LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L3_1_BNROM IS
    PORT (
        coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0); -- Instruction bus
        address : IN unsigned(4 DOWNTO 0));
END L3_1_BNROM;

ARCHITECTURE RTL OF L3_1_BNROM IS

    TYPE ROM_mem IS ARRAY (0 TO 31) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

    CONSTANT ROM_content : ROM_mem :=
    (0=>"0000001011101000"&"0001111000011011",
    1=>"0000000101011000"&"0001010011011100",
    2=>"0000001010111001"&"0001100110000000",
    3=>"0001101100111010"&"0001000000100111",
    4=>"0000011001101001"&"0001010001110001",
    5=>"1111111100110101"&"0001100010100110",
    6=>"0000000101011111"&"0001011001011101",
    7=>"0000101001011110"&"0001010110110110",
    8=>"0000011101001101"&"0001110001001001",
    9=>"0001011100000111"&"0001100001001101",
    10=>"0000001111001011"&"0001011010110100",
    11=>"0000011111111100"&"0001110001111010",
    12=>"0001101011010000"&"0011010001100111",
    13=>"0000010000110100"&"0010101111101001",
    14=>"0000001000100110"&"0001110110100100",
    15=>"0000010110110010"&"0001001000000001",
    16=>"1111110111111011"&"0001100011011001",
    17=>"0000111100101100"&"0001010111011111",
    18=>"0000000111001100"&"0001100011100100",
    19=>"0000001101110011"&"0001101010010010",
    20=>"0000010000111010"&"0010000000011110",
    21=>"1111101110110101"&"0000100101010001",
    22=>"1111111101000111"&"0001110000001000",
    23=>"0000011010010010"&"0001101011000100",
    24=>"0000000101010101"&"0001011111100111",
    25=>"0000101001011001"&"0001100001000000",
    26=>"0000010111100001"&"0001010101110101",
    27=>"0000111001101000"&"0010010101011001",
    28=>"0000100100001000"&"0001010101111100",
    29=>"0001101100111101"&"0001010001111110",
    30=>"0000011000111111"&"0001010101011011",
    31=>"0000001110011100"&"0000110111110000");
    
BEGIN
    coefs <= ROM_content(to_integer(address));
END RTL;