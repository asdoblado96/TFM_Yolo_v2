LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_7_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(8)-1 DOWNTO 0));
END L8_7_WROM;

ARCHITECTURE RTL OF L8_7_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"101000100",
  1=>"001100001",
  2=>"101111011",
  3=>"110000001",
  4=>"001010100",
  5=>"010100100",
  6=>"000011010",
  7=>"101101000",
  8=>"101000000",
  9=>"100011010",
  10=>"100010001",
  11=>"100100001",
  12=>"110111010",
  13=>"000110100",
  14=>"001110010",
  15=>"100011000",
  16=>"111101111",
  17=>"110101101",
  18=>"100110010",
  19=>"111010111",
  20=>"101010111",
  21=>"110000001",
  22=>"111101010",
  23=>"110011101",
  24=>"111001000",
  25=>"110101001",
  26=>"100100001",
  27=>"100110111",
  28=>"101110111",
  29=>"010001011",
  30=>"010010001",
  31=>"001111101",
  32=>"010101001",
  33=>"111010011",
  34=>"100110101",
  35=>"111011010",
  36=>"100111010",
  37=>"000010011",
  38=>"110000000",
  39=>"101001001",
  40=>"100001010",
  41=>"000011110",
  42=>"111110111",
  43=>"100000100",
  44=>"101010001",
  45=>"011001011",
  46=>"111101111",
  47=>"100111100",
  48=>"011111000",
  49=>"011110000",
  50=>"111111111",
  51=>"010111111",
  52=>"011100100",
  53=>"111000111",
  54=>"110111110",
  55=>"111011011",
  56=>"010110011",
  57=>"000000100",
  58=>"001010110",
  59=>"110101010",
  60=>"111101110",
  61=>"111101101",
  62=>"000000110",
  63=>"010000001",
  64=>"111101010",
  65=>"111110001",
  66=>"010100000",
  67=>"111010011",
  68=>"010001000",
  69=>"111010110",
  70=>"111001000",
  71=>"001101011",
  72=>"000101010",
  73=>"101101000",
  74=>"000001000",
  75=>"000111101",
  76=>"110111111",
  77=>"000011100",
  78=>"110010000",
  79=>"101011111",
  80=>"100011110",
  81=>"000000111",
  82=>"000011101",
  83=>"100110101",
  84=>"110000001",
  85=>"000011101",
  86=>"110010011",
  87=>"011101010",
  88=>"100011101",
  89=>"100111010",
  90=>"110001010",
  91=>"000010000",
  92=>"000010001",
  93=>"110000010",
  94=>"100001010",
  95=>"011010111",
  96=>"111110111",
  97=>"010111000",
  98=>"111000010",
  99=>"010010010",
  100=>"110000101",
  101=>"000011001",
  102=>"010100001",
  103=>"010100101",
  104=>"111111101",
  105=>"100011111",
  106=>"010101000",
  107=>"110010000",
  108=>"100101011",
  109=>"010111010",
  110=>"010011111",
  111=>"111111010",
  112=>"110011110",
  113=>"101101101",
  114=>"000010010",
  115=>"010011001",
  116=>"001011000",
  117=>"001101011",
  118=>"010110111",
  119=>"101011000",
  120=>"000011001",
  121=>"101010000",
  122=>"110101110",
  123=>"100101110",
  124=>"110011010",
  125=>"000010101",
  126=>"001011100",
  127=>"100110001",
  128=>"101010100",
  129=>"001000110",
  130=>"101001001",
  131=>"101001001",
  132=>"010100101",
  133=>"111111011",
  134=>"000110100",
  135=>"111101101",
  136=>"100001111",
  137=>"010011010",
  138=>"111011000",
  139=>"010001011",
  140=>"010100100",
  141=>"010111100",
  142=>"000010011",
  143=>"011110010",
  144=>"001110110",
  145=>"100011010",
  146=>"000000101",
  147=>"101001101",
  148=>"001010101",
  149=>"001110111",
  150=>"101101000",
  151=>"111001001",
  152=>"111010011",
  153=>"000111000",
  154=>"000100111",
  155=>"111001111",
  156=>"010100011",
  157=>"010011110",
  158=>"011111100",
  159=>"111011011",
  160=>"101100110",
  161=>"110101111",
  162=>"011001000",
  163=>"010000111",
  164=>"010001001",
  165=>"101011001",
  166=>"100000011",
  167=>"000011010",
  168=>"011010001",
  169=>"101110011",
  170=>"000110010",
  171=>"001111111",
  172=>"101001011",
  173=>"000101010",
  174=>"110111110",
  175=>"000000100",
  176=>"110011110",
  177=>"101110010",
  178=>"111000000",
  179=>"101010000",
  180=>"111100001",
  181=>"101001001",
  182=>"010100001",
  183=>"111101101",
  184=>"100100110",
  185=>"010000010",
  186=>"000111111",
  187=>"000001011",
  188=>"111110111",
  189=>"110101111",
  190=>"000000011",
  191=>"111101000",
  192=>"111001101",
  193=>"011111100",
  194=>"101000111",
  195=>"001100101",
  196=>"000001000",
  197=>"101001111",
  198=>"001100000",
  199=>"111100111",
  200=>"011110011",
  201=>"000011101",
  202=>"000111010",
  203=>"111000001",
  204=>"010111011",
  205=>"111101111",
  206=>"101110111",
  207=>"111000110",
  208=>"001111110",
  209=>"101000101",
  210=>"001101011",
  211=>"101011101",
  212=>"100110000",
  213=>"001010000",
  214=>"111100011",
  215=>"010001011",
  216=>"100111110",
  217=>"010110101",
  218=>"010000100",
  219=>"110000101",
  220=>"000010010",
  221=>"000010100",
  222=>"010000010",
  223=>"111011001",
  224=>"100111000",
  225=>"100001100",
  226=>"000011110",
  227=>"000001001",
  228=>"111010010",
  229=>"011110101",
  230=>"111101010",
  231=>"000000101",
  232=>"101010000",
  233=>"001111010",
  234=>"001101001",
  235=>"000101110",
  236=>"000111001",
  237=>"010000011",
  238=>"010000000",
  239=>"001110000",
  240=>"010110101",
  241=>"001100100",
  242=>"011110101",
  243=>"010000110",
  244=>"011110011",
  245=>"110000001",
  246=>"010000100",
  247=>"101000010",
  248=>"100000100",
  249=>"011000001",
  250=>"011011010",
  251=>"100000100",
  252=>"010101010",
  253=>"100000000",
  254=>"001010010",
  255=>"111000010",
  256=>"101101010",
  257=>"010011000",
  258=>"110001010",
  259=>"001100011",
  260=>"010000011",
  261=>"010011011",
  262=>"001001001",
  263=>"101000111",
  264=>"100110111",
  265=>"011011100",
  266=>"100001000",
  267=>"001110101",
  268=>"010111111",
  269=>"001000110",
  270=>"011101001",
  271=>"101001110",
  272=>"000001100",
  273=>"111000111",
  274=>"100010101",
  275=>"110111011",
  276=>"000000000",
  277=>"000110000",
  278=>"000000001",
  279=>"110101100",
  280=>"110011011",
  281=>"111001111",
  282=>"110111001",
  283=>"100111011",
  284=>"001110111",
  285=>"110010011",
  286=>"010010010",
  287=>"000001100",
  288=>"100011000",
  289=>"001001111",
  290=>"111001000",
  291=>"110000110",
  292=>"000001000",
  293=>"011011101",
  294=>"000001010",
  295=>"101110000",
  296=>"110100110",
  297=>"000111100",
  298=>"100010010",
  299=>"011011110",
  300=>"101001110",
  301=>"010111101",
  302=>"000000011",
  303=>"110010111",
  304=>"001110000",
  305=>"101001110",
  306=>"101111110",
  307=>"010001110",
  308=>"001111111",
  309=>"101111100",
  310=>"011110110",
  311=>"110010110",
  312=>"011001101",
  313=>"000001111",
  314=>"001100101",
  315=>"110100101",
  316=>"010100011",
  317=>"100000111",
  318=>"001110011",
  319=>"111011111",
  320=>"110001011",
  321=>"011111101",
  322=>"011101011",
  323=>"010001000",
  324=>"001110110",
  325=>"010110011",
  326=>"001101000",
  327=>"010011011",
  328=>"101100000",
  329=>"101010111",
  330=>"100101011",
  331=>"000011111",
  332=>"010001010",
  333=>"110010011",
  334=>"010110000",
  335=>"111101100",
  336=>"110101100",
  337=>"001101101",
  338=>"001011111",
  339=>"111010011",
  340=>"010111111",
  341=>"001001111",
  342=>"110001111",
  343=>"000010101",
  344=>"010101100",
  345=>"001010111",
  346=>"110011100",
  347=>"111101100",
  348=>"010001010",
  349=>"100101000",
  350=>"110000000",
  351=>"011010110",
  352=>"011110110",
  353=>"110111001",
  354=>"100101111",
  355=>"111010010",
  356=>"101011010",
  357=>"010010101",
  358=>"111110001",
  359=>"000010000",
  360=>"101010001",
  361=>"101111011",
  362=>"001010000",
  363=>"010110010",
  364=>"111011001",
  365=>"000101101",
  366=>"110010110",
  367=>"011101000",
  368=>"110111111",
  369=>"100000110",
  370=>"001000110",
  371=>"110010010",
  372=>"111100110",
  373=>"010010111",
  374=>"110110010",
  375=>"111100001",
  376=>"001100101",
  377=>"011101001",
  378=>"000110001",
  379=>"101011001",
  380=>"110001010",
  381=>"000100010",
  382=>"000010011",
  383=>"001111101",
  384=>"111000100",
  385=>"100110100",
  386=>"011110111",
  387=>"110101101",
  388=>"000000100",
  389=>"011010110",
  390=>"110101101",
  391=>"010010000",
  392=>"111011000",
  393=>"100101110",
  394=>"010001011",
  395=>"100000111",
  396=>"110100110",
  397=>"110111111",
  398=>"000101100",
  399=>"101111101",
  400=>"011011001",
  401=>"001110000",
  402=>"011101001",
  403=>"111111010",
  404=>"101100000",
  405=>"100000000",
  406=>"011111011",
  407=>"110010101",
  408=>"011010100",
  409=>"100000000",
  410=>"001000101",
  411=>"001100000",
  412=>"111110001",
  413=>"001000100",
  414=>"101101010",
  415=>"010100011",
  416=>"111000101",
  417=>"100000010",
  418=>"100101011",
  419=>"111100001",
  420=>"000000001",
  421=>"010100100",
  422=>"010000111",
  423=>"010100100",
  424=>"011011010",
  425=>"111110100",
  426=>"010110100",
  427=>"000111011",
  428=>"100110100",
  429=>"100001001",
  430=>"101101110",
  431=>"111111011",
  432=>"100100111",
  433=>"111001010",
  434=>"011011100",
  435=>"010001000",
  436=>"101110101",
  437=>"111110000",
  438=>"011001110",
  439=>"100100010",
  440=>"101011111",
  441=>"000000111",
  442=>"000111001",
  443=>"010101001",
  444=>"101100011",
  445=>"010001101",
  446=>"000011111",
  447=>"110111000",
  448=>"101011110",
  449=>"010101100",
  450=>"111101111",
  451=>"111111011",
  452=>"000010100",
  453=>"110001110",
  454=>"111001110",
  455=>"100100010",
  456=>"000001101",
  457=>"001011011",
  458=>"000111110",
  459=>"001100110",
  460=>"000010000",
  461=>"111110011",
  462=>"100100001",
  463=>"101011010",
  464=>"100010110",
  465=>"011111110",
  466=>"101101001",
  467=>"110011011",
  468=>"010111111",
  469=>"111010000",
  470=>"100000111",
  471=>"111000010",
  472=>"011110000",
  473=>"100111000",
  474=>"001011101",
  475=>"001001110",
  476=>"000100110",
  477=>"011110100",
  478=>"110010101",
  479=>"001010110",
  480=>"000011001",
  481=>"001011101",
  482=>"000111101",
  483=>"010100110",
  484=>"001001000",
  485=>"010010011",
  486=>"111011001",
  487=>"111101010",
  488=>"100100001",
  489=>"111010010",
  490=>"110100101",
  491=>"000111010",
  492=>"000001110",
  493=>"100100000",
  494=>"111100110",
  495=>"001101111",
  496=>"000101101",
  497=>"001100101",
  498=>"111001110",
  499=>"101001101",
  500=>"110000010",
  501=>"111010011",
  502=>"010011100",
  503=>"000010010",
  504=>"100011100",
  505=>"010010101",
  506=>"111101110",
  507=>"000100100",
  508=>"000010010",
  509=>"100010011",
  510=>"110010001",
  511=>"101010101",
  512=>"011110110",
  513=>"111010011",
  514=>"100000010",
  515=>"010010001",
  516=>"101111000",
  517=>"110101100",
  518=>"001010111",
  519=>"100111011",
  520=>"101010111",
  521=>"110110001",
  522=>"011011101",
  523=>"110000110",
  524=>"011101111",
  525=>"101111011",
  526=>"001100111",
  527=>"010011000",
  528=>"100000011",
  529=>"011111110",
  530=>"010010001",
  531=>"000001011",
  532=>"000000100",
  533=>"101001010",
  534=>"110011101",
  535=>"001111010",
  536=>"011001011",
  537=>"101001111",
  538=>"011011010",
  539=>"100001111",
  540=>"100110001",
  541=>"011101001",
  542=>"111001000",
  543=>"000100110",
  544=>"000000010",
  545=>"100000100",
  546=>"011010110",
  547=>"111000001",
  548=>"010001011",
  549=>"000110111",
  550=>"101011001",
  551=>"111101110",
  552=>"001000000",
  553=>"001001001",
  554=>"001110110",
  555=>"100100111",
  556=>"010001011",
  557=>"011010011",
  558=>"100011000",
  559=>"000000001",
  560=>"111010011",
  561=>"000011110",
  562=>"011001101",
  563=>"000111001",
  564=>"101011010",
  565=>"101011111",
  566=>"110011011",
  567=>"111001111",
  568=>"000000000",
  569=>"001111000",
  570=>"100101000",
  571=>"010100000",
  572=>"011101011",
  573=>"011011111",
  574=>"011101001",
  575=>"100010100",
  576=>"111111101",
  577=>"110100100",
  578=>"111101000",
  579=>"011110100",
  580=>"111011000",
  581=>"011110000",
  582=>"000100101",
  583=>"000110111",
  584=>"000101000",
  585=>"101100100",
  586=>"101101000",
  587=>"010000100",
  588=>"001100111",
  589=>"101011100",
  590=>"000110011",
  591=>"101010110",
  592=>"100011010",
  593=>"110101001",
  594=>"001000001",
  595=>"000001010",
  596=>"110100001",
  597=>"001010101",
  598=>"001110010",
  599=>"111011110",
  600=>"101100110",
  601=>"110010111",
  602=>"000010000",
  603=>"001000111",
  604=>"111010010",
  605=>"011011101",
  606=>"010010001",
  607=>"000100001",
  608=>"001100011",
  609=>"000001010",
  610=>"111101011",
  611=>"011101010",
  612=>"001000001",
  613=>"010100100",
  614=>"100000111",
  615=>"000000011",
  616=>"000100010",
  617=>"010000101",
  618=>"111001010",
  619=>"100110000",
  620=>"000010100",
  621=>"010100000",
  622=>"110011111",
  623=>"101010100",
  624=>"111010111",
  625=>"010111111",
  626=>"110101111",
  627=>"001000001",
  628=>"000101111",
  629=>"111101100",
  630=>"001110000",
  631=>"101000000",
  632=>"110011001",
  633=>"011011010",
  634=>"001101111",
  635=>"100000011",
  636=>"000101110",
  637=>"110000111",
  638=>"110000111",
  639=>"111111110",
  640=>"011101111",
  641=>"101110101",
  642=>"010001101",
  643=>"000011010",
  644=>"101100011",
  645=>"010100011",
  646=>"011100010",
  647=>"011010010",
  648=>"010010010",
  649=>"010111111",
  650=>"100100111",
  651=>"100001001",
  652=>"111001101",
  653=>"010110011",
  654=>"000000111",
  655=>"100111000",
  656=>"100110111",
  657=>"111101111",
  658=>"010001001",
  659=>"000001110",
  660=>"111001000",
  661=>"011101001",
  662=>"110111101",
  663=>"111000001",
  664=>"101001100",
  665=>"100001011",
  666=>"001100110",
  667=>"111110010",
  668=>"111100110",
  669=>"100101001",
  670=>"010110110",
  671=>"100011100",
  672=>"110001011",
  673=>"100110010",
  674=>"101110110",
  675=>"101000000",
  676=>"100100100",
  677=>"010001010",
  678=>"110100101",
  679=>"001100010",
  680=>"111111001",
  681=>"101101100",
  682=>"000011010",
  683=>"000111101",
  684=>"001101101",
  685=>"001111111",
  686=>"011101110",
  687=>"001000000",
  688=>"001101011",
  689=>"110001011",
  690=>"111010000",
  691=>"111101110",
  692=>"100001011",
  693=>"011011100",
  694=>"011011100",
  695=>"001111110",
  696=>"000000000",
  697=>"111011000",
  698=>"110000000",
  699=>"111000010",
  700=>"010000010",
  701=>"100010000",
  702=>"000100000",
  703=>"011001010",
  704=>"010100110",
  705=>"010101111",
  706=>"100011001",
  707=>"100110001",
  708=>"000000110",
  709=>"000000010",
  710=>"011011110",
  711=>"011011100",
  712=>"101010011",
  713=>"001011110",
  714=>"001110110",
  715=>"001101110",
  716=>"100101100",
  717=>"101110110",
  718=>"011000010",
  719=>"101001111",
  720=>"010000010",
  721=>"101101101",
  722=>"101111101",
  723=>"011000110",
  724=>"100111110",
  725=>"010000100",
  726=>"000000110",
  727=>"111001111",
  728=>"010011010",
  729=>"110111001",
  730=>"111110010",
  731=>"000001111",
  732=>"111110110",
  733=>"111110101",
  734=>"110011010",
  735=>"011101011",
  736=>"010101001",
  737=>"000111001",
  738=>"001100101",
  739=>"100010010",
  740=>"000000000",
  741=>"011001101",
  742=>"010111111",
  743=>"110110011",
  744=>"111000101",
  745=>"101110011",
  746=>"101010001",
  747=>"110000011",
  748=>"101000001",
  749=>"000100001",
  750=>"110011100",
  751=>"111101111",
  752=>"010111111",
  753=>"011101010",
  754=>"100111011",
  755=>"110111111",
  756=>"100001100",
  757=>"011110100",
  758=>"111101100",
  759=>"011010010",
  760=>"010000001",
  761=>"010110110",
  762=>"001111111",
  763=>"011011100",
  764=>"110110111",
  765=>"100001000",
  766=>"010010100",
  767=>"010001101",
  768=>"010010001",
  769=>"011111111",
  770=>"011000011",
  771=>"101111010",
  772=>"101000000",
  773=>"001101101",
  774=>"010000010",
  775=>"101110001",
  776=>"001111110",
  777=>"111110010",
  778=>"110110111",
  779=>"111011101",
  780=>"110101001",
  781=>"000010010",
  782=>"001010001",
  783=>"111011101",
  784=>"101000000",
  785=>"111101101",
  786=>"111001000",
  787=>"111111000",
  788=>"011010011",
  789=>"001011110",
  790=>"111111011",
  791=>"101100010",
  792=>"101101001",
  793=>"001010011",
  794=>"110110110",
  795=>"000000011",
  796=>"010100100",
  797=>"100000001",
  798=>"001100000",
  799=>"100000000",
  800=>"011011010",
  801=>"100001001",
  802=>"001010001",
  803=>"100110011",
  804=>"111001111",
  805=>"011000010",
  806=>"101001100",
  807=>"010111011",
  808=>"000110101",
  809=>"011010110",
  810=>"111011010",
  811=>"000000000",
  812=>"100000100",
  813=>"011010110",
  814=>"101001000",
  815=>"111111111",
  816=>"110000111",
  817=>"001001101",
  818=>"100010111",
  819=>"000110100",
  820=>"111001110",
  821=>"010101011",
  822=>"011100011",
  823=>"111111100",
  824=>"111100101",
  825=>"000110100",
  826=>"111101100",
  827=>"110100010",
  828=>"110000111",
  829=>"110111101",
  830=>"001111111",
  831=>"001100110",
  832=>"000000001",
  833=>"110000010",
  834=>"010001101",
  835=>"000001101",
  836=>"101101010",
  837=>"110011001",
  838=>"010100011",
  839=>"001010000",
  840=>"000000001",
  841=>"011011011",
  842=>"101000011",
  843=>"100001101",
  844=>"101001011",
  845=>"010011100",
  846=>"011101100",
  847=>"111010110",
  848=>"100000000",
  849=>"001010010",
  850=>"001011111",
  851=>"111000111",
  852=>"100011010",
  853=>"111010100",
  854=>"000000011",
  855=>"101011101",
  856=>"000000001",
  857=>"100010101",
  858=>"101111011",
  859=>"000111001",
  860=>"010011010",
  861=>"100001100",
  862=>"110001100",
  863=>"000000111",
  864=>"001100011",
  865=>"111001111",
  866=>"110010101",
  867=>"111001100",
  868=>"101000011",
  869=>"101100101",
  870=>"010010101",
  871=>"100100000",
  872=>"110111101",
  873=>"110000101",
  874=>"000010000",
  875=>"010011000",
  876=>"001100001",
  877=>"000000111",
  878=>"110000001",
  879=>"001001000",
  880=>"011101111",
  881=>"100111111",
  882=>"000101111",
  883=>"010010110",
  884=>"111011001",
  885=>"000001001",
  886=>"110010100",
  887=>"100001011",
  888=>"101100010",
  889=>"110100010",
  890=>"110010000",
  891=>"000100011",
  892=>"000011110",
  893=>"100110010",
  894=>"000100110",
  895=>"000110110",
  896=>"101000001",
  897=>"101101100",
  898=>"001100111",
  899=>"101100100",
  900=>"111101101",
  901=>"100100010",
  902=>"001000000",
  903=>"001101000",
  904=>"100010000",
  905=>"110101100",
  906=>"011011001",
  907=>"111101111",
  908=>"001000011",
  909=>"010011001",
  910=>"110111011",
  911=>"001111011",
  912=>"011111000",
  913=>"010111001",
  914=>"110111001",
  915=>"010111111",
  916=>"100000001",
  917=>"001010100",
  918=>"111010110",
  919=>"011100000",
  920=>"010111101",
  921=>"000000011",
  922=>"111010011",
  923=>"011101001",
  924=>"000001100",
  925=>"110111111",
  926=>"110010000",
  927=>"111111000",
  928=>"010111000",
  929=>"000110101",
  930=>"110000100",
  931=>"000110101",
  932=>"111011101",
  933=>"111111001",
  934=>"000010100",
  935=>"101100011",
  936=>"101101111",
  937=>"111101011",
  938=>"101110011",
  939=>"010010100",
  940=>"110010110",
  941=>"111000100",
  942=>"001010100",
  943=>"100001000",
  944=>"010110101",
  945=>"100111100",
  946=>"110110001",
  947=>"011111010",
  948=>"011100000",
  949=>"011011010",
  950=>"110111111",
  951=>"011010001",
  952=>"111011101",
  953=>"100011100",
  954=>"111010101",
  955=>"110001001",
  956=>"111010100",
  957=>"011100001",
  958=>"100111000",
  959=>"001101001",
  960=>"001100001",
  961=>"010010010",
  962=>"010110100",
  963=>"001001000",
  964=>"101101010",
  965=>"100100101",
  966=>"010101100",
  967=>"110000111",
  968=>"111001100",
  969=>"110100010",
  970=>"111100001",
  971=>"110110011",
  972=>"001001111",
  973=>"111111011",
  974=>"100010001",
  975=>"101000110",
  976=>"011001010",
  977=>"010101010",
  978=>"111111010",
  979=>"010000010",
  980=>"101111111",
  981=>"011001000",
  982=>"001110011",
  983=>"100111110",
  984=>"101001100",
  985=>"100010101",
  986=>"001111011",
  987=>"101011010",
  988=>"111011011",
  989=>"011010001",
  990=>"111011111",
  991=>"101010011",
  992=>"101110110",
  993=>"111101010",
  994=>"001010111",
  995=>"111110010",
  996=>"101011101",
  997=>"100000011",
  998=>"001010000",
  999=>"010001110",
  1000=>"000010010",
  1001=>"001000111",
  1002=>"010001100",
  1003=>"001000111",
  1004=>"010010011",
  1005=>"010001101",
  1006=>"100111011",
  1007=>"110001001",
  1008=>"111101111",
  1009=>"100110001",
  1010=>"111011100",
  1011=>"100001010",
  1012=>"110001101",
  1013=>"001011100",
  1014=>"111010100",
  1015=>"001000111",
  1016=>"001100100",
  1017=>"000110111",
  1018=>"100100111",
  1019=>"100111101",
  1020=>"100101000",
  1021=>"100010111",
  1022=>"101110101",
  1023=>"011000111",
  1024=>"010100101",
  1025=>"011011100",
  1026=>"100010011",
  1027=>"110110111",
  1028=>"000010100",
  1029=>"100000010",
  1030=>"010001100",
  1031=>"000001000",
  1032=>"101110010",
  1033=>"101110111",
  1034=>"101011000",
  1035=>"010111100",
  1036=>"100101100",
  1037=>"111111111",
  1038=>"111111010",
  1039=>"100101100",
  1040=>"010110011",
  1041=>"100010010",
  1042=>"100101001",
  1043=>"001011101",
  1044=>"100100110",
  1045=>"010010010",
  1046=>"001110100",
  1047=>"010111001",
  1048=>"101111100",
  1049=>"011110000",
  1050=>"111100000",
  1051=>"100110001",
  1052=>"010011010",
  1053=>"011111001",
  1054=>"110111100",
  1055=>"010011101",
  1056=>"000111001",
  1057=>"101100111",
  1058=>"011101011",
  1059=>"100100110",
  1060=>"111011110",
  1061=>"001111010",
  1062=>"000100000",
  1063=>"110110011",
  1064=>"001010100",
  1065=>"101101100",
  1066=>"100000101",
  1067=>"110011010",
  1068=>"011001001",
  1069=>"110111001",
  1070=>"000011110",
  1071=>"011000111",
  1072=>"000001101",
  1073=>"100100000",
  1074=>"110001010",
  1075=>"101100101",
  1076=>"111010100",
  1077=>"011011011",
  1078=>"001100011",
  1079=>"111000001",
  1080=>"000000111",
  1081=>"101110000",
  1082=>"001100011",
  1083=>"110110101",
  1084=>"010010101",
  1085=>"000010110",
  1086=>"011100111",
  1087=>"011101000",
  1088=>"100000000",
  1089=>"000000000",
  1090=>"100000010",
  1091=>"100001011",
  1092=>"100000101",
  1093=>"011100110",
  1094=>"010100001",
  1095=>"111110111",
  1096=>"010000011",
  1097=>"000111101",
  1098=>"111101111",
  1099=>"000110101",
  1100=>"010110000",
  1101=>"100001010",
  1102=>"101011100",
  1103=>"101110101",
  1104=>"000000100",
  1105=>"111101011",
  1106=>"000001000",
  1107=>"001010010",
  1108=>"000011010",
  1109=>"001001111",
  1110=>"000101000",
  1111=>"001101101",
  1112=>"101101011",
  1113=>"101101000",
  1114=>"000010111",
  1115=>"110111001",
  1116=>"000000101",
  1117=>"101111010",
  1118=>"011000001",
  1119=>"100000101",
  1120=>"111010001",
  1121=>"101000000",
  1122=>"111111110",
  1123=>"110100111",
  1124=>"010011000",
  1125=>"111101110",
  1126=>"100101010",
  1127=>"000110101",
  1128=>"000111010",
  1129=>"011000100",
  1130=>"000110101",
  1131=>"111101011",
  1132=>"000000011",
  1133=>"001110111",
  1134=>"100000000",
  1135=>"001001010",
  1136=>"111100001",
  1137=>"100111100",
  1138=>"111111110",
  1139=>"100100110",
  1140=>"101010111",
  1141=>"000001000",
  1142=>"110011001",
  1143=>"001111001",
  1144=>"100010101",
  1145=>"011101011",
  1146=>"111100111",
  1147=>"011111000",
  1148=>"011000001",
  1149=>"100000111",
  1150=>"000000000",
  1151=>"011101101",
  1152=>"101000000",
  1153=>"010001100",
  1154=>"001100111",
  1155=>"010001000",
  1156=>"000110000",
  1157=>"001001000",
  1158=>"110001100",
  1159=>"010110001",
  1160=>"110110001",
  1161=>"011111111",
  1162=>"000011000",
  1163=>"001001111",
  1164=>"100000010",
  1165=>"100010100",
  1166=>"110111100",
  1167=>"100110111",
  1168=>"011110100",
  1169=>"111101010",
  1170=>"011011111",
  1171=>"010010110",
  1172=>"010000110",
  1173=>"011001100",
  1174=>"111000000",
  1175=>"110111111",
  1176=>"100001111",
  1177=>"101110111",
  1178=>"000110111",
  1179=>"000011010",
  1180=>"111000010",
  1181=>"100110100",
  1182=>"100111000",
  1183=>"100001011",
  1184=>"011100110",
  1185=>"010111101",
  1186=>"100000011",
  1187=>"110101110",
  1188=>"011011110",
  1189=>"110000111",
  1190=>"010111110",
  1191=>"111110100",
  1192=>"011000011",
  1193=>"111110011",
  1194=>"011010100",
  1195=>"110100000",
  1196=>"111110101",
  1197=>"100111011",
  1198=>"110010110",
  1199=>"100110001",
  1200=>"100011110",
  1201=>"111010111",
  1202=>"001111011",
  1203=>"000110001",
  1204=>"100110110",
  1205=>"110011011",
  1206=>"101100101",
  1207=>"010000110",
  1208=>"100011110",
  1209=>"011011000",
  1210=>"011110110",
  1211=>"000001011",
  1212=>"110010100",
  1213=>"101100001",
  1214=>"100101111",
  1215=>"010110000",
  1216=>"000011001",
  1217=>"111100010",
  1218=>"100100010",
  1219=>"010000010",
  1220=>"001100100",
  1221=>"010010110",
  1222=>"010000101",
  1223=>"010001001",
  1224=>"100000110",
  1225=>"111001001",
  1226=>"010010100",
  1227=>"110010100",
  1228=>"010010000",
  1229=>"011101100",
  1230=>"001001111",
  1231=>"111111100",
  1232=>"110111111",
  1233=>"101000111",
  1234=>"000000110",
  1235=>"110000101",
  1236=>"010111101",
  1237=>"111101000",
  1238=>"001110011",
  1239=>"010101101",
  1240=>"011111001",
  1241=>"100010101",
  1242=>"011101001",
  1243=>"101101010",
  1244=>"011011001",
  1245=>"000000101",
  1246=>"000000011",
  1247=>"111010010",
  1248=>"010000100",
  1249=>"111100111",
  1250=>"111011111",
  1251=>"000000110",
  1252=>"011111101",
  1253=>"011101000",
  1254=>"010111010",
  1255=>"000101000",
  1256=>"101000001",
  1257=>"111111111",
  1258=>"010010011",
  1259=>"000100010",
  1260=>"111100111",
  1261=>"111110101",
  1262=>"000101100",
  1263=>"001111011",
  1264=>"011001111",
  1265=>"111011111",
  1266=>"001011000",
  1267=>"010010110",
  1268=>"100111110",
  1269=>"011100000",
  1270=>"011100001",
  1271=>"110000000",
  1272=>"011101001",
  1273=>"000111011",
  1274=>"101011110",
  1275=>"001000010",
  1276=>"100111111",
  1277=>"000001011",
  1278=>"000010101",
  1279=>"110111000",
  1280=>"011110001",
  1281=>"110010000",
  1282=>"110000101",
  1283=>"001101100",
  1284=>"100111111",
  1285=>"101110100",
  1286=>"001001000",
  1287=>"100011100",
  1288=>"000001111",
  1289=>"011110001",
  1290=>"001010100",
  1291=>"010101000",
  1292=>"110010001",
  1293=>"001011000",
  1294=>"000011100",
  1295=>"111011100",
  1296=>"111100001",
  1297=>"000010001",
  1298=>"000000111",
  1299=>"001011101",
  1300=>"011100010",
  1301=>"011011011",
  1302=>"110000100",
  1303=>"011101101",
  1304=>"000010010",
  1305=>"100111011",
  1306=>"111101101",
  1307=>"011000111",
  1308=>"100100001",
  1309=>"101101001",
  1310=>"011001101",
  1311=>"010000100",
  1312=>"111000110",
  1313=>"100000010",
  1314=>"111110001",
  1315=>"010000001",
  1316=>"100111000",
  1317=>"101100011",
  1318=>"011001111",
  1319=>"100010110",
  1320=>"000111000",
  1321=>"100000100",
  1322=>"010000010",
  1323=>"101111000",
  1324=>"110100101",
  1325=>"000100001",
  1326=>"000011011",
  1327=>"000100111",
  1328=>"001010111",
  1329=>"110101010",
  1330=>"010101001",
  1331=>"000111111",
  1332=>"100000110",
  1333=>"001001001",
  1334=>"000111110",
  1335=>"100000000",
  1336=>"101011111",
  1337=>"100100110",
  1338=>"111100010",
  1339=>"111000101",
  1340=>"001010000",
  1341=>"100100101",
  1342=>"101011010",
  1343=>"000001101",
  1344=>"110011100",
  1345=>"110000100",
  1346=>"100001111",
  1347=>"110001010",
  1348=>"000000111",
  1349=>"010110111",
  1350=>"000010011",
  1351=>"011001010",
  1352=>"001001010",
  1353=>"101001010",
  1354=>"101001001",
  1355=>"000010000",
  1356=>"111100011",
  1357=>"010000010",
  1358=>"111110101",
  1359=>"111110111",
  1360=>"100011110",
  1361=>"101001111",
  1362=>"111100010",
  1363=>"101110101",
  1364=>"110100110",
  1365=>"010001001",
  1366=>"010111010",
  1367=>"000111110",
  1368=>"000011000",
  1369=>"001000010",
  1370=>"001000101",
  1371=>"100001111",
  1372=>"001101100",
  1373=>"110100001",
  1374=>"000010100",
  1375=>"000010111",
  1376=>"000110100",
  1377=>"101111111",
  1378=>"101100110",
  1379=>"000111000",
  1380=>"000000110",
  1381=>"110110010",
  1382=>"111010110",
  1383=>"100011010",
  1384=>"110011000",
  1385=>"000011101",
  1386=>"000010110",
  1387=>"111100110",
  1388=>"001110110",
  1389=>"110011101",
  1390=>"110100101",
  1391=>"111101000",
  1392=>"000111101",
  1393=>"111011010",
  1394=>"111000111",
  1395=>"101110111",
  1396=>"000011111",
  1397=>"000010000",
  1398=>"000000000",
  1399=>"111001000",
  1400=>"110011101",
  1401=>"100011001",
  1402=>"110101010",
  1403=>"110001100",
  1404=>"001010100",
  1405=>"111111101",
  1406=>"010111000",
  1407=>"100000000",
  1408=>"011100010",
  1409=>"001011000",
  1410=>"100011101",
  1411=>"101111100",
  1412=>"100010010",
  1413=>"110011001",
  1414=>"011100101",
  1415=>"011010110",
  1416=>"010001011",
  1417=>"111111110",
  1418=>"100000011",
  1419=>"101101110",
  1420=>"111110111",
  1421=>"100100011",
  1422=>"101100000",
  1423=>"100001000",
  1424=>"010111001",
  1425=>"001000001",
  1426=>"111000110",
  1427=>"010100011",
  1428=>"100111100",
  1429=>"100110101",
  1430=>"111100110",
  1431=>"010000001",
  1432=>"011110110",
  1433=>"010111011",
  1434=>"111111010",
  1435=>"101100010",
  1436=>"100111010",
  1437=>"111101000",
  1438=>"010000000",
  1439=>"110110010",
  1440=>"101101101",
  1441=>"000110100",
  1442=>"101011100",
  1443=>"000000001",
  1444=>"110001101",
  1445=>"111010001",
  1446=>"010000011",
  1447=>"001010001",
  1448=>"011111011",
  1449=>"011011000",
  1450=>"111101001",
  1451=>"111010001",
  1452=>"111010111",
  1453=>"000010000",
  1454=>"011011011",
  1455=>"110111011",
  1456=>"011001110",
  1457=>"101100111",
  1458=>"010100011",
  1459=>"011101001",
  1460=>"101010111",
  1461=>"000100100",
  1462=>"000110010",
  1463=>"111011001",
  1464=>"110011001",
  1465=>"001100011",
  1466=>"010100100",
  1467=>"110000101",
  1468=>"001011111",
  1469=>"011100010",
  1470=>"011101111",
  1471=>"000010100",
  1472=>"100100000",
  1473=>"100111100",
  1474=>"101110110",
  1475=>"111000101",
  1476=>"101000010",
  1477=>"000000100",
  1478=>"001010111",
  1479=>"000111101",
  1480=>"101011111",
  1481=>"010010000",
  1482=>"001100111",
  1483=>"110010011",
  1484=>"100111011",
  1485=>"111100100",
  1486=>"111101001",
  1487=>"111000100",
  1488=>"110100011",
  1489=>"110110111",
  1490=>"011000111",
  1491=>"101010101",
  1492=>"000111110",
  1493=>"100001010",
  1494=>"001111100",
  1495=>"111010111",
  1496=>"110111100",
  1497=>"001100000",
  1498=>"110111101",
  1499=>"100110001",
  1500=>"100001010",
  1501=>"000000110",
  1502=>"000010011",
  1503=>"010001111",
  1504=>"011101000",
  1505=>"011101001",
  1506=>"010111111",
  1507=>"010101011",
  1508=>"100110110",
  1509=>"001111001",
  1510=>"111010000",
  1511=>"010000000",
  1512=>"110101010",
  1513=>"010011000",
  1514=>"100111001",
  1515=>"111110000",
  1516=>"000101111",
  1517=>"011100010",
  1518=>"000111111",
  1519=>"110110000",
  1520=>"101000100",
  1521=>"010010001",
  1522=>"101000011",
  1523=>"001011100",
  1524=>"001000000",
  1525=>"110001110",
  1526=>"011100111",
  1527=>"110010010",
  1528=>"101110001",
  1529=>"001001001",
  1530=>"000010000",
  1531=>"011100001",
  1532=>"001101011",
  1533=>"101011010",
  1534=>"111100110",
  1535=>"111001001",
  1536=>"110111010",
  1537=>"111000101",
  1538=>"111001011",
  1539=>"001101101",
  1540=>"000000001",
  1541=>"100110001",
  1542=>"110010011",
  1543=>"110111011",
  1544=>"011101000",
  1545=>"111001010",
  1546=>"011010010",
  1547=>"111010110",
  1548=>"011100101",
  1549=>"000001011",
  1550=>"111000101",
  1551=>"010000001",
  1552=>"011010000",
  1553=>"001110010",
  1554=>"011101100",
  1555=>"100011001",
  1556=>"010110101",
  1557=>"011010000",
  1558=>"001110101",
  1559=>"011000011",
  1560=>"110111000",
  1561=>"000001001",
  1562=>"111100001",
  1563=>"011000011",
  1564=>"110001110",
  1565=>"001001101",
  1566=>"110011001",
  1567=>"110100111",
  1568=>"111110110",
  1569=>"011100100",
  1570=>"000000101",
  1571=>"110001011",
  1572=>"100001110",
  1573=>"010011110",
  1574=>"010000101",
  1575=>"010110000",
  1576=>"010000101",
  1577=>"011000100",
  1578=>"111000100",
  1579=>"010110100",
  1580=>"001010110",
  1581=>"111111001",
  1582=>"110100011",
  1583=>"011110111",
  1584=>"011100010",
  1585=>"000011101",
  1586=>"000110100",
  1587=>"100011110",
  1588=>"101001110",
  1589=>"001011110",
  1590=>"000011000",
  1591=>"011011000",
  1592=>"000111110",
  1593=>"011000110",
  1594=>"101100011",
  1595=>"111000010",
  1596=>"110111100",
  1597=>"000000101",
  1598=>"101110100",
  1599=>"100010000",
  1600=>"000111110",
  1601=>"010111011",
  1602=>"101001100",
  1603=>"111100011",
  1604=>"110010011",
  1605=>"100000111",
  1606=>"000001010",
  1607=>"001000000",
  1608=>"100000000",
  1609=>"111000000",
  1610=>"011000000",
  1611=>"101011000",
  1612=>"111111101",
  1613=>"101100100",
  1614=>"100001111",
  1615=>"111101010",
  1616=>"111101111",
  1617=>"011010011",
  1618=>"110001011",
  1619=>"111000101",
  1620=>"110000011",
  1621=>"100000010",
  1622=>"110011010",
  1623=>"010101010",
  1624=>"001111100",
  1625=>"000101101",
  1626=>"101110111",
  1627=>"110000100",
  1628=>"000101110",
  1629=>"100000010",
  1630=>"010110010",
  1631=>"010100110",
  1632=>"011000011",
  1633=>"111101101",
  1634=>"110000110",
  1635=>"110010011",
  1636=>"100010111",
  1637=>"101101011",
  1638=>"000101011",
  1639=>"010110110",
  1640=>"000100111",
  1641=>"000110001",
  1642=>"100100000",
  1643=>"100101111",
  1644=>"000111100",
  1645=>"000101000",
  1646=>"000110010",
  1647=>"110011101",
  1648=>"111000011",
  1649=>"000011011",
  1650=>"000101100",
  1651=>"101001001",
  1652=>"111111101",
  1653=>"100000101",
  1654=>"111101110",
  1655=>"001110110",
  1656=>"111001000",
  1657=>"101100101",
  1658=>"110000100",
  1659=>"011000101",
  1660=>"010100111",
  1661=>"110010000",
  1662=>"101011100",
  1663=>"010000000",
  1664=>"111111000",
  1665=>"010011110",
  1666=>"110100001",
  1667=>"010111010",
  1668=>"100011111",
  1669=>"110100010",
  1670=>"001001001",
  1671=>"010011011",
  1672=>"110010010",
  1673=>"010111111",
  1674=>"110000101",
  1675=>"101001110",
  1676=>"011111110",
  1677=>"000000000",
  1678=>"111001011",
  1679=>"111011000",
  1680=>"100110101",
  1681=>"111110011",
  1682=>"000000101",
  1683=>"010100100",
  1684=>"010111000",
  1685=>"110110100",
  1686=>"100101100",
  1687=>"010010011",
  1688=>"100001011",
  1689=>"011111001",
  1690=>"011011011",
  1691=>"001010001",
  1692=>"100111100",
  1693=>"110111000",
  1694=>"111111011",
  1695=>"111111101",
  1696=>"101111101",
  1697=>"110001010",
  1698=>"000010011",
  1699=>"011110100",
  1700=>"010110110",
  1701=>"101111101",
  1702=>"101100111",
  1703=>"111111000",
  1704=>"111101000",
  1705=>"010110001",
  1706=>"111110110",
  1707=>"011100001",
  1708=>"011111111",
  1709=>"000000111",
  1710=>"111100101",
  1711=>"011000010",
  1712=>"010110010",
  1713=>"010110000",
  1714=>"100111001",
  1715=>"101100101",
  1716=>"001001100",
  1717=>"111100111",
  1718=>"011110000",
  1719=>"001001000",
  1720=>"100111011",
  1721=>"001011001",
  1722=>"000110010",
  1723=>"101111101",
  1724=>"001001111",
  1725=>"111000111",
  1726=>"100001100",
  1727=>"100110001",
  1728=>"101010011",
  1729=>"011011110",
  1730=>"010100100",
  1731=>"101101110",
  1732=>"011000001",
  1733=>"010000000",
  1734=>"111110000",
  1735=>"101101111",
  1736=>"000100001",
  1737=>"011101101",
  1738=>"001110100",
  1739=>"010010111",
  1740=>"100001100",
  1741=>"010111000",
  1742=>"001110100",
  1743=>"010000111",
  1744=>"111111001",
  1745=>"101110001",
  1746=>"001111100",
  1747=>"101011011",
  1748=>"001100111",
  1749=>"010101101",
  1750=>"110010101",
  1751=>"010000100",
  1752=>"101101000",
  1753=>"010001011",
  1754=>"101111011",
  1755=>"010110101",
  1756=>"011010001",
  1757=>"001001001",
  1758=>"101110100",
  1759=>"111000100",
  1760=>"111101000",
  1761=>"001100111",
  1762=>"101101101",
  1763=>"110110100",
  1764=>"001110100",
  1765=>"111110000",
  1766=>"010000000",
  1767=>"001011010",
  1768=>"010100011",
  1769=>"000010001",
  1770=>"100001111",
  1771=>"110101100",
  1772=>"011000111",
  1773=>"101010110",
  1774=>"010101010",
  1775=>"100010001",
  1776=>"011100111",
  1777=>"011010111",
  1778=>"010011011",
  1779=>"111100001",
  1780=>"100100000",
  1781=>"101001011",
  1782=>"011101011",
  1783=>"100010000",
  1784=>"011000000",
  1785=>"010001010",
  1786=>"100101010",
  1787=>"010101110",
  1788=>"111001001",
  1789=>"000001111",
  1790=>"010000010",
  1791=>"110110110",
  1792=>"111001111",
  1793=>"001111011",
  1794=>"011111010",
  1795=>"000100001",
  1796=>"001001101",
  1797=>"110000010",
  1798=>"010000100",
  1799=>"110110011",
  1800=>"000101111",
  1801=>"010110100",
  1802=>"001110101",
  1803=>"001100101",
  1804=>"000000000",
  1805=>"010100010",
  1806=>"110111000",
  1807=>"000010010",
  1808=>"001001001",
  1809=>"111100010",
  1810=>"000111111",
  1811=>"110100001",
  1812=>"110111010",
  1813=>"010101000",
  1814=>"010111001",
  1815=>"000000011",
  1816=>"101001101",
  1817=>"110010010",
  1818=>"010010000",
  1819=>"000000101",
  1820=>"110011111",
  1821=>"000001101",
  1822=>"111101011",
  1823=>"000001000",
  1824=>"101001100",
  1825=>"010010000",
  1826=>"011010010",
  1827=>"010111111",
  1828=>"001011011",
  1829=>"111101101",
  1830=>"100010100",
  1831=>"110011010",
  1832=>"001011001",
  1833=>"000000000",
  1834=>"011110001",
  1835=>"101111101",
  1836=>"000001110",
  1837=>"001011101",
  1838=>"101100111",
  1839=>"001110000",
  1840=>"110000101",
  1841=>"100001011",
  1842=>"001000000",
  1843=>"101000001",
  1844=>"111111111",
  1845=>"011010001",
  1846=>"011101000",
  1847=>"111101001",
  1848=>"110010111",
  1849=>"111101011",
  1850=>"000001001",
  1851=>"000111001",
  1852=>"110100111",
  1853=>"101101010",
  1854=>"010000011",
  1855=>"101001110",
  1856=>"010010001",
  1857=>"111110010",
  1858=>"110111101",
  1859=>"110111111",
  1860=>"100011000",
  1861=>"110010000",
  1862=>"111000110",
  1863=>"101111001",
  1864=>"101000110",
  1865=>"100001101",
  1866=>"000000010",
  1867=>"100001011",
  1868=>"100100100",
  1869=>"001000010",
  1870=>"001000101",
  1871=>"110010010",
  1872=>"101001100",
  1873=>"001101100",
  1874=>"011101100",
  1875=>"001010100",
  1876=>"101110010",
  1877=>"000010001",
  1878=>"101001011",
  1879=>"011110000",
  1880=>"111010101",
  1881=>"011001101",
  1882=>"011100111",
  1883=>"100100001",
  1884=>"100001101",
  1885=>"100001001",
  1886=>"001010010",
  1887=>"101000111",
  1888=>"010001110",
  1889=>"110111111",
  1890=>"000110011",
  1891=>"101010110",
  1892=>"111101001",
  1893=>"100101111",
  1894=>"010110100",
  1895=>"110001001",
  1896=>"100001101",
  1897=>"101100011",
  1898=>"001101100",
  1899=>"010110111",
  1900=>"110110110",
  1901=>"000111000",
  1902=>"001000001",
  1903=>"101011000",
  1904=>"001100000",
  1905=>"111101110",
  1906=>"001011001",
  1907=>"110010111",
  1908=>"111101111",
  1909=>"000001111",
  1910=>"111001001",
  1911=>"100001111",
  1912=>"001010101",
  1913=>"000110001",
  1914=>"011010000",
  1915=>"110111010",
  1916=>"111001111",
  1917=>"101011010",
  1918=>"010000000",
  1919=>"011100000",
  1920=>"110001100",
  1921=>"000100011",
  1922=>"000011001",
  1923=>"000111010",
  1924=>"110001010",
  1925=>"110001010",
  1926=>"000000011",
  1927=>"010110100",
  1928=>"111101111",
  1929=>"100110010",
  1930=>"000110011",
  1931=>"111111111",
  1932=>"010001100",
  1933=>"111011110",
  1934=>"100111111",
  1935=>"000100111",
  1936=>"101110100",
  1937=>"111010010",
  1938=>"000000101",
  1939=>"000100000",
  1940=>"011010111",
  1941=>"101110111",
  1942=>"111011110",
  1943=>"100010101",
  1944=>"011001100",
  1945=>"011001111",
  1946=>"101111101",
  1947=>"100011110",
  1948=>"101000001",
  1949=>"001101111",
  1950=>"011001000",
  1951=>"001011010",
  1952=>"101101010",
  1953=>"010101001",
  1954=>"010010101",
  1955=>"111101000",
  1956=>"010011000",
  1957=>"011101010",
  1958=>"011101111",
  1959=>"101100000",
  1960=>"100010111",
  1961=>"100011001",
  1962=>"111101000",
  1963=>"100100001",
  1964=>"110111101",
  1965=>"100011001",
  1966=>"011110101",
  1967=>"011111000",
  1968=>"100001000",
  1969=>"101111110",
  1970=>"110000111",
  1971=>"110110101",
  1972=>"000100111",
  1973=>"001101001",
  1974=>"001011111",
  1975=>"100000100",
  1976=>"000010000",
  1977=>"101111100",
  1978=>"110010001",
  1979=>"100000001",
  1980=>"110011101",
  1981=>"111100001",
  1982=>"000010000",
  1983=>"100101001",
  1984=>"000100000",
  1985=>"111111000",
  1986=>"111010010",
  1987=>"110001100",
  1988=>"010011101",
  1989=>"111001111",
  1990=>"110110111",
  1991=>"100110001",
  1992=>"011100111",
  1993=>"110000101",
  1994=>"101110110",
  1995=>"100110001",
  1996=>"100111100",
  1997=>"100100000",
  1998=>"011011101",
  1999=>"101000010",
  2000=>"110111100",
  2001=>"010101000",
  2002=>"011111111",
  2003=>"100110100",
  2004=>"100111111",
  2005=>"001010010",
  2006=>"100010110",
  2007=>"110101100",
  2008=>"001001110",
  2009=>"011001101",
  2010=>"101010010",
  2011=>"001011011",
  2012=>"111110101",
  2013=>"110110010",
  2014=>"001010010",
  2015=>"110111001",
  2016=>"101001111",
  2017=>"110011000",
  2018=>"000100001",
  2019=>"100010111",
  2020=>"001100111",
  2021=>"000100000",
  2022=>"010110001",
  2023=>"111000001",
  2024=>"100010110",
  2025=>"111010111",
  2026=>"010001100",
  2027=>"000001001",
  2028=>"110100010",
  2029=>"110101110",
  2030=>"101100000",
  2031=>"111101000",
  2032=>"011101101",
  2033=>"010111011",
  2034=>"111011001",
  2035=>"101000011",
  2036=>"100101111",
  2037=>"100001010",
  2038=>"111011011",
  2039=>"010000011",
  2040=>"010010000",
  2041=>"011001000",
  2042=>"001101010",
  2043=>"110100010",
  2044=>"111111101",
  2045=>"010011010",
  2046=>"000111001",
  2047=>"000001101",
  2048=>"111100010",
  2049=>"001001001",
  2050=>"001110001",
  2051=>"011110111",
  2052=>"010010001",
  2053=>"001100101",
  2054=>"011111011",
  2055=>"100000011",
  2056=>"100100101",
  2057=>"100111011",
  2058=>"000101011",
  2059=>"000011010",
  2060=>"100111100",
  2061=>"010000000",
  2062=>"001111001",
  2063=>"110100010",
  2064=>"011011010",
  2065=>"000111111",
  2066=>"111110010",
  2067=>"010100100",
  2068=>"110101000",
  2069=>"100111000",
  2070=>"111111010",
  2071=>"010100000",
  2072=>"011111101",
  2073=>"000110100",
  2074=>"000010111",
  2075=>"111101011",
  2076=>"111100111",
  2077=>"010011100",
  2078=>"011111100",
  2079=>"001000011",
  2080=>"001000010",
  2081=>"110010000",
  2082=>"000011011",
  2083=>"110000000",
  2084=>"001011100",
  2085=>"101101010",
  2086=>"110001111",
  2087=>"011100110",
  2088=>"100110111",
  2089=>"000000111",
  2090=>"110010010",
  2091=>"001011110",
  2092=>"101010101",
  2093=>"101011101",
  2094=>"000110010",
  2095=>"101000110",
  2096=>"011001011",
  2097=>"101010111",
  2098=>"111100110",
  2099=>"011101011",
  2100=>"111000011",
  2101=>"100110011",
  2102=>"101100111",
  2103=>"011011101",
  2104=>"111101101",
  2105=>"010100011",
  2106=>"110110111",
  2107=>"000001110",
  2108=>"010010010",
  2109=>"100110010",
  2110=>"001110100",
  2111=>"100011101",
  2112=>"111011001",
  2113=>"110101001",
  2114=>"101100100",
  2115=>"110110111",
  2116=>"110111000",
  2117=>"100001011",
  2118=>"110110111",
  2119=>"001001000",
  2120=>"100101001",
  2121=>"011101010",
  2122=>"011010110",
  2123=>"011110111",
  2124=>"111100000",
  2125=>"000101100",
  2126=>"101001111",
  2127=>"010010110",
  2128=>"000100001",
  2129=>"111010111",
  2130=>"111110100",
  2131=>"111001000",
  2132=>"100111100",
  2133=>"101101111",
  2134=>"101101000",
  2135=>"010011001",
  2136=>"110001001",
  2137=>"110111001",
  2138=>"010010011",
  2139=>"110010100",
  2140=>"001110001",
  2141=>"110001100",
  2142=>"100110101",
  2143=>"110010111",
  2144=>"000011001",
  2145=>"111011100",
  2146=>"101000000",
  2147=>"000100001",
  2148=>"010000010",
  2149=>"100011101",
  2150=>"111110111",
  2151=>"011100011",
  2152=>"011011111",
  2153=>"111000001",
  2154=>"000100100",
  2155=>"001011100",
  2156=>"101010111",
  2157=>"011100000",
  2158=>"010111000",
  2159=>"011001110",
  2160=>"100100100",
  2161=>"110100000",
  2162=>"100111001",
  2163=>"000111000",
  2164=>"101001000",
  2165=>"000001111",
  2166=>"100000010",
  2167=>"001010010",
  2168=>"100111000",
  2169=>"110000100",
  2170=>"110111100",
  2171=>"100001100",
  2172=>"000100100",
  2173=>"101110011",
  2174=>"100000011",
  2175=>"100011010",
  2176=>"000110010",
  2177=>"010111000",
  2178=>"101100100",
  2179=>"011000010",
  2180=>"101011101",
  2181=>"011000000",
  2182=>"101111101",
  2183=>"111011110",
  2184=>"100001010",
  2185=>"011111000",
  2186=>"101101000",
  2187=>"110000011",
  2188=>"111101110",
  2189=>"010011011",
  2190=>"110000110",
  2191=>"000000100",
  2192=>"111111001",
  2193=>"100001110",
  2194=>"010010000",
  2195=>"001110001",
  2196=>"011100100",
  2197=>"110011001",
  2198=>"111001111",
  2199=>"101100001",
  2200=>"000011001",
  2201=>"010101110",
  2202=>"001100110",
  2203=>"100011100",
  2204=>"010010000",
  2205=>"111100000",
  2206=>"000110010",
  2207=>"111010111",
  2208=>"100010010",
  2209=>"111001001",
  2210=>"111000100",
  2211=>"010010000",
  2212=>"111010110",
  2213=>"110001011",
  2214=>"110110110",
  2215=>"000010111",
  2216=>"010000111",
  2217=>"001010110",
  2218=>"111111011",
  2219=>"111110001",
  2220=>"011001100",
  2221=>"011001000",
  2222=>"000101011",
  2223=>"011101001",
  2224=>"101001011",
  2225=>"110110111",
  2226=>"110000010",
  2227=>"010111110",
  2228=>"001011001",
  2229=>"100100110",
  2230=>"100001101",
  2231=>"011001010",
  2232=>"001100110",
  2233=>"100000011",
  2234=>"001111011",
  2235=>"101001001",
  2236=>"010111101",
  2237=>"001100001",
  2238=>"100101110",
  2239=>"010100010",
  2240=>"010101010",
  2241=>"100001100",
  2242=>"011110011",
  2243=>"100100011",
  2244=>"000011011",
  2245=>"010111011",
  2246=>"000110011",
  2247=>"000000000",
  2248=>"001010010",
  2249=>"110000110",
  2250=>"000100011",
  2251=>"100101110",
  2252=>"111011000",
  2253=>"011011110",
  2254=>"110000100",
  2255=>"111111010",
  2256=>"011000010",
  2257=>"001100111",
  2258=>"111001011",
  2259=>"111000101",
  2260=>"011011101",
  2261=>"000011011",
  2262=>"010110011",
  2263=>"111011110",
  2264=>"011001101",
  2265=>"001001100",
  2266=>"010100111",
  2267=>"011100010",
  2268=>"001010101",
  2269=>"011101011",
  2270=>"001110000",
  2271=>"111000001",
  2272=>"001101101",
  2273=>"001010111",
  2274=>"111010010",
  2275=>"000001000",
  2276=>"000111111",
  2277=>"100000111",
  2278=>"011001000",
  2279=>"110101000",
  2280=>"100111111",
  2281=>"110010000",
  2282=>"000000010",
  2283=>"011010001",
  2284=>"111110100",
  2285=>"001000110",
  2286=>"101001000",
  2287=>"011011101",
  2288=>"001101110",
  2289=>"101101110",
  2290=>"000010001",
  2291=>"000010000",
  2292=>"010001000",
  2293=>"100011101",
  2294=>"001000001",
  2295=>"000101011",
  2296=>"101000010",
  2297=>"010111100",
  2298=>"101111110",
  2299=>"011100110",
  2300=>"100100010",
  2301=>"100010001",
  2302=>"000010000",
  2303=>"010100010",
  2304=>"001110100",
  2305=>"011001100",
  2306=>"100010100",
  2307=>"110000010",
  2308=>"011110010",
  2309=>"001000111",
  2310=>"100001011",
  2311=>"110000011",
  2312=>"001000100",
  2313=>"100110111",
  2314=>"100100010",
  2315=>"000011111",
  2316=>"100000100",
  2317=>"100011110",
  2318=>"110110011",
  2319=>"110001110",
  2320=>"000000110",
  2321=>"000010011",
  2322=>"101010101",
  2323=>"101111101",
  2324=>"010011100",
  2325=>"110100110",
  2326=>"111101000",
  2327=>"110100000",
  2328=>"100000101",
  2329=>"111010101",
  2330=>"111011110",
  2331=>"111111000",
  2332=>"010010110",
  2333=>"011000001",
  2334=>"111100000",
  2335=>"000010110",
  2336=>"011011101",
  2337=>"000011110",
  2338=>"000011110",
  2339=>"011010000",
  2340=>"101101101",
  2341=>"111111000",
  2342=>"000000010",
  2343=>"110010101",
  2344=>"000011111",
  2345=>"100000101",
  2346=>"110000101",
  2347=>"000110100",
  2348=>"101110000",
  2349=>"111010110",
  2350=>"010010010",
  2351=>"110001000",
  2352=>"010100011",
  2353=>"111111110",
  2354=>"011110111",
  2355=>"010000011",
  2356=>"000000111",
  2357=>"101000011",
  2358=>"111101111",
  2359=>"011111000",
  2360=>"101101000",
  2361=>"110100010",
  2362=>"110111011",
  2363=>"001011100",
  2364=>"111010110",
  2365=>"110011000",
  2366=>"001101110",
  2367=>"101001100",
  2368=>"111011011",
  2369=>"100000100",
  2370=>"111110110",
  2371=>"111001000",
  2372=>"010010010",
  2373=>"100110010",
  2374=>"010111001",
  2375=>"110010011",
  2376=>"011111001",
  2377=>"110010001",
  2378=>"110101011",
  2379=>"010100101",
  2380=>"010001000",
  2381=>"110111100",
  2382=>"001101001",
  2383=>"100011110",
  2384=>"000110111",
  2385=>"111111010",
  2386=>"010011010",
  2387=>"011011110",
  2388=>"110001001",
  2389=>"110110011",
  2390=>"111010100",
  2391=>"010001110",
  2392=>"000111010",
  2393=>"111011111",
  2394=>"011011100",
  2395=>"010100101",
  2396=>"111101110",
  2397=>"100011001",
  2398=>"110100110",
  2399=>"101110111",
  2400=>"000011000",
  2401=>"000010010",
  2402=>"000101011",
  2403=>"110011101",
  2404=>"011100101",
  2405=>"110111001",
  2406=>"001010110",
  2407=>"000011110",
  2408=>"010011111",
  2409=>"000100110",
  2410=>"001011010",
  2411=>"111110111",
  2412=>"101001000",
  2413=>"101100001",
  2414=>"011100010",
  2415=>"010001000",
  2416=>"110101100",
  2417=>"001110111",
  2418=>"011000100",
  2419=>"011001100",
  2420=>"010111110",
  2421=>"001000110",
  2422=>"110111111",
  2423=>"011101101",
  2424=>"100011010",
  2425=>"110001000",
  2426=>"110101001",
  2427=>"000111011",
  2428=>"000001110",
  2429=>"000100010",
  2430=>"101100010",
  2431=>"100000111",
  2432=>"101110000",
  2433=>"010000000",
  2434=>"000110101",
  2435=>"000111110",
  2436=>"111000011",
  2437=>"010100010",
  2438=>"110011111",
  2439=>"011101101",
  2440=>"000111001",
  2441=>"001111100",
  2442=>"110101011",
  2443=>"001000001",
  2444=>"111111001",
  2445=>"111001001",
  2446=>"101010011",
  2447=>"010111111",
  2448=>"111001011",
  2449=>"000110000",
  2450=>"100110011",
  2451=>"100011000",
  2452=>"110110101",
  2453=>"001100111",
  2454=>"110110100",
  2455=>"100101101",
  2456=>"101110100",
  2457=>"111100110",
  2458=>"100011010",
  2459=>"011101100",
  2460=>"100111110",
  2461=>"000101000",
  2462=>"010001111",
  2463=>"001101001",
  2464=>"010110100",
  2465=>"000011001",
  2466=>"001110001",
  2467=>"000000010",
  2468=>"001010011",
  2469=>"000010001",
  2470=>"011010010",
  2471=>"010101010",
  2472=>"110101111",
  2473=>"110010001",
  2474=>"111100001",
  2475=>"101111100",
  2476=>"010000110",
  2477=>"010101001",
  2478=>"100011111",
  2479=>"111111000",
  2480=>"010110110",
  2481=>"001011011",
  2482=>"110001001",
  2483=>"010101011",
  2484=>"111001101",
  2485=>"110010101",
  2486=>"111011001",
  2487=>"011011001",
  2488=>"110110101",
  2489=>"000111101",
  2490=>"110010001",
  2491=>"101101111",
  2492=>"110110010",
  2493=>"010101111",
  2494=>"100100111",
  2495=>"110001001",
  2496=>"001000100",
  2497=>"100100110",
  2498=>"000111010",
  2499=>"000100011",
  2500=>"111001011",
  2501=>"111010111",
  2502=>"011011110",
  2503=>"100111000",
  2504=>"010111101",
  2505=>"111101000",
  2506=>"010110100",
  2507=>"110110011",
  2508=>"011001100",
  2509=>"001111101",
  2510=>"010110010",
  2511=>"011110110",
  2512=>"010110111",
  2513=>"101110000",
  2514=>"001000000",
  2515=>"101000000",
  2516=>"101000111",
  2517=>"010000001",
  2518=>"110110111",
  2519=>"000010110",
  2520=>"010110100",
  2521=>"011101000",
  2522=>"010011010",
  2523=>"110011011",
  2524=>"110111010",
  2525=>"010001101",
  2526=>"011100100",
  2527=>"111011000",
  2528=>"100011010",
  2529=>"010111000",
  2530=>"110100010",
  2531=>"110011011",
  2532=>"101000111",
  2533=>"010000111",
  2534=>"100001101",
  2535=>"101001101",
  2536=>"010100000",
  2537=>"000101101",
  2538=>"111111011",
  2539=>"110011111",
  2540=>"010101011",
  2541=>"111011000",
  2542=>"000001011",
  2543=>"100110000",
  2544=>"001001010",
  2545=>"101000100",
  2546=>"100001110",
  2547=>"101110111",
  2548=>"000010101",
  2549=>"111111010",
  2550=>"011101001",
  2551=>"100011111",
  2552=>"001101010",
  2553=>"000001000",
  2554=>"110000111",
  2555=>"011111110",
  2556=>"001110101",
  2557=>"110100110",
  2558=>"000011110",
  2559=>"000100001",
  2560=>"001111010",
  2561=>"101110111",
  2562=>"100110001",
  2563=>"110001111",
  2564=>"110001010",
  2565=>"010000000",
  2566=>"100111011",
  2567=>"111010010",
  2568=>"110100100",
  2569=>"010011110",
  2570=>"010010101",
  2571=>"001000101",
  2572=>"110010101",
  2573=>"110010101",
  2574=>"110101011",
  2575=>"100100101",
  2576=>"110101011",
  2577=>"001001011",
  2578=>"100101011",
  2579=>"011000011",
  2580=>"110101010",
  2581=>"111010000",
  2582=>"010111010",
  2583=>"100010110",
  2584=>"011011101",
  2585=>"110000111",
  2586=>"001101111",
  2587=>"100010001",
  2588=>"010101000",
  2589=>"000000001",
  2590=>"111111001",
  2591=>"011011011",
  2592=>"011001111",
  2593=>"001001101",
  2594=>"100001111",
  2595=>"010001101",
  2596=>"010011010",
  2597=>"110100101",
  2598=>"100010110",
  2599=>"010110110",
  2600=>"110101100",
  2601=>"100111100",
  2602=>"010001110",
  2603=>"011001100",
  2604=>"110110000",
  2605=>"000100110",
  2606=>"000101010",
  2607=>"101100010",
  2608=>"111000101",
  2609=>"100001000",
  2610=>"111101001",
  2611=>"111111110",
  2612=>"100000101",
  2613=>"011010011",
  2614=>"101111010",
  2615=>"101101010",
  2616=>"100011001",
  2617=>"011011000",
  2618=>"101100101",
  2619=>"101110001",
  2620=>"000101000",
  2621=>"001100111",
  2622=>"111001011",
  2623=>"011010010",
  2624=>"011110000",
  2625=>"110001101",
  2626=>"111011100",
  2627=>"010101000",
  2628=>"011100111",
  2629=>"111101001",
  2630=>"100001011",
  2631=>"001111010",
  2632=>"101100010",
  2633=>"011011011",
  2634=>"111100111",
  2635=>"100101010",
  2636=>"111101100",
  2637=>"001101111",
  2638=>"111101011",
  2639=>"001010011",
  2640=>"101011111",
  2641=>"101101000",
  2642=>"010010100",
  2643=>"010111010",
  2644=>"010001000",
  2645=>"010111111",
  2646=>"000001100",
  2647=>"011001110",
  2648=>"110101110",
  2649=>"101001010",
  2650=>"000010000",
  2651=>"100111100",
  2652=>"001010000",
  2653=>"010011000",
  2654=>"001111100",
  2655=>"101111101",
  2656=>"100001110",
  2657=>"011101001",
  2658=>"100010110",
  2659=>"110101110",
  2660=>"101111100",
  2661=>"010110011",
  2662=>"011110001",
  2663=>"011000001",
  2664=>"110111110",
  2665=>"010010101",
  2666=>"011011011",
  2667=>"011110110",
  2668=>"010110011",
  2669=>"011101100",
  2670=>"000111101",
  2671=>"000111111",
  2672=>"110110000",
  2673=>"111000011",
  2674=>"011100111",
  2675=>"100001110",
  2676=>"101001101",
  2677=>"011101101",
  2678=>"100011100",
  2679=>"000000000",
  2680=>"001100101",
  2681=>"010100110",
  2682=>"100110000",
  2683=>"001011010",
  2684=>"100000010",
  2685=>"010100110",
  2686=>"010100011",
  2687=>"010101010",
  2688=>"010101100",
  2689=>"010101111",
  2690=>"100100000",
  2691=>"001001100",
  2692=>"100010000",
  2693=>"111110010",
  2694=>"001101110",
  2695=>"010001101",
  2696=>"101101111",
  2697=>"001111010",
  2698=>"001100110",
  2699=>"001001011",
  2700=>"011010101",
  2701=>"010010001",
  2702=>"100001111",
  2703=>"101011010",
  2704=>"001001010",
  2705=>"010010011",
  2706=>"101011010",
  2707=>"101000001",
  2708=>"110100001",
  2709=>"110111000",
  2710=>"001110110",
  2711=>"111010111",
  2712=>"111111100",
  2713=>"010010010",
  2714=>"000110001",
  2715=>"110101100",
  2716=>"011000110",
  2717=>"001010000",
  2718=>"010010001",
  2719=>"111011100",
  2720=>"011110001",
  2721=>"010001001",
  2722=>"101001101",
  2723=>"100111111",
  2724=>"100011011",
  2725=>"001100100",
  2726=>"001011011",
  2727=>"000011011",
  2728=>"000101101",
  2729=>"100100011",
  2730=>"000110110",
  2731=>"000100101",
  2732=>"010000001",
  2733=>"001011110",
  2734=>"000000101",
  2735=>"011100011",
  2736=>"001000100",
  2737=>"001110101",
  2738=>"011011110",
  2739=>"010100100",
  2740=>"110101100",
  2741=>"111100101",
  2742=>"001011101",
  2743=>"000010110",
  2744=>"100000101",
  2745=>"110110001",
  2746=>"100100100",
  2747=>"101000101",
  2748=>"010111011",
  2749=>"110000101",
  2750=>"011110010",
  2751=>"101111111",
  2752=>"111001110",
  2753=>"100010011",
  2754=>"101100111",
  2755=>"010111101",
  2756=>"111111000",
  2757=>"000010010",
  2758=>"011000000",
  2759=>"010000110",
  2760=>"100111001",
  2761=>"101010111",
  2762=>"001010111",
  2763=>"101011110",
  2764=>"001011101",
  2765=>"001100011",
  2766=>"100101000",
  2767=>"010000110",
  2768=>"110100010",
  2769=>"010000000",
  2770=>"001101110",
  2771=>"011001101",
  2772=>"111110111",
  2773=>"111111000",
  2774=>"100111110",
  2775=>"000101010",
  2776=>"100001101",
  2777=>"111011010",
  2778=>"110110011",
  2779=>"101010011",
  2780=>"010100000",
  2781=>"011000010",
  2782=>"111110011",
  2783=>"001100001",
  2784=>"101110110",
  2785=>"100010111",
  2786=>"110100001",
  2787=>"011100111",
  2788=>"000101001",
  2789=>"000001110",
  2790=>"010001001",
  2791=>"011100111",
  2792=>"001111111",
  2793=>"111110101",
  2794=>"001001000",
  2795=>"010110001",
  2796=>"000010000",
  2797=>"010000001",
  2798=>"111111100",
  2799=>"011101010",
  2800=>"001110101",
  2801=>"000101110",
  2802=>"011010010",
  2803=>"111110100",
  2804=>"000001001",
  2805=>"111001110",
  2806=>"010111100",
  2807=>"001111010",
  2808=>"011111011",
  2809=>"010110101",
  2810=>"101001110",
  2811=>"111011110",
  2812=>"100011100",
  2813=>"111111110",
  2814=>"011111111",
  2815=>"111100111",
  2816=>"110010101",
  2817=>"100110101",
  2818=>"101110111",
  2819=>"011111010",
  2820=>"000100000",
  2821=>"011001111",
  2822=>"011110111",
  2823=>"010011111",
  2824=>"010011110",
  2825=>"111010010",
  2826=>"101100000",
  2827=>"101101110",
  2828=>"111110101",
  2829=>"001011000",
  2830=>"011111010",
  2831=>"011000000",
  2832=>"010000000",
  2833=>"101110101",
  2834=>"110111010",
  2835=>"100110100",
  2836=>"000011111",
  2837=>"111101100",
  2838=>"000101100",
  2839=>"010010110",
  2840=>"110000010",
  2841=>"100011110",
  2842=>"000000111",
  2843=>"001110011",
  2844=>"000111001",
  2845=>"110010011",
  2846=>"000000100",
  2847=>"000010100",
  2848=>"101100000",
  2849=>"001111110",
  2850=>"111100011",
  2851=>"100011101",
  2852=>"100011101",
  2853=>"110000111",
  2854=>"101011111",
  2855=>"001000001",
  2856=>"001101001",
  2857=>"011011001",
  2858=>"110101001",
  2859=>"110011011",
  2860=>"111111000",
  2861=>"001100000",
  2862=>"101000100",
  2863=>"100001011",
  2864=>"100001110",
  2865=>"010100101",
  2866=>"000111101",
  2867=>"101001101",
  2868=>"101111010",
  2869=>"100101110",
  2870=>"110000011",
  2871=>"100101111",
  2872=>"010010101",
  2873=>"011101111",
  2874=>"011100100",
  2875=>"010000111",
  2876=>"000010100",
  2877=>"100001100",
  2878=>"101000000",
  2879=>"011010001",
  2880=>"010100111",
  2881=>"101101001",
  2882=>"010101001",
  2883=>"110010000",
  2884=>"000111011",
  2885=>"010101111",
  2886=>"100101110",
  2887=>"110001010",
  2888=>"101001001",
  2889=>"001111011",
  2890=>"001100011",
  2891=>"111011110",
  2892=>"000100000",
  2893=>"111110111",
  2894=>"110110011",
  2895=>"111000001",
  2896=>"100101001",
  2897=>"100010101",
  2898=>"000000100",
  2899=>"010101011",
  2900=>"100111000",
  2901=>"000001101",
  2902=>"100111001",
  2903=>"110110100",
  2904=>"001111110",
  2905=>"100101100",
  2906=>"001000110",
  2907=>"010000010",
  2908=>"111101011",
  2909=>"101000110",
  2910=>"010111001",
  2911=>"001100101",
  2912=>"000000101",
  2913=>"000001011",
  2914=>"000001100",
  2915=>"110011011",
  2916=>"111011000",
  2917=>"000010010",
  2918=>"010010011",
  2919=>"101101000",
  2920=>"110111101",
  2921=>"000111000",
  2922=>"110101000",
  2923=>"000010111",
  2924=>"111010110",
  2925=>"000111000",
  2926=>"000001001",
  2927=>"100110110",
  2928=>"001011101",
  2929=>"010010110",
  2930=>"111011110",
  2931=>"000000111",
  2932=>"100101010",
  2933=>"000110000",
  2934=>"000100101",
  2935=>"000100010",
  2936=>"100001101",
  2937=>"011110100",
  2938=>"001101110",
  2939=>"100010001",
  2940=>"001110100",
  2941=>"101001101",
  2942=>"111101111",
  2943=>"111010001",
  2944=>"000010111",
  2945=>"101000001",
  2946=>"100000011",
  2947=>"000011001",
  2948=>"000010110",
  2949=>"001010000",
  2950=>"011010111",
  2951=>"000110101",
  2952=>"101101101",
  2953=>"110001100",
  2954=>"101111001",
  2955=>"011011100",
  2956=>"110110110",
  2957=>"111011000",
  2958=>"000010011",
  2959=>"110110001",
  2960=>"000111010",
  2961=>"011010111",
  2962=>"011001111",
  2963=>"001111001",
  2964=>"011111000",
  2965=>"100110011",
  2966=>"010001100",
  2967=>"101010000",
  2968=>"000000110",
  2969=>"011010001",
  2970=>"101010101",
  2971=>"010011110",
  2972=>"010011011",
  2973=>"100010000",
  2974=>"011000001",
  2975=>"101000010",
  2976=>"010010010",
  2977=>"110100000",
  2978=>"000001010",
  2979=>"110100001",
  2980=>"101110101",
  2981=>"000101000",
  2982=>"110000000",
  2983=>"101111001",
  2984=>"101100110",
  2985=>"111010000",
  2986=>"011101000",
  2987=>"100000011",
  2988=>"101001100",
  2989=>"000110000",
  2990=>"101101010",
  2991=>"111110111",
  2992=>"011100010",
  2993=>"010110011",
  2994=>"010000101",
  2995=>"011110111",
  2996=>"010000010",
  2997=>"101000000",
  2998=>"000011111",
  2999=>"011110010",
  3000=>"101101100",
  3001=>"010001000",
  3002=>"000001100",
  3003=>"111100100",
  3004=>"100100000",
  3005=>"010101101",
  3006=>"010101000",
  3007=>"101101001",
  3008=>"000110000",
  3009=>"100010111",
  3010=>"000110010",
  3011=>"100011110",
  3012=>"110011101",
  3013=>"110100110",
  3014=>"110001010",
  3015=>"010010111",
  3016=>"011100101",
  3017=>"010010111",
  3018=>"010100100",
  3019=>"001100001",
  3020=>"000101001",
  3021=>"100000000",
  3022=>"011011000",
  3023=>"101101101",
  3024=>"110000111",
  3025=>"111101101",
  3026=>"110010101",
  3027=>"001110000",
  3028=>"111001111",
  3029=>"000111011",
  3030=>"011111110",
  3031=>"010000101",
  3032=>"001010001",
  3033=>"011100000",
  3034=>"111011111",
  3035=>"000111100",
  3036=>"111111011",
  3037=>"111111100",
  3038=>"001001111",
  3039=>"010101001",
  3040=>"110100010",
  3041=>"100110000",
  3042=>"010001010",
  3043=>"010111001",
  3044=>"111000100",
  3045=>"110000010",
  3046=>"010011011",
  3047=>"011100011",
  3048=>"101011101",
  3049=>"110010000",
  3050=>"001111110",
  3051=>"101001001",
  3052=>"001101010",
  3053=>"010001001",
  3054=>"110110001",
  3055=>"010000100",
  3056=>"000000111",
  3057=>"111001101",
  3058=>"011111111",
  3059=>"111001110",
  3060=>"011111111",
  3061=>"001000000",
  3062=>"100111000",
  3063=>"111101000",
  3064=>"110110101",
  3065=>"010110100",
  3066=>"010100110",
  3067=>"111000100",
  3068=>"001100010",
  3069=>"001111110",
  3070=>"000000101",
  3071=>"010010011",
  3072=>"110101111",
  3073=>"111111100",
  3074=>"001001010",
  3075=>"111001000",
  3076=>"010001101",
  3077=>"101001100",
  3078=>"000000001",
  3079=>"011010000",
  3080=>"101010110",
  3081=>"111110110",
  3082=>"100000111",
  3083=>"001111010",
  3084=>"110110111",
  3085=>"011011011",
  3086=>"011101111",
  3087=>"100010011",
  3088=>"100110001",
  3089=>"111111111",
  3090=>"110011110",
  3091=>"001100101",
  3092=>"011000100",
  3093=>"110001100",
  3094=>"011011001",
  3095=>"110010111",
  3096=>"001101101",
  3097=>"100000001",
  3098=>"110101100",
  3099=>"001101101",
  3100=>"000000100",
  3101=>"111101111",
  3102=>"110010101",
  3103=>"101110000",
  3104=>"111100110",
  3105=>"110101100",
  3106=>"000101001",
  3107=>"101110010",
  3108=>"011000010",
  3109=>"011000001",
  3110=>"011000101",
  3111=>"001110001",
  3112=>"110011110",
  3113=>"000100111",
  3114=>"110101000",
  3115=>"111000101",
  3116=>"000101100",
  3117=>"010010000",
  3118=>"110001111",
  3119=>"001100110",
  3120=>"111111010",
  3121=>"001101110",
  3122=>"010011011",
  3123=>"001100100",
  3124=>"011111100",
  3125=>"000000001",
  3126=>"110110111",
  3127=>"000100000",
  3128=>"010101000",
  3129=>"011110100",
  3130=>"011101100",
  3131=>"010100011",
  3132=>"010000010",
  3133=>"010110111",
  3134=>"010001110",
  3135=>"010010100",
  3136=>"100110000",
  3137=>"101000101",
  3138=>"101000000",
  3139=>"100101000",
  3140=>"010001110",
  3141=>"110011111",
  3142=>"011011101",
  3143=>"001010111",
  3144=>"001100001",
  3145=>"110110110",
  3146=>"001101000",
  3147=>"011100010",
  3148=>"011001010",
  3149=>"110110000",
  3150=>"001110000",
  3151=>"110110111",
  3152=>"100111011",
  3153=>"011000011",
  3154=>"100010111",
  3155=>"101011110",
  3156=>"011100111",
  3157=>"100110101",
  3158=>"011011111",
  3159=>"000010011",
  3160=>"000101110",
  3161=>"001011110",
  3162=>"000010100",
  3163=>"000111011",
  3164=>"010111011",
  3165=>"010000001",
  3166=>"111000010",
  3167=>"111001101",
  3168=>"110110110",
  3169=>"100100010",
  3170=>"000111010",
  3171=>"110011100",
  3172=>"100000000",
  3173=>"111001011",
  3174=>"000000111",
  3175=>"010001001",
  3176=>"000101000",
  3177=>"011101010",
  3178=>"011011000",
  3179=>"001111011",
  3180=>"100100100",
  3181=>"101111000",
  3182=>"011110010",
  3183=>"011011010",
  3184=>"001011011",
  3185=>"111000010",
  3186=>"001001100",
  3187=>"001000110",
  3188=>"111011011",
  3189=>"011001000",
  3190=>"100000100",
  3191=>"111011110",
  3192=>"000000110",
  3193=>"111110010",
  3194=>"011011110",
  3195=>"100110111",
  3196=>"010000010",
  3197=>"001101010",
  3198=>"110100010",
  3199=>"011011101",
  3200=>"101011000",
  3201=>"111100100",
  3202=>"001001001",
  3203=>"010101100",
  3204=>"101100001",
  3205=>"100111101",
  3206=>"001010011",
  3207=>"100001100",
  3208=>"011101010",
  3209=>"111000001",
  3210=>"111110110",
  3211=>"111010110",
  3212=>"110001100",
  3213=>"101000011",
  3214=>"100101000",
  3215=>"000111010",
  3216=>"010001111",
  3217=>"110000010",
  3218=>"111110101",
  3219=>"001100001",
  3220=>"000010101",
  3221=>"110010001",
  3222=>"011000000",
  3223=>"000010111",
  3224=>"101100001",
  3225=>"000011010",
  3226=>"010101100",
  3227=>"000101101",
  3228=>"000011111",
  3229=>"110100110",
  3230=>"011100110",
  3231=>"110011100",
  3232=>"001101011",
  3233=>"011101101",
  3234=>"111011010",
  3235=>"001001000",
  3236=>"100110100",
  3237=>"010010111",
  3238=>"000101001",
  3239=>"011010001",
  3240=>"000000101",
  3241=>"001110010",
  3242=>"001011001",
  3243=>"000000011",
  3244=>"100101001",
  3245=>"000100111",
  3246=>"011101101",
  3247=>"011100010",
  3248=>"001000001",
  3249=>"010100110",
  3250=>"010000110",
  3251=>"111111010",
  3252=>"110100000",
  3253=>"010101000",
  3254=>"001001011",
  3255=>"100100011",
  3256=>"011001010",
  3257=>"000001010",
  3258=>"000101001",
  3259=>"100000000",
  3260=>"010000101",
  3261=>"111111010",
  3262=>"110001111",
  3263=>"010010000",
  3264=>"111000100",
  3265=>"001100111",
  3266=>"000010000",
  3267=>"000110001",
  3268=>"100111111",
  3269=>"110100001",
  3270=>"111100010",
  3271=>"100110111",
  3272=>"101011011",
  3273=>"011101101",
  3274=>"011010110",
  3275=>"001011001",
  3276=>"100010001",
  3277=>"111101000",
  3278=>"001010010",
  3279=>"100111100",
  3280=>"000100000",
  3281=>"011100101",
  3282=>"011001001",
  3283=>"001000110",
  3284=>"010111010",
  3285=>"111110001",
  3286=>"011010000",
  3287=>"001100110",
  3288=>"101100110",
  3289=>"110100101",
  3290=>"110110101",
  3291=>"001000000",
  3292=>"011111000",
  3293=>"000011111",
  3294=>"110111010",
  3295=>"110100001",
  3296=>"000010111",
  3297=>"100010001",
  3298=>"010000101",
  3299=>"110001000",
  3300=>"010011110",
  3301=>"100110011",
  3302=>"110101111",
  3303=>"000110001",
  3304=>"111011100",
  3305=>"010101111",
  3306=>"111101111",
  3307=>"010111000",
  3308=>"101101001",
  3309=>"111111101",
  3310=>"111011101",
  3311=>"101111111",
  3312=>"001011111",
  3313=>"000011010",
  3314=>"110000100",
  3315=>"100010000",
  3316=>"011111011",
  3317=>"111110110",
  3318=>"000111000",
  3319=>"110010111",
  3320=>"010110001",
  3321=>"100111000",
  3322=>"101000010",
  3323=>"100110011",
  3324=>"000110111",
  3325=>"100101100",
  3326=>"011110111",
  3327=>"001001000",
  3328=>"000010111",
  3329=>"001100011",
  3330=>"111011100",
  3331=>"100110001",
  3332=>"010100011",
  3333=>"100010100",
  3334=>"000000100",
  3335=>"010000110",
  3336=>"000110010",
  3337=>"000001110",
  3338=>"011010000",
  3339=>"110110001",
  3340=>"010100010",
  3341=>"100101001",
  3342=>"011100100",
  3343=>"111010101",
  3344=>"110010001",
  3345=>"010101110",
  3346=>"101100100",
  3347=>"101001001",
  3348=>"110100110",
  3349=>"001000100",
  3350=>"011010111",
  3351=>"100100010",
  3352=>"011000000",
  3353=>"100100101",
  3354=>"001100111",
  3355=>"011010000",
  3356=>"000110011",
  3357=>"010110100",
  3358=>"110010110",
  3359=>"100001001",
  3360=>"110011011",
  3361=>"000101000",
  3362=>"000000001",
  3363=>"010011101",
  3364=>"100101001",
  3365=>"000100000",
  3366=>"111110100",
  3367=>"000100011",
  3368=>"111111000",
  3369=>"010100110",
  3370=>"111101001",
  3371=>"101001000",
  3372=>"101011111",
  3373=>"001010011",
  3374=>"111110000",
  3375=>"101001000",
  3376=>"110111000",
  3377=>"110100110",
  3378=>"000101001",
  3379=>"110111000",
  3380=>"111110110",
  3381=>"011000000",
  3382=>"111101101",
  3383=>"110110011",
  3384=>"010010011",
  3385=>"010110010",
  3386=>"011110001",
  3387=>"000001011",
  3388=>"110000100",
  3389=>"000001101",
  3390=>"111110100",
  3391=>"110000010",
  3392=>"101010011",
  3393=>"000101001",
  3394=>"101010001",
  3395=>"001011111",
  3396=>"110101110",
  3397=>"100001000",
  3398=>"110001100",
  3399=>"110010110",
  3400=>"000010101",
  3401=>"001000000",
  3402=>"001100110",
  3403=>"001010101",
  3404=>"010101111",
  3405=>"010011001",
  3406=>"110101110",
  3407=>"111111111",
  3408=>"001000000",
  3409=>"101111011",
  3410=>"011100010",
  3411=>"111100001",
  3412=>"011011011",
  3413=>"111000010",
  3414=>"100111110",
  3415=>"100000010",
  3416=>"011101110",
  3417=>"001111101",
  3418=>"011111000",
  3419=>"100110101",
  3420=>"110101010",
  3421=>"010000010",
  3422=>"110101110",
  3423=>"101100011",
  3424=>"100101001",
  3425=>"101100000",
  3426=>"000001101",
  3427=>"010101001",
  3428=>"100001001",
  3429=>"000100110",
  3430=>"000001010",
  3431=>"010111100",
  3432=>"100111001",
  3433=>"011100100",
  3434=>"110110011",
  3435=>"001100111",
  3436=>"111000001",
  3437=>"011011010",
  3438=>"010000010",
  3439=>"010000011",
  3440=>"001001000",
  3441=>"111001001",
  3442=>"101111111",
  3443=>"101110010",
  3444=>"001010010",
  3445=>"110101111",
  3446=>"111011100",
  3447=>"110110001",
  3448=>"001101010",
  3449=>"001111000",
  3450=>"111100001",
  3451=>"001000110",
  3452=>"101000110",
  3453=>"101010110",
  3454=>"111110100",
  3455=>"100110111",
  3456=>"010000110",
  3457=>"001000010",
  3458=>"110100100",
  3459=>"010101010",
  3460=>"111000010",
  3461=>"000111101",
  3462=>"010010000",
  3463=>"111110101",
  3464=>"111010011",
  3465=>"110111010",
  3466=>"000010000",
  3467=>"100110010",
  3468=>"101000001",
  3469=>"100001110",
  3470=>"100010111",
  3471=>"111100010",
  3472=>"110000101",
  3473=>"111001101",
  3474=>"110110011",
  3475=>"010001100",
  3476=>"001110100",
  3477=>"010000111",
  3478=>"110100110",
  3479=>"101010111",
  3480=>"110011111",
  3481=>"110100010",
  3482=>"110111110",
  3483=>"101100111",
  3484=>"101000110",
  3485=>"100001000",
  3486=>"101100111",
  3487=>"111101101",
  3488=>"100011000",
  3489=>"001100000",
  3490=>"100111100",
  3491=>"101001101",
  3492=>"011100011",
  3493=>"000010101",
  3494=>"101011111",
  3495=>"000010110",
  3496=>"011000010",
  3497=>"000111100",
  3498=>"100111100",
  3499=>"101000100",
  3500=>"110111000",
  3501=>"001100110",
  3502=>"110010011",
  3503=>"100001100",
  3504=>"010100000",
  3505=>"110101110",
  3506=>"011110111",
  3507=>"000010010",
  3508=>"101000111",
  3509=>"010110100",
  3510=>"100101011",
  3511=>"001100010",
  3512=>"101001101",
  3513=>"110111011",
  3514=>"110010100",
  3515=>"111101100",
  3516=>"111010000",
  3517=>"111100100",
  3518=>"001110010",
  3519=>"110110111",
  3520=>"110100011",
  3521=>"010100011",
  3522=>"101111110",
  3523=>"101000001",
  3524=>"011101011",
  3525=>"001011101",
  3526=>"101100010",
  3527=>"100100000",
  3528=>"000100000",
  3529=>"011000110",
  3530=>"101001010",
  3531=>"100010001",
  3532=>"010001101",
  3533=>"111101001",
  3534=>"011001110",
  3535=>"011111000",
  3536=>"111001100",
  3537=>"110100010",
  3538=>"101010001",
  3539=>"101101000",
  3540=>"110111011",
  3541=>"101100001",
  3542=>"010001100",
  3543=>"111100001",
  3544=>"011011100",
  3545=>"100111010",
  3546=>"011000010",
  3547=>"011001000",
  3548=>"000001010",
  3549=>"101100100",
  3550=>"101011001",
  3551=>"101001000",
  3552=>"011001110",
  3553=>"100101100",
  3554=>"011101100",
  3555=>"100100100",
  3556=>"100111011",
  3557=>"110011100",
  3558=>"101101010",
  3559=>"111101101",
  3560=>"101110100",
  3561=>"100000010",
  3562=>"000011000",
  3563=>"000110110",
  3564=>"111111111",
  3565=>"111110101",
  3566=>"100100000",
  3567=>"101010111",
  3568=>"111100110",
  3569=>"110101100",
  3570=>"011001011",
  3571=>"111110010",
  3572=>"000001100",
  3573=>"111010101",
  3574=>"111010111",
  3575=>"000001000",
  3576=>"000110000",
  3577=>"111101010",
  3578=>"001001110",
  3579=>"100011101",
  3580=>"011111001",
  3581=>"111011111",
  3582=>"110110010",
  3583=>"110000000",
  3584=>"111111010",
  3585=>"010011110",
  3586=>"110110000",
  3587=>"101101010",
  3588=>"010010001",
  3589=>"110110111",
  3590=>"010011111",
  3591=>"101101011",
  3592=>"100000101",
  3593=>"001101001",
  3594=>"101111111",
  3595=>"011001010",
  3596=>"010010111",
  3597=>"111000101",
  3598=>"110100000",
  3599=>"010101100",
  3600=>"101010011",
  3601=>"010101010",
  3602=>"011101111",
  3603=>"010100000",
  3604=>"101000100",
  3605=>"100010100",
  3606=>"011000100",
  3607=>"011101110",
  3608=>"011100101",
  3609=>"000010000",
  3610=>"000001100",
  3611=>"110001110",
  3612=>"111111101",
  3613=>"110000100",
  3614=>"000100000",
  3615=>"000001111",
  3616=>"011000001",
  3617=>"101111110",
  3618=>"001000000",
  3619=>"010101100",
  3620=>"011010001",
  3621=>"011011111",
  3622=>"000101100",
  3623=>"110101101",
  3624=>"110100001",
  3625=>"001101111",
  3626=>"111100111",
  3627=>"100001010",
  3628=>"111011011",
  3629=>"011000100",
  3630=>"100011011",
  3631=>"000010111",
  3632=>"001001110",
  3633=>"110011100",
  3634=>"000110010",
  3635=>"000010010",
  3636=>"111100000",
  3637=>"110011111",
  3638=>"101100111",
  3639=>"011010001",
  3640=>"100111011",
  3641=>"011101000",
  3642=>"000001010",
  3643=>"011001001",
  3644=>"000101100",
  3645=>"001111100",
  3646=>"101011100",
  3647=>"001111110",
  3648=>"100011100",
  3649=>"000001001",
  3650=>"001010011",
  3651=>"100000111",
  3652=>"000111011",
  3653=>"000100010",
  3654=>"101001000",
  3655=>"011100001",
  3656=>"111011100",
  3657=>"000010000",
  3658=>"001100001",
  3659=>"001110001",
  3660=>"011001011",
  3661=>"111000100",
  3662=>"010101110",
  3663=>"001101011",
  3664=>"010000000",
  3665=>"001001101",
  3666=>"000101110",
  3667=>"001000111",
  3668=>"100000111",
  3669=>"110000100",
  3670=>"010000001",
  3671=>"010101000",
  3672=>"110010000",
  3673=>"100010000",
  3674=>"100100010",
  3675=>"101011101",
  3676=>"110000101",
  3677=>"010010110",
  3678=>"110010110",
  3679=>"110111100",
  3680=>"111111101",
  3681=>"000010100",
  3682=>"010011101",
  3683=>"001110000",
  3684=>"011101111",
  3685=>"011111011",
  3686=>"000110001",
  3687=>"110111000",
  3688=>"001000110",
  3689=>"100001000",
  3690=>"110101101",
  3691=>"010000000",
  3692=>"100100011",
  3693=>"101011001",
  3694=>"010100110",
  3695=>"011111110",
  3696=>"101101001",
  3697=>"111111100",
  3698=>"101001101",
  3699=>"110111101",
  3700=>"010011100",
  3701=>"101000000",
  3702=>"011100111",
  3703=>"101110100",
  3704=>"000010101",
  3705=>"000101011",
  3706=>"111010000",
  3707=>"111101011",
  3708=>"111111001",
  3709=>"101111101",
  3710=>"011111110",
  3711=>"000111110",
  3712=>"011111111",
  3713=>"101000010",
  3714=>"010101101",
  3715=>"000000011",
  3716=>"000011001",
  3717=>"101100010",
  3718=>"001110010",
  3719=>"011011100",
  3720=>"100101011",
  3721=>"001000110",
  3722=>"001001011",
  3723=>"101000000",
  3724=>"111101000",
  3725=>"110110101",
  3726=>"000101001",
  3727=>"100101100",
  3728=>"010100000",
  3729=>"111011111",
  3730=>"001010101",
  3731=>"111100010",
  3732=>"000111001",
  3733=>"011101101",
  3734=>"010111000",
  3735=>"001111111",
  3736=>"111111011",
  3737=>"011011010",
  3738=>"110100100",
  3739=>"001010010",
  3740=>"000001000",
  3741=>"100110000",
  3742=>"001111011",
  3743=>"111011010",
  3744=>"111000101",
  3745=>"110001100",
  3746=>"100000111",
  3747=>"110101010",
  3748=>"100000100",
  3749=>"010000111",
  3750=>"111001010",
  3751=>"000010000",
  3752=>"001100010",
  3753=>"001100100",
  3754=>"010000110",
  3755=>"010010101",
  3756=>"111011000",
  3757=>"110000000",
  3758=>"001100001",
  3759=>"000101100",
  3760=>"010000110",
  3761=>"011011101",
  3762=>"110111111",
  3763=>"100110001",
  3764=>"000000011",
  3765=>"100100001",
  3766=>"100011100",
  3767=>"100110011",
  3768=>"010111000",
  3769=>"010001110",
  3770=>"001100101",
  3771=>"001001000",
  3772=>"011110010",
  3773=>"100011110",
  3774=>"000110101",
  3775=>"010101111",
  3776=>"111000001",
  3777=>"000000101",
  3778=>"011100111",
  3779=>"110000110",
  3780=>"101010101",
  3781=>"010111110",
  3782=>"110011111",
  3783=>"001100111",
  3784=>"011100110",
  3785=>"110000001",
  3786=>"110000010",
  3787=>"010111010",
  3788=>"011111011",
  3789=>"111011101",
  3790=>"101010110",
  3791=>"000110101",
  3792=>"011100101",
  3793=>"001000111",
  3794=>"000001100",
  3795=>"110111010",
  3796=>"000011011",
  3797=>"000001110",
  3798=>"110111101",
  3799=>"100101011",
  3800=>"000001100",
  3801=>"100110101",
  3802=>"101011110",
  3803=>"100010101",
  3804=>"001110001",
  3805=>"001111001",
  3806=>"011111101",
  3807=>"011100101",
  3808=>"101011001",
  3809=>"001101101",
  3810=>"100000111",
  3811=>"110111100",
  3812=>"111011010",
  3813=>"111011111",
  3814=>"011110000",
  3815=>"100010111",
  3816=>"101010101",
  3817=>"011101100",
  3818=>"101011011",
  3819=>"110000110",
  3820=>"010110110",
  3821=>"100101100",
  3822=>"110011100",
  3823=>"000101000",
  3824=>"000110010",
  3825=>"100111111",
  3826=>"110110001",
  3827=>"100010101",
  3828=>"100001101",
  3829=>"101010111",
  3830=>"010101010",
  3831=>"001000101",
  3832=>"101011101",
  3833=>"010110011",
  3834=>"110001111",
  3835=>"000100101",
  3836=>"000001100",
  3837=>"100000100",
  3838=>"001000000",
  3839=>"100111101",
  3840=>"010110001",
  3841=>"010100011",
  3842=>"010110010",
  3843=>"100101101",
  3844=>"111011010",
  3845=>"001001010",
  3846=>"010110110",
  3847=>"110000000",
  3848=>"101111110",
  3849=>"001011001",
  3850=>"100100000",
  3851=>"101101011",
  3852=>"000011011",
  3853=>"100100001",
  3854=>"011000110",
  3855=>"101000111",
  3856=>"011110100",
  3857=>"000111011",
  3858=>"011111010",
  3859=>"101100000",
  3860=>"011100100",
  3861=>"111100001",
  3862=>"110000101",
  3863=>"011001111",
  3864=>"110000010",
  3865=>"011110111",
  3866=>"001000010",
  3867=>"110111011",
  3868=>"111110111",
  3869=>"001110111",
  3870=>"010110111",
  3871=>"011100000",
  3872=>"111100011",
  3873=>"010110001",
  3874=>"010110001",
  3875=>"111001111",
  3876=>"111110010",
  3877=>"000011000",
  3878=>"011111111",
  3879=>"110010110",
  3880=>"011011010",
  3881=>"000010010",
  3882=>"110011100",
  3883=>"101101100",
  3884=>"110111100",
  3885=>"101000010",
  3886=>"100000010",
  3887=>"111001000",
  3888=>"111010010",
  3889=>"001110100",
  3890=>"010101110",
  3891=>"000000100",
  3892=>"000110010",
  3893=>"110100111",
  3894=>"000001101",
  3895=>"011001110",
  3896=>"110100010",
  3897=>"111010100",
  3898=>"000010100",
  3899=>"111001000",
  3900=>"101000000",
  3901=>"000111010",
  3902=>"111100111",
  3903=>"100001010",
  3904=>"100111010",
  3905=>"011001011",
  3906=>"011001011",
  3907=>"110001001",
  3908=>"110010000",
  3909=>"100110010",
  3910=>"100100001",
  3911=>"110011110",
  3912=>"000010100",
  3913=>"011010110",
  3914=>"110111100",
  3915=>"100000110",
  3916=>"010011010",
  3917=>"000101011",
  3918=>"111001100",
  3919=>"011110101",
  3920=>"011111001",
  3921=>"001100111",
  3922=>"100110010",
  3923=>"100011110",
  3924=>"010011011",
  3925=>"110011111",
  3926=>"110001111",
  3927=>"110100010",
  3928=>"011100111",
  3929=>"001011000",
  3930=>"001111011",
  3931=>"001000101",
  3932=>"100111100",
  3933=>"011010010",
  3934=>"111111001",
  3935=>"101000110",
  3936=>"111110110",
  3937=>"101111100",
  3938=>"011111101",
  3939=>"011010011",
  3940=>"101101101",
  3941=>"010111000",
  3942=>"011011100",
  3943=>"111101110",
  3944=>"010110010",
  3945=>"001110010",
  3946=>"101100010",
  3947=>"010111111",
  3948=>"110011000",
  3949=>"111100001",
  3950=>"110101011",
  3951=>"100100010",
  3952=>"101010001",
  3953=>"111010011",
  3954=>"010000100",
  3955=>"100100011",
  3956=>"100010110",
  3957=>"011100001",
  3958=>"011110010",
  3959=>"000110111",
  3960=>"000010111",
  3961=>"010100111",
  3962=>"101001111",
  3963=>"110001111",
  3964=>"100010010",
  3965=>"010010111",
  3966=>"101001100",
  3967=>"101010000",
  3968=>"111110011",
  3969=>"011011001",
  3970=>"010000110",
  3971=>"000010011",
  3972=>"011101110",
  3973=>"000100000",
  3974=>"000010010",
  3975=>"111100101",
  3976=>"000010111",
  3977=>"110001110",
  3978=>"010010000",
  3979=>"011011011",
  3980=>"110100110",
  3981=>"100101010",
  3982=>"010111100",
  3983=>"110111101",
  3984=>"000111110",
  3985=>"110101010",
  3986=>"110001010",
  3987=>"110101000",
  3988=>"000010000",
  3989=>"111010111",
  3990=>"101100010",
  3991=>"011100101",
  3992=>"101000101",
  3993=>"011101011",
  3994=>"111010010",
  3995=>"010101100",
  3996=>"010011101",
  3997=>"001010000",
  3998=>"101110001",
  3999=>"010001000",
  4000=>"010100010",
  4001=>"110100001",
  4002=>"110011101",
  4003=>"110011100",
  4004=>"001101010",
  4005=>"101100110",
  4006=>"101110111",
  4007=>"001111111",
  4008=>"001000010",
  4009=>"110101011",
  4010=>"000010000",
  4011=>"100111000",
  4012=>"000111110",
  4013=>"000111100",
  4014=>"001110001",
  4015=>"111010110",
  4016=>"001111010",
  4017=>"111001011",
  4018=>"000011111",
  4019=>"000011101",
  4020=>"111010010",
  4021=>"000100110",
  4022=>"101010111",
  4023=>"011000001",
  4024=>"011111110",
  4025=>"111000001",
  4026=>"001010001",
  4027=>"101110010",
  4028=>"010011011",
  4029=>"010010011",
  4030=>"100110101",
  4031=>"011010011",
  4032=>"010101111",
  4033=>"011101100",
  4034=>"011110101",
  4035=>"111111101",
  4036=>"100000100",
  4037=>"100001101",
  4038=>"101110010",
  4039=>"101101010",
  4040=>"000000101",
  4041=>"110010100",
  4042=>"001000110",
  4043=>"111110010",
  4044=>"101110011",
  4045=>"011100010",
  4046=>"111100100",
  4047=>"111111001",
  4048=>"010000010",
  4049=>"001110011",
  4050=>"000101010",
  4051=>"011100010",
  4052=>"001110001",
  4053=>"111001110",
  4054=>"010101000",
  4055=>"000010011",
  4056=>"110110000",
  4057=>"111001010",
  4058=>"000111010",
  4059=>"100111111",
  4060=>"011111011",
  4061=>"011001010",
  4062=>"000111000",
  4063=>"101000011",
  4064=>"000000100",
  4065=>"101110101",
  4066=>"110101110",
  4067=>"010110010",
  4068=>"110000100",
  4069=>"101111011",
  4070=>"110110110",
  4071=>"111011111",
  4072=>"110000000",
  4073=>"111000111",
  4074=>"101100110",
  4075=>"001000011",
  4076=>"000011100",
  4077=>"010011110",
  4078=>"011000011",
  4079=>"000100000",
  4080=>"000100000",
  4081=>"001000010",
  4082=>"011001000",
  4083=>"100011011",
  4084=>"010110000",
  4085=>"100111110",
  4086=>"110110011",
  4087=>"111000010",
  4088=>"101111011",
  4089=>"000001010",
  4090=>"101010101",
  4091=>"000010110",
  4092=>"111110000",
  4093=>"100110000",
  4094=>"000101011",
  4095=>"111101100",
  4096=>"001100010",
  4097=>"000111010",
  4098=>"011011101",
  4099=>"001000110",
  4100=>"010010001",
  4101=>"010011010",
  4102=>"101111010",
  4103=>"111111110",
  4104=>"000100101",
  4105=>"000101011",
  4106=>"101110110",
  4107=>"110010101",
  4108=>"100111000",
  4109=>"111110011",
  4110=>"111110111",
  4111=>"010000011",
  4112=>"010011001",
  4113=>"011000111",
  4114=>"110011011",
  4115=>"001001010",
  4116=>"111001100",
  4117=>"110101111",
  4118=>"000010001",
  4119=>"111100000",
  4120=>"101000011",
  4121=>"101100101",
  4122=>"010111100",
  4123=>"011101000",
  4124=>"111110101",
  4125=>"110111111",
  4126=>"011110011",
  4127=>"000010010",
  4128=>"101111100",
  4129=>"110111101",
  4130=>"010111000",
  4131=>"011100011",
  4132=>"110111010",
  4133=>"011110000",
  4134=>"100010001",
  4135=>"011100110",
  4136=>"110011011",
  4137=>"101110110",
  4138=>"111010010",
  4139=>"010110101",
  4140=>"111001111",
  4141=>"000101011",
  4142=>"111000110",
  4143=>"110100000",
  4144=>"001111100",
  4145=>"111101011",
  4146=>"011101101",
  4147=>"010111010",
  4148=>"010001010",
  4149=>"100111110",
  4150=>"001010110",
  4151=>"011000110",
  4152=>"011111011",
  4153=>"100000110",
  4154=>"111111101",
  4155=>"101010110",
  4156=>"101001110",
  4157=>"000001001",
  4158=>"110110101",
  4159=>"100111000",
  4160=>"001100000",
  4161=>"011100100",
  4162=>"000100000",
  4163=>"011100101",
  4164=>"100001100",
  4165=>"010101111",
  4166=>"000001101",
  4167=>"010010001",
  4168=>"001001011",
  4169=>"011000010",
  4170=>"111101100",
  4171=>"011111111",
  4172=>"101010010",
  4173=>"111011101",
  4174=>"101100001",
  4175=>"111100011",
  4176=>"101111110",
  4177=>"111101101",
  4178=>"100111100",
  4179=>"110110010",
  4180=>"100101000",
  4181=>"000000000",
  4182=>"111010001",
  4183=>"000111100",
  4184=>"111000000",
  4185=>"100011010",
  4186=>"101111110",
  4187=>"111111011",
  4188=>"001011111",
  4189=>"101100011",
  4190=>"111100101",
  4191=>"000010000",
  4192=>"101100111",
  4193=>"100100001",
  4194=>"101010111",
  4195=>"010011110",
  4196=>"100001110",
  4197=>"111001110",
  4198=>"111101000",
  4199=>"000001101",
  4200=>"101111001",
  4201=>"101110110",
  4202=>"001100000",
  4203=>"101010111",
  4204=>"101011011",
  4205=>"111111101",
  4206=>"000000001",
  4207=>"101011001",
  4208=>"010110110",
  4209=>"000010000",
  4210=>"111111001",
  4211=>"000001001",
  4212=>"101000001",
  4213=>"010000110",
  4214=>"001000100",
  4215=>"111111100",
  4216=>"101100000",
  4217=>"111011101",
  4218=>"100010011",
  4219=>"100100100",
  4220=>"101001100",
  4221=>"100000110",
  4222=>"011100010",
  4223=>"101000110",
  4224=>"011001001",
  4225=>"010100010",
  4226=>"000011110",
  4227=>"000110011",
  4228=>"100000010",
  4229=>"001100111",
  4230=>"011010111",
  4231=>"010111000",
  4232=>"111111100",
  4233=>"100101011",
  4234=>"000010101",
  4235=>"000011011",
  4236=>"011100100",
  4237=>"101010101",
  4238=>"111100000",
  4239=>"111010001",
  4240=>"101111101",
  4241=>"111111011",
  4242=>"110011100",
  4243=>"011101000",
  4244=>"010000000",
  4245=>"111110100",
  4246=>"010100010",
  4247=>"101011110",
  4248=>"011111001",
  4249=>"101100001",
  4250=>"000101010",
  4251=>"000010001",
  4252=>"110010000",
  4253=>"001101000",
  4254=>"011111101",
  4255=>"100011011",
  4256=>"011111111",
  4257=>"100101111",
  4258=>"001101100",
  4259=>"111100001",
  4260=>"111101100",
  4261=>"101010110",
  4262=>"101001100",
  4263=>"100100111",
  4264=>"010010011",
  4265=>"010101010",
  4266=>"000000100",
  4267=>"111100101",
  4268=>"110110100",
  4269=>"011010001",
  4270=>"010111000",
  4271=>"001000011",
  4272=>"011100110",
  4273=>"000101111",
  4274=>"110100111",
  4275=>"101110000",
  4276=>"001111111",
  4277=>"101101100",
  4278=>"010011100",
  4279=>"101110101",
  4280=>"000001010",
  4281=>"110110011",
  4282=>"100010010",
  4283=>"101011111",
  4284=>"001010011",
  4285=>"100101111",
  4286=>"010000100",
  4287=>"111101011",
  4288=>"001001111",
  4289=>"000101111",
  4290=>"100100000",
  4291=>"111110010",
  4292=>"011110010",
  4293=>"000001110",
  4294=>"110111111",
  4295=>"110110111",
  4296=>"101011010",
  4297=>"111001011",
  4298=>"010101001",
  4299=>"001010111",
  4300=>"010111011",
  4301=>"001101110",
  4302=>"011111100",
  4303=>"111011100",
  4304=>"010010011",
  4305=>"100101011",
  4306=>"101010010",
  4307=>"111011001",
  4308=>"000110110",
  4309=>"110010011",
  4310=>"101010010",
  4311=>"100010000",
  4312=>"111000010",
  4313=>"010010011",
  4314=>"011110000",
  4315=>"011000001",
  4316=>"110100111",
  4317=>"111101101",
  4318=>"001111001",
  4319=>"000110000",
  4320=>"101100001",
  4321=>"111101010",
  4322=>"100111000",
  4323=>"111011100",
  4324=>"011011101",
  4325=>"100001100",
  4326=>"100100101",
  4327=>"010111010",
  4328=>"000000011",
  4329=>"010100010",
  4330=>"011100011",
  4331=>"111110111",
  4332=>"101000010",
  4333=>"110010110",
  4334=>"011011100",
  4335=>"000110000",
  4336=>"110001101",
  4337=>"101101111",
  4338=>"101011001",
  4339=>"001000111",
  4340=>"001011110",
  4341=>"111001100",
  4342=>"111110101",
  4343=>"010100000",
  4344=>"001010110",
  4345=>"110011101",
  4346=>"001110101",
  4347=>"001000110",
  4348=>"110100011",
  4349=>"000111100",
  4350=>"001101100",
  4351=>"001010011",
  4352=>"100011111",
  4353=>"001101100",
  4354=>"111111100",
  4355=>"010100001",
  4356=>"000101010",
  4357=>"010000110",
  4358=>"001110001",
  4359=>"100101001",
  4360=>"100110000",
  4361=>"000111011",
  4362=>"010101010",
  4363=>"101010001",
  4364=>"011000011",
  4365=>"100110010",
  4366=>"010110000",
  4367=>"001100111",
  4368=>"101001100",
  4369=>"101000010",
  4370=>"110100110",
  4371=>"011100110",
  4372=>"010101111",
  4373=>"001011011",
  4374=>"011010111",
  4375=>"111110001",
  4376=>"101101001",
  4377=>"001110000",
  4378=>"111010010",
  4379=>"011001111",
  4380=>"000000110",
  4381=>"000010101",
  4382=>"100010100",
  4383=>"100011011",
  4384=>"111010111",
  4385=>"110100000",
  4386=>"000110100",
  4387=>"011011111",
  4388=>"000100000",
  4389=>"001010000",
  4390=>"101110110",
  4391=>"110010111",
  4392=>"111001100",
  4393=>"101011010",
  4394=>"110100111",
  4395=>"001100001",
  4396=>"101101101",
  4397=>"000001100",
  4398=>"101111111",
  4399=>"001111000",
  4400=>"110001110",
  4401=>"000101001",
  4402=>"100011010",
  4403=>"011010110",
  4404=>"010111100",
  4405=>"100001100",
  4406=>"010100011",
  4407=>"111000010",
  4408=>"001010010",
  4409=>"011101011",
  4410=>"010000010",
  4411=>"000111000",
  4412=>"000111110",
  4413=>"101101110",
  4414=>"010100100",
  4415=>"100101011",
  4416=>"011011101",
  4417=>"000101001",
  4418=>"110000001",
  4419=>"001011110",
  4420=>"100010101",
  4421=>"011110111",
  4422=>"000011110",
  4423=>"001000111",
  4424=>"100001001",
  4425=>"100111110",
  4426=>"111100010",
  4427=>"001010000",
  4428=>"111000111",
  4429=>"011111111",
  4430=>"110110010",
  4431=>"011110100",
  4432=>"010000001",
  4433=>"100000110",
  4434=>"100110110",
  4435=>"100000011",
  4436=>"101000010",
  4437=>"000101011",
  4438=>"110110010",
  4439=>"010111101",
  4440=>"111010111",
  4441=>"001101000",
  4442=>"100011000",
  4443=>"101100010",
  4444=>"001110101",
  4445=>"111011000",
  4446=>"011110000",
  4447=>"101001100",
  4448=>"011111000",
  4449=>"001111111",
  4450=>"000111011",
  4451=>"001111111",
  4452=>"110001011",
  4453=>"110100110",
  4454=>"000111101",
  4455=>"010111011",
  4456=>"011000011",
  4457=>"001111111",
  4458=>"001111110",
  4459=>"101100001",
  4460=>"111000001",
  4461=>"100001000",
  4462=>"101010111",
  4463=>"011011111",
  4464=>"110110001",
  4465=>"001101001",
  4466=>"000010010",
  4467=>"110000001",
  4468=>"000011101",
  4469=>"110001101",
  4470=>"001100001",
  4471=>"110000100",
  4472=>"001110100",
  4473=>"011000100",
  4474=>"001010001",
  4475=>"011100011",
  4476=>"111001101",
  4477=>"111111111",
  4478=>"111101011",
  4479=>"101001001",
  4480=>"110001111",
  4481=>"001001111",
  4482=>"101110100",
  4483=>"000100001",
  4484=>"100100101",
  4485=>"000000100",
  4486=>"110011011",
  4487=>"010010001",
  4488=>"000011011",
  4489=>"111111110",
  4490=>"100101100",
  4491=>"011001001",
  4492=>"100101100",
  4493=>"111100110",
  4494=>"001100101",
  4495=>"100001101",
  4496=>"001110110",
  4497=>"100110110",
  4498=>"010001010",
  4499=>"110111000",
  4500=>"101110010",
  4501=>"000011110",
  4502=>"000000000",
  4503=>"101011010",
  4504=>"011110101",
  4505=>"111101011",
  4506=>"110110111",
  4507=>"010001111",
  4508=>"011100011",
  4509=>"100010111",
  4510=>"000100001",
  4511=>"110010110",
  4512=>"000011100",
  4513=>"100111011",
  4514=>"011111001",
  4515=>"010110110",
  4516=>"000100110",
  4517=>"001011000",
  4518=>"110010100",
  4519=>"000011101",
  4520=>"110111101",
  4521=>"011110000",
  4522=>"111111000",
  4523=>"110010110",
  4524=>"111100110",
  4525=>"000001101",
  4526=>"110101011",
  4527=>"110100010",
  4528=>"011010000",
  4529=>"001111010",
  4530=>"001111111",
  4531=>"001000000",
  4532=>"110010111",
  4533=>"111111100",
  4534=>"111000110",
  4535=>"011011000",
  4536=>"111111010",
  4537=>"111000011",
  4538=>"001110010",
  4539=>"110000010",
  4540=>"101100101",
  4541=>"011001101",
  4542=>"001000100",
  4543=>"010000000",
  4544=>"101001100",
  4545=>"100000010",
  4546=>"010111110",
  4547=>"010000010",
  4548=>"011010101",
  4549=>"111100110",
  4550=>"110101111",
  4551=>"100110100",
  4552=>"100000001",
  4553=>"000100100",
  4554=>"101011011",
  4555=>"111101010",
  4556=>"111011000",
  4557=>"110011000",
  4558=>"100111111",
  4559=>"011100001",
  4560=>"111111000",
  4561=>"001001011",
  4562=>"110111100",
  4563=>"100100101",
  4564=>"101110110",
  4565=>"100001110",
  4566=>"000001101",
  4567=>"111100101",
  4568=>"011011111",
  4569=>"101000110",
  4570=>"111000001",
  4571=>"101001000",
  4572=>"010011011",
  4573=>"001111001",
  4574=>"111000011",
  4575=>"001111110",
  4576=>"011010110",
  4577=>"110010100",
  4578=>"110110001",
  4579=>"100011011",
  4580=>"011100000",
  4581=>"000001010",
  4582=>"011010001",
  4583=>"001110001",
  4584=>"101000010",
  4585=>"111001100",
  4586=>"000111010",
  4587=>"101100000",
  4588=>"000000001",
  4589=>"101001100",
  4590=>"000100011",
  4591=>"101010011",
  4592=>"010111110",
  4593=>"010100011",
  4594=>"111001000",
  4595=>"000100101",
  4596=>"111100110",
  4597=>"110111111",
  4598=>"111000000",
  4599=>"101010001",
  4600=>"000110111",
  4601=>"110010000",
  4602=>"100110000",
  4603=>"100010000",
  4604=>"101011110",
  4605=>"010101101",
  4606=>"111100101",
  4607=>"101111101",
  4608=>"010010100",
  4609=>"000011111",
  4610=>"100010010",
  4611=>"001010000",
  4612=>"011000100",
  4613=>"101101111",
  4614=>"111100001",
  4615=>"010111000",
  4616=>"101000010",
  4617=>"010101110",
  4618=>"100111101",
  4619=>"110011011",
  4620=>"001000000",
  4621=>"010011110",
  4622=>"111000010",
  4623=>"110110010",
  4624=>"000110001",
  4625=>"011100011",
  4626=>"101100110",
  4627=>"101000000",
  4628=>"010010001",
  4629=>"011001001",
  4630=>"110010010",
  4631=>"001110011",
  4632=>"110110001",
  4633=>"100010100",
  4634=>"001100000",
  4635=>"011001100",
  4636=>"100100010",
  4637=>"110101110",
  4638=>"110011100",
  4639=>"110101111",
  4640=>"001010101",
  4641=>"001000000",
  4642=>"000010110",
  4643=>"101100011",
  4644=>"101011101",
  4645=>"010101011",
  4646=>"010001011",
  4647=>"010001111",
  4648=>"111001111",
  4649=>"100000010",
  4650=>"111111011",
  4651=>"111101111",
  4652=>"011010110",
  4653=>"100110101",
  4654=>"000010101",
  4655=>"111110011",
  4656=>"000100110",
  4657=>"011111110",
  4658=>"010111001",
  4659=>"011000110",
  4660=>"010011000",
  4661=>"000111101",
  4662=>"100111010",
  4663=>"000111101",
  4664=>"000001101",
  4665=>"111111000",
  4666=>"001010001",
  4667=>"000001010",
  4668=>"010101000",
  4669=>"000000000",
  4670=>"001011010",
  4671=>"101100001",
  4672=>"111010111",
  4673=>"001110010",
  4674=>"001000101",
  4675=>"001100101",
  4676=>"101000001",
  4677=>"011111100",
  4678=>"101001111",
  4679=>"010010011",
  4680=>"011101100",
  4681=>"011100001",
  4682=>"101110111",
  4683=>"011101111",
  4684=>"010011010",
  4685=>"111011100",
  4686=>"000001101",
  4687=>"011011111",
  4688=>"110000101",
  4689=>"000110101",
  4690=>"101111110",
  4691=>"011110110",
  4692=>"100111111",
  4693=>"000001110",
  4694=>"000000000",
  4695=>"000011010",
  4696=>"101110110",
  4697=>"011100010",
  4698=>"100100000",
  4699=>"100101110",
  4700=>"100110100",
  4701=>"000010111",
  4702=>"111100000",
  4703=>"111000000",
  4704=>"000001111",
  4705=>"000110110",
  4706=>"110000100",
  4707=>"011011010",
  4708=>"001100101",
  4709=>"101010111",
  4710=>"111011001",
  4711=>"000010101",
  4712=>"000010000",
  4713=>"110011001",
  4714=>"101000001",
  4715=>"101110000",
  4716=>"100110001",
  4717=>"100100011",
  4718=>"110101110",
  4719=>"011101101",
  4720=>"100110101",
  4721=>"000001010",
  4722=>"000011000",
  4723=>"001010111",
  4724=>"111001101",
  4725=>"011100111",
  4726=>"010000000",
  4727=>"000111110",
  4728=>"001010101",
  4729=>"110110100",
  4730=>"001011111",
  4731=>"010111000",
  4732=>"110010001",
  4733=>"010111001",
  4734=>"011100110",
  4735=>"110100001",
  4736=>"011010111",
  4737=>"111001111",
  4738=>"010100101",
  4739=>"101111011",
  4740=>"110000010",
  4741=>"110110101",
  4742=>"111110111",
  4743=>"001101011",
  4744=>"000110100",
  4745=>"000100010",
  4746=>"001011000",
  4747=>"000111100",
  4748=>"000101111",
  4749=>"001011000",
  4750=>"110011110",
  4751=>"001011000",
  4752=>"100010010",
  4753=>"101001101",
  4754=>"001111101",
  4755=>"100111111",
  4756=>"111111010",
  4757=>"100011100",
  4758=>"010000100",
  4759=>"100011101",
  4760=>"010001010",
  4761=>"111001010",
  4762=>"010011000",
  4763=>"101010110",
  4764=>"000000000",
  4765=>"100100000",
  4766=>"100001110",
  4767=>"100011101",
  4768=>"100000001",
  4769=>"101100000",
  4770=>"111110001",
  4771=>"100011000",
  4772=>"010011111",
  4773=>"001011100",
  4774=>"001101011",
  4775=>"000000000",
  4776=>"000000011",
  4777=>"100001101",
  4778=>"010011101",
  4779=>"010110001",
  4780=>"010001000",
  4781=>"101100000",
  4782=>"110100101",
  4783=>"000001110",
  4784=>"001110010",
  4785=>"110100011",
  4786=>"000011001",
  4787=>"011000110",
  4788=>"111010000",
  4789=>"010101001",
  4790=>"110011001",
  4791=>"111111010",
  4792=>"001100001",
  4793=>"010100100",
  4794=>"110101011",
  4795=>"110100001",
  4796=>"000111101",
  4797=>"101000000",
  4798=>"011100001",
  4799=>"110011100",
  4800=>"100001111",
  4801=>"110110110",
  4802=>"111100011",
  4803=>"010101000",
  4804=>"011110010",
  4805=>"001101001",
  4806=>"111100001",
  4807=>"100001101",
  4808=>"000011100",
  4809=>"000111000",
  4810=>"100000000",
  4811=>"001000101",
  4812=>"100000010",
  4813=>"011011010",
  4814=>"101011100",
  4815=>"110100011",
  4816=>"100000101",
  4817=>"101110111",
  4818=>"011001100",
  4819=>"011111010",
  4820=>"110101100",
  4821=>"110101111",
  4822=>"000001000",
  4823=>"011000100",
  4824=>"000110011",
  4825=>"000001110",
  4826=>"000100011",
  4827=>"011111011",
  4828=>"101101111",
  4829=>"010001100",
  4830=>"110000010",
  4831=>"010101011",
  4832=>"111111000",
  4833=>"110000010",
  4834=>"110010111",
  4835=>"010010101",
  4836=>"001110011",
  4837=>"100000011",
  4838=>"000011110",
  4839=>"111110001",
  4840=>"110101100",
  4841=>"010111111",
  4842=>"011001010",
  4843=>"011111000",
  4844=>"001000100",
  4845=>"110011001",
  4846=>"100010110",
  4847=>"110101000",
  4848=>"100100111",
  4849=>"110011000",
  4850=>"000110000",
  4851=>"101110000",
  4852=>"001011011",
  4853=>"001111110",
  4854=>"100000010",
  4855=>"111000101",
  4856=>"111011101",
  4857=>"000010011",
  4858=>"011011000",
  4859=>"001010110",
  4860=>"000000010",
  4861=>"010100111",
  4862=>"000100000",
  4863=>"110101001",
  4864=>"001100001",
  4865=>"011110001",
  4866=>"010101001",
  4867=>"100110001",
  4868=>"111110011",
  4869=>"100001000",
  4870=>"101111010",
  4871=>"101010111",
  4872=>"011000011",
  4873=>"001111111",
  4874=>"010100000",
  4875=>"001000010",
  4876=>"101000111",
  4877=>"010101011",
  4878=>"110011100",
  4879=>"110110011",
  4880=>"011001111",
  4881=>"001010110",
  4882=>"010101100",
  4883=>"011000000",
  4884=>"110110001",
  4885=>"011010101",
  4886=>"111010100",
  4887=>"111010000",
  4888=>"010001001",
  4889=>"100011001",
  4890=>"110111000",
  4891=>"101111011",
  4892=>"110101110",
  4893=>"010100110",
  4894=>"100010100",
  4895=>"001101110",
  4896=>"001111011",
  4897=>"000010111",
  4898=>"010101110",
  4899=>"011000001",
  4900=>"110001100",
  4901=>"101000100",
  4902=>"010001001",
  4903=>"111110010",
  4904=>"111010110",
  4905=>"101000001",
  4906=>"101101100",
  4907=>"111001110",
  4908=>"110001100",
  4909=>"011110001",
  4910=>"111110110",
  4911=>"010111000",
  4912=>"011000011",
  4913=>"011100100",
  4914=>"101011000",
  4915=>"010110000",
  4916=>"111111111",
  4917=>"001111101",
  4918=>"011001111",
  4919=>"000111010",
  4920=>"101011101",
  4921=>"001111101",
  4922=>"101101010",
  4923=>"111110011",
  4924=>"111000010",
  4925=>"110101011",
  4926=>"000110110",
  4927=>"110011001",
  4928=>"101100001",
  4929=>"110110010",
  4930=>"001011011",
  4931=>"001110001",
  4932=>"100111011",
  4933=>"000000011",
  4934=>"001101101",
  4935=>"001010010",
  4936=>"110010101",
  4937=>"110110101",
  4938=>"101010011",
  4939=>"011110100",
  4940=>"111010111",
  4941=>"000001001",
  4942=>"000010101",
  4943=>"010011101",
  4944=>"110101001",
  4945=>"000111110",
  4946=>"000110110",
  4947=>"100000110",
  4948=>"010010111",
  4949=>"001000101",
  4950=>"101000010",
  4951=>"010101111",
  4952=>"000001100",
  4953=>"110111011",
  4954=>"001110100",
  4955=>"101001111",
  4956=>"001101010",
  4957=>"111101011",
  4958=>"000011000",
  4959=>"111000010",
  4960=>"101011110",
  4961=>"101110101",
  4962=>"101111010",
  4963=>"000110100",
  4964=>"001011001",
  4965=>"000011000",
  4966=>"110010000",
  4967=>"010100000",
  4968=>"001110111",
  4969=>"010110011",
  4970=>"010101010",
  4971=>"101011111",
  4972=>"100100111",
  4973=>"010000101",
  4974=>"101010111",
  4975=>"111011101",
  4976=>"001001000",
  4977=>"110110000",
  4978=>"110011110",
  4979=>"000011011",
  4980=>"100100010",
  4981=>"010000001",
  4982=>"001001111",
  4983=>"011011011",
  4984=>"000110001",
  4985=>"100100011",
  4986=>"011101010",
  4987=>"001111011",
  4988=>"000000000",
  4989=>"101000001",
  4990=>"110111110",
  4991=>"100010001",
  4992=>"111000101",
  4993=>"001100010",
  4994=>"110100100",
  4995=>"010101111",
  4996=>"110011011",
  4997=>"111110101",
  4998=>"100011000",
  4999=>"110111110",
  5000=>"010100001",
  5001=>"100000001",
  5002=>"000100111",
  5003=>"001111011",
  5004=>"000110110",
  5005=>"000001001",
  5006=>"101100001",
  5007=>"100101100",
  5008=>"100111110",
  5009=>"111100011",
  5010=>"001010100",
  5011=>"001111110",
  5012=>"010111101",
  5013=>"011000101",
  5014=>"100000000",
  5015=>"001011101",
  5016=>"010011010",
  5017=>"010011110",
  5018=>"001100011",
  5019=>"100001110",
  5020=>"100111010",
  5021=>"100000110",
  5022=>"110110101",
  5023=>"010100001",
  5024=>"101001000",
  5025=>"111000001",
  5026=>"000011110",
  5027=>"010001001",
  5028=>"011000001",
  5029=>"100110111",
  5030=>"010000101",
  5031=>"100011000",
  5032=>"000010001",
  5033=>"010000110",
  5034=>"011101110",
  5035=>"111101011",
  5036=>"001111001",
  5037=>"011110010",
  5038=>"001011111",
  5039=>"110011010",
  5040=>"111100010",
  5041=>"011010000",
  5042=>"011101001",
  5043=>"111010110",
  5044=>"011011001",
  5045=>"010011011",
  5046=>"100110000",
  5047=>"001100100",
  5048=>"101110110",
  5049=>"011011011",
  5050=>"000010010",
  5051=>"001100011",
  5052=>"110010010",
  5053=>"101111101",
  5054=>"000010001",
  5055=>"000100001",
  5056=>"111100111",
  5057=>"111010001",
  5058=>"111111011",
  5059=>"011010010",
  5060=>"110001011",
  5061=>"000001011",
  5062=>"000110001",
  5063=>"111100001",
  5064=>"001011011",
  5065=>"001101111",
  5066=>"001110010",
  5067=>"111110111",
  5068=>"100110101",
  5069=>"000000101",
  5070=>"010100010",
  5071=>"010000001",
  5072=>"111000100",
  5073=>"000100010",
  5074=>"000011010",
  5075=>"100111100",
  5076=>"111000111",
  5077=>"101011001",
  5078=>"111011001",
  5079=>"010111111",
  5080=>"101010111",
  5081=>"101001100",
  5082=>"111100001",
  5083=>"100000000",
  5084=>"000000000",
  5085=>"000100010",
  5086=>"100111101",
  5087=>"010111111",
  5088=>"100001011",
  5089=>"110111001",
  5090=>"110100111",
  5091=>"110000111",
  5092=>"110001110",
  5093=>"110111001",
  5094=>"101010001",
  5095=>"110001010",
  5096=>"001111001",
  5097=>"010101100",
  5098=>"001100101",
  5099=>"111100100",
  5100=>"101110100",
  5101=>"000101101",
  5102=>"110011110",
  5103=>"010011100",
  5104=>"011001000",
  5105=>"110100101",
  5106=>"101100111",
  5107=>"111111011",
  5108=>"001001110",
  5109=>"110000001",
  5110=>"000111111",
  5111=>"001001101",
  5112=>"001110001",
  5113=>"000011111",
  5114=>"100010111",
  5115=>"010000101",
  5116=>"000110010",
  5117=>"101000101",
  5118=>"000101101",
  5119=>"111111110",
  5120=>"101110110",
  5121=>"000011001",
  5122=>"100011011",
  5123=>"001111011",
  5124=>"010101000",
  5125=>"100001010",
  5126=>"111100010",
  5127=>"100110101",
  5128=>"111000110",
  5129=>"000111100",
  5130=>"000000110",
  5131=>"000011101",
  5132=>"001101100",
  5133=>"101001010",
  5134=>"011000100",
  5135=>"000001100",
  5136=>"010101001",
  5137=>"000010010",
  5138=>"101101000",
  5139=>"110101010",
  5140=>"100100011",
  5141=>"100011111",
  5142=>"100110110",
  5143=>"111011000",
  5144=>"010010110",
  5145=>"011000001",
  5146=>"111110110",
  5147=>"111001010",
  5148=>"001001010",
  5149=>"000011111",
  5150=>"011000000",
  5151=>"111111100",
  5152=>"110010010",
  5153=>"010011100",
  5154=>"011100010",
  5155=>"000101101",
  5156=>"001110110",
  5157=>"011110101",
  5158=>"010011100",
  5159=>"100001010",
  5160=>"111100111",
  5161=>"110011101",
  5162=>"100101011",
  5163=>"111000100",
  5164=>"000000011",
  5165=>"000101011",
  5166=>"000001000",
  5167=>"010101100",
  5168=>"010111011",
  5169=>"110001111",
  5170=>"011100001",
  5171=>"101000000",
  5172=>"101111101",
  5173=>"011111001",
  5174=>"100100000",
  5175=>"100011010",
  5176=>"000000000",
  5177=>"100111101",
  5178=>"110010010",
  5179=>"100001010",
  5180=>"110110011",
  5181=>"011000011",
  5182=>"110110100",
  5183=>"000110010",
  5184=>"000001100",
  5185=>"000001001",
  5186=>"101011011",
  5187=>"100110011",
  5188=>"011001001",
  5189=>"010000010",
  5190=>"101011001",
  5191=>"110010000",
  5192=>"110110101",
  5193=>"000011011",
  5194=>"010101001",
  5195=>"010100001",
  5196=>"010111000",
  5197=>"001101100",
  5198=>"101010111",
  5199=>"111110111",
  5200=>"101000111",
  5201=>"111100010",
  5202=>"101000111",
  5203=>"011101101",
  5204=>"111000100",
  5205=>"001010100",
  5206=>"100101001",
  5207=>"100001110",
  5208=>"010011111",
  5209=>"001011010",
  5210=>"010101010",
  5211=>"111010111",
  5212=>"010000001",
  5213=>"000001100",
  5214=>"101101101",
  5215=>"111101111",
  5216=>"000110000",
  5217=>"111011000",
  5218=>"101001111",
  5219=>"000101101",
  5220=>"001001100",
  5221=>"101110000",
  5222=>"100001101",
  5223=>"010010100",
  5224=>"010111001",
  5225=>"111101110",
  5226=>"010000010",
  5227=>"111000110",
  5228=>"100011001",
  5229=>"001000111",
  5230=>"001000100",
  5231=>"000011101",
  5232=>"101010011",
  5233=>"011011001",
  5234=>"010100010",
  5235=>"101001010",
  5236=>"000010101",
  5237=>"001011111",
  5238=>"011111110",
  5239=>"100010010",
  5240=>"100011001",
  5241=>"100100011",
  5242=>"111001001",
  5243=>"110100010",
  5244=>"011111010",
  5245=>"001001111",
  5246=>"011000000",
  5247=>"111011011",
  5248=>"111111011",
  5249=>"110000001",
  5250=>"010001011",
  5251=>"111010000",
  5252=>"110111001",
  5253=>"010111001",
  5254=>"101000010",
  5255=>"011111100",
  5256=>"110011010",
  5257=>"100100011",
  5258=>"110000101",
  5259=>"010000101",
  5260=>"111110011",
  5261=>"100010100",
  5262=>"001110101",
  5263=>"111001101",
  5264=>"100000010",
  5265=>"110110011",
  5266=>"111001001",
  5267=>"010101111",
  5268=>"110001101",
  5269=>"010111110",
  5270=>"000000011",
  5271=>"100010000",
  5272=>"000111100",
  5273=>"111111001",
  5274=>"110010110",
  5275=>"001000011",
  5276=>"000110010",
  5277=>"111010100",
  5278=>"010000100",
  5279=>"010101110",
  5280=>"001001010",
  5281=>"101011011",
  5282=>"010110100",
  5283=>"110110100",
  5284=>"110010111",
  5285=>"001001100",
  5286=>"111100100",
  5287=>"001110110",
  5288=>"011111100",
  5289=>"011001000",
  5290=>"101101010",
  5291=>"100101000",
  5292=>"001100011",
  5293=>"111001101",
  5294=>"011100111",
  5295=>"111011110",
  5296=>"001100001",
  5297=>"010001111",
  5298=>"111000000",
  5299=>"001010100",
  5300=>"111000100",
  5301=>"011000000",
  5302=>"001110111",
  5303=>"110010100",
  5304=>"110000000",
  5305=>"100011001",
  5306=>"010010110",
  5307=>"010000110",
  5308=>"001010001",
  5309=>"100100001",
  5310=>"101100011",
  5311=>"011001100",
  5312=>"111011111",
  5313=>"001111111",
  5314=>"000010110",
  5315=>"111100000",
  5316=>"001001111",
  5317=>"000101000",
  5318=>"000000101",
  5319=>"001001101",
  5320=>"101111011",
  5321=>"110000001",
  5322=>"011100101",
  5323=>"100000000",
  5324=>"101101111",
  5325=>"111011010",
  5326=>"001010000",
  5327=>"111001001",
  5328=>"100111101",
  5329=>"010001000",
  5330=>"011101010",
  5331=>"000100010",
  5332=>"001111001",
  5333=>"101000000",
  5334=>"000000100",
  5335=>"000111100",
  5336=>"000100100",
  5337=>"010011000",
  5338=>"010100101",
  5339=>"111000100",
  5340=>"011110000",
  5341=>"110000110",
  5342=>"010100100",
  5343=>"111100110",
  5344=>"110011000",
  5345=>"000001111",
  5346=>"000000101",
  5347=>"101101011",
  5348=>"000000001",
  5349=>"111111100",
  5350=>"010011010",
  5351=>"010010000",
  5352=>"000100010",
  5353=>"011000110",
  5354=>"100010010",
  5355=>"010111011",
  5356=>"101011100",
  5357=>"010000111",
  5358=>"111100010",
  5359=>"100110101",
  5360=>"111111101",
  5361=>"010111110",
  5362=>"010010000",
  5363=>"100111011",
  5364=>"001100100",
  5365=>"101101100",
  5366=>"001110111",
  5367=>"100000000",
  5368=>"111011010",
  5369=>"110010011",
  5370=>"011000111",
  5371=>"101111000",
  5372=>"000101001",
  5373=>"010001100",
  5374=>"101011010",
  5375=>"111011011",
  5376=>"010101100",
  5377=>"111001011",
  5378=>"111001011",
  5379=>"001001011",
  5380=>"111110111",
  5381=>"001011010",
  5382=>"001011010",
  5383=>"011011010",
  5384=>"101000001",
  5385=>"101011101",
  5386=>"110010101",
  5387=>"110101100",
  5388=>"110000010",
  5389=>"000101111",
  5390=>"100000011",
  5391=>"011101110",
  5392=>"011010111",
  5393=>"000101001",
  5394=>"111111110",
  5395=>"101001100",
  5396=>"110100110",
  5397=>"101011100",
  5398=>"111011111",
  5399=>"010100110",
  5400=>"010100010",
  5401=>"111011011",
  5402=>"100111000",
  5403=>"000011100",
  5404=>"101001010",
  5405=>"111010110",
  5406=>"111100101",
  5407=>"011110101",
  5408=>"001011000",
  5409=>"010001011",
  5410=>"000100110",
  5411=>"100000110",
  5412=>"010101111",
  5413=>"111100010",
  5414=>"011000111",
  5415=>"011001010",
  5416=>"011011001",
  5417=>"101111111",
  5418=>"001011111",
  5419=>"001101100",
  5420=>"101010000",
  5421=>"111101111",
  5422=>"000100101",
  5423=>"010100011",
  5424=>"000010011",
  5425=>"100000000",
  5426=>"111101111",
  5427=>"000010100",
  5428=>"001000010",
  5429=>"010000001",
  5430=>"011100011",
  5431=>"111100000",
  5432=>"000110000",
  5433=>"000011110",
  5434=>"011101111",
  5435=>"100010000",
  5436=>"111011011",
  5437=>"110010110",
  5438=>"110110111",
  5439=>"010010101",
  5440=>"101011110",
  5441=>"100001001",
  5442=>"111111101",
  5443=>"100111100",
  5444=>"011110110",
  5445=>"111000110",
  5446=>"100000100",
  5447=>"010000111",
  5448=>"110001110",
  5449=>"111000111",
  5450=>"001001101",
  5451=>"101110101",
  5452=>"111111110",
  5453=>"101100010",
  5454=>"001001011",
  5455=>"101000111",
  5456=>"101001110",
  5457=>"100001001",
  5458=>"001110000",
  5459=>"101110111",
  5460=>"010111001",
  5461=>"100100000",
  5462=>"010110110",
  5463=>"101010111",
  5464=>"010000001",
  5465=>"101101010",
  5466=>"111010011",
  5467=>"000110111",
  5468=>"001101101",
  5469=>"101101101",
  5470=>"010100001",
  5471=>"010000000",
  5472=>"110101001",
  5473=>"100101100",
  5474=>"010100110",
  5475=>"000000101",
  5476=>"110010000",
  5477=>"101100100",
  5478=>"110000110",
  5479=>"000001010",
  5480=>"001011101",
  5481=>"100000000",
  5482=>"111100110",
  5483=>"001010110",
  5484=>"100101111",
  5485=>"100101111",
  5486=>"000110111",
  5487=>"001000011",
  5488=>"000101101",
  5489=>"100111010",
  5490=>"001001101",
  5491=>"111100110",
  5492=>"000001101",
  5493=>"010110010",
  5494=>"001000001",
  5495=>"011100010",
  5496=>"011100100",
  5497=>"110011100",
  5498=>"010000101",
  5499=>"001101011",
  5500=>"011000010",
  5501=>"011100110",
  5502=>"100011101",
  5503=>"001000011",
  5504=>"100010100",
  5505=>"111000001",
  5506=>"100101111",
  5507=>"110101001",
  5508=>"011000011",
  5509=>"010010110",
  5510=>"000101011",
  5511=>"010110001",
  5512=>"100010101",
  5513=>"100001001",
  5514=>"111110001",
  5515=>"010010000",
  5516=>"110011111",
  5517=>"100001001",
  5518=>"000000001",
  5519=>"100101011",
  5520=>"011101110",
  5521=>"010010000",
  5522=>"000011010",
  5523=>"111110001",
  5524=>"000010110",
  5525=>"110001001",
  5526=>"111111101",
  5527=>"101001111",
  5528=>"010000110",
  5529=>"111000111",
  5530=>"101010000",
  5531=>"010001100",
  5532=>"111001000",
  5533=>"000100101",
  5534=>"101011111",
  5535=>"010111000",
  5536=>"000100001",
  5537=>"100010001",
  5538=>"101011100",
  5539=>"110100011",
  5540=>"100111101",
  5541=>"101000001",
  5542=>"100111011",
  5543=>"010011101",
  5544=>"010111111",
  5545=>"111110110",
  5546=>"000010000",
  5547=>"010010010",
  5548=>"011111000",
  5549=>"111100100",
  5550=>"010000101",
  5551=>"000110001",
  5552=>"100011011",
  5553=>"010101011",
  5554=>"010010101",
  5555=>"101100100",
  5556=>"100011100",
  5557=>"001010011",
  5558=>"100100100",
  5559=>"010011010",
  5560=>"100101111",
  5561=>"000001010",
  5562=>"011000101",
  5563=>"111110001",
  5564=>"110111010",
  5565=>"000001111",
  5566=>"010111100",
  5567=>"101001111",
  5568=>"101100101",
  5569=>"100101101",
  5570=>"110000111",
  5571=>"001001010",
  5572=>"000101011",
  5573=>"011111101",
  5574=>"011001000",
  5575=>"101000000",
  5576=>"001000010",
  5577=>"110101100",
  5578=>"001001001",
  5579=>"111001111",
  5580=>"011011001",
  5581=>"010001011",
  5582=>"000010110",
  5583=>"111111110",
  5584=>"111011100",
  5585=>"011111011",
  5586=>"010110010",
  5587=>"001001010",
  5588=>"101000100",
  5589=>"100010101",
  5590=>"000000010",
  5591=>"100001001",
  5592=>"100001000",
  5593=>"000011010",
  5594=>"010110001",
  5595=>"101100100",
  5596=>"011011101",
  5597=>"001010100",
  5598=>"010100000",
  5599=>"111100010",
  5600=>"100000111",
  5601=>"000001100",
  5602=>"011101101",
  5603=>"000000011",
  5604=>"110101110",
  5605=>"100000111",
  5606=>"001011111",
  5607=>"001100010",
  5608=>"111110010",
  5609=>"011101000",
  5610=>"010000101",
  5611=>"001000001",
  5612=>"001110111",
  5613=>"001101001",
  5614=>"000000010",
  5615=>"101100110",
  5616=>"011100100",
  5617=>"000000011",
  5618=>"101101010",
  5619=>"100010001",
  5620=>"010100101",
  5621=>"011011001",
  5622=>"001000101",
  5623=>"101011001",
  5624=>"010101001",
  5625=>"001000110",
  5626=>"101000011",
  5627=>"101001001",
  5628=>"100011111",
  5629=>"000111001",
  5630=>"111001001",
  5631=>"101110101",
  5632=>"010001111",
  5633=>"010001011",
  5634=>"110111010",
  5635=>"011001101",
  5636=>"110110101",
  5637=>"000010000",
  5638=>"001101001",
  5639=>"001101010",
  5640=>"010101100",
  5641=>"010011101",
  5642=>"010011000",
  5643=>"110011111",
  5644=>"001010111",
  5645=>"110101001",
  5646=>"111010011",
  5647=>"110101010",
  5648=>"110010100",
  5649=>"101000100",
  5650=>"100001000",
  5651=>"111000111",
  5652=>"100010001",
  5653=>"100100110",
  5654=>"111100111",
  5655=>"011011010",
  5656=>"111010100",
  5657=>"101010011",
  5658=>"101101101",
  5659=>"000100011",
  5660=>"000000000",
  5661=>"111101001",
  5662=>"110101011",
  5663=>"000010001",
  5664=>"111100100",
  5665=>"101100101",
  5666=>"000001000",
  5667=>"101000001",
  5668=>"101000101",
  5669=>"000101011",
  5670=>"111011110",
  5671=>"000011100",
  5672=>"010100001",
  5673=>"100001000",
  5674=>"000000000",
  5675=>"001000001",
  5676=>"101011001",
  5677=>"000100011",
  5678=>"001010110",
  5679=>"001101111",
  5680=>"110001000",
  5681=>"101010001",
  5682=>"001111011",
  5683=>"000000010",
  5684=>"000010101",
  5685=>"101010111",
  5686=>"000001110",
  5687=>"000000110",
  5688=>"100101010",
  5689=>"000000101",
  5690=>"101010011",
  5691=>"100100011",
  5692=>"100010010",
  5693=>"011011111",
  5694=>"010101111",
  5695=>"010100110",
  5696=>"011101100",
  5697=>"001000000",
  5698=>"010000111",
  5699=>"010010011",
  5700=>"100011111",
  5701=>"101011110",
  5702=>"101100011",
  5703=>"100100100",
  5704=>"110010000",
  5705=>"011010000",
  5706=>"110011101",
  5707=>"011001000",
  5708=>"101100101",
  5709=>"101000001",
  5710=>"100101010",
  5711=>"010111101",
  5712=>"010111011",
  5713=>"010110000",
  5714=>"110110101",
  5715=>"000000111",
  5716=>"000000011",
  5717=>"110000011",
  5718=>"110111111",
  5719=>"101110110",
  5720=>"010001111",
  5721=>"001000110",
  5722=>"001000101",
  5723=>"000000100",
  5724=>"001011000",
  5725=>"100000101",
  5726=>"101110010",
  5727=>"100110010",
  5728=>"010010111",
  5729=>"110101101",
  5730=>"111000011",
  5731=>"000001111",
  5732=>"000101010",
  5733=>"100101101",
  5734=>"111001011",
  5735=>"011101001",
  5736=>"101111101",
  5737=>"010101000",
  5738=>"010011110",
  5739=>"100011010",
  5740=>"100000101",
  5741=>"011100100",
  5742=>"110100110",
  5743=>"101100111",
  5744=>"101001001",
  5745=>"111101000",
  5746=>"000011001",
  5747=>"000011000",
  5748=>"010000000",
  5749=>"100000110",
  5750=>"010000110",
  5751=>"001000011",
  5752=>"011101010",
  5753=>"100011110",
  5754=>"001110111",
  5755=>"000000000",
  5756=>"000001000",
  5757=>"110011011",
  5758=>"101001100",
  5759=>"101011101",
  5760=>"111001011",
  5761=>"100111100",
  5762=>"000001010",
  5763=>"010111001",
  5764=>"111110010",
  5765=>"100101111",
  5766=>"001110001",
  5767=>"100101111",
  5768=>"100110011",
  5769=>"101111001",
  5770=>"101100110",
  5771=>"000100010",
  5772=>"000100011",
  5773=>"001000101",
  5774=>"001010100",
  5775=>"100010110",
  5776=>"110010011",
  5777=>"111010001",
  5778=>"011110110",
  5779=>"010100110",
  5780=>"000101111",
  5781=>"110000011",
  5782=>"111000011",
  5783=>"010100110",
  5784=>"110111110",
  5785=>"000101101",
  5786=>"011101111",
  5787=>"001111110",
  5788=>"100000001",
  5789=>"100101111",
  5790=>"110001001",
  5791=>"000110111",
  5792=>"000100111",
  5793=>"011001111",
  5794=>"001001011",
  5795=>"101111101",
  5796=>"001110011",
  5797=>"110111111",
  5798=>"001000011",
  5799=>"000000100",
  5800=>"000100000",
  5801=>"110000011",
  5802=>"100001100",
  5803=>"000001001",
  5804=>"100000111",
  5805=>"000111000",
  5806=>"110111000",
  5807=>"011000000",
  5808=>"100100101",
  5809=>"001111111",
  5810=>"111100000",
  5811=>"011100100",
  5812=>"010101100",
  5813=>"111101000",
  5814=>"010101100",
  5815=>"110001100",
  5816=>"011000000",
  5817=>"110110101",
  5818=>"001000000",
  5819=>"001101010",
  5820=>"101110001",
  5821=>"100100110",
  5822=>"001110100",
  5823=>"011010111",
  5824=>"011001001",
  5825=>"111011000",
  5826=>"000110011",
  5827=>"001011101",
  5828=>"001010110",
  5829=>"011001110",
  5830=>"101010010",
  5831=>"101101001",
  5832=>"101101000",
  5833=>"000001000",
  5834=>"111010001",
  5835=>"000100001",
  5836=>"100001011",
  5837=>"100111011",
  5838=>"100011101",
  5839=>"011100001",
  5840=>"001110001",
  5841=>"011111110",
  5842=>"111110111",
  5843=>"101101101",
  5844=>"101101000",
  5845=>"000111011",
  5846=>"000010111",
  5847=>"111011101",
  5848=>"001010100",
  5849=>"001111001",
  5850=>"000110000",
  5851=>"011110001",
  5852=>"110101000",
  5853=>"000110000",
  5854=>"011100010",
  5855=>"100100111",
  5856=>"100000010",
  5857=>"011100011",
  5858=>"100101011",
  5859=>"011000010",
  5860=>"100110110",
  5861=>"010111010",
  5862=>"111100111",
  5863=>"000111010",
  5864=>"001111101",
  5865=>"010110100",
  5866=>"011110100",
  5867=>"001110001",
  5868=>"100001110",
  5869=>"111010111",
  5870=>"100110100",
  5871=>"100000110",
  5872=>"111101111",
  5873=>"101100111",
  5874=>"010010101",
  5875=>"101010000",
  5876=>"111011111",
  5877=>"011010010",
  5878=>"100000010",
  5879=>"001111010",
  5880=>"010011101",
  5881=>"001000111",
  5882=>"010010100",
  5883=>"011110010",
  5884=>"010111001",
  5885=>"010110000",
  5886=>"010100100",
  5887=>"101001010",
  5888=>"001010000",
  5889=>"011100001",
  5890=>"011111011",
  5891=>"111010011",
  5892=>"000101000",
  5893=>"001110010",
  5894=>"010011101",
  5895=>"001111100",
  5896=>"100010110",
  5897=>"101111110",
  5898=>"101010101",
  5899=>"100101000",
  5900=>"000011010",
  5901=>"111000010",
  5902=>"110001001",
  5903=>"110000100",
  5904=>"100101100",
  5905=>"011001110",
  5906=>"000000010",
  5907=>"101000000",
  5908=>"111101110",
  5909=>"001011111",
  5910=>"010011001",
  5911=>"011001000",
  5912=>"011000101",
  5913=>"000000100",
  5914=>"101101001",
  5915=>"010011000",
  5916=>"011010111",
  5917=>"011001001",
  5918=>"110010101",
  5919=>"111111010",
  5920=>"110010100",
  5921=>"111111100",
  5922=>"011000001",
  5923=>"011111010",
  5924=>"000010001",
  5925=>"111101010",
  5926=>"001010100",
  5927=>"011000110",
  5928=>"110101000",
  5929=>"001000101",
  5930=>"000110110",
  5931=>"111101110",
  5932=>"100100111",
  5933=>"111111110",
  5934=>"100010011",
  5935=>"111101101",
  5936=>"001010111",
  5937=>"110000010",
  5938=>"001000001",
  5939=>"000010110",
  5940=>"011100111",
  5941=>"111010011",
  5942=>"101111111",
  5943=>"001010100",
  5944=>"011010111",
  5945=>"101011110",
  5946=>"101100011",
  5947=>"111111001",
  5948=>"110100100",
  5949=>"111110111",
  5950=>"010101101",
  5951=>"111011101",
  5952=>"100011111",
  5953=>"111111100",
  5954=>"101000101",
  5955=>"111101111",
  5956=>"100001110",
  5957=>"111110000",
  5958=>"110100010",
  5959=>"110001101",
  5960=>"101111111",
  5961=>"001111010",
  5962=>"000111100",
  5963=>"010000000",
  5964=>"000100110",
  5965=>"010000110",
  5966=>"110100011",
  5967=>"101101100",
  5968=>"010101110",
  5969=>"001001111",
  5970=>"011111000",
  5971=>"001010111",
  5972=>"000011001",
  5973=>"101101010",
  5974=>"001001111",
  5975=>"000101011",
  5976=>"001101111",
  5977=>"000100111",
  5978=>"010010010",
  5979=>"010110010",
  5980=>"010110000",
  5981=>"101001111",
  5982=>"111110110",
  5983=>"011010010",
  5984=>"101111101",
  5985=>"001111000",
  5986=>"000001011",
  5987=>"110100110",
  5988=>"100011010",
  5989=>"111010001",
  5990=>"010101100",
  5991=>"000011010",
  5992=>"010111101",
  5993=>"101010001",
  5994=>"001001111",
  5995=>"001101110",
  5996=>"100011110",
  5997=>"011111101",
  5998=>"010110000",
  5999=>"110101100",
  6000=>"100111100",
  6001=>"000011000",
  6002=>"111110101",
  6003=>"011100111",
  6004=>"010000111",
  6005=>"000101010",
  6006=>"100010011",
  6007=>"010000011",
  6008=>"001011001",
  6009=>"011101010",
  6010=>"010111011",
  6011=>"000111010",
  6012=>"001001110",
  6013=>"111100000",
  6014=>"010010111",
  6015=>"101011110",
  6016=>"001101010",
  6017=>"101110101",
  6018=>"010011110",
  6019=>"110111001",
  6020=>"000010101",
  6021=>"100110011",
  6022=>"101011000",
  6023=>"111110100",
  6024=>"011101001",
  6025=>"000101110",
  6026=>"010111110",
  6027=>"011010111",
  6028=>"110101101",
  6029=>"010001101",
  6030=>"011011100",
  6031=>"101101000",
  6032=>"000001001",
  6033=>"001111111",
  6034=>"001001100",
  6035=>"001011000",
  6036=>"011011100",
  6037=>"101001010",
  6038=>"000010110",
  6039=>"100111010",
  6040=>"111001100",
  6041=>"111111011",
  6042=>"010111001",
  6043=>"100000100",
  6044=>"101010110",
  6045=>"101010111",
  6046=>"101000000",
  6047=>"001111101",
  6048=>"111001000",
  6049=>"101000001",
  6050=>"010010110",
  6051=>"100101000",
  6052=>"001100110",
  6053=>"100110110",
  6054=>"011010000",
  6055=>"011110101",
  6056=>"100100101",
  6057=>"111111100",
  6058=>"111010011",
  6059=>"000111110",
  6060=>"010010110",
  6061=>"000101011",
  6062=>"011011110",
  6063=>"000101011",
  6064=>"100100011",
  6065=>"111001111",
  6066=>"010111110",
  6067=>"101010111",
  6068=>"000000011",
  6069=>"000101101",
  6070=>"010101110",
  6071=>"000010101",
  6072=>"010101010",
  6073=>"110100101",
  6074=>"010110000",
  6075=>"001001100",
  6076=>"001101010",
  6077=>"010000101",
  6078=>"000011101",
  6079=>"011000001",
  6080=>"001000110",
  6081=>"011011001",
  6082=>"001111011",
  6083=>"101000000",
  6084=>"101100001",
  6085=>"001000101",
  6086=>"001001001",
  6087=>"000011000",
  6088=>"101011010",
  6089=>"000011011",
  6090=>"101100010",
  6091=>"011000001",
  6092=>"010011100",
  6093=>"100000010",
  6094=>"101001111",
  6095=>"110011101",
  6096=>"010111101",
  6097=>"111011011",
  6098=>"100100011",
  6099=>"000010101",
  6100=>"111001100",
  6101=>"111111110",
  6102=>"110110110",
  6103=>"000111110",
  6104=>"011101000",
  6105=>"000100111",
  6106=>"011001101",
  6107=>"011100100",
  6108=>"011000110",
  6109=>"100101111",
  6110=>"001011110",
  6111=>"011000011",
  6112=>"010111110",
  6113=>"001000010",
  6114=>"000101110",
  6115=>"000111011",
  6116=>"100110101",
  6117=>"000100110",
  6118=>"110010010",
  6119=>"011111101",
  6120=>"110101101",
  6121=>"101101100",
  6122=>"001011000",
  6123=>"100110111",
  6124=>"100101111",
  6125=>"010000010",
  6126=>"010010100",
  6127=>"100011101",
  6128=>"001101111",
  6129=>"011000101",
  6130=>"110111101",
  6131=>"111010110",
  6132=>"011011111",
  6133=>"101111010",
  6134=>"111001000",
  6135=>"000011011",
  6136=>"100001001",
  6137=>"000101000",
  6138=>"100011101",
  6139=>"001100001",
  6140=>"111001010",
  6141=>"000100011",
  6142=>"000101001",
  6143=>"000110110",
  6144=>"111111000",
  6145=>"010010001",
  6146=>"010101001",
  6147=>"111111100",
  6148=>"101100101",
  6149=>"010111110",
  6150=>"010100011",
  6151=>"001101000",
  6152=>"101010000",
  6153=>"001011101",
  6154=>"001100101",
  6155=>"110100111",
  6156=>"011000010",
  6157=>"111111010",
  6158=>"000011010",
  6159=>"001011011",
  6160=>"101110011",
  6161=>"111111001",
  6162=>"101100001",
  6163=>"111101011",
  6164=>"100011010",
  6165=>"011110110",
  6166=>"101101011",
  6167=>"001111101",
  6168=>"111011000",
  6169=>"001100011",
  6170=>"011001111",
  6171=>"100101100",
  6172=>"111110000",
  6173=>"111011101",
  6174=>"101010111",
  6175=>"001110111",
  6176=>"110001011",
  6177=>"001001101",
  6178=>"001000001",
  6179=>"011010011",
  6180=>"010011100",
  6181=>"111111000",
  6182=>"011000100",
  6183=>"111111111",
  6184=>"101100101",
  6185=>"001111011",
  6186=>"011110000",
  6187=>"000110111",
  6188=>"000111111",
  6189=>"111000011",
  6190=>"100100000",
  6191=>"101110111",
  6192=>"000111100",
  6193=>"100100111",
  6194=>"000101100",
  6195=>"111100000",
  6196=>"110001011",
  6197=>"011011100",
  6198=>"001101111",
  6199=>"111011111",
  6200=>"010100001",
  6201=>"010110110",
  6202=>"100111111",
  6203=>"110000010",
  6204=>"111000011",
  6205=>"111101110",
  6206=>"111001101",
  6207=>"101110100",
  6208=>"110101111",
  6209=>"010100110",
  6210=>"000100100",
  6211=>"001000010",
  6212=>"100110010",
  6213=>"100100001",
  6214=>"110010010",
  6215=>"010001001",
  6216=>"100001000",
  6217=>"100100111",
  6218=>"011000111",
  6219=>"000011111",
  6220=>"111000010",
  6221=>"011010001",
  6222=>"111111111",
  6223=>"010000000",
  6224=>"001001010",
  6225=>"000000111",
  6226=>"001111000",
  6227=>"000010011",
  6228=>"001000001",
  6229=>"111111101",
  6230=>"101100011",
  6231=>"011001111",
  6232=>"100000101",
  6233=>"110000001",
  6234=>"011000111",
  6235=>"011111101",
  6236=>"110001011",
  6237=>"000101001",
  6238=>"101111001",
  6239=>"101101101",
  6240=>"111101010",
  6241=>"011000111",
  6242=>"010011110",
  6243=>"011011001",
  6244=>"010010010",
  6245=>"000010110",
  6246=>"110111101",
  6247=>"001111100",
  6248=>"111001011",
  6249=>"100111111",
  6250=>"001000100",
  6251=>"011110111",
  6252=>"100001001",
  6253=>"010101110",
  6254=>"000000011",
  6255=>"011001000",
  6256=>"010110111",
  6257=>"001011100",
  6258=>"101110001",
  6259=>"000100010",
  6260=>"001010111",
  6261=>"111110100",
  6262=>"001101010",
  6263=>"001110101",
  6264=>"100010001",
  6265=>"100000000",
  6266=>"101011110",
  6267=>"000100010",
  6268=>"101000111",
  6269=>"111000101",
  6270=>"011011110",
  6271=>"001100101",
  6272=>"100001100",
  6273=>"100111101",
  6274=>"110101111",
  6275=>"101000011",
  6276=>"000000100",
  6277=>"000000010",
  6278=>"000010001",
  6279=>"110011101",
  6280=>"000011010",
  6281=>"110011011",
  6282=>"001100011",
  6283=>"100110111",
  6284=>"100110011",
  6285=>"001100101",
  6286=>"111101100",
  6287=>"000110010",
  6288=>"001010000",
  6289=>"000111100",
  6290=>"100110100",
  6291=>"010000001",
  6292=>"000110001",
  6293=>"100100110",
  6294=>"011010101",
  6295=>"100011101",
  6296=>"110101111",
  6297=>"010100111",
  6298=>"101110101",
  6299=>"010001001",
  6300=>"111011101",
  6301=>"010000101",
  6302=>"100010111",
  6303=>"011011110",
  6304=>"111000110",
  6305=>"001101010",
  6306=>"001011110",
  6307=>"010100110",
  6308=>"100011101",
  6309=>"000000000",
  6310=>"101011111",
  6311=>"100000000",
  6312=>"010000011",
  6313=>"110111111",
  6314=>"110000111",
  6315=>"011001101",
  6316=>"001001110",
  6317=>"000000111",
  6318=>"000001010",
  6319=>"111001111",
  6320=>"001111000",
  6321=>"010011100",
  6322=>"000110000",
  6323=>"101111101",
  6324=>"010111011",
  6325=>"001010000",
  6326=>"111111110",
  6327=>"001000010",
  6328=>"000100100",
  6329=>"011001010",
  6330=>"000110010",
  6331=>"100100110",
  6332=>"001110111",
  6333=>"000001110",
  6334=>"100010011",
  6335=>"110001110",
  6336=>"011011101",
  6337=>"101101100",
  6338=>"010110110",
  6339=>"010010000",
  6340=>"101011111",
  6341=>"000010001",
  6342=>"101100101",
  6343=>"010110011",
  6344=>"111111111",
  6345=>"111101001",
  6346=>"101101100",
  6347=>"011000111",
  6348=>"001010111",
  6349=>"110000011",
  6350=>"111001000",
  6351=>"101100110",
  6352=>"100010010",
  6353=>"010101100",
  6354=>"011001010",
  6355=>"011010101",
  6356=>"101011010",
  6357=>"100110011",
  6358=>"000101011",
  6359=>"011110111",
  6360=>"011001100",
  6361=>"110100111",
  6362=>"110001111",
  6363=>"110110111",
  6364=>"001011000",
  6365=>"111001101",
  6366=>"101101101",
  6367=>"111011001",
  6368=>"011001001",
  6369=>"110111111",
  6370=>"010111001",
  6371=>"101001011",
  6372=>"011111110",
  6373=>"000101010",
  6374=>"100111110",
  6375=>"101001010",
  6376=>"101000000",
  6377=>"110001100",
  6378=>"100110100",
  6379=>"000101101",
  6380=>"010111101",
  6381=>"001111011",
  6382=>"111111101",
  6383=>"101100111",
  6384=>"110000100",
  6385=>"100011000",
  6386=>"000101000",
  6387=>"000001010",
  6388=>"000011100",
  6389=>"000110000",
  6390=>"100110011",
  6391=>"110001110",
  6392=>"101011000",
  6393=>"001100101",
  6394=>"101000001",
  6395=>"101001111",
  6396=>"111010101",
  6397=>"011010110",
  6398=>"011111111",
  6399=>"001111111",
  6400=>"111110011",
  6401=>"000110100",
  6402=>"111011100",
  6403=>"011110100",
  6404=>"100111010",
  6405=>"100001101",
  6406=>"101110001",
  6407=>"101000010",
  6408=>"001010000",
  6409=>"111001111",
  6410=>"100101101",
  6411=>"111111011",
  6412=>"111101000",
  6413=>"011010010",
  6414=>"001110000",
  6415=>"011111110",
  6416=>"101100110",
  6417=>"101001101",
  6418=>"010011110",
  6419=>"010101000",
  6420=>"001111000",
  6421=>"010111110",
  6422=>"110001010",
  6423=>"100110100",
  6424=>"011000100",
  6425=>"110110010",
  6426=>"000010101",
  6427=>"010100110",
  6428=>"000110110",
  6429=>"111111001",
  6430=>"010110000",
  6431=>"001011100",
  6432=>"110110111",
  6433=>"110011111",
  6434=>"101010101",
  6435=>"010010011",
  6436=>"000000011",
  6437=>"001110000",
  6438=>"111100100",
  6439=>"110110000",
  6440=>"010010100",
  6441=>"000010111",
  6442=>"100001010",
  6443=>"101010010",
  6444=>"101101111",
  6445=>"100010000",
  6446=>"000101111",
  6447=>"010111000",
  6448=>"011110001",
  6449=>"000101001",
  6450=>"110100001",
  6451=>"110110010",
  6452=>"110000101",
  6453=>"010010110",
  6454=>"110111111",
  6455=>"011010100",
  6456=>"001011101",
  6457=>"010110001",
  6458=>"000100000",
  6459=>"001100011",
  6460=>"010001010",
  6461=>"001000001",
  6462=>"110010010",
  6463=>"111001111",
  6464=>"010001000",
  6465=>"010111111",
  6466=>"001001010",
  6467=>"011110001",
  6468=>"011001100",
  6469=>"100100111",
  6470=>"000000100",
  6471=>"011001001",
  6472=>"000000000",
  6473=>"110101011",
  6474=>"000101101",
  6475=>"010011010",
  6476=>"100000110",
  6477=>"011110011",
  6478=>"101110101",
  6479=>"111111011",
  6480=>"010111101",
  6481=>"111100001",
  6482=>"101011110",
  6483=>"011000110",
  6484=>"111010000",
  6485=>"010001010",
  6486=>"110111101",
  6487=>"011001100",
  6488=>"000100011",
  6489=>"110001111",
  6490=>"000010011",
  6491=>"010111000",
  6492=>"100101010",
  6493=>"001100001",
  6494=>"011101000",
  6495=>"111011001",
  6496=>"001101101",
  6497=>"110110100",
  6498=>"101000011",
  6499=>"000000110",
  6500=>"010011100",
  6501=>"110010100",
  6502=>"101110110",
  6503=>"000000111",
  6504=>"000000001",
  6505=>"010110000",
  6506=>"001110001",
  6507=>"010100010",
  6508=>"011010011",
  6509=>"100100111",
  6510=>"011101001",
  6511=>"000110010",
  6512=>"111011110",
  6513=>"111101101",
  6514=>"001010001",
  6515=>"110100010",
  6516=>"001010010",
  6517=>"101111111",
  6518=>"101110000",
  6519=>"101101011",
  6520=>"010110000",
  6521=>"101011011",
  6522=>"010010101",
  6523=>"000010101",
  6524=>"001101011",
  6525=>"100000110",
  6526=>"000111000",
  6527=>"001100111",
  6528=>"101011101",
  6529=>"011011001",
  6530=>"010110101",
  6531=>"111001101",
  6532=>"001000110",
  6533=>"101000101",
  6534=>"100110001",
  6535=>"000100011",
  6536=>"110010101",
  6537=>"110110011",
  6538=>"110000001",
  6539=>"101000100",
  6540=>"101010111",
  6541=>"110110011",
  6542=>"001001010",
  6543=>"011000000",
  6544=>"111111100",
  6545=>"000011000",
  6546=>"001000001",
  6547=>"111101110",
  6548=>"010001111",
  6549=>"110101011",
  6550=>"000010000",
  6551=>"010010100",
  6552=>"100010000",
  6553=>"101001000",
  6554=>"110011101",
  6555=>"000111100",
  6556=>"001000011",
  6557=>"010101110",
  6558=>"100000110",
  6559=>"010110001",
  6560=>"101100101",
  6561=>"000100110",
  6562=>"000001101",
  6563=>"001100001",
  6564=>"110001011",
  6565=>"100011101",
  6566=>"110001001",
  6567=>"001011011",
  6568=>"100010000",
  6569=>"110100101",
  6570=>"001010010",
  6571=>"000010110",
  6572=>"100111001",
  6573=>"100110110",
  6574=>"000000001",
  6575=>"101111110",
  6576=>"101111111",
  6577=>"011011010",
  6578=>"001111101",
  6579=>"000110010",
  6580=>"000101000",
  6581=>"000010111",
  6582=>"100000010",
  6583=>"100000100",
  6584=>"001100101",
  6585=>"011110100",
  6586=>"011011000",
  6587=>"010101110",
  6588=>"110110000",
  6589=>"111110000",
  6590=>"111100011",
  6591=>"110101011",
  6592=>"110011111",
  6593=>"111111111",
  6594=>"011110110",
  6595=>"100110111",
  6596=>"010000111",
  6597=>"000001010",
  6598=>"011001001",
  6599=>"111101101",
  6600=>"110101111",
  6601=>"111001010",
  6602=>"000101111",
  6603=>"000100000",
  6604=>"111111011",
  6605=>"110111011",
  6606=>"000111000",
  6607=>"010101000",
  6608=>"110101110",
  6609=>"011010011",
  6610=>"010001010",
  6611=>"110011010",
  6612=>"101000100",
  6613=>"111000111",
  6614=>"101111110",
  6615=>"111111101",
  6616=>"001001111",
  6617=>"000011100",
  6618=>"111011010",
  6619=>"101111011",
  6620=>"100111101",
  6621=>"001001010",
  6622=>"111010011",
  6623=>"000110000",
  6624=>"000110010",
  6625=>"000010001",
  6626=>"101001001",
  6627=>"001110001",
  6628=>"001101001",
  6629=>"011001100",
  6630=>"101001011",
  6631=>"111000111",
  6632=>"110000100",
  6633=>"101101000",
  6634=>"001111011",
  6635=>"111011100",
  6636=>"011100000",
  6637=>"010011000",
  6638=>"110100111",
  6639=>"110111111",
  6640=>"001100001",
  6641=>"100001100",
  6642=>"011111111",
  6643=>"010100010",
  6644=>"001011000",
  6645=>"000000111",
  6646=>"110010000",
  6647=>"010000000",
  6648=>"001011110",
  6649=>"010000000",
  6650=>"001011101",
  6651=>"010110001",
  6652=>"001000010",
  6653=>"001110001",
  6654=>"100110000",
  6655=>"000011100",
  6656=>"010110011",
  6657=>"010001100",
  6658=>"111110010",
  6659=>"011010001",
  6660=>"110110001",
  6661=>"110001001",
  6662=>"100110111",
  6663=>"100101011",
  6664=>"111111100",
  6665=>"000111010",
  6666=>"000001101",
  6667=>"010000110",
  6668=>"110111110",
  6669=>"110101000",
  6670=>"101100001",
  6671=>"101010100",
  6672=>"000110110",
  6673=>"011011010",
  6674=>"111101011",
  6675=>"111110100",
  6676=>"001011001",
  6677=>"010000101",
  6678=>"111001000",
  6679=>"101100110",
  6680=>"010000110",
  6681=>"111010011",
  6682=>"001101101",
  6683=>"111010101",
  6684=>"010001110",
  6685=>"010110001",
  6686=>"011011111",
  6687=>"011110001",
  6688=>"001001000",
  6689=>"110111101",
  6690=>"011100110",
  6691=>"101101111",
  6692=>"101001010",
  6693=>"001100000",
  6694=>"100000111",
  6695=>"100001101",
  6696=>"001101001",
  6697=>"110000110",
  6698=>"100000101",
  6699=>"101101000",
  6700=>"011100100",
  6701=>"010011101",
  6702=>"101001001",
  6703=>"100110101",
  6704=>"100000110",
  6705=>"100011110",
  6706=>"001011111",
  6707=>"000100001",
  6708=>"010010111",
  6709=>"111111110",
  6710=>"110011011",
  6711=>"110001100",
  6712=>"100110001",
  6713=>"011110000",
  6714=>"111100111",
  6715=>"100011110",
  6716=>"010000000",
  6717=>"101100011",
  6718=>"011100111",
  6719=>"000110010",
  6720=>"111100011",
  6721=>"100000000",
  6722=>"010000010",
  6723=>"000111110",
  6724=>"100100011",
  6725=>"000111111",
  6726=>"001000001",
  6727=>"001110110",
  6728=>"010100011",
  6729=>"111111110",
  6730=>"111101111",
  6731=>"100110010",
  6732=>"110011011",
  6733=>"111000101",
  6734=>"101011010",
  6735=>"000110101",
  6736=>"100001100",
  6737=>"011101101",
  6738=>"101011101",
  6739=>"100111010",
  6740=>"011110000",
  6741=>"010111000",
  6742=>"101001111",
  6743=>"000011000",
  6744=>"000010101",
  6745=>"000100010",
  6746=>"000110101",
  6747=>"100111100",
  6748=>"000001111",
  6749=>"001000011",
  6750=>"111101110",
  6751=>"000010110",
  6752=>"110111001",
  6753=>"010000100",
  6754=>"101011101",
  6755=>"101110011",
  6756=>"010011100",
  6757=>"111001110",
  6758=>"100110010",
  6759=>"001000000",
  6760=>"010110011",
  6761=>"101101001",
  6762=>"101000010",
  6763=>"001001010",
  6764=>"011100101",
  6765=>"011010100",
  6766=>"000110001",
  6767=>"110110111",
  6768=>"000110111",
  6769=>"110111010",
  6770=>"100001101",
  6771=>"110110111",
  6772=>"011100011",
  6773=>"000111111",
  6774=>"101001111",
  6775=>"010010110",
  6776=>"110100011",
  6777=>"100101101",
  6778=>"011110011",
  6779=>"111000110",
  6780=>"011000000",
  6781=>"010001110",
  6782=>"011000100",
  6783=>"110001000",
  6784=>"001111011",
  6785=>"110110010",
  6786=>"001001001",
  6787=>"100010101",
  6788=>"100101110",
  6789=>"111000010",
  6790=>"101010101",
  6791=>"110001101",
  6792=>"011101111",
  6793=>"100001111",
  6794=>"100100101",
  6795=>"110101100",
  6796=>"110000111",
  6797=>"111101011",
  6798=>"110100100",
  6799=>"000000101",
  6800=>"000111001",
  6801=>"011110001",
  6802=>"001110001",
  6803=>"100000001",
  6804=>"101111001",
  6805=>"101010001",
  6806=>"111001000",
  6807=>"000001010",
  6808=>"101011000",
  6809=>"011010011",
  6810=>"100101011",
  6811=>"111101011",
  6812=>"100011010",
  6813=>"111010101",
  6814=>"000001110",
  6815=>"101011000",
  6816=>"010100011",
  6817=>"110010101",
  6818=>"001001011",
  6819=>"110101001",
  6820=>"011100001",
  6821=>"001001011",
  6822=>"100010110",
  6823=>"101001101",
  6824=>"001111100",
  6825=>"110111101",
  6826=>"100001011",
  6827=>"111011001",
  6828=>"100000001",
  6829=>"000100000",
  6830=>"111011011",
  6831=>"010010010",
  6832=>"101010110",
  6833=>"001111101",
  6834=>"111110111",
  6835=>"101010000",
  6836=>"001001011",
  6837=>"111111001",
  6838=>"010010000",
  6839=>"101101110",
  6840=>"110001011",
  6841=>"110001111",
  6842=>"010010101",
  6843=>"101110001",
  6844=>"111000101",
  6845=>"111111101",
  6846=>"000000010",
  6847=>"001110111",
  6848=>"001011100",
  6849=>"000101111",
  6850=>"011011001",
  6851=>"110101101",
  6852=>"010010010",
  6853=>"100101010",
  6854=>"001001001",
  6855=>"000101001",
  6856=>"110011000",
  6857=>"010111011",
  6858=>"001011011",
  6859=>"010101010",
  6860=>"000100011",
  6861=>"101111110",
  6862=>"010111110",
  6863=>"010010001",
  6864=>"001001110",
  6865=>"101100100",
  6866=>"111010010",
  6867=>"101011111",
  6868=>"011000100",
  6869=>"000010101",
  6870=>"011001000",
  6871=>"000011110",
  6872=>"110000100",
  6873=>"110111110",
  6874=>"001010001",
  6875=>"001001011",
  6876=>"101011110",
  6877=>"000100111",
  6878=>"100011011",
  6879=>"100000100",
  6880=>"100111110",
  6881=>"010000110",
  6882=>"011000111",
  6883=>"000111011",
  6884=>"100111010",
  6885=>"001000000",
  6886=>"100111100",
  6887=>"000110001",
  6888=>"000101011",
  6889=>"100010101",
  6890=>"110000001",
  6891=>"111101111",
  6892=>"011101001",
  6893=>"100110110",
  6894=>"011100010",
  6895=>"101110010",
  6896=>"110111111",
  6897=>"111011111",
  6898=>"110111101",
  6899=>"100100010",
  6900=>"011100011",
  6901=>"100110110",
  6902=>"000001100",
  6903=>"011010000",
  6904=>"010011111",
  6905=>"101000111",
  6906=>"010001010",
  6907=>"111101011",
  6908=>"000000101",
  6909=>"010010000",
  6910=>"100001110",
  6911=>"101001001",
  6912=>"100111111",
  6913=>"001000000",
  6914=>"001110001",
  6915=>"110100100",
  6916=>"110000110",
  6917=>"101001011",
  6918=>"011111111",
  6919=>"111101001",
  6920=>"100000001",
  6921=>"101111101",
  6922=>"100101010",
  6923=>"001101001",
  6924=>"001001101",
  6925=>"011110110",
  6926=>"110111011",
  6927=>"110000111",
  6928=>"101001001",
  6929=>"010001101",
  6930=>"000010000",
  6931=>"101000000",
  6932=>"001111101",
  6933=>"111001110",
  6934=>"110011001",
  6935=>"010110011",
  6936=>"111111101",
  6937=>"011111110",
  6938=>"100111101",
  6939=>"111100110",
  6940=>"100010101",
  6941=>"101111000",
  6942=>"011110000",
  6943=>"111001000",
  6944=>"001011111",
  6945=>"110011110",
  6946=>"111010110",
  6947=>"101011100",
  6948=>"110111000",
  6949=>"000110101",
  6950=>"001110010",
  6951=>"000101111",
  6952=>"111011011",
  6953=>"011010011",
  6954=>"011110101",
  6955=>"010001111",
  6956=>"110000001",
  6957=>"010010100",
  6958=>"011000001",
  6959=>"010101111",
  6960=>"010001000",
  6961=>"011001101",
  6962=>"111101100",
  6963=>"101101101",
  6964=>"111001011",
  6965=>"010000100",
  6966=>"110100100",
  6967=>"110010011",
  6968=>"101111011",
  6969=>"111011000",
  6970=>"100110011",
  6971=>"000010000",
  6972=>"111101000",
  6973=>"110001100",
  6974=>"110010111",
  6975=>"110001011",
  6976=>"110111100",
  6977=>"001010111",
  6978=>"101000110",
  6979=>"001001101",
  6980=>"001110100",
  6981=>"101010001",
  6982=>"110001110",
  6983=>"101000000",
  6984=>"110000110",
  6985=>"101101100",
  6986=>"101110100",
  6987=>"111000011",
  6988=>"001111001",
  6989=>"111100110",
  6990=>"111100100",
  6991=>"110000100",
  6992=>"000001001",
  6993=>"011000100",
  6994=>"011111011",
  6995=>"111000000",
  6996=>"110100011",
  6997=>"101101110",
  6998=>"001001011",
  6999=>"010110010",
  7000=>"001010100",
  7001=>"011011010",
  7002=>"101110000",
  7003=>"011000001",
  7004=>"001101111",
  7005=>"000010011",
  7006=>"110111100",
  7007=>"000111010",
  7008=>"111001101",
  7009=>"001110011",
  7010=>"000000111",
  7011=>"010010010",
  7012=>"010111011",
  7013=>"011010000",
  7014=>"010011100",
  7015=>"110000101",
  7016=>"000011001",
  7017=>"101101111",
  7018=>"111001000",
  7019=>"100011001",
  7020=>"101000001",
  7021=>"101011101",
  7022=>"111011011",
  7023=>"000010101",
  7024=>"000001001",
  7025=>"100100001",
  7026=>"011011001",
  7027=>"111100000",
  7028=>"011011111",
  7029=>"111111011",
  7030=>"110100101",
  7031=>"001011001",
  7032=>"100101101",
  7033=>"011110011",
  7034=>"001101111",
  7035=>"110000000",
  7036=>"011100001",
  7037=>"111011111",
  7038=>"100011011",
  7039=>"111011100",
  7040=>"110101001",
  7041=>"100110101",
  7042=>"000010011",
  7043=>"110110001",
  7044=>"100110101",
  7045=>"100110000",
  7046=>"100111100",
  7047=>"101001010",
  7048=>"111111110",
  7049=>"111011110",
  7050=>"010111011",
  7051=>"101010001",
  7052=>"010110000",
  7053=>"011011000",
  7054=>"101100001",
  7055=>"111011001",
  7056=>"001000100",
  7057=>"010011001",
  7058=>"011010001",
  7059=>"110000011",
  7060=>"111011010",
  7061=>"111001011",
  7062=>"011000010",
  7063=>"010001011",
  7064=>"110010100",
  7065=>"101011001",
  7066=>"000110110",
  7067=>"110110110",
  7068=>"110011011",
  7069=>"111000110",
  7070=>"010110001",
  7071=>"010000100",
  7072=>"101101111",
  7073=>"111110011",
  7074=>"011110011",
  7075=>"100001101",
  7076=>"010011111",
  7077=>"100111011",
  7078=>"110100100",
  7079=>"001000111",
  7080=>"101110101",
  7081=>"110000110",
  7082=>"001001110",
  7083=>"000011100",
  7084=>"111100111",
  7085=>"100010110",
  7086=>"011000101",
  7087=>"000101001",
  7088=>"000100101",
  7089=>"011000011",
  7090=>"000011111",
  7091=>"010011111",
  7092=>"111001110",
  7093=>"011000110",
  7094=>"101100100",
  7095=>"110001010",
  7096=>"011101101",
  7097=>"111001110",
  7098=>"010110110",
  7099=>"001011001",
  7100=>"111111101",
  7101=>"001101110",
  7102=>"000111000",
  7103=>"000001001",
  7104=>"001110101",
  7105=>"000110100",
  7106=>"000001001",
  7107=>"110001110",
  7108=>"100111100",
  7109=>"001000101",
  7110=>"110110110",
  7111=>"100111111",
  7112=>"000110110",
  7113=>"011001001",
  7114=>"101101001",
  7115=>"010101010",
  7116=>"010111110",
  7117=>"101010011",
  7118=>"000100000",
  7119=>"100101101",
  7120=>"000101111",
  7121=>"000101001",
  7122=>"001011010",
  7123=>"000100111",
  7124=>"011111000",
  7125=>"110000100",
  7126=>"110101101",
  7127=>"000011101",
  7128=>"000001101",
  7129=>"000000110",
  7130=>"110101101",
  7131=>"111100110",
  7132=>"101101111",
  7133=>"111010010",
  7134=>"001110000",
  7135=>"001001110",
  7136=>"100101101",
  7137=>"011111000",
  7138=>"011111001",
  7139=>"101111011",
  7140=>"110011101",
  7141=>"000111010",
  7142=>"000010011",
  7143=>"010011001",
  7144=>"001000010",
  7145=>"011000101",
  7146=>"001010011",
  7147=>"000010111",
  7148=>"000100110",
  7149=>"111000001",
  7150=>"111111100",
  7151=>"101101000",
  7152=>"001100000",
  7153=>"101110100",
  7154=>"000110111",
  7155=>"111100001",
  7156=>"111010000",
  7157=>"011111110",
  7158=>"001111111",
  7159=>"001111100",
  7160=>"011010100",
  7161=>"001100101",
  7162=>"010110111",
  7163=>"111110001",
  7164=>"011000010",
  7165=>"000000100",
  7166=>"001100000",
  7167=>"010010100",
  7168=>"100011111",
  7169=>"100001010",
  7170=>"100010110",
  7171=>"100001110",
  7172=>"000100000",
  7173=>"010011010",
  7174=>"101000110",
  7175=>"100000001",
  7176=>"000111100",
  7177=>"001000100",
  7178=>"101010010",
  7179=>"111101101",
  7180=>"001110110",
  7181=>"111001011",
  7182=>"010010101",
  7183=>"110001001",
  7184=>"001010001",
  7185=>"000100011",
  7186=>"101011000",
  7187=>"001101011",
  7188=>"110011101",
  7189=>"010000010",
  7190=>"100001101",
  7191=>"000000111",
  7192=>"110110101",
  7193=>"000100000",
  7194=>"101010111",
  7195=>"111100110",
  7196=>"010100111",
  7197=>"000110000",
  7198=>"111001110",
  7199=>"011010001",
  7200=>"101001000",
  7201=>"110100100",
  7202=>"110001001",
  7203=>"100100011",
  7204=>"001111110",
  7205=>"100010000",
  7206=>"001000011",
  7207=>"100101111",
  7208=>"010001010",
  7209=>"001011110",
  7210=>"111001100",
  7211=>"001010011",
  7212=>"010101000",
  7213=>"101110100",
  7214=>"010101001",
  7215=>"111011111",
  7216=>"011001111",
  7217=>"100111110",
  7218=>"101111011",
  7219=>"110011000",
  7220=>"011101101",
  7221=>"100000010",
  7222=>"111001110",
  7223=>"010010011",
  7224=>"111110100",
  7225=>"001011000",
  7226=>"111000110",
  7227=>"010011000",
  7228=>"001111100",
  7229=>"001001101",
  7230=>"010001111",
  7231=>"001110000",
  7232=>"100100001",
  7233=>"100111110",
  7234=>"000100110",
  7235=>"001001101",
  7236=>"010001010",
  7237=>"000011000",
  7238=>"110010100",
  7239=>"011010100",
  7240=>"101100010",
  7241=>"001000001",
  7242=>"110101111",
  7243=>"111000111",
  7244=>"000000110",
  7245=>"010010001",
  7246=>"001010011",
  7247=>"010111001",
  7248=>"000100111",
  7249=>"110100000",
  7250=>"100010000",
  7251=>"100111011",
  7252=>"001001111",
  7253=>"000111100",
  7254=>"111110010",
  7255=>"101110101",
  7256=>"000011001",
  7257=>"111101000",
  7258=>"001110000",
  7259=>"000111011",
  7260=>"111111000",
  7261=>"110011001",
  7262=>"011000101",
  7263=>"000000111",
  7264=>"000011100",
  7265=>"000101111",
  7266=>"111010110",
  7267=>"110110100",
  7268=>"110001010",
  7269=>"101110100",
  7270=>"010011101",
  7271=>"101011011",
  7272=>"111011001",
  7273=>"101100111",
  7274=>"100000001",
  7275=>"011110010",
  7276=>"011101110",
  7277=>"110100111",
  7278=>"001001100",
  7279=>"011010101",
  7280=>"100010011",
  7281=>"111111011",
  7282=>"111010010",
  7283=>"011001111",
  7284=>"110011000",
  7285=>"010111010",
  7286=>"000001000",
  7287=>"110010101",
  7288=>"001000111",
  7289=>"011000010",
  7290=>"010010100",
  7291=>"110110000",
  7292=>"110111100",
  7293=>"001111100",
  7294=>"011000010",
  7295=>"100100101",
  7296=>"000101000",
  7297=>"010111000",
  7298=>"011010000",
  7299=>"110100110",
  7300=>"001100110",
  7301=>"010111001",
  7302=>"111001111",
  7303=>"100011101",
  7304=>"110111001",
  7305=>"011100001",
  7306=>"001111111",
  7307=>"001000110",
  7308=>"101000011",
  7309=>"100000100",
  7310=>"001010100",
  7311=>"010000010",
  7312=>"110100000",
  7313=>"100111101",
  7314=>"001101111",
  7315=>"010000000",
  7316=>"101001101",
  7317=>"101111111",
  7318=>"111110001",
  7319=>"011001011",
  7320=>"110011000",
  7321=>"101101010",
  7322=>"000001111",
  7323=>"010010011",
  7324=>"101110101",
  7325=>"111111111",
  7326=>"110001100",
  7327=>"010110110",
  7328=>"001010100",
  7329=>"100001100",
  7330=>"101000101",
  7331=>"000010010",
  7332=>"110101111",
  7333=>"100101000",
  7334=>"000100111",
  7335=>"011011101",
  7336=>"001010110",
  7337=>"011001111",
  7338=>"011111100",
  7339=>"010000010",
  7340=>"000101011",
  7341=>"001101101",
  7342=>"001011000",
  7343=>"100001011",
  7344=>"000001110",
  7345=>"111011010",
  7346=>"110110001",
  7347=>"000110010",
  7348=>"110101000",
  7349=>"000000101",
  7350=>"010111011",
  7351=>"110010000",
  7352=>"010111100",
  7353=>"100101100",
  7354=>"101001100",
  7355=>"101111111",
  7356=>"011000000",
  7357=>"001100000",
  7358=>"010011101",
  7359=>"000001110",
  7360=>"001111001",
  7361=>"010000101",
  7362=>"000000101",
  7363=>"001000011",
  7364=>"000100110",
  7365=>"011001000",
  7366=>"110101010",
  7367=>"010010110",
  7368=>"010111011",
  7369=>"100100010",
  7370=>"001001111",
  7371=>"011111100",
  7372=>"111101100",
  7373=>"111010001",
  7374=>"100100101",
  7375=>"010110000",
  7376=>"001000100",
  7377=>"101000101",
  7378=>"011100010",
  7379=>"001100001",
  7380=>"100001010",
  7381=>"011101100",
  7382=>"010010110",
  7383=>"101101001",
  7384=>"000111111",
  7385=>"001001011",
  7386=>"000100000",
  7387=>"001100001",
  7388=>"000110111",
  7389=>"000111000",
  7390=>"110011111",
  7391=>"111101101",
  7392=>"110000100",
  7393=>"100111010",
  7394=>"010000110",
  7395=>"100000100",
  7396=>"001010100",
  7397=>"101000001",
  7398=>"100111111",
  7399=>"100110011",
  7400=>"110101111",
  7401=>"100100000",
  7402=>"011100010",
  7403=>"101010111",
  7404=>"011110000",
  7405=>"110011110",
  7406=>"000000010",
  7407=>"000110000",
  7408=>"011100000",
  7409=>"000000011",
  7410=>"101101001",
  7411=>"110101100",
  7412=>"011111100",
  7413=>"011010101",
  7414=>"110000000",
  7415=>"011010101",
  7416=>"001000011",
  7417=>"000001100",
  7418=>"111010101",
  7419=>"010110001",
  7420=>"101111111",
  7421=>"100000100",
  7422=>"000001001",
  7423=>"111100011",
  7424=>"111110110",
  7425=>"111111010",
  7426=>"000111100",
  7427=>"110001111",
  7428=>"111010110",
  7429=>"010010000",
  7430=>"001010011",
  7431=>"010010010",
  7432=>"011010000",
  7433=>"111011110",
  7434=>"010010111",
  7435=>"011000110",
  7436=>"011000011",
  7437=>"101000110",
  7438=>"111111101",
  7439=>"011101110",
  7440=>"011000111",
  7441=>"000100100",
  7442=>"010000100",
  7443=>"010001010",
  7444=>"011110010",
  7445=>"101011111",
  7446=>"100111100",
  7447=>"001010010",
  7448=>"001010101",
  7449=>"011001010",
  7450=>"000001010",
  7451=>"011001011",
  7452=>"001010111",
  7453=>"101101000",
  7454=>"000010011",
  7455=>"100001000",
  7456=>"010001100",
  7457=>"010110101",
  7458=>"101111100",
  7459=>"000010011",
  7460=>"110000000",
  7461=>"010010100",
  7462=>"100101011",
  7463=>"101100010",
  7464=>"011010110",
  7465=>"101100010",
  7466=>"101000010",
  7467=>"101010110",
  7468=>"001100000",
  7469=>"101001101",
  7470=>"111101001",
  7471=>"010111100",
  7472=>"010100010",
  7473=>"010011101",
  7474=>"101010110",
  7475=>"101101010",
  7476=>"101011010",
  7477=>"111001010",
  7478=>"111000100",
  7479=>"010001010",
  7480=>"111110001",
  7481=>"110001000",
  7482=>"000101010",
  7483=>"011101000",
  7484=>"111010101",
  7485=>"100110111",
  7486=>"111111100",
  7487=>"011111101",
  7488=>"011100100",
  7489=>"000011110",
  7490=>"000010011",
  7491=>"101001000",
  7492=>"000100110",
  7493=>"101101001",
  7494=>"110111111",
  7495=>"010000100",
  7496=>"001011110",
  7497=>"101010001",
  7498=>"101111100",
  7499=>"010000100",
  7500=>"111011111",
  7501=>"011011101",
  7502=>"011011100",
  7503=>"101001100",
  7504=>"101111010",
  7505=>"100010100",
  7506=>"010110111",
  7507=>"011001011",
  7508=>"110011101",
  7509=>"001011100",
  7510=>"000101010",
  7511=>"001101011",
  7512=>"101010001",
  7513=>"101001001",
  7514=>"101010111",
  7515=>"000001010",
  7516=>"111011110",
  7517=>"110111111",
  7518=>"010001111",
  7519=>"010100111",
  7520=>"100110000",
  7521=>"000111010",
  7522=>"100011110",
  7523=>"001100000",
  7524=>"000001100",
  7525=>"001001011",
  7526=>"010011011",
  7527=>"001010100",
  7528=>"011000001",
  7529=>"011100001",
  7530=>"100110111",
  7531=>"000110100",
  7532=>"111001101",
  7533=>"000001001",
  7534=>"000101111",
  7535=>"001000001",
  7536=>"100101110",
  7537=>"000111001",
  7538=>"101001010",
  7539=>"111101110",
  7540=>"001110011",
  7541=>"111111000",
  7542=>"001000111",
  7543=>"111000001",
  7544=>"001101101",
  7545=>"101110010",
  7546=>"010001101",
  7547=>"010110111",
  7548=>"001010101",
  7549=>"111011010",
  7550=>"011011011",
  7551=>"000010011",
  7552=>"000010010",
  7553=>"000001011",
  7554=>"010000001",
  7555=>"101111000",
  7556=>"110111010",
  7557=>"101100011",
  7558=>"010001011",
  7559=>"111010111",
  7560=>"011010000",
  7561=>"000010100",
  7562=>"000000101",
  7563=>"010011110",
  7564=>"110000011",
  7565=>"001010010",
  7566=>"011000001",
  7567=>"001101000",
  7568=>"010001010",
  7569=>"000000000",
  7570=>"110110100",
  7571=>"011101101",
  7572=>"001101110",
  7573=>"000100101",
  7574=>"110000011",
  7575=>"101111010",
  7576=>"100001000",
  7577=>"010010001",
  7578=>"000111001",
  7579=>"011110110",
  7580=>"101111001",
  7581=>"101001101",
  7582=>"000010011",
  7583=>"111111111",
  7584=>"011100001",
  7585=>"000011101",
  7586=>"000111011",
  7587=>"000111100",
  7588=>"111111101",
  7589=>"001000111",
  7590=>"011001010",
  7591=>"010101000",
  7592=>"001110100",
  7593=>"110001100",
  7594=>"110101110",
  7595=>"001010111",
  7596=>"101101111",
  7597=>"111001011",
  7598=>"111000000",
  7599=>"011000001",
  7600=>"101100000",
  7601=>"000100100",
  7602=>"100011011",
  7603=>"001010100",
  7604=>"011111011",
  7605=>"000001100",
  7606=>"000010000",
  7607=>"110000101",
  7608=>"111101110",
  7609=>"000101111",
  7610=>"011011010",
  7611=>"000011101",
  7612=>"100100001",
  7613=>"000000101",
  7614=>"110101001",
  7615=>"110110010",
  7616=>"100100101",
  7617=>"000011110",
  7618=>"110110110",
  7619=>"011010000",
  7620=>"100000010",
  7621=>"110101011",
  7622=>"101011010",
  7623=>"001101110",
  7624=>"001011011",
  7625=>"000001100",
  7626=>"000100000",
  7627=>"110010000",
  7628=>"111000110",
  7629=>"000110100",
  7630=>"100000010",
  7631=>"110010100",
  7632=>"011010101",
  7633=>"000111100",
  7634=>"110110001",
  7635=>"101010010",
  7636=>"011101111",
  7637=>"100101000",
  7638=>"011100101",
  7639=>"011001011",
  7640=>"000011010",
  7641=>"010100101",
  7642=>"110111011",
  7643=>"000101000",
  7644=>"010010111",
  7645=>"101010011",
  7646=>"101110010",
  7647=>"111011101",
  7648=>"010100011",
  7649=>"110111100",
  7650=>"101111101",
  7651=>"001010001",
  7652=>"110001010",
  7653=>"100111100",
  7654=>"100011001",
  7655=>"001001001",
  7656=>"001011010",
  7657=>"100010001",
  7658=>"101110100",
  7659=>"001011101",
  7660=>"001110010",
  7661=>"000011000",
  7662=>"000100101",
  7663=>"001000010",
  7664=>"011000101",
  7665=>"000001101",
  7666=>"100110101",
  7667=>"001011000",
  7668=>"010000111",
  7669=>"100100001",
  7670=>"111010001",
  7671=>"011001001",
  7672=>"100101110",
  7673=>"010000101",
  7674=>"000101101",
  7675=>"100010110",
  7676=>"110110111",
  7677=>"111100000",
  7678=>"111111111",
  7679=>"110001111",
  7680=>"000000100",
  7681=>"101010101",
  7682=>"011010001",
  7683=>"010001100",
  7684=>"010111011",
  7685=>"001011001",
  7686=>"011000000",
  7687=>"011010100",
  7688=>"001110100",
  7689=>"000011110",
  7690=>"000110011",
  7691=>"110011111",
  7692=>"101011011",
  7693=>"011011010",
  7694=>"000001101",
  7695=>"101001001",
  7696=>"000110010",
  7697=>"001100001",
  7698=>"000001101",
  7699=>"111010100",
  7700=>"110000000",
  7701=>"000110010",
  7702=>"111001111",
  7703=>"000000000",
  7704=>"100011000",
  7705=>"110001001",
  7706=>"001001001",
  7707=>"100111000",
  7708=>"100000010",
  7709=>"101111000",
  7710=>"101111011",
  7711=>"111011111",
  7712=>"010111000",
  7713=>"101001011",
  7714=>"011110111",
  7715=>"000101010",
  7716=>"111011111",
  7717=>"101101010",
  7718=>"010101101",
  7719=>"101111111",
  7720=>"011011001",
  7721=>"111011001",
  7722=>"100110111",
  7723=>"101011010",
  7724=>"101111001",
  7725=>"100100101",
  7726=>"001001110",
  7727=>"110110100",
  7728=>"000001000",
  7729=>"100100000",
  7730=>"100010111",
  7731=>"011111110",
  7732=>"001111001",
  7733=>"010110110",
  7734=>"001000011",
  7735=>"110111010",
  7736=>"010101010",
  7737=>"000110001",
  7738=>"111100100",
  7739=>"111110110",
  7740=>"011001011",
  7741=>"101010000",
  7742=>"111110001",
  7743=>"000100110",
  7744=>"111001000",
  7745=>"111001110",
  7746=>"000011100",
  7747=>"111101110",
  7748=>"011110111",
  7749=>"100010110",
  7750=>"001011111",
  7751=>"101011100",
  7752=>"011110011",
  7753=>"100001111",
  7754=>"010000101",
  7755=>"110110011",
  7756=>"011010111",
  7757=>"000100110",
  7758=>"011000001",
  7759=>"101010010",
  7760=>"001100100",
  7761=>"010000010",
  7762=>"000001011",
  7763=>"100101111",
  7764=>"011001000",
  7765=>"001111000",
  7766=>"000110010",
  7767=>"100011011",
  7768=>"100011010",
  7769=>"000000100",
  7770=>"101010001",
  7771=>"101101101",
  7772=>"100001010",
  7773=>"100011000",
  7774=>"000000011",
  7775=>"010110110",
  7776=>"000100000",
  7777=>"100011101",
  7778=>"001101100",
  7779=>"110011010",
  7780=>"110001110",
  7781=>"010011011",
  7782=>"100001111",
  7783=>"110111101",
  7784=>"011100001",
  7785=>"000100100",
  7786=>"111011011",
  7787=>"111101010",
  7788=>"001000000",
  7789=>"100010011",
  7790=>"101001011",
  7791=>"000010110",
  7792=>"101111011",
  7793=>"000011000",
  7794=>"111001101",
  7795=>"010111110",
  7796=>"100010010",
  7797=>"001110010",
  7798=>"110010110",
  7799=>"001111100",
  7800=>"010111000",
  7801=>"000011100",
  7802=>"010000010",
  7803=>"111000101",
  7804=>"011001011",
  7805=>"000110110",
  7806=>"110001111",
  7807=>"000110010",
  7808=>"001000001",
  7809=>"001110101",
  7810=>"111010111",
  7811=>"101000011",
  7812=>"001010101",
  7813=>"000010100",
  7814=>"001011001",
  7815=>"010110110",
  7816=>"101110111",
  7817=>"110100100",
  7818=>"100011010",
  7819=>"101000101",
  7820=>"101100001",
  7821=>"011000101",
  7822=>"110111110",
  7823=>"110110011",
  7824=>"000110111",
  7825=>"100111010",
  7826=>"100111001",
  7827=>"001101010",
  7828=>"111000000",
  7829=>"001000011",
  7830=>"010101111",
  7831=>"001111101",
  7832=>"100000011",
  7833=>"000000000",
  7834=>"011101010",
  7835=>"101111010",
  7836=>"101001000",
  7837=>"110010100",
  7838=>"100001110",
  7839=>"100110111",
  7840=>"101100010",
  7841=>"001101101",
  7842=>"101101000",
  7843=>"010111011",
  7844=>"110001101",
  7845=>"101111011",
  7846=>"111111100",
  7847=>"111000101",
  7848=>"101111010",
  7849=>"111100110",
  7850=>"011000101",
  7851=>"010000000",
  7852=>"111101101",
  7853=>"011100001",
  7854=>"100001110",
  7855=>"110001101",
  7856=>"011100010",
  7857=>"101111100",
  7858=>"011010111",
  7859=>"111011111",
  7860=>"001101111",
  7861=>"101101110",
  7862=>"110101001",
  7863=>"101110010",
  7864=>"011100101",
  7865=>"010111110",
  7866=>"111111011",
  7867=>"010000111",
  7868=>"101111001",
  7869=>"000000110",
  7870=>"101001100",
  7871=>"000111111",
  7872=>"001000010",
  7873=>"001011000",
  7874=>"100001101",
  7875=>"111011100",
  7876=>"101111101",
  7877=>"110101010",
  7878=>"100110011",
  7879=>"110110000",
  7880=>"001000001",
  7881=>"100001001",
  7882=>"011001000",
  7883=>"101001101",
  7884=>"001101000",
  7885=>"011000111",
  7886=>"010010011",
  7887=>"000000001",
  7888=>"010001100",
  7889=>"011001010",
  7890=>"101100110",
  7891=>"001101001",
  7892=>"001011110",
  7893=>"000010111",
  7894=>"101001001",
  7895=>"000101010",
  7896=>"110110100",
  7897=>"001101011",
  7898=>"010000111",
  7899=>"001110100",
  7900=>"110100010",
  7901=>"110111011",
  7902=>"101010011",
  7903=>"000000100",
  7904=>"010011000",
  7905=>"001010001",
  7906=>"101001111",
  7907=>"111111000",
  7908=>"100101011",
  7909=>"111101100",
  7910=>"001010111",
  7911=>"111101011",
  7912=>"000011000",
  7913=>"111101101",
  7914=>"000010011",
  7915=>"100001010",
  7916=>"011000101",
  7917=>"101000101",
  7918=>"111011011",
  7919=>"101010100",
  7920=>"001110110",
  7921=>"011111100",
  7922=>"000010100",
  7923=>"000110111",
  7924=>"101000001",
  7925=>"111001000",
  7926=>"101110111",
  7927=>"101000001",
  7928=>"011011111",
  7929=>"110001010",
  7930=>"001110100",
  7931=>"001100101",
  7932=>"000000101",
  7933=>"110111110",
  7934=>"101101100",
  7935=>"111100010",
  7936=>"111000010",
  7937=>"101000100",
  7938=>"111110111",
  7939=>"000001011",
  7940=>"101000001",
  7941=>"001111110",
  7942=>"110010111",
  7943=>"111011001",
  7944=>"100000101",
  7945=>"111000010",
  7946=>"111001100",
  7947=>"111101101",
  7948=>"100111000",
  7949=>"000111001",
  7950=>"000111001",
  7951=>"100110110",
  7952=>"101111111",
  7953=>"111011000",
  7954=>"101111011",
  7955=>"100101011",
  7956=>"000111010",
  7957=>"000001011",
  7958=>"010101001",
  7959=>"011110010",
  7960=>"000000110",
  7961=>"101001000",
  7962=>"000010100",
  7963=>"111111100",
  7964=>"111001010",
  7965=>"100011110",
  7966=>"101100101",
  7967=>"011011000",
  7968=>"000101100",
  7969=>"110101000",
  7970=>"100110000",
  7971=>"000110100",
  7972=>"000000100",
  7973=>"111100111",
  7974=>"101111100",
  7975=>"110001111",
  7976=>"110100001",
  7977=>"000111100",
  7978=>"000000000",
  7979=>"100101111",
  7980=>"010100100",
  7981=>"011101110",
  7982=>"111001000",
  7983=>"110000110",
  7984=>"010000111",
  7985=>"100100001",
  7986=>"101101111",
  7987=>"011000111",
  7988=>"000101001",
  7989=>"011000100",
  7990=>"110111000",
  7991=>"000111110",
  7992=>"110111100",
  7993=>"110000100",
  7994=>"000001101",
  7995=>"100101001",
  7996=>"001001110",
  7997=>"110101110",
  7998=>"010110111",
  7999=>"110000000",
  8000=>"101111000",
  8001=>"100110011",
  8002=>"111001001",
  8003=>"100100111",
  8004=>"000011001",
  8005=>"010001101",
  8006=>"010101001",
  8007=>"011010111",
  8008=>"000111111",
  8009=>"100011100",
  8010=>"110111101",
  8011=>"001011000",
  8012=>"011000011",
  8013=>"000110111",
  8014=>"101011110",
  8015=>"101010010",
  8016=>"100001110",
  8017=>"111111101",
  8018=>"000001001",
  8019=>"111001010",
  8020=>"100001101",
  8021=>"111111000",
  8022=>"010100000",
  8023=>"111101101",
  8024=>"001101111",
  8025=>"110111000",
  8026=>"001110100",
  8027=>"000001001",
  8028=>"101110111",
  8029=>"000100001",
  8030=>"010100001",
  8031=>"000111110",
  8032=>"100110011",
  8033=>"100110110",
  8034=>"001101111",
  8035=>"010111111",
  8036=>"110011101",
  8037=>"000001000",
  8038=>"111101110",
  8039=>"001101000",
  8040=>"100000101",
  8041=>"101111000",
  8042=>"111000010",
  8043=>"111100011",
  8044=>"100111001",
  8045=>"011011101",
  8046=>"000100101",
  8047=>"100001110",
  8048=>"001000100",
  8049=>"100111001",
  8050=>"001110000",
  8051=>"101100000",
  8052=>"101101011",
  8053=>"110000100",
  8054=>"001011000",
  8055=>"011100000",
  8056=>"000110101",
  8057=>"001001111",
  8058=>"010001010",
  8059=>"011111101",
  8060=>"001101001",
  8061=>"001100110",
  8062=>"011100010",
  8063=>"011111111",
  8064=>"010010100",
  8065=>"101011110",
  8066=>"011100010",
  8067=>"101110000",
  8068=>"110111110",
  8069=>"111101011",
  8070=>"101000101",
  8071=>"000000111",
  8072=>"011111001",
  8073=>"111011010",
  8074=>"010010000",
  8075=>"110010011",
  8076=>"110111000",
  8077=>"101110110",
  8078=>"000010100",
  8079=>"001100010",
  8080=>"111111011",
  8081=>"100101011",
  8082=>"101100001",
  8083=>"111111011",
  8084=>"000110001",
  8085=>"010100110",
  8086=>"111100101",
  8087=>"101111100",
  8088=>"011111111",
  8089=>"000101010",
  8090=>"110011100",
  8091=>"101001111",
  8092=>"111001010",
  8093=>"000111011",
  8094=>"111001011",
  8095=>"011101011",
  8096=>"001111101",
  8097=>"101100001",
  8098=>"111110100",
  8099=>"011001100",
  8100=>"111111101",
  8101=>"010000101",
  8102=>"110000101",
  8103=>"001101111",
  8104=>"011000001",
  8105=>"001010110",
  8106=>"011110100",
  8107=>"001111101",
  8108=>"011110011",
  8109=>"111010000",
  8110=>"000001000",
  8111=>"111111011",
  8112=>"010011010",
  8113=>"111001110",
  8114=>"010110000",
  8115=>"011001100",
  8116=>"110010111",
  8117=>"100110001",
  8118=>"110111001",
  8119=>"000110011",
  8120=>"111000001",
  8121=>"010001101",
  8122=>"001011111",
  8123=>"010100001",
  8124=>"110000111",
  8125=>"010000001",
  8126=>"000100000",
  8127=>"011101111",
  8128=>"100010111",
  8129=>"010101011",
  8130=>"010110111",
  8131=>"010011101",
  8132=>"011001010",
  8133=>"001011111",
  8134=>"100010111",
  8135=>"001111111",
  8136=>"111100110",
  8137=>"101000111",
  8138=>"111101001",
  8139=>"001011110",
  8140=>"011001101",
  8141=>"111000111",
  8142=>"101100000",
  8143=>"101100101",
  8144=>"001011100",
  8145=>"100010001",
  8146=>"000001001",
  8147=>"100000010",
  8148=>"111001000",
  8149=>"100000010",
  8150=>"111101010",
  8151=>"010111010",
  8152=>"110001000",
  8153=>"000011110",
  8154=>"100011010",
  8155=>"011001100",
  8156=>"001001011",
  8157=>"000001001",
  8158=>"011100111",
  8159=>"000110011",
  8160=>"001100010",
  8161=>"101111001",
  8162=>"110100110",
  8163=>"000110100",
  8164=>"100001100",
  8165=>"001100110",
  8166=>"001101100",
  8167=>"111001010",
  8168=>"111011111",
  8169=>"011101010",
  8170=>"100010101",
  8171=>"100001111",
  8172=>"110100000",
  8173=>"001001001",
  8174=>"001100001",
  8175=>"111011111",
  8176=>"100010111",
  8177=>"110100000",
  8178=>"101111111",
  8179=>"001110111",
  8180=>"010001001",
  8181=>"001000100",
  8182=>"110110010",
  8183=>"100111010",
  8184=>"110001000",
  8185=>"101110000",
  8186=>"011100111",
  8187=>"110000000",
  8188=>"011100011",
  8189=>"111001101",
  8190=>"011111110",
  8191=>"011000010",
  8192=>"110011010",
  8193=>"110110011",
  8194=>"110010100",
  8195=>"110100001",
  8196=>"000000110",
  8197=>"111010101",
  8198=>"011110100",
  8199=>"111100110",
  8200=>"011001000",
  8201=>"111110001",
  8202=>"101100011",
  8203=>"000010001",
  8204=>"111001111",
  8205=>"000101001",
  8206=>"110011000",
  8207=>"001110000",
  8208=>"000000010",
  8209=>"101010000",
  8210=>"110000100",
  8211=>"000001111",
  8212=>"000101000",
  8213=>"101101011",
  8214=>"000101010",
  8215=>"101101011",
  8216=>"100000001",
  8217=>"000010001",
  8218=>"000101000",
  8219=>"100001111",
  8220=>"011000011",
  8221=>"110001101",
  8222=>"001010000",
  8223=>"001100101",
  8224=>"110100111",
  8225=>"001011001",
  8226=>"111011111",
  8227=>"001101011",
  8228=>"110001000",
  8229=>"011101110",
  8230=>"001100100",
  8231=>"000111111",
  8232=>"101011111",
  8233=>"000110110",
  8234=>"111110101",
  8235=>"111010010",
  8236=>"111100110",
  8237=>"001110111",
  8238=>"110001010",
  8239=>"010101001",
  8240=>"111101011",
  8241=>"100111111",
  8242=>"011100101",
  8243=>"110101010",
  8244=>"101011100",
  8245=>"110111101",
  8246=>"001010010",
  8247=>"011011101",
  8248=>"101111100",
  8249=>"100000100",
  8250=>"101001101",
  8251=>"101011010",
  8252=>"111111001",
  8253=>"110011111",
  8254=>"111001011",
  8255=>"100010110",
  8256=>"100010010",
  8257=>"011011010",
  8258=>"010110100",
  8259=>"101010101",
  8260=>"111101100",
  8261=>"100100000",
  8262=>"011111111",
  8263=>"111100001",
  8264=>"110110011",
  8265=>"111100010",
  8266=>"001100011",
  8267=>"111001110",
  8268=>"011001010",
  8269=>"100101101",
  8270=>"111010100",
  8271=>"110100111",
  8272=>"111101111",
  8273=>"000001000",
  8274=>"101011111",
  8275=>"010101000",
  8276=>"110111111",
  8277=>"100000100",
  8278=>"100001011",
  8279=>"001001011",
  8280=>"011111111",
  8281=>"110010000",
  8282=>"110110101",
  8283=>"110111000",
  8284=>"100100100",
  8285=>"000101011",
  8286=>"100010000",
  8287=>"110110000",
  8288=>"111110001",
  8289=>"010001000",
  8290=>"000011101",
  8291=>"010011001",
  8292=>"010111010",
  8293=>"001111101",
  8294=>"101111111",
  8295=>"010001101",
  8296=>"101100111",
  8297=>"110000011",
  8298=>"000100101",
  8299=>"101110111",
  8300=>"101101100",
  8301=>"101100010",
  8302=>"110010010",
  8303=>"001101011",
  8304=>"010111000",
  8305=>"001011100",
  8306=>"001010110",
  8307=>"101110001",
  8308=>"000001011",
  8309=>"100011101",
  8310=>"111111111",
  8311=>"011110111",
  8312=>"001010010",
  8313=>"010010111",
  8314=>"110111001",
  8315=>"000010000",
  8316=>"010011001",
  8317=>"000010001",
  8318=>"010001111",
  8319=>"011010000",
  8320=>"010100000",
  8321=>"100100110",
  8322=>"011110010",
  8323=>"000100100",
  8324=>"011010101",
  8325=>"011000001",
  8326=>"011000111",
  8327=>"111000110",
  8328=>"100010011",
  8329=>"000010011",
  8330=>"011001001",
  8331=>"100101110",
  8332=>"010101011",
  8333=>"110101010",
  8334=>"011000010",
  8335=>"010110000",
  8336=>"010011100",
  8337=>"001111001",
  8338=>"111001001",
  8339=>"100011101",
  8340=>"111101010",
  8341=>"101111100",
  8342=>"010010010",
  8343=>"000101011",
  8344=>"111011011",
  8345=>"000011000",
  8346=>"100101001",
  8347=>"001001111",
  8348=>"111000100",
  8349=>"010101000",
  8350=>"100101001",
  8351=>"100010000",
  8352=>"001100001",
  8353=>"101000101",
  8354=>"110010110",
  8355=>"111000101",
  8356=>"100100001",
  8357=>"001000011",
  8358=>"101010101",
  8359=>"010110100",
  8360=>"001111100",
  8361=>"100110010",
  8362=>"110111111",
  8363=>"001010000",
  8364=>"010110110",
  8365=>"000100100",
  8366=>"111110000",
  8367=>"110110111",
  8368=>"001010100",
  8369=>"100100010",
  8370=>"101110111",
  8371=>"100101000",
  8372=>"011111011",
  8373=>"000001111",
  8374=>"100010100",
  8375=>"110101110",
  8376=>"010100000",
  8377=>"000100010",
  8378=>"111100100",
  8379=>"010100110",
  8380=>"001101000",
  8381=>"101110000",
  8382=>"111001001",
  8383=>"101111011",
  8384=>"011101101",
  8385=>"110000010",
  8386=>"111110011",
  8387=>"010110100",
  8388=>"011000011",
  8389=>"000110011",
  8390=>"010001000",
  8391=>"000110101",
  8392=>"100000110",
  8393=>"101111010",
  8394=>"111001101",
  8395=>"111001010",
  8396=>"100110110",
  8397=>"000100100",
  8398=>"101010001",
  8399=>"011000001",
  8400=>"101001010",
  8401=>"011101010",
  8402=>"110000000",
  8403=>"011011111",
  8404=>"101100001",
  8405=>"110001111",
  8406=>"110010011",
  8407=>"010111010",
  8408=>"000101100",
  8409=>"001001111",
  8410=>"000100000",
  8411=>"000010111",
  8412=>"100011101",
  8413=>"111011110",
  8414=>"001100111",
  8415=>"010111110",
  8416=>"110000000",
  8417=>"001000010",
  8418=>"110110011",
  8419=>"010101010",
  8420=>"010101110",
  8421=>"000101011",
  8422=>"000010000",
  8423=>"011101011",
  8424=>"100001000",
  8425=>"011101001",
  8426=>"010000011",
  8427=>"100100001",
  8428=>"011010000",
  8429=>"011001000",
  8430=>"010000000",
  8431=>"001100000",
  8432=>"011000101",
  8433=>"010101101",
  8434=>"000001011",
  8435=>"100110111",
  8436=>"001100110",
  8437=>"111010000",
  8438=>"000100001",
  8439=>"010000010",
  8440=>"111011111",
  8441=>"100101110",
  8442=>"000110000",
  8443=>"110011100",
  8444=>"101011111",
  8445=>"111110011",
  8446=>"111111111",
  8447=>"110111100",
  8448=>"100110111",
  8449=>"101110001",
  8450=>"000010111",
  8451=>"010110100",
  8452=>"011010111",
  8453=>"011100000",
  8454=>"111011100",
  8455=>"101100100",
  8456=>"100001011",
  8457=>"000011000",
  8458=>"011000101",
  8459=>"010100100",
  8460=>"111101111",
  8461=>"011000001",
  8462=>"000011000",
  8463=>"111101001",
  8464=>"010110000",
  8465=>"111100101",
  8466=>"001111111",
  8467=>"000000111",
  8468=>"000111111",
  8469=>"100001000",
  8470=>"011000000",
  8471=>"000100000",
  8472=>"111101011",
  8473=>"111111101",
  8474=>"100000001",
  8475=>"111100101",
  8476=>"100011111",
  8477=>"100001000",
  8478=>"111110111",
  8479=>"110110110",
  8480=>"111100111",
  8481=>"001110000",
  8482=>"110010100",
  8483=>"100010011",
  8484=>"100010000",
  8485=>"010110000",
  8486=>"111111111",
  8487=>"110011111",
  8488=>"111101000",
  8489=>"100010001",
  8490=>"101101000",
  8491=>"100011010",
  8492=>"111100010",
  8493=>"111111111",
  8494=>"010100100",
  8495=>"100010001",
  8496=>"011000111",
  8497=>"100011000",
  8498=>"100111100",
  8499=>"001010011",
  8500=>"111100111",
  8501=>"010100000",
  8502=>"100000111",
  8503=>"001101110",
  8504=>"101111110",
  8505=>"110100011",
  8506=>"000011110",
  8507=>"001000010",
  8508=>"101010111",
  8509=>"001000111",
  8510=>"111110100",
  8511=>"111001111",
  8512=>"001011110",
  8513=>"111100001",
  8514=>"001101001",
  8515=>"000101011",
  8516=>"001000011",
  8517=>"000010000",
  8518=>"000001000",
  8519=>"011100110",
  8520=>"100110011",
  8521=>"000100000",
  8522=>"110100100",
  8523=>"111100100",
  8524=>"001010011",
  8525=>"010111010",
  8526=>"000111110",
  8527=>"001010011",
  8528=>"010100001",
  8529=>"101111000",
  8530=>"100001010",
  8531=>"110111100",
  8532=>"010101000",
  8533=>"101000010",
  8534=>"010101111",
  8535=>"000001000",
  8536=>"111011001",
  8537=>"011110001",
  8538=>"000110100",
  8539=>"111001100",
  8540=>"100111100",
  8541=>"000111111",
  8542=>"010111011",
  8543=>"011100111",
  8544=>"010101011",
  8545=>"110101110",
  8546=>"010101000",
  8547=>"110001101",
  8548=>"101010011",
  8549=>"000100111",
  8550=>"101011000",
  8551=>"000110110",
  8552=>"001001111",
  8553=>"011111000",
  8554=>"111010110",
  8555=>"111110001",
  8556=>"010110011",
  8557=>"011111000",
  8558=>"010001000",
  8559=>"100000100",
  8560=>"110111011",
  8561=>"100110001",
  8562=>"110000110",
  8563=>"001100001",
  8564=>"000111010",
  8565=>"010001010",
  8566=>"110001000",
  8567=>"111111111",
  8568=>"110011011",
  8569=>"000110011",
  8570=>"001100111",
  8571=>"110001101",
  8572=>"000101000",
  8573=>"110011100",
  8574=>"101011101",
  8575=>"010011110",
  8576=>"000000111",
  8577=>"010110000",
  8578=>"000111101",
  8579=>"010100010",
  8580=>"001010111",
  8581=>"001001111",
  8582=>"011001100",
  8583=>"000010000",
  8584=>"101000000",
  8585=>"000001000",
  8586=>"000001111",
  8587=>"111010010",
  8588=>"001111100",
  8589=>"001110000",
  8590=>"110000011",
  8591=>"001110000",
  8592=>"111010100",
  8593=>"000000111",
  8594=>"010001110",
  8595=>"011110001",
  8596=>"000101000",
  8597=>"000100001",
  8598=>"000010000",
  8599=>"111001101",
  8600=>"000001100",
  8601=>"011000000",
  8602=>"000010010",
  8603=>"100011010",
  8604=>"010001000",
  8605=>"001001110",
  8606=>"111010110",
  8607=>"001000010",
  8608=>"011101101",
  8609=>"001000111",
  8610=>"100100110",
  8611=>"101100001",
  8612=>"110100011",
  8613=>"001000101",
  8614=>"110111001",
  8615=>"111001110",
  8616=>"001011011",
  8617=>"011001111",
  8618=>"011110001",
  8619=>"111101111",
  8620=>"110000010",
  8621=>"100010011",
  8622=>"010001101",
  8623=>"110010001",
  8624=>"110011110",
  8625=>"111000001",
  8626=>"000011001",
  8627=>"011111010",
  8628=>"101101101",
  8629=>"000011011",
  8630=>"001010010",
  8631=>"111101101",
  8632=>"000010111",
  8633=>"010100110",
  8634=>"011011000",
  8635=>"100111101",
  8636=>"000000101",
  8637=>"011000011",
  8638=>"111101001",
  8639=>"100110001",
  8640=>"010000000",
  8641=>"001001101",
  8642=>"000000110",
  8643=>"101011101",
  8644=>"001010101",
  8645=>"001110100",
  8646=>"000110011",
  8647=>"101000000",
  8648=>"111011010",
  8649=>"011100111",
  8650=>"001001100",
  8651=>"011110000",
  8652=>"100001011",
  8653=>"011001001",
  8654=>"100000111",
  8655=>"000111101",
  8656=>"011000100",
  8657=>"011001010",
  8658=>"011000110",
  8659=>"000100110",
  8660=>"001110011",
  8661=>"110100100",
  8662=>"111111011",
  8663=>"110111100",
  8664=>"101001101",
  8665=>"110011101",
  8666=>"111010001",
  8667=>"011100110",
  8668=>"010100011",
  8669=>"001101001",
  8670=>"010101100",
  8671=>"001010111",
  8672=>"010011111",
  8673=>"010001000",
  8674=>"100001000",
  8675=>"000000011",
  8676=>"111010011",
  8677=>"001001001",
  8678=>"000111110",
  8679=>"000111001",
  8680=>"100001011",
  8681=>"100101000",
  8682=>"101001001",
  8683=>"010100111",
  8684=>"011011001",
  8685=>"111011011",
  8686=>"011111011",
  8687=>"100000101",
  8688=>"100001010",
  8689=>"111111011",
  8690=>"110100011",
  8691=>"111011000",
  8692=>"011100010",
  8693=>"011110011",
  8694=>"110000011",
  8695=>"001000100",
  8696=>"000000101",
  8697=>"011001011",
  8698=>"001001000",
  8699=>"101101010",
  8700=>"000011110",
  8701=>"001011101",
  8702=>"000110110",
  8703=>"110100000",
  8704=>"010001011",
  8705=>"101111110",
  8706=>"101001101",
  8707=>"011011001",
  8708=>"100001001",
  8709=>"010001010",
  8710=>"100000110",
  8711=>"011110000",
  8712=>"011110001",
  8713=>"000001001",
  8714=>"111001010",
  8715=>"000000001",
  8716=>"001110010",
  8717=>"100100010",
  8718=>"110100010",
  8719=>"110101001",
  8720=>"010001101",
  8721=>"001010111",
  8722=>"101100100",
  8723=>"111000100",
  8724=>"011000110",
  8725=>"111000100",
  8726=>"001111111",
  8727=>"010110001",
  8728=>"000010011",
  8729=>"011111111",
  8730=>"011000110",
  8731=>"101011101",
  8732=>"010100100",
  8733=>"111010111",
  8734=>"001011101",
  8735=>"100001111",
  8736=>"001011001",
  8737=>"000001111",
  8738=>"101000100",
  8739=>"110011011",
  8740=>"001111101",
  8741=>"000011011",
  8742=>"011111111",
  8743=>"010111000",
  8744=>"100110010",
  8745=>"100101010",
  8746=>"011111011",
  8747=>"010110010",
  8748=>"010110101",
  8749=>"011100111",
  8750=>"000000000",
  8751=>"111011111",
  8752=>"101001111",
  8753=>"011001101",
  8754=>"001010001",
  8755=>"100000011",
  8756=>"111110110",
  8757=>"101000010",
  8758=>"000001101",
  8759=>"011100101",
  8760=>"001010001",
  8761=>"011111001",
  8762=>"101100001",
  8763=>"000000110",
  8764=>"111100010",
  8765=>"111011001",
  8766=>"110101101",
  8767=>"011011111",
  8768=>"011010100",
  8769=>"011010110",
  8770=>"001000111",
  8771=>"010111001",
  8772=>"101011111",
  8773=>"000010001",
  8774=>"001000000",
  8775=>"001101100",
  8776=>"010001011",
  8777=>"111111010",
  8778=>"100001001",
  8779=>"000000100",
  8780=>"111001110",
  8781=>"101010001",
  8782=>"011100010",
  8783=>"000111010",
  8784=>"111011001",
  8785=>"000110010",
  8786=>"111110000",
  8787=>"000000011",
  8788=>"011100011",
  8789=>"000110000",
  8790=>"000101100",
  8791=>"100100100",
  8792=>"011100111",
  8793=>"111000001",
  8794=>"000001100",
  8795=>"101001111",
  8796=>"000100111",
  8797=>"000000010",
  8798=>"011110111",
  8799=>"010011111",
  8800=>"100001010",
  8801=>"110001000",
  8802=>"100111011",
  8803=>"010110111",
  8804=>"000111110",
  8805=>"100101101",
  8806=>"100000010",
  8807=>"100001111",
  8808=>"111111110",
  8809=>"100100011",
  8810=>"001100011",
  8811=>"110001000",
  8812=>"000000100",
  8813=>"001100101",
  8814=>"101010011",
  8815=>"001110110",
  8816=>"000001100",
  8817=>"010010100",
  8818=>"100011001",
  8819=>"110110111",
  8820=>"111011000",
  8821=>"110111100",
  8822=>"100001001",
  8823=>"100001011",
  8824=>"111001010",
  8825=>"010111010",
  8826=>"100111110",
  8827=>"111010010",
  8828=>"010000001",
  8829=>"001001000",
  8830=>"000011101",
  8831=>"101001100",
  8832=>"111101000",
  8833=>"110011001",
  8834=>"010011010",
  8835=>"110000100",
  8836=>"000100000",
  8837=>"100001010",
  8838=>"000011100",
  8839=>"100011101",
  8840=>"111100111",
  8841=>"111011100",
  8842=>"110011110",
  8843=>"001110111",
  8844=>"011000010",
  8845=>"010000110",
  8846=>"101000101",
  8847=>"001000001",
  8848=>"111110001",
  8849=>"100110111",
  8850=>"110100011",
  8851=>"110111101",
  8852=>"101000101",
  8853=>"100110100",
  8854=>"011101010",
  8855=>"110110111",
  8856=>"100000110",
  8857=>"011110000",
  8858=>"011000101",
  8859=>"111101110",
  8860=>"011001111",
  8861=>"000011010",
  8862=>"111000001",
  8863=>"011001001",
  8864=>"001011111",
  8865=>"110101110",
  8866=>"101101011",
  8867=>"000101111",
  8868=>"111111010",
  8869=>"000100010",
  8870=>"001000001",
  8871=>"111001001",
  8872=>"011011000",
  8873=>"101010000",
  8874=>"001101011",
  8875=>"001100010",
  8876=>"010010010",
  8877=>"000100001",
  8878=>"111011001",
  8879=>"010010001",
  8880=>"001100111",
  8881=>"000001110",
  8882=>"101001111",
  8883=>"111110000",
  8884=>"100000110",
  8885=>"010101111",
  8886=>"010100001",
  8887=>"101000011",
  8888=>"111001010",
  8889=>"110101010",
  8890=>"000101100",
  8891=>"110101011",
  8892=>"001000001",
  8893=>"101010000",
  8894=>"011001100",
  8895=>"111110010",
  8896=>"011101001",
  8897=>"000111101",
  8898=>"001011000",
  8899=>"010111011",
  8900=>"110111100",
  8901=>"110010000",
  8902=>"100010000",
  8903=>"000101010",
  8904=>"111010100",
  8905=>"100010101",
  8906=>"110011001",
  8907=>"000000000",
  8908=>"010001111",
  8909=>"101110001",
  8910=>"110111111",
  8911=>"010101010",
  8912=>"001100100",
  8913=>"100100111",
  8914=>"001001000",
  8915=>"011011011",
  8916=>"111000100",
  8917=>"011100000",
  8918=>"011011000",
  8919=>"100011011",
  8920=>"101001101",
  8921=>"110101100",
  8922=>"110001111",
  8923=>"100010011",
  8924=>"111000000",
  8925=>"001001111",
  8926=>"111101111",
  8927=>"000100010",
  8928=>"010001000",
  8929=>"101000111",
  8930=>"100001111",
  8931=>"010000110",
  8932=>"001010000",
  8933=>"101010101",
  8934=>"000000001",
  8935=>"001111000",
  8936=>"000101111",
  8937=>"101001110",
  8938=>"110000101",
  8939=>"110010111",
  8940=>"110010011",
  8941=>"010000111",
  8942=>"111100100",
  8943=>"001111100",
  8944=>"000110111",
  8945=>"010101110",
  8946=>"110000100",
  8947=>"001100100",
  8948=>"000111101",
  8949=>"111110011",
  8950=>"110101111",
  8951=>"011110101",
  8952=>"100000111",
  8953=>"001001111",
  8954=>"011001011",
  8955=>"110001001",
  8956=>"000011001",
  8957=>"110100110",
  8958=>"010001001",
  8959=>"100110010",
  8960=>"100110010",
  8961=>"000111111",
  8962=>"000011110",
  8963=>"011000101",
  8964=>"100001000",
  8965=>"011000010",
  8966=>"000100111",
  8967=>"100101000",
  8968=>"000000101",
  8969=>"011100101",
  8970=>"000111110",
  8971=>"111001100",
  8972=>"111100011",
  8973=>"010100101",
  8974=>"101101011",
  8975=>"010000111",
  8976=>"010110100",
  8977=>"100101011",
  8978=>"000110010",
  8979=>"111110010",
  8980=>"111010110",
  8981=>"000100101",
  8982=>"101011111",
  8983=>"000011010",
  8984=>"111101101",
  8985=>"000011011",
  8986=>"000001010",
  8987=>"001100111",
  8988=>"110110001",
  8989=>"111100011",
  8990=>"011101011",
  8991=>"101010010",
  8992=>"011010110",
  8993=>"111111011",
  8994=>"111100010",
  8995=>"111101000",
  8996=>"001111000",
  8997=>"010001001",
  8998=>"000000110",
  8999=>"001111010",
  9000=>"101010011",
  9001=>"011101001",
  9002=>"001111101",
  9003=>"010111111",
  9004=>"000000001",
  9005=>"101001111",
  9006=>"101011000",
  9007=>"101001100",
  9008=>"001100100",
  9009=>"100011001",
  9010=>"010110111",
  9011=>"110000000",
  9012=>"011111111",
  9013=>"100001110",
  9014=>"010111010",
  9015=>"110110001",
  9016=>"001001101",
  9017=>"001001010",
  9018=>"100110010",
  9019=>"001111101",
  9020=>"011101001",
  9021=>"111000101",
  9022=>"101101000",
  9023=>"011110110",
  9024=>"111111010",
  9025=>"111111011",
  9026=>"100111001",
  9027=>"110111100",
  9028=>"110100011",
  9029=>"111111100",
  9030=>"101001100",
  9031=>"100010100",
  9032=>"110011000",
  9033=>"010111000",
  9034=>"101010101",
  9035=>"001101100",
  9036=>"110010110",
  9037=>"110110110",
  9038=>"111111011",
  9039=>"110001111",
  9040=>"011001000",
  9041=>"010110010",
  9042=>"010011000",
  9043=>"010000000",
  9044=>"011100100",
  9045=>"001110010",
  9046=>"100000011",
  9047=>"000111110",
  9048=>"100111110",
  9049=>"010110011",
  9050=>"000101000",
  9051=>"101100011",
  9052=>"101111111",
  9053=>"000001110",
  9054=>"111111111",
  9055=>"110010000",
  9056=>"010010100",
  9057=>"110101001",
  9058=>"110010101",
  9059=>"000011101",
  9060=>"010110001",
  9061=>"011101000",
  9062=>"011010001",
  9063=>"100111111",
  9064=>"111011010",
  9065=>"100001111",
  9066=>"100110101",
  9067=>"111010000",
  9068=>"100100111",
  9069=>"100001011",
  9070=>"110110001",
  9071=>"100001111",
  9072=>"111101111",
  9073=>"001111010",
  9074=>"001001001",
  9075=>"011011111",
  9076=>"011011110",
  9077=>"110110110",
  9078=>"111101001",
  9079=>"010011100",
  9080=>"011101110",
  9081=>"010000110",
  9082=>"001110100",
  9083=>"000100101",
  9084=>"001000000",
  9085=>"001000001",
  9086=>"101110011",
  9087=>"011001110",
  9088=>"001011011",
  9089=>"000111110",
  9090=>"111001010",
  9091=>"001001001",
  9092=>"100110110",
  9093=>"011111011",
  9094=>"101111011",
  9095=>"011011100",
  9096=>"011000111",
  9097=>"101110001",
  9098=>"001000001",
  9099=>"001101001",
  9100=>"101101010",
  9101=>"111000000",
  9102=>"001011101",
  9103=>"110101100",
  9104=>"111001101",
  9105=>"110001100",
  9106=>"101010000",
  9107=>"000001001",
  9108=>"111101111",
  9109=>"010000010",
  9110=>"011011111",
  9111=>"110010001",
  9112=>"111100110",
  9113=>"110001010",
  9114=>"011011010",
  9115=>"110010001",
  9116=>"100100000",
  9117=>"010110010",
  9118=>"100000010",
  9119=>"110000100",
  9120=>"111011011",
  9121=>"011111001",
  9122=>"000100110",
  9123=>"011001100",
  9124=>"111010110",
  9125=>"100001000",
  9126=>"000101101",
  9127=>"010111001",
  9128=>"111011010",
  9129=>"010000000",
  9130=>"001111100",
  9131=>"000000101",
  9132=>"111111001",
  9133=>"000110001",
  9134=>"111000000",
  9135=>"101110010",
  9136=>"111101110",
  9137=>"100000000",
  9138=>"011010011",
  9139=>"001100110",
  9140=>"010100100",
  9141=>"001101010",
  9142=>"011001101",
  9143=>"011110001",
  9144=>"101000101",
  9145=>"000011011",
  9146=>"010111111",
  9147=>"001010011",
  9148=>"111010011",
  9149=>"111110110",
  9150=>"110010010",
  9151=>"100011111",
  9152=>"010110110",
  9153=>"001100101",
  9154=>"100011000",
  9155=>"101000000",
  9156=>"010000010",
  9157=>"111010010",
  9158=>"100111101",
  9159=>"100001110",
  9160=>"110011000",
  9161=>"100110010",
  9162=>"100101101",
  9163=>"011101100",
  9164=>"101010110",
  9165=>"101001000",
  9166=>"100111110",
  9167=>"011101101",
  9168=>"101111101",
  9169=>"110111101",
  9170=>"100101100",
  9171=>"110000100",
  9172=>"111110001",
  9173=>"000010111",
  9174=>"011000011",
  9175=>"000010101",
  9176=>"111001001",
  9177=>"001011100",
  9178=>"110111101",
  9179=>"111011111",
  9180=>"110001001",
  9181=>"000010000",
  9182=>"011000001",
  9183=>"001100011",
  9184=>"111111101",
  9185=>"010010100",
  9186=>"011110111",
  9187=>"110111001",
  9188=>"011011010",
  9189=>"011000111",
  9190=>"000100111",
  9191=>"100001011",
  9192=>"111100001",
  9193=>"000000001",
  9194=>"111111101",
  9195=>"110001101",
  9196=>"011101000",
  9197=>"110100010",
  9198=>"110010111",
  9199=>"110010110",
  9200=>"000100110",
  9201=>"010001010",
  9202=>"110000010",
  9203=>"000000100",
  9204=>"010010010",
  9205=>"000011111",
  9206=>"001011000",
  9207=>"100101101",
  9208=>"111001011",
  9209=>"011011100",
  9210=>"000100101",
  9211=>"110111111",
  9212=>"001010111",
  9213=>"110000101",
  9214=>"011111110",
  9215=>"110100001",
  9216=>"101010111",
  9217=>"011011011",
  9218=>"110000001",
  9219=>"010001010",
  9220=>"100111111",
  9221=>"101010101",
  9222=>"001100000",
  9223=>"000110010",
  9224=>"001110001",
  9225=>"010100001",
  9226=>"101000000",
  9227=>"111111100",
  9228=>"111101101",
  9229=>"100101100",
  9230=>"111100010",
  9231=>"011000011",
  9232=>"011010101",
  9233=>"100001100",
  9234=>"000101000",
  9235=>"100111000",
  9236=>"001010010",
  9237=>"010001100",
  9238=>"011010110",
  9239=>"000110110",
  9240=>"101111000",
  9241=>"010101110",
  9242=>"110100000",
  9243=>"010101110",
  9244=>"010011010",
  9245=>"110000001",
  9246=>"001011001",
  9247=>"100011001",
  9248=>"000000101",
  9249=>"001010101",
  9250=>"011010010",
  9251=>"101111111",
  9252=>"111010000",
  9253=>"011100110",
  9254=>"001010101",
  9255=>"110110110",
  9256=>"010001010",
  9257=>"000101110",
  9258=>"101011110",
  9259=>"110111100",
  9260=>"101010011",
  9261=>"100011111",
  9262=>"110111111",
  9263=>"100100010",
  9264=>"111010010",
  9265=>"110000111",
  9266=>"111000110",
  9267=>"111011101",
  9268=>"000000000",
  9269=>"100011000",
  9270=>"011000000",
  9271=>"111011111",
  9272=>"110000000",
  9273=>"000001010",
  9274=>"001110101",
  9275=>"010100111",
  9276=>"010101100",
  9277=>"110001101",
  9278=>"011110111",
  9279=>"011101001",
  9280=>"000111111",
  9281=>"110011000",
  9282=>"111011001",
  9283=>"011100111",
  9284=>"111001010",
  9285=>"001000101",
  9286=>"010011011",
  9287=>"010111100",
  9288=>"011100100",
  9289=>"101111110",
  9290=>"011010110",
  9291=>"001111111",
  9292=>"100010111",
  9293=>"000010001",
  9294=>"110000110",
  9295=>"101101101",
  9296=>"111101011",
  9297=>"001111000",
  9298=>"101011100",
  9299=>"110010100",
  9300=>"110110011",
  9301=>"110110011",
  9302=>"010000111",
  9303=>"111010000",
  9304=>"001000000",
  9305=>"101100101",
  9306=>"000000111",
  9307=>"010100010",
  9308=>"001101110",
  9309=>"110111111",
  9310=>"010101010",
  9311=>"110011101",
  9312=>"001101001",
  9313=>"101000010",
  9314=>"010001000",
  9315=>"000111100",
  9316=>"000100111",
  9317=>"110110100",
  9318=>"000110010",
  9319=>"001111100",
  9320=>"010111101",
  9321=>"001110110",
  9322=>"011100011",
  9323=>"010010111",
  9324=>"010010010",
  9325=>"111011111",
  9326=>"011100101",
  9327=>"111100110",
  9328=>"100010100",
  9329=>"111101011",
  9330=>"000001100",
  9331=>"110010110",
  9332=>"110000010",
  9333=>"111100101",
  9334=>"111111110",
  9335=>"010011010",
  9336=>"010000000",
  9337=>"010100100",
  9338=>"001100100",
  9339=>"101101010",
  9340=>"010000100",
  9341=>"011000001",
  9342=>"111110111",
  9343=>"110110000",
  9344=>"000100010",
  9345=>"110100011",
  9346=>"001100000",
  9347=>"001010111",
  9348=>"110111000",
  9349=>"000010111",
  9350=>"011110001",
  9351=>"010100100",
  9352=>"101110000",
  9353=>"001100111",
  9354=>"101100001",
  9355=>"101010110",
  9356=>"010000101",
  9357=>"011001100",
  9358=>"100000100",
  9359=>"001001111",
  9360=>"111110011",
  9361=>"010000001",
  9362=>"100100101",
  9363=>"010110101",
  9364=>"010010000",
  9365=>"111101100",
  9366=>"011101100",
  9367=>"011000100",
  9368=>"011010001",
  9369=>"000000100",
  9370=>"111100110",
  9371=>"111011100",
  9372=>"001000010",
  9373=>"011101111",
  9374=>"000001010",
  9375=>"110111010",
  9376=>"100000110",
  9377=>"110010001",
  9378=>"000011010",
  9379=>"000001101",
  9380=>"001011001",
  9381=>"101110110",
  9382=>"001010110",
  9383=>"011010000",
  9384=>"110110100",
  9385=>"100011100",
  9386=>"010101101",
  9387=>"100000001",
  9388=>"110111010",
  9389=>"110101101",
  9390=>"110011110",
  9391=>"101011110",
  9392=>"010100011",
  9393=>"111101111",
  9394=>"010100000",
  9395=>"011101001",
  9396=>"001101110",
  9397=>"000111000",
  9398=>"100000011",
  9399=>"111101001",
  9400=>"001010110",
  9401=>"001111001",
  9402=>"101011010",
  9403=>"101101010",
  9404=>"101101011",
  9405=>"011000011",
  9406=>"000011011",
  9407=>"100011010",
  9408=>"000010011",
  9409=>"010000100",
  9410=>"001001111",
  9411=>"110100101",
  9412=>"101001111",
  9413=>"101000111",
  9414=>"000101011",
  9415=>"010010101",
  9416=>"010110111",
  9417=>"011101000",
  9418=>"000011010",
  9419=>"010110011",
  9420=>"011100000",
  9421=>"000001000",
  9422=>"001011111",
  9423=>"110110010",
  9424=>"101110001",
  9425=>"101010101",
  9426=>"011010110",
  9427=>"110010110",
  9428=>"110011010",
  9429=>"010000101",
  9430=>"010011101",
  9431=>"101000011",
  9432=>"111000010",
  9433=>"101000100",
  9434=>"100100001",
  9435=>"011010011",
  9436=>"010000011",
  9437=>"111101111",
  9438=>"101110001",
  9439=>"000001010",
  9440=>"010011101",
  9441=>"011001010",
  9442=>"010100001",
  9443=>"001111000",
  9444=>"010110100",
  9445=>"100111011",
  9446=>"110111001",
  9447=>"011010110",
  9448=>"100001111",
  9449=>"000000110",
  9450=>"001100010",
  9451=>"100000010",
  9452=>"000000111",
  9453=>"101000110",
  9454=>"110111010",
  9455=>"001110111",
  9456=>"010010110",
  9457=>"111001000",
  9458=>"011001011",
  9459=>"011001000",
  9460=>"010110111",
  9461=>"101000110",
  9462=>"011000000",
  9463=>"100000111",
  9464=>"101001100",
  9465=>"010100101",
  9466=>"001011001",
  9467=>"010011101",
  9468=>"110001011",
  9469=>"010110110",
  9470=>"101010110",
  9471=>"000001001",
  9472=>"101110111",
  9473=>"111001110",
  9474=>"101110010",
  9475=>"111110110",
  9476=>"111001010",
  9477=>"100001001",
  9478=>"100100010",
  9479=>"101100011",
  9480=>"010111001",
  9481=>"001110100",
  9482=>"010001111",
  9483=>"000100011",
  9484=>"001010101",
  9485=>"011010011",
  9486=>"100011110",
  9487=>"100100111",
  9488=>"000001110",
  9489=>"011110110",
  9490=>"101110111",
  9491=>"100110000",
  9492=>"001001010",
  9493=>"110100110",
  9494=>"111011101",
  9495=>"010010101",
  9496=>"100110001",
  9497=>"010110101",
  9498=>"110000100",
  9499=>"100010010",
  9500=>"110000001",
  9501=>"000010000",
  9502=>"010111101",
  9503=>"010010101",
  9504=>"001001001",
  9505=>"001101000",
  9506=>"111000110",
  9507=>"110010001",
  9508=>"000111110",
  9509=>"010110000",
  9510=>"111010000",
  9511=>"100011001",
  9512=>"010000011",
  9513=>"001101010",
  9514=>"010101011",
  9515=>"101001101",
  9516=>"111010011",
  9517=>"100110010",
  9518=>"110100110",
  9519=>"011110010",
  9520=>"000010010",
  9521=>"011110101",
  9522=>"010011001",
  9523=>"111111111",
  9524=>"110100001",
  9525=>"001000010",
  9526=>"011110011",
  9527=>"101011111",
  9528=>"001011011",
  9529=>"100000110",
  9530=>"100111101",
  9531=>"010100011",
  9532=>"001001100",
  9533=>"111000100",
  9534=>"000100010",
  9535=>"111111110",
  9536=>"100101100",
  9537=>"000000001",
  9538=>"011010101",
  9539=>"101110110",
  9540=>"111110011",
  9541=>"100111001",
  9542=>"011100111",
  9543=>"100001011",
  9544=>"000001001",
  9545=>"011110011",
  9546=>"100011110",
  9547=>"011000000",
  9548=>"001110101",
  9549=>"001111111",
  9550=>"010000011",
  9551=>"011110011",
  9552=>"110011010",
  9553=>"100110111",
  9554=>"000110100",
  9555=>"010001000",
  9556=>"010010111",
  9557=>"111010111",
  9558=>"110011001",
  9559=>"100011010",
  9560=>"100101111",
  9561=>"111110110",
  9562=>"010011010",
  9563=>"010101100",
  9564=>"011111000",
  9565=>"011101011",
  9566=>"110101100",
  9567=>"110111011",
  9568=>"101111110",
  9569=>"111001101",
  9570=>"010101101",
  9571=>"110001001",
  9572=>"101100101",
  9573=>"000110000",
  9574=>"100101000",
  9575=>"011111011",
  9576=>"001000101",
  9577=>"000000100",
  9578=>"111111110",
  9579=>"011111110",
  9580=>"100011100",
  9581=>"110001110",
  9582=>"110001001",
  9583=>"110111000",
  9584=>"010110011",
  9585=>"110000110",
  9586=>"010010011",
  9587=>"100100000",
  9588=>"001101010",
  9589=>"110110001",
  9590=>"000001111",
  9591=>"100110110",
  9592=>"101100000",
  9593=>"010101001",
  9594=>"001011011",
  9595=>"110010111",
  9596=>"010110110",
  9597=>"000000010",
  9598=>"010100101",
  9599=>"000101000",
  9600=>"111111010",
  9601=>"101000011",
  9602=>"110010011",
  9603=>"111001010",
  9604=>"010000000",
  9605=>"110001001",
  9606=>"110111010",
  9607=>"000000000",
  9608=>"101111001",
  9609=>"011100110",
  9610=>"100101011",
  9611=>"010000011",
  9612=>"111111100",
  9613=>"101010000",
  9614=>"011111011",
  9615=>"101001010",
  9616=>"001011111",
  9617=>"000001000",
  9618=>"100001101",
  9619=>"111011111",
  9620=>"111111100",
  9621=>"000011100",
  9622=>"000010010",
  9623=>"101001010",
  9624=>"111001101",
  9625=>"101001011",
  9626=>"110111100",
  9627=>"000101001",
  9628=>"000011011",
  9629=>"011101110",
  9630=>"101101101",
  9631=>"010010110",
  9632=>"000001111",
  9633=>"011001010",
  9634=>"100110010",
  9635=>"000100100",
  9636=>"101110100",
  9637=>"000001110",
  9638=>"010000000",
  9639=>"101010111",
  9640=>"010000110",
  9641=>"001001001",
  9642=>"000010010",
  9643=>"011001011",
  9644=>"001111100",
  9645=>"010010111",
  9646=>"111100100",
  9647=>"001011101",
  9648=>"001100001",
  9649=>"011011100",
  9650=>"010000000",
  9651=>"001111010",
  9652=>"111111000",
  9653=>"010010100",
  9654=>"001011000",
  9655=>"101110110",
  9656=>"011000111",
  9657=>"101000111",
  9658=>"010011011",
  9659=>"100000000",
  9660=>"111011111",
  9661=>"110000110",
  9662=>"101011111",
  9663=>"110100101",
  9664=>"101001010",
  9665=>"010101011",
  9666=>"100111111",
  9667=>"110000001",
  9668=>"110000110",
  9669=>"010110000",
  9670=>"110011100",
  9671=>"001000011",
  9672=>"011010011",
  9673=>"111001010",
  9674=>"001000001",
  9675=>"100101011",
  9676=>"000001100",
  9677=>"111010100",
  9678=>"011111010",
  9679=>"101100100",
  9680=>"101011011",
  9681=>"011110111",
  9682=>"010010001",
  9683=>"000100100",
  9684=>"010111111",
  9685=>"001100011",
  9686=>"110101101",
  9687=>"011000001",
  9688=>"001101010",
  9689=>"001101011",
  9690=>"111111010",
  9691=>"101001011",
  9692=>"111000100",
  9693=>"101000011",
  9694=>"001110010",
  9695=>"110110110",
  9696=>"010110011",
  9697=>"100111100",
  9698=>"100110101",
  9699=>"111001010",
  9700=>"100011000",
  9701=>"000011000",
  9702=>"001000000",
  9703=>"110000001",
  9704=>"101101000",
  9705=>"111111100",
  9706=>"100010000",
  9707=>"101001101",
  9708=>"000111011",
  9709=>"011000111",
  9710=>"111000110",
  9711=>"110101111",
  9712=>"000000110",
  9713=>"001111110",
  9714=>"110111000",
  9715=>"101110010",
  9716=>"000010010",
  9717=>"000110111",
  9718=>"111011101",
  9719=>"100000011",
  9720=>"000011100",
  9721=>"110000001",
  9722=>"000100101",
  9723=>"001110001",
  9724=>"111011100",
  9725=>"110111100",
  9726=>"000001000",
  9727=>"010100110",
  9728=>"100111001",
  9729=>"000010000",
  9730=>"100011100",
  9731=>"101111010",
  9732=>"111010110",
  9733=>"000001000",
  9734=>"010010110",
  9735=>"110000010",
  9736=>"001000100",
  9737=>"111100011",
  9738=>"111100111",
  9739=>"111100100",
  9740=>"101111011",
  9741=>"111000101",
  9742=>"110111011",
  9743=>"010101001",
  9744=>"101100000",
  9745=>"100000010",
  9746=>"000111001",
  9747=>"110001001",
  9748=>"110101000",
  9749=>"110110101",
  9750=>"011000111",
  9751=>"000101011",
  9752=>"110111111",
  9753=>"000101111",
  9754=>"000100111",
  9755=>"010010111",
  9756=>"010010010",
  9757=>"010010010",
  9758=>"101101100",
  9759=>"000011011",
  9760=>"101000001",
  9761=>"101101001",
  9762=>"000010011",
  9763=>"101101001",
  9764=>"010000101",
  9765=>"111110001",
  9766=>"101111000",
  9767=>"010110110",
  9768=>"010010110",
  9769=>"101111001",
  9770=>"110000001",
  9771=>"101011100",
  9772=>"110010101",
  9773=>"110001100",
  9774=>"110001001",
  9775=>"101101101",
  9776=>"011000001",
  9777=>"001001110",
  9778=>"101000111",
  9779=>"101010110",
  9780=>"010100000",
  9781=>"000100000",
  9782=>"101010110",
  9783=>"011000101",
  9784=>"010000111",
  9785=>"101000000",
  9786=>"010011011",
  9787=>"110011001",
  9788=>"010111111",
  9789=>"101001010",
  9790=>"000101100",
  9791=>"111011110",
  9792=>"100000001",
  9793=>"001101001",
  9794=>"110001110",
  9795=>"011111100",
  9796=>"000001000",
  9797=>"000100011",
  9798=>"101011101",
  9799=>"111011100",
  9800=>"000000101",
  9801=>"000001000",
  9802=>"100010111",
  9803=>"101101010",
  9804=>"110010001",
  9805=>"001001001",
  9806=>"101111010",
  9807=>"010001010",
  9808=>"001101010",
  9809=>"001001111",
  9810=>"100010011",
  9811=>"001100101",
  9812=>"110111011",
  9813=>"011000101",
  9814=>"010010111",
  9815=>"011101011",
  9816=>"011011110",
  9817=>"001000110",
  9818=>"100101100",
  9819=>"011110011",
  9820=>"010011110",
  9821=>"000001010",
  9822=>"000011111",
  9823=>"110111111",
  9824=>"010011001",
  9825=>"101100010",
  9826=>"001111000",
  9827=>"000111001",
  9828=>"000000001",
  9829=>"001110110",
  9830=>"010111101",
  9831=>"100111000",
  9832=>"011000011",
  9833=>"010010011",
  9834=>"101100110",
  9835=>"000011110",
  9836=>"000011101",
  9837=>"100011001",
  9838=>"101011111",
  9839=>"110111000",
  9840=>"110110100",
  9841=>"101110001",
  9842=>"100110011",
  9843=>"010011100",
  9844=>"001011001",
  9845=>"011101001",
  9846=>"010010001",
  9847=>"011111001",
  9848=>"000101100",
  9849=>"000011001",
  9850=>"101000000",
  9851=>"011111110",
  9852=>"101110011",
  9853=>"000100111",
  9854=>"010011000",
  9855=>"101011111",
  9856=>"110111111",
  9857=>"001001010",
  9858=>"111011001",
  9859=>"100000110",
  9860=>"001100110",
  9861=>"010001011",
  9862=>"111011100",
  9863=>"010111010",
  9864=>"111111000",
  9865=>"010100101",
  9866=>"000001011",
  9867=>"101011110",
  9868=>"011010111",
  9869=>"101111110",
  9870=>"111010011",
  9871=>"101011001",
  9872=>"110010101",
  9873=>"101101010",
  9874=>"011010011",
  9875=>"110011010",
  9876=>"001010100",
  9877=>"011001010",
  9878=>"010010111",
  9879=>"010101110",
  9880=>"101000111",
  9881=>"111101101",
  9882=>"111101111",
  9883=>"011011010",
  9884=>"101111011",
  9885=>"111001011",
  9886=>"101100011",
  9887=>"000011001",
  9888=>"000011000",
  9889=>"101000011",
  9890=>"000000100",
  9891=>"101010100",
  9892=>"100101001",
  9893=>"001001101",
  9894=>"100110100",
  9895=>"010100000",
  9896=>"110001010",
  9897=>"101011001",
  9898=>"101011110",
  9899=>"011100111",
  9900=>"110111100",
  9901=>"011011011",
  9902=>"010110011",
  9903=>"100000100",
  9904=>"010100011",
  9905=>"001000101",
  9906=>"000001011",
  9907=>"100101100",
  9908=>"000110111",
  9909=>"101101000",
  9910=>"111111100",
  9911=>"100100000",
  9912=>"001111010",
  9913=>"111101110",
  9914=>"111100101",
  9915=>"001011111",
  9916=>"110000010",
  9917=>"110001010",
  9918=>"001111100",
  9919=>"001110011",
  9920=>"001110100",
  9921=>"100011101",
  9922=>"011001010",
  9923=>"101000100",
  9924=>"001100101",
  9925=>"110111101",
  9926=>"001000001",
  9927=>"101010100",
  9928=>"101100110",
  9929=>"101101011",
  9930=>"101011011",
  9931=>"111111101",
  9932=>"101111000",
  9933=>"010100011",
  9934=>"011000111",
  9935=>"101111011",
  9936=>"010001000",
  9937=>"100100010",
  9938=>"010100110",
  9939=>"101011100",
  9940=>"010011101",
  9941=>"001000001",
  9942=>"101101111",
  9943=>"111111100",
  9944=>"000000111",
  9945=>"010111001",
  9946=>"001011111",
  9947=>"101011110",
  9948=>"011111011",
  9949=>"111001101",
  9950=>"100101101",
  9951=>"110110110",
  9952=>"011011000",
  9953=>"010101001",
  9954=>"111011100",
  9955=>"000000011",
  9956=>"011011110",
  9957=>"010010000",
  9958=>"101001011",
  9959=>"000000010",
  9960=>"001011110",
  9961=>"011011111",
  9962=>"011001101",
  9963=>"111111111",
  9964=>"010110000",
  9965=>"111101000",
  9966=>"100100001",
  9967=>"001011100",
  9968=>"010000010",
  9969=>"100101000",
  9970=>"000010010",
  9971=>"101111010",
  9972=>"101000010",
  9973=>"000011100",
  9974=>"111100011",
  9975=>"101101111",
  9976=>"101100001",
  9977=>"100001101",
  9978=>"101111010",
  9979=>"111100100",
  9980=>"101101100",
  9981=>"101010100",
  9982=>"111100101",
  9983=>"110100101",
  9984=>"010100110",
  9985=>"001010011",
  9986=>"110110011",
  9987=>"101101100",
  9988=>"011001111",
  9989=>"011111010",
  9990=>"011111100",
  9991=>"000100000",
  9992=>"010111111",
  9993=>"001111111",
  9994=>"111110000",
  9995=>"011010011",
  9996=>"000111100",
  9997=>"010100111",
  9998=>"000111111",
  9999=>"110111010",
  10000=>"110110010",
  10001=>"100100101",
  10002=>"111010111",
  10003=>"010010111",
  10004=>"101101000",
  10005=>"000010100",
  10006=>"110000111",
  10007=>"100101001",
  10008=>"101101011",
  10009=>"001111111",
  10010=>"000000110",
  10011=>"110000001",
  10012=>"000101001",
  10013=>"011011100",
  10014=>"101011000",
  10015=>"100101000",
  10016=>"111111000",
  10017=>"001001001",
  10018=>"111000110",
  10019=>"111010101",
  10020=>"000100000",
  10021=>"000101010",
  10022=>"010100001",
  10023=>"100111100",
  10024=>"111010101",
  10025=>"111001010",
  10026=>"110011100",
  10027=>"010111010",
  10028=>"001111010",
  10029=>"000001110",
  10030=>"111110101",
  10031=>"100011010",
  10032=>"110011101",
  10033=>"100111011",
  10034=>"000010100",
  10035=>"101101101",
  10036=>"010000001",
  10037=>"000111100",
  10038=>"010001001",
  10039=>"001011010",
  10040=>"101000101",
  10041=>"001001110",
  10042=>"000001010",
  10043=>"010101111",
  10044=>"101101101",
  10045=>"001011000",
  10046=>"110000001",
  10047=>"110110001",
  10048=>"010000000",
  10049=>"100010101",
  10050=>"011101100",
  10051=>"010000011",
  10052=>"001101011",
  10053=>"011010101",
  10054=>"101110001",
  10055=>"001010001",
  10056=>"011000001",
  10057=>"111011111",
  10058=>"011001011",
  10059=>"100001101",
  10060=>"110110000",
  10061=>"111010101",
  10062=>"110000001",
  10063=>"010111011",
  10064=>"001001111",
  10065=>"000101000",
  10066=>"100100100",
  10067=>"000011011",
  10068=>"000110011",
  10069=>"010010101",
  10070=>"011100111",
  10071=>"000100001",
  10072=>"100100011",
  10073=>"001110100",
  10074=>"101010110",
  10075=>"110101100",
  10076=>"001110011",
  10077=>"111100110",
  10078=>"110011101",
  10079=>"001010101",
  10080=>"000101101",
  10081=>"011010110",
  10082=>"001001010",
  10083=>"010011001",
  10084=>"101111101",
  10085=>"111001100",
  10086=>"111001100",
  10087=>"001101100",
  10088=>"111010001",
  10089=>"100111101",
  10090=>"110010111",
  10091=>"101001101",
  10092=>"011100101",
  10093=>"111110011",
  10094=>"001100000",
  10095=>"000001101",
  10096=>"101111110",
  10097=>"001000101",
  10098=>"111100001",
  10099=>"111111111",
  10100=>"000011000",
  10101=>"110001001",
  10102=>"111001101",
  10103=>"101110110",
  10104=>"000001111",
  10105=>"000011010",
  10106=>"111000001",
  10107=>"111111111",
  10108=>"111011001",
  10109=>"000100011",
  10110=>"101011000",
  10111=>"011000110",
  10112=>"011101010",
  10113=>"000110111",
  10114=>"000011001",
  10115=>"110001111",
  10116=>"111101101",
  10117=>"010010001",
  10118=>"001111101",
  10119=>"011010001",
  10120=>"101110010",
  10121=>"010000011",
  10122=>"000100000",
  10123=>"011101101",
  10124=>"010010100",
  10125=>"000001101",
  10126=>"010000101",
  10127=>"110001011",
  10128=>"001110001",
  10129=>"110110010",
  10130=>"000111110",
  10131=>"011000100",
  10132=>"000101000",
  10133=>"001010001",
  10134=>"000100001",
  10135=>"001000100",
  10136=>"100001111",
  10137=>"000010001",
  10138=>"000010101",
  10139=>"101010101",
  10140=>"101001000",
  10141=>"111001001",
  10142=>"110010010",
  10143=>"111011111",
  10144=>"000101011",
  10145=>"001011001",
  10146=>"101001001",
  10147=>"111101100",
  10148=>"100011010",
  10149=>"000111011",
  10150=>"000100100",
  10151=>"111011010",
  10152=>"110000011",
  10153=>"011000000",
  10154=>"111101001",
  10155=>"011001000",
  10156=>"000000010",
  10157=>"010001100",
  10158=>"010011100",
  10159=>"011101110",
  10160=>"111011000",
  10161=>"010000101",
  10162=>"011101111",
  10163=>"000001001",
  10164=>"101011111",
  10165=>"110000010",
  10166=>"001110001",
  10167=>"001110111",
  10168=>"001010010",
  10169=>"110101110",
  10170=>"110001110",
  10171=>"101100000",
  10172=>"110100010",
  10173=>"110100010",
  10174=>"010110101",
  10175=>"000001001",
  10176=>"101010111",
  10177=>"101000011",
  10178=>"001010000",
  10179=>"100111011",
  10180=>"101110011",
  10181=>"000101100",
  10182=>"010000010",
  10183=>"010000100",
  10184=>"100010110",
  10185=>"001101101",
  10186=>"001100101",
  10187=>"001100111",
  10188=>"100010000",
  10189=>"101000011",
  10190=>"010010100",
  10191=>"101110000",
  10192=>"010101010",
  10193=>"100111111",
  10194=>"000100110",
  10195=>"110111000",
  10196=>"110000000",
  10197=>"011100111",
  10198=>"001001110",
  10199=>"101100001",
  10200=>"111001001",
  10201=>"000100110",
  10202=>"110001101",
  10203=>"000011100",
  10204=>"011000101",
  10205=>"101011111",
  10206=>"010001001",
  10207=>"110000110",
  10208=>"011111000",
  10209=>"100111111",
  10210=>"101101100",
  10211=>"111001101",
  10212=>"001100011",
  10213=>"111111101",
  10214=>"000101110",
  10215=>"110001010",
  10216=>"011011100",
  10217=>"011001100",
  10218=>"011100010",
  10219=>"101101100",
  10220=>"011101010",
  10221=>"110110111",
  10222=>"110110111",
  10223=>"011001110",
  10224=>"001110100",
  10225=>"100111101",
  10226=>"001100110",
  10227=>"110100110",
  10228=>"011111101",
  10229=>"011000100",
  10230=>"111011011",
  10231=>"110011100",
  10232=>"111010011",
  10233=>"011111110",
  10234=>"101100100",
  10235=>"100110011",
  10236=>"101000111",
  10237=>"101100010",
  10238=>"111100110",
  10239=>"101100100",
  10240=>"100110100",
  10241=>"111010010",
  10242=>"100101011",
  10243=>"011110111",
  10244=>"100110101",
  10245=>"101011001",
  10246=>"001010001",
  10247=>"000010010",
  10248=>"010001110",
  10249=>"011001111",
  10250=>"010010001",
  10251=>"001110001",
  10252=>"010001010",
  10253=>"011010000",
  10254=>"000011001",
  10255=>"001001000",
  10256=>"011001011",
  10257=>"011101101",
  10258=>"010110101",
  10259=>"001111100",
  10260=>"001111100",
  10261=>"100010010",
  10262=>"110111100",
  10263=>"010001001",
  10264=>"010000110",
  10265=>"001001011",
  10266=>"100100010",
  10267=>"000110001",
  10268=>"000000000",
  10269=>"010111101",
  10270=>"101010010",
  10271=>"110000000",
  10272=>"101000001",
  10273=>"110111110",
  10274=>"100111111",
  10275=>"000101100",
  10276=>"011010001",
  10277=>"011011101",
  10278=>"001011001",
  10279=>"100100011",
  10280=>"010010001",
  10281=>"000110011",
  10282=>"010000000",
  10283=>"110000110",
  10284=>"111011110",
  10285=>"011010001",
  10286=>"110001000",
  10287=>"001011110",
  10288=>"100101001",
  10289=>"111000101",
  10290=>"000110010",
  10291=>"111001110",
  10292=>"001010000",
  10293=>"110001000",
  10294=>"110111100",
  10295=>"110100000",
  10296=>"000101001",
  10297=>"110000001",
  10298=>"000001110",
  10299=>"100110111",
  10300=>"111111010",
  10301=>"000011101",
  10302=>"011100001",
  10303=>"011110000",
  10304=>"010000000",
  10305=>"010101111",
  10306=>"111001011",
  10307=>"100111001",
  10308=>"010110110",
  10309=>"110011001",
  10310=>"001110111",
  10311=>"110111001",
  10312=>"010001010",
  10313=>"010011101",
  10314=>"001000000",
  10315=>"000000010",
  10316=>"000011111",
  10317=>"010001100",
  10318=>"000000001",
  10319=>"101001000",
  10320=>"000000110",
  10321=>"000101010",
  10322=>"101101001",
  10323=>"010100011",
  10324=>"010100101",
  10325=>"000101000",
  10326=>"011111011",
  10327=>"001010000",
  10328=>"101111001",
  10329=>"110111110",
  10330=>"111100101",
  10331=>"111001110",
  10332=>"011010010",
  10333=>"001001101",
  10334=>"110111100",
  10335=>"010110111",
  10336=>"111001011",
  10337=>"001001000",
  10338=>"001010011",
  10339=>"011011000",
  10340=>"001010001",
  10341=>"101010010",
  10342=>"100011111",
  10343=>"001110000",
  10344=>"000001100",
  10345=>"010001110",
  10346=>"010101111",
  10347=>"010001101",
  10348=>"000110000",
  10349=>"111010111",
  10350=>"010110000",
  10351=>"011010010",
  10352=>"110111100",
  10353=>"010101100",
  10354=>"101010010",
  10355=>"100110111",
  10356=>"011111110",
  10357=>"110111110",
  10358=>"110110001",
  10359=>"101000001",
  10360=>"001010011",
  10361=>"100010001",
  10362=>"000100011",
  10363=>"100101010",
  10364=>"001111010",
  10365=>"100001100",
  10366=>"110100101",
  10367=>"000010010",
  10368=>"110000010",
  10369=>"001100111",
  10370=>"010001010",
  10371=>"111011110",
  10372=>"111000100",
  10373=>"000000000",
  10374=>"010101110",
  10375=>"111110111",
  10376=>"111111100",
  10377=>"001110111",
  10378=>"110100111",
  10379=>"101110100",
  10380=>"000100100",
  10381=>"100011111",
  10382=>"001100101",
  10383=>"011111100",
  10384=>"010100110",
  10385=>"011010110",
  10386=>"000000010",
  10387=>"011000101",
  10388=>"000011010",
  10389=>"011001101",
  10390=>"101010110",
  10391=>"000101110",
  10392=>"010001111",
  10393=>"000000000",
  10394=>"010101010",
  10395=>"111101101",
  10396=>"000011001",
  10397=>"101011001",
  10398=>"100110110",
  10399=>"001011001",
  10400=>"110111111",
  10401=>"001010110",
  10402=>"111111101",
  10403=>"000001010",
  10404=>"000100110",
  10405=>"000011011",
  10406=>"101110110",
  10407=>"100011010",
  10408=>"011010001",
  10409=>"101101011",
  10410=>"010100010",
  10411=>"011011000",
  10412=>"001000100",
  10413=>"100011111",
  10414=>"000001111",
  10415=>"011010111",
  10416=>"101000011",
  10417=>"111101110",
  10418=>"011100101",
  10419=>"111010011",
  10420=>"001001111",
  10421=>"100011111",
  10422=>"100110001",
  10423=>"111001110",
  10424=>"111011110",
  10425=>"000010000",
  10426=>"110101010",
  10427=>"010001000",
  10428=>"101100110",
  10429=>"001011101",
  10430=>"111010011",
  10431=>"110000000",
  10432=>"101100000",
  10433=>"101110011",
  10434=>"111111100",
  10435=>"010011011",
  10436=>"011000001",
  10437=>"000000110",
  10438=>"110111001",
  10439=>"110011000",
  10440=>"000111010",
  10441=>"000001101",
  10442=>"000110100",
  10443=>"111110001",
  10444=>"010000110",
  10445=>"100111111",
  10446=>"001110011",
  10447=>"010010100",
  10448=>"111100001",
  10449=>"110000010",
  10450=>"100101111",
  10451=>"001011100",
  10452=>"011110100",
  10453=>"011101100",
  10454=>"101000001",
  10455=>"000100111",
  10456=>"001011000",
  10457=>"100010010",
  10458=>"000101011",
  10459=>"011110100",
  10460=>"101101110",
  10461=>"011011110",
  10462=>"010001011",
  10463=>"010100101",
  10464=>"000100000",
  10465=>"001001001",
  10466=>"101111101",
  10467=>"111000111",
  10468=>"001000101",
  10469=>"001000001",
  10470=>"000011111",
  10471=>"111010000",
  10472=>"000011000",
  10473=>"001011001",
  10474=>"010010100",
  10475=>"100010111",
  10476=>"100000101",
  10477=>"100010101",
  10478=>"010001110",
  10479=>"101111111",
  10480=>"010101010",
  10481=>"000000010",
  10482=>"011100001",
  10483=>"111000111",
  10484=>"000001100",
  10485=>"110011001",
  10486=>"001101111",
  10487=>"001100010",
  10488=>"001000101",
  10489=>"010011010",
  10490=>"101100100",
  10491=>"101000111",
  10492=>"100101000",
  10493=>"011001000",
  10494=>"001101111",
  10495=>"110011001",
  10496=>"010011000",
  10497=>"001001110",
  10498=>"001111111",
  10499=>"111111011",
  10500=>"011011001",
  10501=>"010010110",
  10502=>"011110110",
  10503=>"000101011",
  10504=>"110111101",
  10505=>"000010000",
  10506=>"100100100",
  10507=>"100100100",
  10508=>"011011000",
  10509=>"101011011",
  10510=>"000100011",
  10511=>"110011100",
  10512=>"011010111",
  10513=>"011000000",
  10514=>"111010010",
  10515=>"011100011",
  10516=>"001011111",
  10517=>"100010001",
  10518=>"011110011",
  10519=>"100000100",
  10520=>"010010010",
  10521=>"110101010",
  10522=>"100010000",
  10523=>"100010010",
  10524=>"011011101",
  10525=>"001110111",
  10526=>"001001100",
  10527=>"010010001",
  10528=>"100100100",
  10529=>"111010100",
  10530=>"110101001",
  10531=>"000100001",
  10532=>"111110100",
  10533=>"110000100",
  10534=>"001110111",
  10535=>"111000101",
  10536=>"010001110",
  10537=>"101000001",
  10538=>"000101010",
  10539=>"111010000",
  10540=>"111111100",
  10541=>"000000011",
  10542=>"000110010",
  10543=>"110110111",
  10544=>"101110000",
  10545=>"010001110",
  10546=>"100111010",
  10547=>"010001010",
  10548=>"001111111",
  10549=>"000000010",
  10550=>"000100001",
  10551=>"100001010",
  10552=>"101010100",
  10553=>"010000010",
  10554=>"110001110",
  10555=>"011110000",
  10556=>"111101111",
  10557=>"101111110",
  10558=>"001001000",
  10559=>"111001101",
  10560=>"110100000",
  10561=>"110001101",
  10562=>"011000100",
  10563=>"000101010",
  10564=>"001100000",
  10565=>"101010111",
  10566=>"100100101",
  10567=>"101111010",
  10568=>"000110111",
  10569=>"011101000",
  10570=>"100011010",
  10571=>"110100001",
  10572=>"011011100",
  10573=>"011101011",
  10574=>"110010010",
  10575=>"110100000",
  10576=>"001110001",
  10577=>"000000001",
  10578=>"111100010",
  10579=>"001110001",
  10580=>"110111000",
  10581=>"011001101",
  10582=>"011100111",
  10583=>"000001111",
  10584=>"001110100",
  10585=>"011000011",
  10586=>"010001011",
  10587=>"100011111",
  10588=>"001111110",
  10589=>"111001101",
  10590=>"101001001",
  10591=>"000111100",
  10592=>"100100010",
  10593=>"101110010",
  10594=>"000001000",
  10595=>"001110010",
  10596=>"011110110",
  10597=>"111110111",
  10598=>"011001001",
  10599=>"100110100",
  10600=>"101111111",
  10601=>"000110000",
  10602=>"110001010",
  10603=>"111101011",
  10604=>"110111100",
  10605=>"111100100",
  10606=>"000000111",
  10607=>"111011100",
  10608=>"101000110",
  10609=>"101010000",
  10610=>"000110001",
  10611=>"010011011",
  10612=>"100101110",
  10613=>"101001010",
  10614=>"000000111",
  10615=>"111000100",
  10616=>"011101010",
  10617=>"101000111",
  10618=>"000010110",
  10619=>"100010001",
  10620=>"000010100",
  10621=>"000101011",
  10622=>"001100011",
  10623=>"110011001",
  10624=>"101101000",
  10625=>"011111110",
  10626=>"011101011",
  10627=>"011101000",
  10628=>"010010010",
  10629=>"100111100",
  10630=>"111010111",
  10631=>"000101111",
  10632=>"000101100",
  10633=>"111001111",
  10634=>"100011100",
  10635=>"001000100",
  10636=>"100110010",
  10637=>"101010101",
  10638=>"010011001",
  10639=>"011101001",
  10640=>"011110000",
  10641=>"110101000",
  10642=>"110001010",
  10643=>"010000110",
  10644=>"100010010",
  10645=>"110111011",
  10646=>"001001100",
  10647=>"101100101",
  10648=>"011000100",
  10649=>"110110101",
  10650=>"100010010",
  10651=>"101000101",
  10652=>"100101101",
  10653=>"011100110",
  10654=>"100010101",
  10655=>"100110100",
  10656=>"110100011",
  10657=>"110100110",
  10658=>"010000001",
  10659=>"011111000",
  10660=>"011100101",
  10661=>"001001100",
  10662=>"110010110",
  10663=>"111111011",
  10664=>"101101000",
  10665=>"010010101",
  10666=>"010001011",
  10667=>"000010101",
  10668=>"110110011",
  10669=>"110011101",
  10670=>"111111111",
  10671=>"011100100",
  10672=>"000111101",
  10673=>"010010000",
  10674=>"111010011",
  10675=>"011110010",
  10676=>"010100111",
  10677=>"011010000",
  10678=>"100111111",
  10679=>"111111010",
  10680=>"001101010",
  10681=>"110010000",
  10682=>"011111000",
  10683=>"011011100",
  10684=>"110110011",
  10685=>"110111010",
  10686=>"111110101",
  10687=>"110111000",
  10688=>"011001001",
  10689=>"000100000",
  10690=>"110100101",
  10691=>"110111110",
  10692=>"111111110",
  10693=>"000000110",
  10694=>"111000111",
  10695=>"010101101",
  10696=>"101101111",
  10697=>"101000000",
  10698=>"000110100",
  10699=>"100110001",
  10700=>"101100100",
  10701=>"111010101",
  10702=>"000010001",
  10703=>"110110101",
  10704=>"100001100",
  10705=>"101111111",
  10706=>"100111000",
  10707=>"111011011",
  10708=>"010111110",
  10709=>"101100101",
  10710=>"100111101",
  10711=>"011000100",
  10712=>"011001011",
  10713=>"010000000",
  10714=>"011100001",
  10715=>"111110001",
  10716=>"001010000",
  10717=>"101110011",
  10718=>"100001101",
  10719=>"010100110",
  10720=>"100011011",
  10721=>"101011011",
  10722=>"010011010",
  10723=>"011001111",
  10724=>"100010011",
  10725=>"001011011",
  10726=>"101110101",
  10727=>"100110010",
  10728=>"100110011",
  10729=>"010111011",
  10730=>"110010111",
  10731=>"011011010",
  10732=>"101111001",
  10733=>"011111011",
  10734=>"010010101",
  10735=>"111111111",
  10736=>"101001100",
  10737=>"000010001",
  10738=>"110100000",
  10739=>"001111111",
  10740=>"000111110",
  10741=>"101100011",
  10742=>"101011011",
  10743=>"100100000",
  10744=>"101100000",
  10745=>"001010100",
  10746=>"101001000",
  10747=>"001010010",
  10748=>"001001001",
  10749=>"111100100",
  10750=>"010110100",
  10751=>"010010001",
  10752=>"100111011",
  10753=>"000110011",
  10754=>"110011001",
  10755=>"000100110",
  10756=>"001010011",
  10757=>"011010111",
  10758=>"010110000",
  10759=>"000010110",
  10760=>"100111000",
  10761=>"111101100",
  10762=>"001011101",
  10763=>"011000001",
  10764=>"010101100",
  10765=>"000001011",
  10766=>"001101011",
  10767=>"100010001",
  10768=>"111100010",
  10769=>"101011110",
  10770=>"001010001",
  10771=>"110000000",
  10772=>"001000001",
  10773=>"100000001",
  10774=>"010001000",
  10775=>"000111011",
  10776=>"011011110",
  10777=>"101100111",
  10778=>"110001010",
  10779=>"000101111",
  10780=>"101101000",
  10781=>"111110111",
  10782=>"011010011",
  10783=>"001010110",
  10784=>"000100010",
  10785=>"101111010",
  10786=>"111001101",
  10787=>"010100101",
  10788=>"000001000",
  10789=>"111101101",
  10790=>"101001110",
  10791=>"011001100",
  10792=>"010100000",
  10793=>"001110101",
  10794=>"101111010",
  10795=>"000111000",
  10796=>"000000000",
  10797=>"001011110",
  10798=>"001110101",
  10799=>"101110011",
  10800=>"000100000",
  10801=>"100001000",
  10802=>"101010001",
  10803=>"001011010",
  10804=>"111011000",
  10805=>"110110100",
  10806=>"101111011",
  10807=>"100110010",
  10808=>"010011010",
  10809=>"100001110",
  10810=>"001011000",
  10811=>"011110111",
  10812=>"000100001",
  10813=>"100011101",
  10814=>"110100000",
  10815=>"000010011",
  10816=>"000100000",
  10817=>"000001110",
  10818=>"111101001",
  10819=>"111001010",
  10820=>"100001010",
  10821=>"011011100",
  10822=>"101011101",
  10823=>"110011110",
  10824=>"010101100",
  10825=>"111101011",
  10826=>"111010010",
  10827=>"001001111",
  10828=>"011001110",
  10829=>"101010000",
  10830=>"111100100",
  10831=>"000100111",
  10832=>"111011010",
  10833=>"101110100",
  10834=>"101000001",
  10835=>"111000100",
  10836=>"000100001",
  10837=>"110010001",
  10838=>"001101011",
  10839=>"110100001",
  10840=>"010010010",
  10841=>"100011100",
  10842=>"010010111",
  10843=>"011111010",
  10844=>"000111111",
  10845=>"010101010",
  10846=>"000011110",
  10847=>"111101101",
  10848=>"001110011",
  10849=>"011000111",
  10850=>"010010000",
  10851=>"001001100",
  10852=>"110111100",
  10853=>"100100010",
  10854=>"000010011",
  10855=>"100001010",
  10856=>"001101110",
  10857=>"001101010",
  10858=>"001010000",
  10859=>"010000011",
  10860=>"011001100",
  10861=>"100010010",
  10862=>"001000010",
  10863=>"110011100",
  10864=>"010111110",
  10865=>"111000100",
  10866=>"111100000",
  10867=>"011001110",
  10868=>"010000110",
  10869=>"101111010",
  10870=>"100000000",
  10871=>"100011111",
  10872=>"000110000",
  10873=>"010010100",
  10874=>"101001010",
  10875=>"010100100",
  10876=>"001001111",
  10877=>"001100010",
  10878=>"101001011",
  10879=>"011110111",
  10880=>"000111010",
  10881=>"111111111",
  10882=>"111100101",
  10883=>"111000101",
  10884=>"010000110",
  10885=>"001001000",
  10886=>"011010001",
  10887=>"110101001",
  10888=>"101111101",
  10889=>"000111001",
  10890=>"110100110",
  10891=>"110100110",
  10892=>"100000010",
  10893=>"110011000",
  10894=>"111101011",
  10895=>"101101110",
  10896=>"111101010",
  10897=>"101011111",
  10898=>"011000010",
  10899=>"111100101",
  10900=>"110100110",
  10901=>"000110101",
  10902=>"101000111",
  10903=>"001111111",
  10904=>"100001101",
  10905=>"100011111",
  10906=>"001111001",
  10907=>"001011110",
  10908=>"111001011",
  10909=>"010110001",
  10910=>"110010111",
  10911=>"001101001",
  10912=>"001110101",
  10913=>"010001001",
  10914=>"011000001",
  10915=>"100110001",
  10916=>"010010111",
  10917=>"000000011",
  10918=>"111000011",
  10919=>"101101111",
  10920=>"011101111",
  10921=>"010100010",
  10922=>"100000110",
  10923=>"010110001",
  10924=>"101111000",
  10925=>"011000100",
  10926=>"010010010",
  10927=>"100000010",
  10928=>"010010011",
  10929=>"000111001",
  10930=>"001000010",
  10931=>"000001101",
  10932=>"000011110",
  10933=>"111110001",
  10934=>"010011001",
  10935=>"100101100",
  10936=>"110011001",
  10937=>"000111001",
  10938=>"001111000",
  10939=>"101011000",
  10940=>"100111110",
  10941=>"000000100",
  10942=>"100000110",
  10943=>"011110110",
  10944=>"101010010",
  10945=>"110110111",
  10946=>"111110100",
  10947=>"101001101",
  10948=>"111000010",
  10949=>"110101001",
  10950=>"010111010",
  10951=>"011111011",
  10952=>"101010011",
  10953=>"111111101",
  10954=>"000101101",
  10955=>"011101101",
  10956=>"111010111",
  10957=>"011111010",
  10958=>"111110010",
  10959=>"111110010",
  10960=>"110001100",
  10961=>"101000111",
  10962=>"111010111",
  10963=>"111000011",
  10964=>"000100100",
  10965=>"100111001",
  10966=>"110010011",
  10967=>"100001001",
  10968=>"110000000",
  10969=>"010000010",
  10970=>"110000111",
  10971=>"001011110",
  10972=>"001100011",
  10973=>"111100111",
  10974=>"000110100",
  10975=>"110110001",
  10976=>"100000011",
  10977=>"000011111",
  10978=>"001001101",
  10979=>"000000000",
  10980=>"111001111",
  10981=>"100000010",
  10982=>"011111110",
  10983=>"011110011",
  10984=>"011101000",
  10985=>"111110111",
  10986=>"100010111",
  10987=>"011110010",
  10988=>"010000010",
  10989=>"010011010",
  10990=>"101101010",
  10991=>"011001000",
  10992=>"101011010",
  10993=>"001000011",
  10994=>"000010101",
  10995=>"111110001",
  10996=>"111101101",
  10997=>"001011100",
  10998=>"010101101",
  10999=>"001100001",
  11000=>"001100011",
  11001=>"010111111",
  11002=>"110011100",
  11003=>"001101100",
  11004=>"111111100",
  11005=>"100011101",
  11006=>"110100000",
  11007=>"011011001",
  11008=>"111000001",
  11009=>"001111101",
  11010=>"011011101",
  11011=>"100011011",
  11012=>"000000111",
  11013=>"110010001",
  11014=>"001110001",
  11015=>"111111110",
  11016=>"110101011",
  11017=>"000011001",
  11018=>"001000011",
  11019=>"000000010",
  11020=>"001101000",
  11021=>"000111011",
  11022=>"110001101",
  11023=>"011011011",
  11024=>"010101010",
  11025=>"110100010",
  11026=>"101110011",
  11027=>"101100000",
  11028=>"100000110",
  11029=>"100011100",
  11030=>"100100001",
  11031=>"111000100",
  11032=>"010110010",
  11033=>"000100111",
  11034=>"001000111",
  11035=>"100110011",
  11036=>"010011101",
  11037=>"111000001",
  11038=>"101111110",
  11039=>"110001000",
  11040=>"010010010",
  11041=>"101011001",
  11042=>"110000010",
  11043=>"001011010",
  11044=>"010100000",
  11045=>"011110111",
  11046=>"100000100",
  11047=>"011101001",
  11048=>"110011111",
  11049=>"010111011",
  11050=>"100111010",
  11051=>"110111110",
  11052=>"101000001",
  11053=>"000111101",
  11054=>"111110010",
  11055=>"101000101",
  11056=>"010010110",
  11057=>"111111101",
  11058=>"001011000",
  11059=>"000000000",
  11060=>"001100111",
  11061=>"001010010",
  11062=>"000010111",
  11063=>"001010010",
  11064=>"101110110",
  11065=>"101100111",
  11066=>"010011001",
  11067=>"001001110",
  11068=>"010000000",
  11069=>"000000110",
  11070=>"110011101",
  11071=>"000100111",
  11072=>"111101100",
  11073=>"100011111",
  11074=>"011000110",
  11075=>"110110000",
  11076=>"011011011",
  11077=>"000000010",
  11078=>"001101110",
  11079=>"100011011",
  11080=>"101111010",
  11081=>"001000001",
  11082=>"111011000",
  11083=>"001101010",
  11084=>"010010000",
  11085=>"000100000",
  11086=>"000110010",
  11087=>"100001011",
  11088=>"010101100",
  11089=>"110000101",
  11090=>"001001000",
  11091=>"011001011",
  11092=>"010011110",
  11093=>"000101110",
  11094=>"000010001",
  11095=>"110111100",
  11096=>"111101011",
  11097=>"111000110",
  11098=>"110011101",
  11099=>"111101101",
  11100=>"011110011",
  11101=>"110110111",
  11102=>"111001010",
  11103=>"010011011",
  11104=>"100001111",
  11105=>"010011110",
  11106=>"101011000",
  11107=>"000110101",
  11108=>"111000111",
  11109=>"001000111",
  11110=>"011110100",
  11111=>"000100110",
  11112=>"001110101",
  11113=>"111101110",
  11114=>"110111010",
  11115=>"011111101",
  11116=>"011011101",
  11117=>"011010100",
  11118=>"101110001",
  11119=>"000100111",
  11120=>"100000111",
  11121=>"010001010",
  11122=>"101111100",
  11123=>"001110000",
  11124=>"010011001",
  11125=>"000011000",
  11126=>"101001101",
  11127=>"011011001",
  11128=>"111010000",
  11129=>"001001000",
  11130=>"100001011",
  11131=>"000101111",
  11132=>"101101001",
  11133=>"001000100",
  11134=>"000100000",
  11135=>"100100110",
  11136=>"101110111",
  11137=>"101001000",
  11138=>"100011110",
  11139=>"011100001",
  11140=>"110011110",
  11141=>"001100010",
  11142=>"000000011",
  11143=>"001010111",
  11144=>"001110010",
  11145=>"001100011",
  11146=>"001111110",
  11147=>"101100100",
  11148=>"100000111",
  11149=>"111000111",
  11150=>"000000000",
  11151=>"010110111",
  11152=>"011011001",
  11153=>"010101001",
  11154=>"110111001",
  11155=>"111010100",
  11156=>"001100000",
  11157=>"101110111",
  11158=>"111101011",
  11159=>"000111000",
  11160=>"010111111",
  11161=>"100110000",
  11162=>"100000100",
  11163=>"101111010",
  11164=>"111011100",
  11165=>"000101100",
  11166=>"000110010",
  11167=>"101001011",
  11168=>"101111001",
  11169=>"110100011",
  11170=>"000111011",
  11171=>"010101100",
  11172=>"010110100",
  11173=>"010100100",
  11174=>"010000110",
  11175=>"110011010",
  11176=>"011010001",
  11177=>"101010000",
  11178=>"000000001",
  11179=>"111100111",
  11180=>"000111101",
  11181=>"101010110",
  11182=>"111111011",
  11183=>"000000100",
  11184=>"110011000",
  11185=>"000111010",
  11186=>"011000110",
  11187=>"011011111",
  11188=>"000110101",
  11189=>"100010001",
  11190=>"010110101",
  11191=>"111000001",
  11192=>"011010110",
  11193=>"111011111",
  11194=>"011101100",
  11195=>"110101101",
  11196=>"100000110",
  11197=>"001000000",
  11198=>"100100010",
  11199=>"000000100",
  11200=>"010000111",
  11201=>"100000100",
  11202=>"000101011",
  11203=>"110010010",
  11204=>"101100111",
  11205=>"101011000",
  11206=>"111001010",
  11207=>"100011100",
  11208=>"111000100",
  11209=>"110101111",
  11210=>"000100100",
  11211=>"000011110",
  11212=>"011110100",
  11213=>"100111101",
  11214=>"110101011",
  11215=>"011111011",
  11216=>"000100010",
  11217=>"100100111",
  11218=>"101100011",
  11219=>"100111011",
  11220=>"111101101",
  11221=>"001111000",
  11222=>"010000011",
  11223=>"100110101",
  11224=>"000000100",
  11225=>"100001000",
  11226=>"110010111",
  11227=>"000010001",
  11228=>"001010101",
  11229=>"110000010",
  11230=>"010001000",
  11231=>"000010000",
  11232=>"001100001",
  11233=>"101111111",
  11234=>"000111111",
  11235=>"011100000",
  11236=>"000000110",
  11237=>"000110101",
  11238=>"000010101",
  11239=>"011000000",
  11240=>"101101100",
  11241=>"101110010",
  11242=>"100010010",
  11243=>"001000100",
  11244=>"001101110",
  11245=>"001000010",
  11246=>"110010001",
  11247=>"101111000",
  11248=>"001100000",
  11249=>"010011001",
  11250=>"101011110",
  11251=>"101001101",
  11252=>"010110111",
  11253=>"011000100",
  11254=>"111011111",
  11255=>"100101100",
  11256=>"110100101",
  11257=>"111011111",
  11258=>"110011101",
  11259=>"001101011",
  11260=>"000100100",
  11261=>"000000101",
  11262=>"010000100",
  11263=>"011110011",
  11264=>"000011010",
  11265=>"100010011",
  11266=>"100110000",
  11267=>"110011110",
  11268=>"101111000",
  11269=>"110111101",
  11270=>"110101000",
  11271=>"010110010",
  11272=>"010000000",
  11273=>"001010111",
  11274=>"011101110",
  11275=>"010000111",
  11276=>"011011111",
  11277=>"010111100",
  11278=>"001001111",
  11279=>"111011111",
  11280=>"011100101",
  11281=>"001110010",
  11282=>"111000101",
  11283=>"011101111",
  11284=>"110010101",
  11285=>"100001101",
  11286=>"000110100",
  11287=>"011111101",
  11288=>"110111100",
  11289=>"101111101",
  11290=>"001010110",
  11291=>"100000101",
  11292=>"110110010",
  11293=>"101110111",
  11294=>"110111110",
  11295=>"110111011",
  11296=>"100100000",
  11297=>"001011000",
  11298=>"000001000",
  11299=>"000100000",
  11300=>"100110101",
  11301=>"101100110",
  11302=>"111000010",
  11303=>"000001000",
  11304=>"011001100",
  11305=>"101011111",
  11306=>"001111010",
  11307=>"100101110",
  11308=>"110110100",
  11309=>"000001001",
  11310=>"101011010",
  11311=>"101011110",
  11312=>"111101111",
  11313=>"010111110",
  11314=>"011011010",
  11315=>"110001001",
  11316=>"010110011",
  11317=>"000101010",
  11318=>"110000100",
  11319=>"101100001",
  11320=>"000111011",
  11321=>"011110111",
  11322=>"011111111",
  11323=>"101111011",
  11324=>"101111010",
  11325=>"110111000",
  11326=>"110010000",
  11327=>"011100111",
  11328=>"000010110",
  11329=>"111111110",
  11330=>"110001001",
  11331=>"011100011",
  11332=>"000000110",
  11333=>"000010100",
  11334=>"100001000",
  11335=>"000011111",
  11336=>"010001010",
  11337=>"001101110",
  11338=>"110111100",
  11339=>"111111111",
  11340=>"000111011",
  11341=>"000001101",
  11342=>"001000000",
  11343=>"000101101",
  11344=>"001010100",
  11345=>"101110001",
  11346=>"110001111",
  11347=>"001000001",
  11348=>"010000010",
  11349=>"101001111",
  11350=>"011010110",
  11351=>"011011110",
  11352=>"100000010",
  11353=>"111110010",
  11354=>"111111001",
  11355=>"100111010",
  11356=>"011111011",
  11357=>"111110110",
  11358=>"010111010",
  11359=>"111101111",
  11360=>"010110000",
  11361=>"011111111",
  11362=>"010100100",
  11363=>"111111110",
  11364=>"100111011",
  11365=>"100010101",
  11366=>"100011011",
  11367=>"111111111",
  11368=>"111011100",
  11369=>"111101011",
  11370=>"010001000",
  11371=>"000011001",
  11372=>"111111111",
  11373=>"100100000",
  11374=>"011001010",
  11375=>"011111111",
  11376=>"100110010",
  11377=>"111111001",
  11378=>"111010011",
  11379=>"111010101",
  11380=>"010100110",
  11381=>"001000011",
  11382=>"011000011",
  11383=>"001110001",
  11384=>"111001111",
  11385=>"110101010",
  11386=>"000011111",
  11387=>"000011110",
  11388=>"001001110",
  11389=>"011000000",
  11390=>"111110111",
  11391=>"001010010",
  11392=>"001111110",
  11393=>"101100101",
  11394=>"101110111",
  11395=>"111110100",
  11396=>"000010011",
  11397=>"100101010",
  11398=>"001011000",
  11399=>"100111000",
  11400=>"110111111",
  11401=>"101111100",
  11402=>"111001111",
  11403=>"001111110",
  11404=>"101010100",
  11405=>"111100100",
  11406=>"110000010",
  11407=>"110101111",
  11408=>"101000101",
  11409=>"110010010",
  11410=>"011010111",
  11411=>"100100101",
  11412=>"011101010",
  11413=>"011001011",
  11414=>"110001110",
  11415=>"000011100",
  11416=>"111110110",
  11417=>"011000111",
  11418=>"000010111",
  11419=>"010001110",
  11420=>"111011001",
  11421=>"111101001",
  11422=>"011011001",
  11423=>"110001010",
  11424=>"111100000",
  11425=>"111000100",
  11426=>"000000011",
  11427=>"011111001",
  11428=>"100010110",
  11429=>"111110100",
  11430=>"010001101",
  11431=>"011011000",
  11432=>"000111100",
  11433=>"101111101",
  11434=>"111001001",
  11435=>"000000010",
  11436=>"100010110",
  11437=>"011011001",
  11438=>"011001101",
  11439=>"111000001",
  11440=>"111011100",
  11441=>"111101111",
  11442=>"011001110",
  11443=>"111111110",
  11444=>"110101101",
  11445=>"100101100",
  11446=>"101101110",
  11447=>"000111111",
  11448=>"101111111",
  11449=>"011010111",
  11450=>"110010010",
  11451=>"101100010",
  11452=>"000001010",
  11453=>"010111010",
  11454=>"010011011",
  11455=>"001000101",
  11456=>"100000001",
  11457=>"001001111",
  11458=>"110010111",
  11459=>"111011111",
  11460=>"101101110",
  11461=>"011110010",
  11462=>"101011000",
  11463=>"111010000",
  11464=>"011000000",
  11465=>"000110100",
  11466=>"000001001",
  11467=>"010110111",
  11468=>"110101000",
  11469=>"111101011",
  11470=>"000010010",
  11471=>"001111011",
  11472=>"111011111",
  11473=>"110100010",
  11474=>"101100110",
  11475=>"111011011",
  11476=>"110001110",
  11477=>"101010011",
  11478=>"000000100",
  11479=>"111000001",
  11480=>"001011101",
  11481=>"001101111",
  11482=>"110110000",
  11483=>"100100000",
  11484=>"110010110",
  11485=>"101010100",
  11486=>"100000000",
  11487=>"111111110",
  11488=>"101011000",
  11489=>"100111101",
  11490=>"110101000",
  11491=>"111011001",
  11492=>"000111110",
  11493=>"111111111",
  11494=>"100010011",
  11495=>"010111000",
  11496=>"100011010",
  11497=>"100111001",
  11498=>"001110001",
  11499=>"101001010",
  11500=>"100001001",
  11501=>"101111100",
  11502=>"111101111",
  11503=>"111111111",
  11504=>"011110101",
  11505=>"100001111",
  11506=>"111111111",
  11507=>"101000100",
  11508=>"010010010",
  11509=>"100011001",
  11510=>"100100100",
  11511=>"111111111",
  11512=>"000111001",
  11513=>"111010100",
  11514=>"011011101",
  11515=>"011111011",
  11516=>"011111100",
  11517=>"111011101",
  11518=>"101000100",
  11519=>"111010101",
  11520=>"001000000",
  11521=>"100010101",
  11522=>"100111011",
  11523=>"111111100",
  11524=>"001001110",
  11525=>"110100100",
  11526=>"111111111",
  11527=>"000000101",
  11528=>"101100011",
  11529=>"111100111",
  11530=>"111111100",
  11531=>"101111011",
  11532=>"011110111",
  11533=>"101111111",
  11534=>"001001100",
  11535=>"111011011",
  11536=>"000000101",
  11537=>"010010100",
  11538=>"001011111",
  11539=>"010101101",
  11540=>"101011101",
  11541=>"101011011",
  11542=>"110011111",
  11543=>"110000111",
  11544=>"000000001",
  11545=>"011000111",
  11546=>"010001010",
  11547=>"000000101",
  11548=>"010011010",
  11549=>"001010011",
  11550=>"000110001",
  11551=>"111000110",
  11552=>"111110101",
  11553=>"110010110",
  11554=>"111010011",
  11555=>"110111111",
  11556=>"101100000",
  11557=>"000100000",
  11558=>"000001111",
  11559=>"001000010",
  11560=>"101110001",
  11561=>"000111000",
  11562=>"111100000",
  11563=>"110000110",
  11564=>"100001101",
  11565=>"001111011",
  11566=>"011111011",
  11567=>"100101011",
  11568=>"110111101",
  11569=>"000000000",
  11570=>"011100000",
  11571=>"111110111",
  11572=>"111101011",
  11573=>"010011010",
  11574=>"110011000",
  11575=>"001111000",
  11576=>"111110110",
  11577=>"011001100",
  11578=>"111001101",
  11579=>"110101111",
  11580=>"111101110",
  11581=>"011101000",
  11582=>"000110111",
  11583=>"110000010",
  11584=>"111010010",
  11585=>"111111011",
  11586=>"010011010",
  11587=>"010011010",
  11588=>"001111011",
  11589=>"100001000",
  11590=>"111101111",
  11591=>"011110111",
  11592=>"010100001",
  11593=>"111011110",
  11594=>"101001010",
  11595=>"100111101",
  11596=>"100011000",
  11597=>"110110000",
  11598=>"010110000",
  11599=>"011011001",
  11600=>"011011000",
  11601=>"111001011",
  11602=>"100010110",
  11603=>"111111110",
  11604=>"111111111",
  11605=>"010111110",
  11606=>"111000000",
  11607=>"011011111",
  11608=>"000110011",
  11609=>"111110111",
  11610=>"011110111",
  11611=>"000111111",
  11612=>"000101010",
  11613=>"001101111",
  11614=>"111110011",
  11615=>"111111111",
  11616=>"111010110",
  11617=>"000111110",
  11618=>"101110111",
  11619=>"100110101",
  11620=>"100011110",
  11621=>"101000100",
  11622=>"001110111",
  11623=>"010100000",
  11624=>"110011000",
  11625=>"010100110",
  11626=>"111101101",
  11627=>"111011000",
  11628=>"011011001",
  11629=>"000100110",
  11630=>"110101100",
  11631=>"011101110",
  11632=>"011111111",
  11633=>"011100010",
  11634=>"111111111",
  11635=>"000100001",
  11636=>"001000111",
  11637=>"111010110",
  11638=>"010011110",
  11639=>"011100100",
  11640=>"011110011",
  11641=>"011100100",
  11642=>"101101001",
  11643=>"010110100",
  11644=>"010111101",
  11645=>"110000101",
  11646=>"000110100",
  11647=>"100100101",
  11648=>"101101111",
  11649=>"001110101",
  11650=>"000001000",
  11651=>"100000111",
  11652=>"011001000",
  11653=>"101111010",
  11654=>"011101100",
  11655=>"001111011",
  11656=>"111010110",
  11657=>"011110101",
  11658=>"100110100",
  11659=>"000001100",
  11660=>"101110101",
  11661=>"000110101",
  11662=>"000100001",
  11663=>"000100111",
  11664=>"110000100",
  11665=>"111000010",
  11666=>"111000001",
  11667=>"011100011",
  11668=>"111111111",
  11669=>"101110011",
  11670=>"011000111",
  11671=>"000000001",
  11672=>"001001000",
  11673=>"111111100",
  11674=>"011011010",
  11675=>"010110100",
  11676=>"000000100",
  11677=>"111111111",
  11678=>"011000010",
  11679=>"110101101",
  11680=>"001001001",
  11681=>"111011111",
  11682=>"000010110",
  11683=>"111111101",
  11684=>"001100001",
  11685=>"101111001",
  11686=>"000111110",
  11687=>"100001001",
  11688=>"110000110",
  11689=>"101001001",
  11690=>"110000111",
  11691=>"010011111",
  11692=>"111010111",
  11693=>"100101101",
  11694=>"011110011",
  11695=>"110010010",
  11696=>"010001011",
  11697=>"110111011",
  11698=>"001101100",
  11699=>"011110100",
  11700=>"010010010",
  11701=>"111000110",
  11702=>"110101110",
  11703=>"111111000",
  11704=>"001000000",
  11705=>"111010111",
  11706=>"111110001",
  11707=>"110111011",
  11708=>"000000010",
  11709=>"000010000",
  11710=>"111110111",
  11711=>"001000111",
  11712=>"010001110",
  11713=>"111110110",
  11714=>"001011001",
  11715=>"010100100",
  11716=>"101001100",
  11717=>"010001100",
  11718=>"011011111",
  11719=>"000001001",
  11720=>"111000000",
  11721=>"111001001",
  11722=>"010111010",
  11723=>"010110110",
  11724=>"111001111",
  11725=>"000111010",
  11726=>"101011001",
  11727=>"001101111",
  11728=>"010000001",
  11729=>"000100111",
  11730=>"011110100",
  11731=>"001001110",
  11732=>"100111011",
  11733=>"101001110",
  11734=>"000011000",
  11735=>"100101010",
  11736=>"111010011",
  11737=>"111110001",
  11738=>"111101100",
  11739=>"001001110",
  11740=>"100001111",
  11741=>"000111111",
  11742=>"110111001",
  11743=>"110111111",
  11744=>"111101111",
  11745=>"010011000",
  11746=>"010011111",
  11747=>"111000010",
  11748=>"110111111",
  11749=>"000110111",
  11750=>"010111001",
  11751=>"001100110",
  11752=>"111101100",
  11753=>"011100000",
  11754=>"111111110",
  11755=>"001010100",
  11756=>"001101001",
  11757=>"001000000",
  11758=>"110011010",
  11759=>"101110101",
  11760=>"001111110",
  11761=>"010100101",
  11762=>"110101100",
  11763=>"000111011",
  11764=>"100000000",
  11765=>"001011001",
  11766=>"010011100",
  11767=>"101000001",
  11768=>"110101110",
  11769=>"101100111",
  11770=>"111101111",
  11771=>"100111110",
  11772=>"101111010",
  11773=>"001000111",
  11774=>"100110000",
  11775=>"000101101",
  11776=>"001011110",
  11777=>"011000101",
  11778=>"110111011",
  11779=>"001011111",
  11780=>"111100001",
  11781=>"000011111",
  11782=>"000001110",
  11783=>"110001111",
  11784=>"011011110",
  11785=>"011001001",
  11786=>"000111101",
  11787=>"100111111",
  11788=>"001111001",
  11789=>"000111000",
  11790=>"001001111",
  11791=>"101010100",
  11792=>"010001011",
  11793=>"100000101",
  11794=>"100010001",
  11795=>"101101001",
  11796=>"011001010",
  11797=>"110010010",
  11798=>"100010011",
  11799=>"111100001",
  11800=>"010001110",
  11801=>"100110111",
  11802=>"001110111",
  11803=>"110111111",
  11804=>"100111010",
  11805=>"010010111",
  11806=>"000001011",
  11807=>"100000100",
  11808=>"000011011",
  11809=>"110100100",
  11810=>"111001110",
  11811=>"100011000",
  11812=>"010101001",
  11813=>"101010100",
  11814=>"011110001",
  11815=>"000110011",
  11816=>"111100110",
  11817=>"110000101",
  11818=>"101110011",
  11819=>"010111100",
  11820=>"110110000",
  11821=>"011111101",
  11822=>"101000100",
  11823=>"101010111",
  11824=>"100111100",
  11825=>"010001000",
  11826=>"011001000",
  11827=>"111000111",
  11828=>"111111111",
  11829=>"101100101",
  11830=>"111001101",
  11831=>"101110101",
  11832=>"100000110",
  11833=>"001100000",
  11834=>"011111111",
  11835=>"110111111",
  11836=>"110010111",
  11837=>"011111111",
  11838=>"010111000",
  11839=>"010101000",
  11840=>"111011111",
  11841=>"100000101",
  11842=>"001110011",
  11843=>"110001100",
  11844=>"000110001",
  11845=>"011011101",
  11846=>"011100111",
  11847=>"100110000",
  11848=>"011110010",
  11849=>"100100000",
  11850=>"001010010",
  11851=>"111111111",
  11852=>"010010101",
  11853=>"101011001",
  11854=>"001100001",
  11855=>"000100110",
  11856=>"111000101",
  11857=>"111110000",
  11858=>"111110111",
  11859=>"111110111",
  11860=>"110111011",
  11861=>"100111111",
  11862=>"000111101",
  11863=>"001011111",
  11864=>"100011011",
  11865=>"010011011",
  11866=>"011110111",
  11867=>"110111011",
  11868=>"000110010",
  11869=>"101000111",
  11870=>"111110101",
  11871=>"101000001",
  11872=>"011111101",
  11873=>"011111101",
  11874=>"110001010",
  11875=>"111100000",
  11876=>"010011111",
  11877=>"111001011",
  11878=>"101011100",
  11879=>"111111010",
  11880=>"110101101",
  11881=>"000010111",
  11882=>"111000111",
  11883=>"011011111",
  11884=>"011100101",
  11885=>"000011101",
  11886=>"111010000",
  11887=>"111011111",
  11888=>"111010000",
  11889=>"010001111",
  11890=>"010000011",
  11891=>"000111101",
  11892=>"111011000",
  11893=>"010110110",
  11894=>"011011111",
  11895=>"100111011",
  11896=>"111111110",
  11897=>"001001011",
  11898=>"100001110",
  11899=>"011001001",
  11900=>"100111011",
  11901=>"101011111",
  11902=>"101100011",
  11903=>"100010101",
  11904=>"001110011",
  11905=>"000011110",
  11906=>"000000110",
  11907=>"100111110",
  11908=>"100100110",
  11909=>"111110111",
  11910=>"001011100",
  11911=>"101001010",
  11912=>"100010000",
  11913=>"000000011",
  11914=>"001000000",
  11915=>"111010110",
  11916=>"111011110",
  11917=>"011101111",
  11918=>"010001111",
  11919=>"100101001",
  11920=>"010010110",
  11921=>"001001001",
  11922=>"011100100",
  11923=>"111010110",
  11924=>"111110001",
  11925=>"001010100",
  11926=>"001010000",
  11927=>"011000000",
  11928=>"011100111",
  11929=>"110010110",
  11930=>"000111100",
  11931=>"101010010",
  11932=>"001011111",
  11933=>"100100100",
  11934=>"111111101",
  11935=>"000110111",
  11936=>"011110110",
  11937=>"101001110",
  11938=>"100010000",
  11939=>"111111100",
  11940=>"111101001",
  11941=>"111000010",
  11942=>"011010000",
  11943=>"111111100",
  11944=>"111110111",
  11945=>"100100111",
  11946=>"001000001",
  11947=>"110110111",
  11948=>"110110111",
  11949=>"100011100",
  11950=>"000010111",
  11951=>"100110101",
  11952=>"011010111",
  11953=>"101000111",
  11954=>"100000110",
  11955=>"000010001",
  11956=>"101001001",
  11957=>"010100000",
  11958=>"110101010",
  11959=>"011001101",
  11960=>"111110110",
  11961=>"011101000",
  11962=>"101110010",
  11963=>"111100111",
  11964=>"101101101",
  11965=>"010011011",
  11966=>"101011011",
  11967=>"000111011",
  11968=>"000010101",
  11969=>"100110110",
  11970=>"011100111",
  11971=>"011011111",
  11972=>"111011001",
  11973=>"111111111",
  11974=>"100100010",
  11975=>"001111101",
  11976=>"000000010",
  11977=>"101100101",
  11978=>"101101001",
  11979=>"111111110",
  11980=>"011000011",
  11981=>"001101000",
  11982=>"011010101",
  11983=>"000011111",
  11984=>"011110111",
  11985=>"001111110",
  11986=>"110111111",
  11987=>"111110110",
  11988=>"100110011",
  11989=>"110101110",
  11990=>"111000100",
  11991=>"011001110",
  11992=>"111000011",
  11993=>"110100110",
  11994=>"111011000",
  11995=>"001001111",
  11996=>"111111010",
  11997=>"000110011",
  11998=>"110100111",
  11999=>"011000010",
  12000=>"100011111",
  12001=>"010010010",
  12002=>"100101010",
  12003=>"000110010",
  12004=>"111111000",
  12005=>"000100011",
  12006=>"101110111",
  12007=>"010010111",
  12008=>"001100001",
  12009=>"100100000",
  12010=>"011100001",
  12011=>"001011011",
  12012=>"111110110",
  12013=>"010010010",
  12014=>"010010110",
  12015=>"101101000",
  12016=>"011010100",
  12017=>"101010110",
  12018=>"010110101",
  12019=>"000100100",
  12020=>"000100000",
  12021=>"101100000",
  12022=>"000010110",
  12023=>"000010110",
  12024=>"010011010",
  12025=>"111001111",
  12026=>"001010100",
  12027=>"111011100",
  12028=>"100000100",
  12029=>"000001111",
  12030=>"011110010",
  12031=>"101101000",
  12032=>"011111010",
  12033=>"110001011",
  12034=>"010000111",
  12035=>"111111000",
  12036=>"001101101",
  12037=>"100011111",
  12038=>"111100010",
  12039=>"001011000",
  12040=>"101111101",
  12041=>"111101111",
  12042=>"101000101",
  12043=>"110011110",
  12044=>"000011100",
  12045=>"010110100",
  12046=>"100010111",
  12047=>"100111000",
  12048=>"111001001",
  12049=>"111111111",
  12050=>"001000110",
  12051=>"000101100",
  12052=>"000111110",
  12053=>"101010100",
  12054=>"010000010",
  12055=>"100111011",
  12056=>"011011010",
  12057=>"011111111",
  12058=>"110111111",
  12059=>"010000101",
  12060=>"110110011",
  12061=>"010000010",
  12062=>"010001111",
  12063=>"001000110",
  12064=>"011100000",
  12065=>"110010000",
  12066=>"001010000",
  12067=>"001100011",
  12068=>"101011110",
  12069=>"011101111",
  12070=>"001100100",
  12071=>"111011111",
  12072=>"111010100",
  12073=>"000010000",
  12074=>"110111000",
  12075=>"110001011",
  12076=>"111100111",
  12077=>"110111111",
  12078=>"011001111",
  12079=>"111101101",
  12080=>"111011111",
  12081=>"011110110",
  12082=>"111111011",
  12083=>"001010111",
  12084=>"000000110",
  12085=>"011010100",
  12086=>"111011000",
  12087=>"110001001",
  12088=>"000010011",
  12089=>"000000011",
  12090=>"111011110",
  12091=>"001000011",
  12092=>"111111011",
  12093=>"011111111",
  12094=>"000011110",
  12095=>"000101110",
  12096=>"111010001",
  12097=>"100001000",
  12098=>"000000100",
  12099=>"010001111",
  12100=>"011011111",
  12101=>"000101110",
  12102=>"000101101",
  12103=>"101011010",
  12104=>"101111000",
  12105=>"101111000",
  12106=>"100011111",
  12107=>"101111010",
  12108=>"010000001",
  12109=>"011011111",
  12110=>"010001111",
  12111=>"000001110",
  12112=>"001101111",
  12113=>"111001011",
  12114=>"100111111",
  12115=>"001100111",
  12116=>"000001010",
  12117=>"001111001",
  12118=>"111101010",
  12119=>"111011111",
  12120=>"110110010",
  12121=>"110110000",
  12122=>"110001111",
  12123=>"100101111",
  12124=>"000010000",
  12125=>"101000001",
  12126=>"000100001",
  12127=>"110111111",
  12128=>"100000011",
  12129=>"001010011",
  12130=>"111010111",
  12131=>"001000010",
  12132=>"101011111",
  12133=>"011100110",
  12134=>"001001000",
  12135=>"110000101",
  12136=>"010000101",
  12137=>"011011100",
  12138=>"100111111",
  12139=>"110100111",
  12140=>"000100011",
  12141=>"011001001",
  12142=>"000101010",
  12143=>"011010010",
  12144=>"101101100",
  12145=>"010011011",
  12146=>"000010010",
  12147=>"111001101",
  12148=>"011001111",
  12149=>"111011110",
  12150=>"111000000",
  12151=>"111010100",
  12152=>"111101000",
  12153=>"110110111",
  12154=>"111100000",
  12155=>"000110110",
  12156=>"011111111",
  12157=>"011110101",
  12158=>"001011011",
  12159=>"000100001",
  12160=>"001100000",
  12161=>"101010000",
  12162=>"001101000",
  12163=>"110110001",
  12164=>"111101100",
  12165=>"100001000",
  12166=>"111001111",
  12167=>"101010010",
  12168=>"000111000",
  12169=>"101001001",
  12170=>"111111100",
  12171=>"001001011",
  12172=>"101010010",
  12173=>"001000100",
  12174=>"000101010",
  12175=>"010010000",
  12176=>"001000011",
  12177=>"010101101",
  12178=>"001101111",
  12179=>"011110011",
  12180=>"011000111",
  12181=>"001100100",
  12182=>"001111101",
  12183=>"001011011",
  12184=>"111101100",
  12185=>"000100111",
  12186=>"001110111",
  12187=>"111110100",
  12188=>"111101000",
  12189=>"001101111",
  12190=>"110001010",
  12191=>"010100010",
  12192=>"011101001",
  12193=>"011000000",
  12194=>"110110111",
  12195=>"000111010",
  12196=>"101000011",
  12197=>"101000110",
  12198=>"000110111",
  12199=>"000110001",
  12200=>"000000111",
  12201=>"010111100",
  12202=>"011101011",
  12203=>"111100111",
  12204=>"111011110",
  12205=>"000000000",
  12206=>"010100111",
  12207=>"000001101",
  12208=>"100111101",
  12209=>"111010010",
  12210=>"010000000",
  12211=>"011110001",
  12212=>"010000011",
  12213=>"010001001",
  12214=>"110010101",
  12215=>"010111100",
  12216=>"101100111",
  12217=>"011010111",
  12218=>"100001110",
  12219=>"010111011",
  12220=>"010000011",
  12221=>"001100101",
  12222=>"000111001",
  12223=>"111111101",
  12224=>"011111110",
  12225=>"110100000",
  12226=>"110111011",
  12227=>"001011111",
  12228=>"111001011",
  12229=>"100000010",
  12230=>"101000000",
  12231=>"101000101",
  12232=>"111111101",
  12233=>"111001001",
  12234=>"100001111",
  12235=>"011110010",
  12236=>"000010110",
  12237=>"001001111",
  12238=>"001110000",
  12239=>"001111000",
  12240=>"111100111",
  12241=>"001110101",
  12242=>"101101111",
  12243=>"110101111",
  12244=>"111111010",
  12245=>"111010100",
  12246=>"101111110",
  12247=>"101100111",
  12248=>"110111111",
  12249=>"010101110",
  12250=>"101110011",
  12251=>"100111100",
  12252=>"001010100",
  12253=>"010101101",
  12254=>"111100001",
  12255=>"111100110",
  12256=>"001111100",
  12257=>"111110100",
  12258=>"100000001",
  12259=>"110100110",
  12260=>"110011111",
  12261=>"111010110",
  12262=>"110110110",
  12263=>"110010000",
  12264=>"011100110",
  12265=>"110111000",
  12266=>"010110111",
  12267=>"110001111",
  12268=>"110110001",
  12269=>"111010011",
  12270=>"001010001",
  12271=>"110110001",
  12272=>"000101100",
  12273=>"101111011",
  12274=>"101111111",
  12275=>"100001000",
  12276=>"101000011",
  12277=>"101111110",
  12278=>"000010111",
  12279=>"111001101",
  12280=>"111011100",
  12281=>"111000001",
  12282=>"111101000",
  12283=>"100000011",
  12284=>"110101111",
  12285=>"110100110",
  12286=>"010000101",
  12287=>"010011011",
  12288=>"000001010",
  12289=>"001110111",
  12290=>"010100001",
  12291=>"110111011",
  12292=>"111101110",
  12293=>"010011010",
  12294=>"100011111",
  12295=>"110010010",
  12296=>"100010010",
  12297=>"000010100",
  12298=>"101011000",
  12299=>"100101000",
  12300=>"110011001",
  12301=>"100010110",
  12302=>"100101011",
  12303=>"100011011",
  12304=>"000000001",
  12305=>"101110000",
  12306=>"010000001",
  12307=>"011100100",
  12308=>"000100000",
  12309=>"111110101",
  12310=>"001111110",
  12311=>"100101000",
  12312=>"110111101",
  12313=>"101000001",
  12314=>"010001100",
  12315=>"110100101",
  12316=>"110110011",
  12317=>"001001010",
  12318=>"000011101",
  12319=>"000111000",
  12320=>"011010111",
  12321=>"101100011",
  12322=>"111110110",
  12323=>"010011001",
  12324=>"111001000",
  12325=>"011101110",
  12326=>"111100010",
  12327=>"000100000",
  12328=>"011010010",
  12329=>"000001000",
  12330=>"010000101",
  12331=>"110011111",
  12332=>"100011000",
  12333=>"001011001",
  12334=>"111000100",
  12335=>"000000101",
  12336=>"100111101",
  12337=>"001001001",
  12338=>"100111111",
  12339=>"010001001",
  12340=>"011100000",
  12341=>"011001111",
  12342=>"010010010",
  12343=>"111001111",
  12344=>"001000100",
  12345=>"100001001",
  12346=>"110000110",
  12347=>"011010110",
  12348=>"001011110",
  12349=>"000000001",
  12350=>"010110101",
  12351=>"100101101",
  12352=>"101111011",
  12353=>"110101011",
  12354=>"010000000",
  12355=>"011101000",
  12356=>"111111111",
  12357=>"011000001",
  12358=>"011010110",
  12359=>"001111000",
  12360=>"001110111",
  12361=>"011000000",
  12362=>"100111000",
  12363=>"101100101",
  12364=>"011100011",
  12365=>"110010101",
  12366=>"010111001",
  12367=>"101101011",
  12368=>"000110110",
  12369=>"001100000",
  12370=>"110101011",
  12371=>"000100000",
  12372=>"010110111",
  12373=>"001000111",
  12374=>"001101010",
  12375=>"010101111",
  12376=>"001111111",
  12377=>"011111111",
  12378=>"001111111",
  12379=>"101010011",
  12380=>"101110110",
  12381=>"111011001",
  12382=>"110111001",
  12383=>"100101010",
  12384=>"100110101",
  12385=>"100000101",
  12386=>"011000010",
  12387=>"001010010",
  12388=>"110100111",
  12389=>"101000001",
  12390=>"010011000",
  12391=>"010010111",
  12392=>"010000001",
  12393=>"000010100",
  12394=>"011101110",
  12395=>"111011001",
  12396=>"010000100",
  12397=>"111011111",
  12398=>"111000000",
  12399=>"101110100",
  12400=>"011111000",
  12401=>"101000001",
  12402=>"111000110",
  12403=>"010110001",
  12404=>"000001011",
  12405=>"100001000",
  12406=>"010001111",
  12407=>"101100010",
  12408=>"100101011",
  12409=>"011001111",
  12410=>"000001010",
  12411=>"101110010",
  12412=>"101001011",
  12413=>"100101001",
  12414=>"101011101",
  12415=>"000101010",
  12416=>"001110010",
  12417=>"111111110",
  12418=>"010110101",
  12419=>"111111011",
  12420=>"010111001",
  12421=>"100011110",
  12422=>"111000111",
  12423=>"010111110",
  12424=>"010110111",
  12425=>"011100010",
  12426=>"111110000",
  12427=>"010000111",
  12428=>"111100011",
  12429=>"100101111",
  12430=>"000101110",
  12431=>"100101001",
  12432=>"111000110",
  12433=>"110010001",
  12434=>"010010101",
  12435=>"111000000",
  12436=>"110101000",
  12437=>"011101110",
  12438=>"111000010",
  12439=>"111110000",
  12440=>"001111011",
  12441=>"010001011",
  12442=>"011100101",
  12443=>"010111011",
  12444=>"001101011",
  12445=>"100110000",
  12446=>"100111100",
  12447=>"110010000",
  12448=>"111011011",
  12449=>"010000100",
  12450=>"100111101",
  12451=>"000011010",
  12452=>"011111100",
  12453=>"010100100",
  12454=>"101001011",
  12455=>"000000011",
  12456=>"101111100",
  12457=>"010111011",
  12458=>"001001111",
  12459=>"110001010",
  12460=>"110100001",
  12461=>"101110010",
  12462=>"101111111",
  12463=>"101110011",
  12464=>"101111010",
  12465=>"000100110",
  12466=>"010000100",
  12467=>"001101011",
  12468=>"000100001",
  12469=>"100111111",
  12470=>"111110110",
  12471=>"100100001",
  12472=>"111000111",
  12473=>"011000000",
  12474=>"000110101",
  12475=>"101011001",
  12476=>"111010001",
  12477=>"100110001",
  12478=>"000100110",
  12479=>"000010100",
  12480=>"000011010",
  12481=>"111110100",
  12482=>"000000010",
  12483=>"010110111",
  12484=>"000101010",
  12485=>"011111000",
  12486=>"011100111",
  12487=>"111000110",
  12488=>"001011100",
  12489=>"101110101",
  12490=>"110001001",
  12491=>"011011000",
  12492=>"111011101",
  12493=>"011101101",
  12494=>"101111010",
  12495=>"100010101",
  12496=>"101111000",
  12497=>"000100111",
  12498=>"011011111",
  12499=>"011101110",
  12500=>"011010110",
  12501=>"111111100",
  12502=>"111000001",
  12503=>"011000011",
  12504=>"010011011",
  12505=>"000110111",
  12506=>"010111001",
  12507=>"010000110",
  12508=>"101000011",
  12509=>"111111100",
  12510=>"011001101",
  12511=>"000000010",
  12512=>"010111000",
  12513=>"011000001",
  12514=>"000100111",
  12515=>"010001001",
  12516=>"011110001",
  12517=>"000000101",
  12518=>"101100111",
  12519=>"101010100",
  12520=>"000111100",
  12521=>"101101011",
  12522=>"111000001",
  12523=>"100100010",
  12524=>"100001100",
  12525=>"011000111",
  12526=>"000100100",
  12527=>"000111111",
  12528=>"011110011",
  12529=>"111010010",
  12530=>"111011000",
  12531=>"110001001",
  12532=>"111110000",
  12533=>"000100001",
  12534=>"111001111",
  12535=>"000100011",
  12536=>"101010000",
  12537=>"111100000",
  12538=>"110110011",
  12539=>"000110000",
  12540=>"000001010",
  12541=>"011110010",
  12542=>"111001011",
  12543=>"101110000",
  12544=>"000010110",
  12545=>"011001101",
  12546=>"110011010",
  12547=>"010100111",
  12548=>"100101010",
  12549=>"100110101",
  12550=>"100100110",
  12551=>"001010001",
  12552=>"010010100",
  12553=>"100010001",
  12554=>"000101111",
  12555=>"110001111",
  12556=>"001010101",
  12557=>"010100011",
  12558=>"101011001",
  12559=>"010110100",
  12560=>"010111011",
  12561=>"110100010",
  12562=>"111110110",
  12563=>"010010011",
  12564=>"110011000",
  12565=>"111010101",
  12566=>"010010110",
  12567=>"101110111",
  12568=>"000101000",
  12569=>"101000000",
  12570=>"100110011",
  12571=>"111000111",
  12572=>"001100000",
  12573=>"110000001",
  12574=>"001000001",
  12575=>"010001000",
  12576=>"000101010",
  12577=>"000110000",
  12578=>"110010100",
  12579=>"110100001",
  12580=>"000011100",
  12581=>"111100010",
  12582=>"011100001",
  12583=>"010110001",
  12584=>"110011110",
  12585=>"000011110",
  12586=>"010000001",
  12587=>"101111101",
  12588=>"110101100",
  12589=>"001111011",
  12590=>"001110100",
  12591=>"110111001",
  12592=>"100010110",
  12593=>"110000000",
  12594=>"011001001",
  12595=>"000001111",
  12596=>"110001110",
  12597=>"110010110",
  12598=>"100101000",
  12599=>"111110110",
  12600=>"011000111",
  12601=>"101011011",
  12602=>"010011100",
  12603=>"110010101",
  12604=>"100100000",
  12605=>"110110010",
  12606=>"110000101",
  12607=>"100010010",
  12608=>"110010001",
  12609=>"011000111",
  12610=>"000100000",
  12611=>"011111010",
  12612=>"001011011",
  12613=>"011010110",
  12614=>"010100011",
  12615=>"011001000",
  12616=>"110110100",
  12617=>"111101011",
  12618=>"101101011",
  12619=>"000001101",
  12620=>"011001101",
  12621=>"100001010",
  12622=>"001000110",
  12623=>"010110111",
  12624=>"111001011",
  12625=>"111100101",
  12626=>"101100000",
  12627=>"010101110",
  12628=>"011011011",
  12629=>"001011111",
  12630=>"000000001",
  12631=>"000011010",
  12632=>"101100010",
  12633=>"000000011",
  12634=>"000000111",
  12635=>"001100011",
  12636=>"110111110",
  12637=>"011101110",
  12638=>"111011001",
  12639=>"011100111",
  12640=>"011111011",
  12641=>"010011010",
  12642=>"000001111",
  12643=>"011000111",
  12644=>"001000111",
  12645=>"001101101",
  12646=>"000010111",
  12647=>"010011101",
  12648=>"111101010",
  12649=>"000111000",
  12650=>"101000010",
  12651=>"100110110",
  12652=>"011010110",
  12653=>"000111110",
  12654=>"001101011",
  12655=>"000010000",
  12656=>"011000111",
  12657=>"011010000",
  12658=>"100111010",
  12659=>"010000011",
  12660=>"011110111",
  12661=>"000001100",
  12662=>"100100001",
  12663=>"100000100",
  12664=>"101100011",
  12665=>"001111111",
  12666=>"000111100",
  12667=>"011110011",
  12668=>"100101011",
  12669=>"010110001",
  12670=>"001001101",
  12671=>"000000010",
  12672=>"101000000",
  12673=>"101101110",
  12674=>"000111010",
  12675=>"000010001",
  12676=>"111100011",
  12677=>"001110001",
  12678=>"111001001",
  12679=>"111100001",
  12680=>"101011001",
  12681=>"010100100",
  12682=>"010110100",
  12683=>"101101011",
  12684=>"010100001",
  12685=>"010010101",
  12686=>"011100000",
  12687=>"010111110",
  12688=>"010011101",
  12689=>"101100000",
  12690=>"111001001",
  12691=>"000011001",
  12692=>"011110001",
  12693=>"111101000",
  12694=>"000101000",
  12695=>"011111110",
  12696=>"110000100",
  12697=>"101111000",
  12698=>"001110000",
  12699=>"101000111",
  12700=>"111010111",
  12701=>"000100111",
  12702=>"000101100",
  12703=>"111000000",
  12704=>"101111011",
  12705=>"011010000",
  12706=>"101010010",
  12707=>"101100100",
  12708=>"101010010",
  12709=>"001111011",
  12710=>"000001001",
  12711=>"001000010",
  12712=>"100111011",
  12713=>"001100010",
  12714=>"100100100",
  12715=>"100010010",
  12716=>"100100101",
  12717=>"100101010",
  12718=>"000010100",
  12719=>"110000000",
  12720=>"000111010",
  12721=>"101100100",
  12722=>"011110111",
  12723=>"101000000",
  12724=>"110000101",
  12725=>"000010101",
  12726=>"011011100",
  12727=>"011000001",
  12728=>"100001010",
  12729=>"110000000",
  12730=>"101000010",
  12731=>"100100011",
  12732=>"101011100",
  12733=>"111011110",
  12734=>"101000000",
  12735=>"111110001",
  12736=>"100001001",
  12737=>"110011001",
  12738=>"110100110",
  12739=>"101111001",
  12740=>"000100111",
  12741=>"111001001",
  12742=>"101001111",
  12743=>"001010000",
  12744=>"010011010",
  12745=>"110010110",
  12746=>"111011110",
  12747=>"111001101",
  12748=>"000100001",
  12749=>"011100001",
  12750=>"001000111",
  12751=>"100001101",
  12752=>"101111110",
  12753=>"001101101",
  12754=>"001011000",
  12755=>"101101111",
  12756=>"010010110",
  12757=>"111110011",
  12758=>"010011101",
  12759=>"111010101",
  12760=>"110011110",
  12761=>"101101010",
  12762=>"001100001",
  12763=>"111001100",
  12764=>"110010010",
  12765=>"101000110",
  12766=>"101110011",
  12767=>"110000001",
  12768=>"001000001",
  12769=>"010010101",
  12770=>"001110001",
  12771=>"101010100",
  12772=>"000010100",
  12773=>"000000110",
  12774=>"001101111",
  12775=>"010101111",
  12776=>"001001001",
  12777=>"010000010",
  12778=>"001011001",
  12779=>"100001100",
  12780=>"000100001",
  12781=>"110100100",
  12782=>"000000000",
  12783=>"101000100",
  12784=>"010101011",
  12785=>"110110001",
  12786=>"110110101",
  12787=>"011100101",
  12788=>"101110110",
  12789=>"011010011",
  12790=>"101011001",
  12791=>"100011110",
  12792=>"101110010",
  12793=>"010000011",
  12794=>"110100100",
  12795=>"011111110",
  12796=>"111000001",
  12797=>"111100111",
  12798=>"110000111",
  12799=>"001000000",
  12800=>"110111101",
  12801=>"110110110",
  12802=>"000011101",
  12803=>"001101110",
  12804=>"000110011",
  12805=>"001110011",
  12806=>"001110100",
  12807=>"110100010",
  12808=>"001010110",
  12809=>"111100111",
  12810=>"111001000",
  12811=>"101100111",
  12812=>"100100010",
  12813=>"110001010",
  12814=>"000000001",
  12815=>"010000110",
  12816=>"110101010",
  12817=>"001001000",
  12818=>"111000001",
  12819=>"110001000",
  12820=>"111010110",
  12821=>"111101011",
  12822=>"000111010",
  12823=>"011010000",
  12824=>"001111101",
  12825=>"011011000",
  12826=>"000100010",
  12827=>"010000010",
  12828=>"000011101",
  12829=>"011111101",
  12830=>"000000001",
  12831=>"110111010",
  12832=>"001110101",
  12833=>"001011111",
  12834=>"111001100",
  12835=>"000111001",
  12836=>"011010111",
  12837=>"000100111",
  12838=>"101100011",
  12839=>"000100111",
  12840=>"001100000",
  12841=>"111000000",
  12842=>"010010101",
  12843=>"101101000",
  12844=>"000110101",
  12845=>"101001111",
  12846=>"110111111",
  12847=>"110101111",
  12848=>"110001011",
  12849=>"101000100",
  12850=>"011100010",
  12851=>"100011100",
  12852=>"011011000",
  12853=>"110111011",
  12854=>"111111011",
  12855=>"010010001",
  12856=>"000111111",
  12857=>"011110111",
  12858=>"111010100",
  12859=>"101111111",
  12860=>"100101111",
  12861=>"001010100",
  12862=>"000101010",
  12863=>"011000010",
  12864=>"111010110",
  12865=>"011101101",
  12866=>"111101110",
  12867=>"111100100",
  12868=>"000000110",
  12869=>"010011100",
  12870=>"000000001",
  12871=>"000000110",
  12872=>"100010001",
  12873=>"000111101",
  12874=>"011111100",
  12875=>"111010111",
  12876=>"100100111",
  12877=>"000001101",
  12878=>"101111000",
  12879=>"000010110",
  12880=>"101110110",
  12881=>"110010000",
  12882=>"111001011",
  12883=>"000001101",
  12884=>"100010101",
  12885=>"000111000",
  12886=>"010010111",
  12887=>"011110000",
  12888=>"110010010",
  12889=>"101110110",
  12890=>"001011011",
  12891=>"011000010",
  12892=>"100110011",
  12893=>"101100101",
  12894=>"111001010",
  12895=>"101110011",
  12896=>"000010011",
  12897=>"000010100",
  12898=>"001111011",
  12899=>"011001101",
  12900=>"111011001",
  12901=>"001000101",
  12902=>"100100000",
  12903=>"011010101",
  12904=>"110110111",
  12905=>"111010100",
  12906=>"011001110",
  12907=>"110110101",
  12908=>"001111101",
  12909=>"101001100",
  12910=>"001001110",
  12911=>"111111111",
  12912=>"001101001",
  12913=>"010001111",
  12914=>"101101101",
  12915=>"010100010",
  12916=>"011000001",
  12917=>"000111011",
  12918=>"100001110",
  12919=>"001000000",
  12920=>"111011111",
  12921=>"010010000",
  12922=>"010011101",
  12923=>"100000001",
  12924=>"010100101",
  12925=>"101001110",
  12926=>"110001111",
  12927=>"111111100",
  12928=>"000001100",
  12929=>"101110100",
  12930=>"111001010",
  12931=>"011001001",
  12932=>"100111100",
  12933=>"100000010",
  12934=>"111010111",
  12935=>"001001100",
  12936=>"011111010",
  12937=>"001100000",
  12938=>"110100011",
  12939=>"111000111",
  12940=>"011010110",
  12941=>"001101010",
  12942=>"110011000",
  12943=>"011110110",
  12944=>"011100110",
  12945=>"011100010",
  12946=>"010000101",
  12947=>"011001001",
  12948=>"011001100",
  12949=>"000100000",
  12950=>"010010000",
  12951=>"001100101",
  12952=>"001111110",
  12953=>"000000110",
  12954=>"000000101",
  12955=>"010000000",
  12956=>"000000010",
  12957=>"100111101",
  12958=>"011101001",
  12959=>"001100100",
  12960=>"011110000",
  12961=>"000000100",
  12962=>"001010010",
  12963=>"001111000",
  12964=>"100011100",
  12965=>"101111111",
  12966=>"101010001",
  12967=>"010111000",
  12968=>"011011000",
  12969=>"010110000",
  12970=>"010010111",
  12971=>"001101010",
  12972=>"010011010",
  12973=>"101101011",
  12974=>"000000000",
  12975=>"010010000",
  12976=>"011100101",
  12977=>"110010001",
  12978=>"110011001",
  12979=>"101110111",
  12980=>"111111110",
  12981=>"001011010",
  12982=>"001001111",
  12983=>"011010100",
  12984=>"010110010",
  12985=>"001010110",
  12986=>"110100000",
  12987=>"000000000",
  12988=>"100111110",
  12989=>"011010000",
  12990=>"111111001",
  12991=>"111100000",
  12992=>"111101100",
  12993=>"011111010",
  12994=>"101110111",
  12995=>"011001001",
  12996=>"010100111",
  12997=>"001101001",
  12998=>"011101110",
  12999=>"000000000",
  13000=>"000001011",
  13001=>"011101010",
  13002=>"111100001",
  13003=>"111010100",
  13004=>"001001001",
  13005=>"111011111",
  13006=>"111110110",
  13007=>"100111100",
  13008=>"111110011",
  13009=>"110000011",
  13010=>"011100000",
  13011=>"110011000",
  13012=>"100011100",
  13013=>"100011001",
  13014=>"110110111",
  13015=>"001011001",
  13016=>"110000000",
  13017=>"100111100",
  13018=>"100010001",
  13019=>"100101100",
  13020=>"110101110",
  13021=>"111001010",
  13022=>"101101111",
  13023=>"010000111",
  13024=>"011100111",
  13025=>"011101111",
  13026=>"000010111",
  13027=>"000110000",
  13028=>"010001101",
  13029=>"010001010",
  13030=>"110101000",
  13031=>"000010111",
  13032=>"001110011",
  13033=>"101000111",
  13034=>"011101000",
  13035=>"101010100",
  13036=>"011000110",
  13037=>"000100010",
  13038=>"101011010",
  13039=>"001010001",
  13040=>"000101111",
  13041=>"011011000",
  13042=>"100011101",
  13043=>"101011101",
  13044=>"101110010",
  13045=>"100011000",
  13046=>"010111000",
  13047=>"111110001",
  13048=>"001101111",
  13049=>"001001110",
  13050=>"000010001",
  13051=>"110001010",
  13052=>"101111110",
  13053=>"001101011",
  13054=>"000010010",
  13055=>"111110100",
  13056=>"101110000",
  13057=>"010010011",
  13058=>"000110111",
  13059=>"100001110",
  13060=>"001100110",
  13061=>"010100011",
  13062=>"111000100",
  13063=>"110110101",
  13064=>"110000011",
  13065=>"101011011",
  13066=>"010101110",
  13067=>"100100100",
  13068=>"010000111",
  13069=>"111001011",
  13070=>"101000001",
  13071=>"100100111",
  13072=>"000100110",
  13073=>"001000101",
  13074=>"001101011",
  13075=>"111011110",
  13076=>"101110110",
  13077=>"110111111",
  13078=>"011010110",
  13079=>"101111101",
  13080=>"100000111",
  13081=>"001010011",
  13082=>"000000000",
  13083=>"001101001",
  13084=>"011001111",
  13085=>"010000110",
  13086=>"001001101",
  13087=>"000010100",
  13088=>"100011110",
  13089=>"110110010",
  13090=>"011010010",
  13091=>"010101100",
  13092=>"110101100",
  13093=>"110100000",
  13094=>"111110100",
  13095=>"101111010",
  13096=>"101100111",
  13097=>"000101011",
  13098=>"010101100",
  13099=>"001100011",
  13100=>"110001101",
  13101=>"011001000",
  13102=>"110001011",
  13103=>"111010101",
  13104=>"010000000",
  13105=>"010010010",
  13106=>"101111000",
  13107=>"000110100",
  13108=>"010000000",
  13109=>"101111111",
  13110=>"110101010",
  13111=>"000011101",
  13112=>"110110000",
  13113=>"011010010",
  13114=>"000001110",
  13115=>"111111101",
  13116=>"000000011",
  13117=>"011001000",
  13118=>"001100011",
  13119=>"011110101",
  13120=>"110100101",
  13121=>"100100010",
  13122=>"111111010",
  13123=>"110011101",
  13124=>"011000010",
  13125=>"111101111",
  13126=>"100011101",
  13127=>"000011010",
  13128=>"000011101",
  13129=>"010011011",
  13130=>"000110110",
  13131=>"110000111",
  13132=>"001111010",
  13133=>"000111110",
  13134=>"110111110",
  13135=>"111011011",
  13136=>"101001100",
  13137=>"011011000",
  13138=>"010010100",
  13139=>"001001010",
  13140=>"100100101",
  13141=>"011011110",
  13142=>"010001000",
  13143=>"011000100",
  13144=>"111100010",
  13145=>"101001011",
  13146=>"001011100",
  13147=>"011010001",
  13148=>"010111111",
  13149=>"001100101",
  13150=>"100010111",
  13151=>"000110101",
  13152=>"111001010",
  13153=>"011001010",
  13154=>"000000011",
  13155=>"010000110",
  13156=>"110001010",
  13157=>"111101101",
  13158=>"111100100",
  13159=>"001001000",
  13160=>"101101011",
  13161=>"010111001",
  13162=>"000010010",
  13163=>"101000010",
  13164=>"100101100",
  13165=>"001000011",
  13166=>"110011110",
  13167=>"000001110",
  13168=>"011101010",
  13169=>"101011110",
  13170=>"110110101",
  13171=>"111100111",
  13172=>"100100111",
  13173=>"111100000",
  13174=>"110001100",
  13175=>"111000101",
  13176=>"011000110",
  13177=>"001010111",
  13178=>"110110100",
  13179=>"000100000",
  13180=>"000010100",
  13181=>"010101101",
  13182=>"011010110",
  13183=>"101010101",
  13184=>"011010111",
  13185=>"001000110",
  13186=>"100000110",
  13187=>"000101011",
  13188=>"101010010",
  13189=>"110010001",
  13190=>"000000111",
  13191=>"101001011",
  13192=>"001111111",
  13193=>"001111011",
  13194=>"111001100",
  13195=>"101111000",
  13196=>"011101010",
  13197=>"010011011",
  13198=>"111100001",
  13199=>"001111101",
  13200=>"010010100",
  13201=>"101001100",
  13202=>"010100000",
  13203=>"010010100",
  13204=>"010001001",
  13205=>"100110100",
  13206=>"000100001",
  13207=>"000100010",
  13208=>"101100011",
  13209=>"010000101",
  13210=>"100111010",
  13211=>"010110100",
  13212=>"110101110",
  13213=>"010101100",
  13214=>"100111100",
  13215=>"000001110",
  13216=>"110111011",
  13217=>"100010001",
  13218=>"100111111",
  13219=>"011000000",
  13220=>"100110000",
  13221=>"101000110",
  13222=>"000100011",
  13223=>"011111011",
  13224=>"011000000",
  13225=>"010100011",
  13226=>"110000110",
  13227=>"101000010",
  13228=>"001111011",
  13229=>"101011100",
  13230=>"111110100",
  13231=>"001111110",
  13232=>"111111011",
  13233=>"111101100",
  13234=>"110001111",
  13235=>"100110101",
  13236=>"000001100",
  13237=>"101101111",
  13238=>"000111010",
  13239=>"001111011",
  13240=>"100110000",
  13241=>"100000000",
  13242=>"101010111",
  13243=>"000000000",
  13244=>"101011010",
  13245=>"101010001",
  13246=>"010110111",
  13247=>"001011000",
  13248=>"110000000",
  13249=>"000101010",
  13250=>"010010100",
  13251=>"100001010",
  13252=>"110111111",
  13253=>"111100000",
  13254=>"010101001",
  13255=>"010000001",
  13256=>"101111110",
  13257=>"011000011",
  13258=>"100101000",
  13259=>"010010100",
  13260=>"101101101",
  13261=>"011101100",
  13262=>"100111011",
  13263=>"111010100",
  13264=>"100101000",
  13265=>"001010011",
  13266=>"111110011",
  13267=>"010000100",
  13268=>"111001011",
  13269=>"111010001",
  13270=>"111001010",
  13271=>"110010110",
  13272=>"110000010",
  13273=>"110000011",
  13274=>"100000001",
  13275=>"000110111",
  13276=>"001011100",
  13277=>"011110010",
  13278=>"001111100",
  13279=>"010100001",
  13280=>"100101010",
  13281=>"110100111",
  13282=>"100100001",
  13283=>"001010010",
  13284=>"100000000",
  13285=>"011100001",
  13286=>"101001001",
  13287=>"010010111",
  13288=>"100011101",
  13289=>"010000111",
  13290=>"110011000",
  13291=>"111011110",
  13292=>"010011000",
  13293=>"101000000",
  13294=>"011111000",
  13295=>"000110100",
  13296=>"000101111",
  13297=>"000101101",
  13298=>"011111010",
  13299=>"001010110",
  13300=>"101010111",
  13301=>"000101101",
  13302=>"100011111",
  13303=>"110000010",
  13304=>"001111100",
  13305=>"111000111",
  13306=>"011101101",
  13307=>"001011100",
  13308=>"110000111",
  13309=>"100111000",
  13310=>"111101111",
  13311=>"001101100",
  13312=>"001100011",
  13313=>"101001101",
  13314=>"110111101",
  13315=>"000001001",
  13316=>"001000101",
  13317=>"111000100",
  13318=>"011001010",
  13319=>"100100111",
  13320=>"100011000",
  13321=>"110010010",
  13322=>"011010110",
  13323=>"000111101",
  13324=>"101101101",
  13325=>"011010010",
  13326=>"011111101",
  13327=>"001000111",
  13328=>"110110111",
  13329=>"001100001",
  13330=>"100011111",
  13331=>"000000111",
  13332=>"111100011",
  13333=>"101001100",
  13334=>"000011101",
  13335=>"010000010",
  13336=>"010100110",
  13337=>"001110000",
  13338=>"110111000",
  13339=>"100011000",
  13340=>"110001110",
  13341=>"001010110",
  13342=>"000101100",
  13343=>"100110010",
  13344=>"100010100",
  13345=>"011110110",
  13346=>"001011110",
  13347=>"110011011",
  13348=>"001000010",
  13349=>"011100111",
  13350=>"111011010",
  13351=>"001000001",
  13352=>"000110110",
  13353=>"110000000",
  13354=>"110110101",
  13355=>"101010110",
  13356=>"101010101",
  13357=>"001010011",
  13358=>"001000100",
  13359=>"101001100",
  13360=>"001100110",
  13361=>"111101101",
  13362=>"010011111",
  13363=>"010101100",
  13364=>"110110110",
  13365=>"000010110",
  13366=>"000001110",
  13367=>"000000011",
  13368=>"100111100",
  13369=>"010101101",
  13370=>"011100100",
  13371=>"110101010",
  13372=>"111000000",
  13373=>"001010101",
  13374=>"100000110",
  13375=>"000010100",
  13376=>"011100101",
  13377=>"001010010",
  13378=>"110100000",
  13379=>"000110110",
  13380=>"110111010",
  13381=>"101110110",
  13382=>"111100000",
  13383=>"001000011",
  13384=>"011101010",
  13385=>"111011001",
  13386=>"001000010",
  13387=>"101111001",
  13388=>"100000000",
  13389=>"111001010",
  13390=>"110100011",
  13391=>"100111000",
  13392=>"001101111",
  13393=>"000111100",
  13394=>"010100000",
  13395=>"100001111",
  13396=>"000100100",
  13397=>"110011010",
  13398=>"011011111",
  13399=>"111100001",
  13400=>"101101101",
  13401=>"101110000",
  13402=>"000110110",
  13403=>"111100110",
  13404=>"010001111",
  13405=>"001100111",
  13406=>"011111101",
  13407=>"110101111",
  13408=>"011101111",
  13409=>"111110000",
  13410=>"010001010",
  13411=>"011000000",
  13412=>"010011011",
  13413=>"111111110",
  13414=>"000111010",
  13415=>"100100110",
  13416=>"111100111",
  13417=>"111101011",
  13418=>"011011100",
  13419=>"001010111",
  13420=>"010000000",
  13421=>"101001100",
  13422=>"101100011",
  13423=>"100100011",
  13424=>"000011011",
  13425=>"010000001",
  13426=>"000000100",
  13427=>"001110000",
  13428=>"101101110",
  13429=>"110101000",
  13430=>"000001111",
  13431=>"001001010",
  13432=>"101101111",
  13433=>"010100011",
  13434=>"001101011",
  13435=>"010011001",
  13436=>"001111011",
  13437=>"111011110",
  13438=>"001001110",
  13439=>"111101000",
  13440=>"100111011",
  13441=>"010100101",
  13442=>"000010100",
  13443=>"100000000",
  13444=>"011110001",
  13445=>"100010011",
  13446=>"011111111",
  13447=>"011010010",
  13448=>"000001110",
  13449=>"111101110",
  13450=>"001001011",
  13451=>"111111110",
  13452=>"001000011",
  13453=>"110011001",
  13454=>"110101000",
  13455=>"000000001",
  13456=>"000000001",
  13457=>"110111100",
  13458=>"100010011",
  13459=>"010000010",
  13460=>"000001010",
  13461=>"111110011",
  13462=>"010000111",
  13463=>"111001000",
  13464=>"100001100",
  13465=>"001011110",
  13466=>"001001101",
  13467=>"101000000",
  13468=>"100011001",
  13469=>"110100110",
  13470=>"000001000",
  13471=>"011001011",
  13472=>"010000001",
  13473=>"011000101",
  13474=>"000010100",
  13475=>"111001100",
  13476=>"010110000",
  13477=>"101010010",
  13478=>"111000110",
  13479=>"101110000",
  13480=>"111011010",
  13481=>"000100101",
  13482=>"100111110",
  13483=>"001010011",
  13484=>"111001001",
  13485=>"000100001",
  13486=>"010111100",
  13487=>"100100101",
  13488=>"011011010",
  13489=>"010000001",
  13490=>"000111111",
  13491=>"101000110",
  13492=>"111011011",
  13493=>"010100110",
  13494=>"010110101",
  13495=>"111010100",
  13496=>"100010000",
  13497=>"101000001",
  13498=>"011111111",
  13499=>"011100010",
  13500=>"011001001",
  13501=>"111111010",
  13502=>"011001101",
  13503=>"001010001",
  13504=>"111101111",
  13505=>"001010010",
  13506=>"101010001",
  13507=>"100101111",
  13508=>"100001010",
  13509=>"101000010",
  13510=>"001101011",
  13511=>"111101010",
  13512=>"011010000",
  13513=>"100100100",
  13514=>"001010111",
  13515=>"100100011",
  13516=>"101111110",
  13517=>"000110010",
  13518=>"111001111",
  13519=>"100010000",
  13520=>"000000001",
  13521=>"101100110",
  13522=>"000010110",
  13523=>"001101100",
  13524=>"010001100",
  13525=>"011100101",
  13526=>"010010111",
  13527=>"111010101",
  13528=>"100100100",
  13529=>"111100001",
  13530=>"001010000",
  13531=>"110011101",
  13532=>"101001111",
  13533=>"111101011",
  13534=>"001010001",
  13535=>"010011011",
  13536=>"000000010",
  13537=>"101010100",
  13538=>"000010001",
  13539=>"011011001",
  13540=>"111011011",
  13541=>"001010110",
  13542=>"000110010",
  13543=>"100100110",
  13544=>"010101111",
  13545=>"010011010",
  13546=>"011000000",
  13547=>"001110111",
  13548=>"100001001",
  13549=>"110011000",
  13550=>"010111001",
  13551=>"100011101",
  13552=>"101000010",
  13553=>"010000010",
  13554=>"100010110",
  13555=>"001011111",
  13556=>"100000110",
  13557=>"000000101",
  13558=>"001111011",
  13559=>"100101010",
  13560=>"011110110",
  13561=>"001101010",
  13562=>"011110000",
  13563=>"110010101",
  13564=>"011001001",
  13565=>"110010010",
  13566=>"011110110",
  13567=>"000111010",
  13568=>"111110000",
  13569=>"100001101",
  13570=>"011010111",
  13571=>"101001111",
  13572=>"011010111",
  13573=>"011010101",
  13574=>"000011001",
  13575=>"011110100",
  13576=>"110011111",
  13577=>"011100001",
  13578=>"111111111",
  13579=>"000100000",
  13580=>"000000100",
  13581=>"101110101",
  13582=>"100011001",
  13583=>"011101000",
  13584=>"001101011",
  13585=>"011001100",
  13586=>"010110111",
  13587=>"110010100",
  13588=>"010101000",
  13589=>"000100001",
  13590=>"000000000",
  13591=>"101000000",
  13592=>"011011100",
  13593=>"101101001",
  13594=>"100110001",
  13595=>"111110100",
  13596=>"111111001",
  13597=>"000010010",
  13598=>"111101000",
  13599=>"011101000",
  13600=>"000110011",
  13601=>"101001001",
  13602=>"111001110",
  13603=>"100000100",
  13604=>"000100110",
  13605=>"001111101",
  13606=>"101011110",
  13607=>"010000011",
  13608=>"001011101",
  13609=>"110000001",
  13610=>"001001011",
  13611=>"101110111",
  13612=>"110101110",
  13613=>"101100110",
  13614=>"010011110",
  13615=>"011101010",
  13616=>"001001010",
  13617=>"011111001",
  13618=>"101101100",
  13619=>"011010100",
  13620=>"100001111",
  13621=>"100111101",
  13622=>"110111100",
  13623=>"100110001",
  13624=>"000011000",
  13625=>"101100100",
  13626=>"010000110",
  13627=>"010100011",
  13628=>"010000100",
  13629=>"010000111",
  13630=>"100101010",
  13631=>"000001011",
  13632=>"001110001",
  13633=>"110110100",
  13634=>"100011010",
  13635=>"011000000",
  13636=>"100000010",
  13637=>"100000100",
  13638=>"011011000",
  13639=>"000101010",
  13640=>"111100011",
  13641=>"010001001",
  13642=>"100011011",
  13643=>"011000111",
  13644=>"011101010",
  13645=>"010110110",
  13646=>"010001000",
  13647=>"101001001",
  13648=>"100000001",
  13649=>"101011011",
  13650=>"111000010",
  13651=>"101101000",
  13652=>"000010101",
  13653=>"001101100",
  13654=>"110001111",
  13655=>"101010000",
  13656=>"110100001",
  13657=>"011110100",
  13658=>"000100100",
  13659=>"100100001",
  13660=>"011101111",
  13661=>"101010010",
  13662=>"110001100",
  13663=>"100010000",
  13664=>"101000000",
  13665=>"011110111",
  13666=>"001000110",
  13667=>"111010010",
  13668=>"010101100",
  13669=>"010100111",
  13670=>"110000010",
  13671=>"011001011",
  13672=>"110110100",
  13673=>"100111110",
  13674=>"001010001",
  13675=>"111111001",
  13676=>"000110010",
  13677=>"111110001",
  13678=>"100000001",
  13679=>"001110111",
  13680=>"011010100",
  13681=>"010111000",
  13682=>"000101011",
  13683=>"011011100",
  13684=>"011000101",
  13685=>"000101011",
  13686=>"100110011",
  13687=>"111111001",
  13688=>"111111100",
  13689=>"000111010",
  13690=>"111100000",
  13691=>"000110101",
  13692=>"101001001",
  13693=>"110001110",
  13694=>"010001010",
  13695=>"111111011",
  13696=>"010111011",
  13697=>"010010110",
  13698=>"000110001",
  13699=>"101100101",
  13700=>"111110001",
  13701=>"000001011",
  13702=>"000100111",
  13703=>"110101001",
  13704=>"100100000",
  13705=>"010001001",
  13706=>"110110110",
  13707=>"101001111",
  13708=>"110011110",
  13709=>"000010000",
  13710=>"100001011",
  13711=>"100011100",
  13712=>"000111011",
  13713=>"000000000",
  13714=>"110110110",
  13715=>"000110001",
  13716=>"011100111",
  13717=>"000100111",
  13718=>"100010011",
  13719=>"100101110",
  13720=>"111011101",
  13721=>"110111011",
  13722=>"110010111",
  13723=>"001000111",
  13724=>"101011010",
  13725=>"111001011",
  13726=>"000111101",
  13727=>"100110110",
  13728=>"101011101",
  13729=>"011011000",
  13730=>"101110110",
  13731=>"111010000",
  13732=>"110001000",
  13733=>"100010101",
  13734=>"111111110",
  13735=>"000000101",
  13736=>"110010010",
  13737=>"011000110",
  13738=>"001110101",
  13739=>"000111000",
  13740=>"000010010",
  13741=>"011010001",
  13742=>"000000000",
  13743=>"000101000",
  13744=>"000100000",
  13745=>"100111100",
  13746=>"110110011",
  13747=>"111001111",
  13748=>"111110001",
  13749=>"001010100",
  13750=>"010011000",
  13751=>"110010110",
  13752=>"101111111",
  13753=>"111101110",
  13754=>"111111101",
  13755=>"101001100",
  13756=>"100101101",
  13757=>"010101101",
  13758=>"010110010",
  13759=>"000010010",
  13760=>"000001010",
  13761=>"111110111",
  13762=>"001110110",
  13763=>"101100001",
  13764=>"100100000",
  13765=>"101000111",
  13766=>"000100011",
  13767=>"010010000",
  13768=>"011001001",
  13769=>"000011111",
  13770=>"111001010",
  13771=>"001100111",
  13772=>"101110011",
  13773=>"100110000",
  13774=>"100010111",
  13775=>"000100111",
  13776=>"110010110",
  13777=>"001100001",
  13778=>"011111010",
  13779=>"101101011",
  13780=>"110111111",
  13781=>"110010110",
  13782=>"101100010",
  13783=>"011100000",
  13784=>"100111101",
  13785=>"001111010",
  13786=>"101111111",
  13787=>"001110000",
  13788=>"100111010",
  13789=>"000010011",
  13790=>"000111111",
  13791=>"111110001",
  13792=>"010100110",
  13793=>"010011000",
  13794=>"110010000",
  13795=>"001011111",
  13796=>"010111111",
  13797=>"100011000",
  13798=>"101110110",
  13799=>"001111100",
  13800=>"100010010",
  13801=>"000110111",
  13802=>"000001000",
  13803=>"100010001",
  13804=>"111101100",
  13805=>"110110001",
  13806=>"101001101",
  13807=>"101110000",
  13808=>"011111111",
  13809=>"111011011",
  13810=>"101010010",
  13811=>"010110101",
  13812=>"001100000",
  13813=>"010110100",
  13814=>"011011101",
  13815=>"111100000",
  13816=>"111110111",
  13817=>"010011100",
  13818=>"001101101",
  13819=>"111100111",
  13820=>"110110111",
  13821=>"111001000",
  13822=>"011010110",
  13823=>"100111000",
  13824=>"000010110",
  13825=>"000000100",
  13826=>"011011101",
  13827=>"010010100",
  13828=>"110000010",
  13829=>"111110100",
  13830=>"110010010",
  13831=>"100101000",
  13832=>"000100000",
  13833=>"000100001",
  13834=>"011111111",
  13835=>"001110100",
  13836=>"011010100",
  13837=>"111101010",
  13838=>"100000001",
  13839=>"100000101",
  13840=>"010011001",
  13841=>"011001111",
  13842=>"000000100",
  13843=>"101001110",
  13844=>"001000101",
  13845=>"000001011",
  13846=>"110100010",
  13847=>"110000100",
  13848=>"010011100",
  13849=>"100000110",
  13850=>"001001001",
  13851=>"000000110",
  13852=>"110000000",
  13853=>"110000100",
  13854=>"111100110",
  13855=>"110101100",
  13856=>"000001100",
  13857=>"001111101",
  13858=>"100110011",
  13859=>"111010000",
  13860=>"000100000",
  13861=>"110010011",
  13862=>"110100000",
  13863=>"110110001",
  13864=>"101111000",
  13865=>"111010101",
  13866=>"110111000",
  13867=>"111101101",
  13868=>"001010000",
  13869=>"110010111",
  13870=>"010111000",
  13871=>"110001110",
  13872=>"000010100",
  13873=>"001101100",
  13874=>"101111011",
  13875=>"100001111",
  13876=>"011010110",
  13877=>"001101110",
  13878=>"000011100",
  13879=>"110111011",
  13880=>"000111001",
  13881=>"101001011",
  13882=>"111001010",
  13883=>"010101010",
  13884=>"101101100",
  13885=>"001000011",
  13886=>"010000101",
  13887=>"001101101",
  13888=>"110101110",
  13889=>"000000110",
  13890=>"000110011",
  13891=>"011000111",
  13892=>"010010000",
  13893=>"011010010",
  13894=>"101000011",
  13895=>"100110110",
  13896=>"011010000",
  13897=>"001001010",
  13898=>"111001100",
  13899=>"000001101",
  13900=>"111110001",
  13901=>"000000010",
  13902=>"011011110",
  13903=>"011001011",
  13904=>"001100011",
  13905=>"011100110",
  13906=>"000010000",
  13907=>"000110111",
  13908=>"010000100",
  13909=>"010000010",
  13910=>"010011000",
  13911=>"100000101",
  13912=>"101000101",
  13913=>"100010101",
  13914=>"001101001",
  13915=>"010010000",
  13916=>"011011011",
  13917=>"111000100",
  13918=>"101101101",
  13919=>"001101100",
  13920=>"010001011",
  13921=>"111101100",
  13922=>"000101101",
  13923=>"111111110",
  13924=>"101011010",
  13925=>"000100101",
  13926=>"101011000",
  13927=>"001111110",
  13928=>"000000101",
  13929=>"000111110",
  13930=>"111110001",
  13931=>"001101100",
  13932=>"000100001",
  13933=>"111011000",
  13934=>"011011110",
  13935=>"110010111",
  13936=>"110110100",
  13937=>"000111110",
  13938=>"110101110",
  13939=>"001101101",
  13940=>"111110100",
  13941=>"001000001",
  13942=>"011101101",
  13943=>"111000000",
  13944=>"011011000",
  13945=>"010000110",
  13946=>"101010010",
  13947=>"111001101",
  13948=>"000000100",
  13949=>"100110010",
  13950=>"011101110",
  13951=>"101110100",
  13952=>"011110101",
  13953=>"011001000",
  13954=>"101010010",
  13955=>"001001100",
  13956=>"001000111",
  13957=>"010000000",
  13958=>"111110111",
  13959=>"110010111",
  13960=>"011100111",
  13961=>"010011101",
  13962=>"010100110",
  13963=>"000101101",
  13964=>"100100111",
  13965=>"110111010",
  13966=>"001000111",
  13967=>"011010111",
  13968=>"100001010",
  13969=>"111000011",
  13970=>"000010110",
  13971=>"101010000",
  13972=>"100000011",
  13973=>"110101100",
  13974=>"011111001",
  13975=>"001100110",
  13976=>"111011001",
  13977=>"101001111",
  13978=>"111000010",
  13979=>"000000000",
  13980=>"001111100",
  13981=>"110110110",
  13982=>"111100010",
  13983=>"010110000",
  13984=>"000100101",
  13985=>"111101100",
  13986=>"000001000",
  13987=>"111000111",
  13988=>"011000010",
  13989=>"100101111",
  13990=>"001100101",
  13991=>"100000011",
  13992=>"110110011",
  13993=>"000010111",
  13994=>"001100011",
  13995=>"000110110",
  13996=>"011000110",
  13997=>"001111101",
  13998=>"011111001",
  13999=>"100110101",
  14000=>"110101100",
  14001=>"001100011",
  14002=>"000110010",
  14003=>"000100000",
  14004=>"111011111",
  14005=>"101100110",
  14006=>"011000101",
  14007=>"111001100",
  14008=>"110110000",
  14009=>"110100110",
  14010=>"101000000",
  14011=>"001011101",
  14012=>"111000011",
  14013=>"001110000",
  14014=>"111011100",
  14015=>"101011111",
  14016=>"001101100",
  14017=>"010001100",
  14018=>"101100001",
  14019=>"011000111",
  14020=>"011011001",
  14021=>"110101011",
  14022=>"001010011",
  14023=>"001110010",
  14024=>"010100000",
  14025=>"010111101",
  14026=>"001001101",
  14027=>"000111010",
  14028=>"010011111",
  14029=>"001001100",
  14030=>"100111100",
  14031=>"010100010",
  14032=>"001100100",
  14033=>"100110100",
  14034=>"101010000",
  14035=>"001011010",
  14036=>"000010010",
  14037=>"001101011",
  14038=>"010101111",
  14039=>"101000110",
  14040=>"011100001",
  14041=>"110000001",
  14042=>"011001100",
  14043=>"001001001",
  14044=>"100101101",
  14045=>"011101000",
  14046=>"101001010",
  14047=>"110000110",
  14048=>"001001001",
  14049=>"100001111",
  14050=>"111000111",
  14051=>"100011010",
  14052=>"110010011",
  14053=>"011011110",
  14054=>"111110101",
  14055=>"001011100",
  14056=>"010010011",
  14057=>"011001000",
  14058=>"101011011",
  14059=>"110111111",
  14060=>"001010000",
  14061=>"110000111",
  14062=>"111010000",
  14063=>"000111111",
  14064=>"111100111",
  14065=>"101110010",
  14066=>"110110110",
  14067=>"011010100",
  14068=>"010110111",
  14069=>"001011111",
  14070=>"111100000",
  14071=>"100010100",
  14072=>"100000011",
  14073=>"101010110",
  14074=>"100101011",
  14075=>"000111100",
  14076=>"001100101",
  14077=>"111111000",
  14078=>"101111001",
  14079=>"110101100",
  14080=>"101110010",
  14081=>"001001101",
  14082=>"100100000",
  14083=>"100000101",
  14084=>"001010110",
  14085=>"110101001",
  14086=>"000001100",
  14087=>"111100101",
  14088=>"101010011",
  14089=>"011011000",
  14090=>"100010010",
  14091=>"101011011",
  14092=>"000001111",
  14093=>"111111001",
  14094=>"000011101",
  14095=>"110011010",
  14096=>"111011000",
  14097=>"010111001",
  14098=>"110011111",
  14099=>"101010110",
  14100=>"111010010",
  14101=>"010010001",
  14102=>"111110110",
  14103=>"011001001",
  14104=>"011111010",
  14105=>"010110001",
  14106=>"101111111",
  14107=>"111101011",
  14108=>"110110010",
  14109=>"111101000",
  14110=>"100100011",
  14111=>"011010101",
  14112=>"101000111",
  14113=>"011110000",
  14114=>"100010110",
  14115=>"100101001",
  14116=>"111011000",
  14117=>"111001000",
  14118=>"101001001",
  14119=>"110111111",
  14120=>"001101001",
  14121=>"000110010",
  14122=>"101101100",
  14123=>"110001011",
  14124=>"011001011",
  14125=>"001101111",
  14126=>"011010011",
  14127=>"010000110",
  14128=>"100010010",
  14129=>"100000011",
  14130=>"110000101",
  14131=>"100110000",
  14132=>"000100000",
  14133=>"001100001",
  14134=>"000011011",
  14135=>"100001001",
  14136=>"100111101",
  14137=>"010100010",
  14138=>"000100101",
  14139=>"011011110",
  14140=>"111001101",
  14141=>"000010000",
  14142=>"101000010",
  14143=>"101010110",
  14144=>"011000111",
  14145=>"100000111",
  14146=>"011011010",
  14147=>"010101010",
  14148=>"000011111",
  14149=>"111110001",
  14150=>"101000000",
  14151=>"001111100",
  14152=>"110111101",
  14153=>"011011110",
  14154=>"001001001",
  14155=>"101010100",
  14156=>"101010011",
  14157=>"000001111",
  14158=>"110000011",
  14159=>"110100001",
  14160=>"010011000",
  14161=>"101111010",
  14162=>"010101000",
  14163=>"011000001",
  14164=>"001011111",
  14165=>"100110011",
  14166=>"010011110",
  14167=>"100001000",
  14168=>"001100001",
  14169=>"100001101",
  14170=>"110111100",
  14171=>"000001001",
  14172=>"011100000",
  14173=>"111001111",
  14174=>"011011100",
  14175=>"001010111",
  14176=>"111111110",
  14177=>"000111011",
  14178=>"000111111",
  14179=>"011100101",
  14180=>"011100010",
  14181=>"000111001",
  14182=>"110110010",
  14183=>"001000101",
  14184=>"100001100",
  14185=>"010001001",
  14186=>"001100000",
  14187=>"101011110",
  14188=>"001010111",
  14189=>"111001010",
  14190=>"010100010",
  14191=>"001111100",
  14192=>"110000010",
  14193=>"011001111",
  14194=>"010001111",
  14195=>"101000010",
  14196=>"110101111",
  14197=>"111101001",
  14198=>"111000100",
  14199=>"110000010",
  14200=>"011110011",
  14201=>"110111000",
  14202=>"011111000",
  14203=>"010011011",
  14204=>"000010010",
  14205=>"010100101",
  14206=>"100101010",
  14207=>"101111011",
  14208=>"111101001",
  14209=>"010100101",
  14210=>"000100110",
  14211=>"001001110",
  14212=>"010101110",
  14213=>"010100001",
  14214=>"000011001",
  14215=>"011001011",
  14216=>"011111110",
  14217=>"000001011",
  14218=>"001101101",
  14219=>"010001011",
  14220=>"100101100",
  14221=>"101011000",
  14222=>"100010001",
  14223=>"101011110",
  14224=>"010000001",
  14225=>"010000110",
  14226=>"100000100",
  14227=>"011101111",
  14228=>"010011000",
  14229=>"110111111",
  14230=>"111101101",
  14231=>"011100000",
  14232=>"100010001",
  14233=>"010110000",
  14234=>"001100001",
  14235=>"000111011",
  14236=>"100110111",
  14237=>"100011101",
  14238=>"000011110",
  14239=>"111001000",
  14240=>"010000000",
  14241=>"100001111",
  14242=>"110000110",
  14243=>"101011011",
  14244=>"100000100",
  14245=>"101000001",
  14246=>"001111110",
  14247=>"000000001",
  14248=>"010100100",
  14249=>"011010101",
  14250=>"101001001",
  14251=>"110000100",
  14252=>"001000010",
  14253=>"111010011",
  14254=>"101111101",
  14255=>"111011010",
  14256=>"100001011",
  14257=>"110110100",
  14258=>"001011001",
  14259=>"000000111",
  14260=>"111011011",
  14261=>"010100100",
  14262=>"110011000",
  14263=>"111100100",
  14264=>"010101101",
  14265=>"000111010",
  14266=>"100000100",
  14267=>"011000101",
  14268=>"001011010",
  14269=>"010110101",
  14270=>"100001110",
  14271=>"000110011",
  14272=>"011111101",
  14273=>"000000001",
  14274=>"101001010",
  14275=>"101101100",
  14276=>"111010100",
  14277=>"001101000",
  14278=>"111000001",
  14279=>"100111101",
  14280=>"101101110",
  14281=>"000001000",
  14282=>"110100100",
  14283=>"110000000",
  14284=>"010001001",
  14285=>"111000000",
  14286=>"110101110",
  14287=>"111010110",
  14288=>"001101100",
  14289=>"000000010",
  14290=>"001001100",
  14291=>"100000000",
  14292=>"010011001",
  14293=>"000110110",
  14294=>"000100111",
  14295=>"001101101",
  14296=>"111100111",
  14297=>"100011100",
  14298=>"100010000",
  14299=>"101010010",
  14300=>"100110101",
  14301=>"011101100",
  14302=>"110011100",
  14303=>"010111011",
  14304=>"000000101",
  14305=>"010111010",
  14306=>"111001110",
  14307=>"001100101",
  14308=>"011101110",
  14309=>"100010100",
  14310=>"000100100",
  14311=>"110011010",
  14312=>"100000100",
  14313=>"111000010",
  14314=>"100000000",
  14315=>"001100110",
  14316=>"000100010",
  14317=>"100111001",
  14318=>"011100011",
  14319=>"010111101",
  14320=>"100001001",
  14321=>"000111101",
  14322=>"001100010",
  14323=>"101100001",
  14324=>"101110110",
  14325=>"001000001",
  14326=>"000110011",
  14327=>"011110101",
  14328=>"111011100",
  14329=>"000110100",
  14330=>"001101110",
  14331=>"000101101",
  14332=>"001000011",
  14333=>"101011010",
  14334=>"101000000",
  14335=>"011111101",
  14336=>"001000111",
  14337=>"111110101",
  14338=>"100010000",
  14339=>"100111000",
  14340=>"111111000",
  14341=>"100101001",
  14342=>"000000110",
  14343=>"110100011",
  14344=>"110010100",
  14345=>"001010000",
  14346=>"000011101",
  14347=>"101001000",
  14348=>"100011010",
  14349=>"000110000",
  14350=>"010001111",
  14351=>"000000010",
  14352=>"110000101",
  14353=>"110100101",
  14354=>"101110011",
  14355=>"010110101",
  14356=>"011101011",
  14357=>"010100100",
  14358=>"101011000",
  14359=>"100010000",
  14360=>"110011010",
  14361=>"100010101",
  14362=>"000001100",
  14363=>"100001011",
  14364=>"101001001",
  14365=>"011000110",
  14366=>"000001101",
  14367=>"101001101",
  14368=>"101111001",
  14369=>"010101001",
  14370=>"001010000",
  14371=>"011110110",
  14372=>"001011111",
  14373=>"010011010",
  14374=>"001110010",
  14375=>"110000100",
  14376=>"001111010",
  14377=>"010101011",
  14378=>"100111100",
  14379=>"011011111",
  14380=>"100100010",
  14381=>"001010010",
  14382=>"010011011",
  14383=>"110001001",
  14384=>"111100100",
  14385=>"111110101",
  14386=>"001100001",
  14387=>"111101101",
  14388=>"111100110",
  14389=>"000011110",
  14390=>"000000011",
  14391=>"011001101",
  14392=>"000100010",
  14393=>"001010100",
  14394=>"000011010",
  14395=>"001000011",
  14396=>"001110000",
  14397=>"000110111",
  14398=>"010101011",
  14399=>"001100111",
  14400=>"101001110",
  14401=>"100111010",
  14402=>"000000001",
  14403=>"011011000",
  14404=>"011000001",
  14405=>"001010110",
  14406=>"111010000",
  14407=>"000001010",
  14408=>"100001010",
  14409=>"001110010",
  14410=>"100100011",
  14411=>"100111001",
  14412=>"101111110",
  14413=>"010111010",
  14414=>"110010110",
  14415=>"010001100",
  14416=>"100101011",
  14417=>"100000011",
  14418=>"010011000",
  14419=>"011101100",
  14420=>"110000101",
  14421=>"111010000",
  14422=>"010100011",
  14423=>"100001010",
  14424=>"001101000",
  14425=>"101101001",
  14426=>"001000111",
  14427=>"110110101",
  14428=>"110010101",
  14429=>"101010110",
  14430=>"100111111",
  14431=>"010111110",
  14432=>"001111001",
  14433=>"111010000",
  14434=>"000101101",
  14435=>"000101000",
  14436=>"001001111",
  14437=>"101100101",
  14438=>"111000100",
  14439=>"010100000",
  14440=>"101010011",
  14441=>"011111100",
  14442=>"001111000",
  14443=>"011011101",
  14444=>"111111010",
  14445=>"011110000",
  14446=>"100010111",
  14447=>"011000111",
  14448=>"001111100",
  14449=>"100101000",
  14450=>"100010010",
  14451=>"010001001",
  14452=>"011110110",
  14453=>"101111000",
  14454=>"001111010",
  14455=>"010100011",
  14456=>"001101010",
  14457=>"001001000",
  14458=>"110110010",
  14459=>"010000100",
  14460=>"110000010",
  14461=>"100010111",
  14462=>"101111011",
  14463=>"111001110",
  14464=>"011011101",
  14465=>"101011100",
  14466=>"000001000",
  14467=>"100110111",
  14468=>"110100010",
  14469=>"010001000",
  14470=>"011000101",
  14471=>"100111100",
  14472=>"011010101",
  14473=>"101000111",
  14474=>"110000100",
  14475=>"111101110",
  14476=>"001101000",
  14477=>"101100110",
  14478=>"011011111",
  14479=>"000100011",
  14480=>"000000101",
  14481=>"011110100",
  14482=>"011010001",
  14483=>"101010100",
  14484=>"101101111",
  14485=>"111010000",
  14486=>"001110001",
  14487=>"011110000",
  14488=>"011010000",
  14489=>"000000100",
  14490=>"011101100",
  14491=>"110010001",
  14492=>"111111000",
  14493=>"111010011",
  14494=>"111000010",
  14495=>"011001111",
  14496=>"101011101",
  14497=>"110001100",
  14498=>"010011111",
  14499=>"111111011",
  14500=>"010001111",
  14501=>"110111110",
  14502=>"110010101",
  14503=>"101010011",
  14504=>"011111110",
  14505=>"010010011",
  14506=>"010010011",
  14507=>"001000100",
  14508=>"100011010",
  14509=>"100010111",
  14510=>"111100110",
  14511=>"111001010",
  14512=>"111111101",
  14513=>"110100011",
  14514=>"011100011",
  14515=>"001110010",
  14516=>"110011001",
  14517=>"001010100",
  14518=>"011011110",
  14519=>"010000011",
  14520=>"110101100",
  14521=>"100100001",
  14522=>"010110111",
  14523=>"000110011",
  14524=>"111101010",
  14525=>"010100011",
  14526=>"011011111",
  14527=>"111100000",
  14528=>"011001111",
  14529=>"111100100",
  14530=>"110111000",
  14531=>"010101111",
  14532=>"110000000",
  14533=>"110100100",
  14534=>"101100000",
  14535=>"111100011",
  14536=>"011000111",
  14537=>"111110000",
  14538=>"111011001",
  14539=>"110111001",
  14540=>"111111010",
  14541=>"100011100",
  14542=>"011000110",
  14543=>"000010001",
  14544=>"110000000",
  14545=>"011100011",
  14546=>"100010110",
  14547=>"000111000",
  14548=>"110010101",
  14549=>"010111001",
  14550=>"011011111",
  14551=>"011110110",
  14552=>"111101001",
  14553=>"101111000",
  14554=>"011001101",
  14555=>"011110101",
  14556=>"111010001",
  14557=>"001111110",
  14558=>"010000101",
  14559=>"001110101",
  14560=>"000011001",
  14561=>"101001011",
  14562=>"000000100",
  14563=>"111101011",
  14564=>"011011110",
  14565=>"000000001",
  14566=>"101000111",
  14567=>"000110111",
  14568=>"111001000",
  14569=>"111011011",
  14570=>"000111000",
  14571=>"000001001",
  14572=>"110100010",
  14573=>"100000000",
  14574=>"101010010",
  14575=>"111111010",
  14576=>"111111100",
  14577=>"001001000",
  14578=>"100100110",
  14579=>"111000110",
  14580=>"110011101",
  14581=>"100010010",
  14582=>"000100001",
  14583=>"000000100",
  14584=>"000001111",
  14585=>"110000010",
  14586=>"101011101",
  14587=>"100100011",
  14588=>"111111110",
  14589=>"001100000",
  14590=>"111111111",
  14591=>"010110000",
  14592=>"000010000",
  14593=>"101000110",
  14594=>"101111001",
  14595=>"000000111",
  14596=>"100000101",
  14597=>"010011000",
  14598=>"111000001",
  14599=>"101101100",
  14600=>"000110011",
  14601=>"101000111",
  14602=>"101001111",
  14603=>"110111110",
  14604=>"000010100",
  14605=>"111001110",
  14606=>"101111111",
  14607=>"110111110",
  14608=>"101000101",
  14609=>"100110110",
  14610=>"001000110",
  14611=>"001110100",
  14612=>"110110110",
  14613=>"111000010",
  14614=>"101110000",
  14615=>"010110000",
  14616=>"111110101",
  14617=>"100010011",
  14618=>"001110100",
  14619=>"000010110",
  14620=>"110010011",
  14621=>"101011101",
  14622=>"001101001",
  14623=>"111101100",
  14624=>"110110001",
  14625=>"001100001",
  14626=>"000011101",
  14627=>"110110100",
  14628=>"011111100",
  14629=>"010111100",
  14630=>"110100001",
  14631=>"000101001",
  14632=>"110111011",
  14633=>"111100011",
  14634=>"001001010",
  14635=>"010100100",
  14636=>"111110010",
  14637=>"111000000",
  14638=>"001111111",
  14639=>"101110000",
  14640=>"111111101",
  14641=>"000010010",
  14642=>"011001001",
  14643=>"110100001",
  14644=>"001100011",
  14645=>"001100111",
  14646=>"010001000",
  14647=>"101001100",
  14648=>"010000101",
  14649=>"011000001",
  14650=>"010000101",
  14651=>"001001101",
  14652=>"101111001",
  14653=>"100111110",
  14654=>"000110101",
  14655=>"011011101",
  14656=>"001000111",
  14657=>"111111110",
  14658=>"010000101",
  14659=>"100011100",
  14660=>"101011100",
  14661=>"101010110",
  14662=>"011000011",
  14663=>"000110101",
  14664=>"000010000",
  14665=>"010001100",
  14666=>"100110100",
  14667=>"010010110",
  14668=>"010100100",
  14669=>"101101011",
  14670=>"011010000",
  14671=>"111111100",
  14672=>"010000011",
  14673=>"010110001",
  14674=>"111011010",
  14675=>"101111000",
  14676=>"101000100",
  14677=>"111100110",
  14678=>"010110001",
  14679=>"111001110",
  14680=>"001000111",
  14681=>"000010111",
  14682=>"010111010",
  14683=>"111100111",
  14684=>"110011101",
  14685=>"100001000",
  14686=>"111001101",
  14687=>"000101011",
  14688=>"001110100",
  14689=>"100001100",
  14690=>"000001110",
  14691=>"001101111",
  14692=>"111001110",
  14693=>"010001101",
  14694=>"111111010",
  14695=>"100001000",
  14696=>"010000110",
  14697=>"000000001",
  14698=>"011000001",
  14699=>"000110110",
  14700=>"111010100",
  14701=>"101100001",
  14702=>"110010101",
  14703=>"101000100",
  14704=>"110011111",
  14705=>"001010001",
  14706=>"010000110",
  14707=>"111011010",
  14708=>"011011000",
  14709=>"011001010",
  14710=>"000101000",
  14711=>"110111010",
  14712=>"000111100",
  14713=>"000011011",
  14714=>"111011010",
  14715=>"000111100",
  14716=>"010111100",
  14717=>"001001010",
  14718=>"110000111",
  14719=>"000011101",
  14720=>"001111110",
  14721=>"001101101",
  14722=>"010001010",
  14723=>"100100011",
  14724=>"001011111",
  14725=>"000010110",
  14726=>"011111100",
  14727=>"010111100",
  14728=>"111010111",
  14729=>"110110011",
  14730=>"110011010",
  14731=>"000100000",
  14732=>"001000001",
  14733=>"000000010",
  14734=>"110001101",
  14735=>"000010010",
  14736=>"001110101",
  14737=>"000000010",
  14738=>"000011011",
  14739=>"111001000",
  14740=>"011000111",
  14741=>"000101001",
  14742=>"001101111",
  14743=>"011101011",
  14744=>"010000010",
  14745=>"000001101",
  14746=>"011100000",
  14747=>"110010010",
  14748=>"100110110",
  14749=>"111111011",
  14750=>"010111010",
  14751=>"100101110",
  14752=>"011000011",
  14753=>"001100101",
  14754=>"011100000",
  14755=>"100001000",
  14756=>"110110101",
  14757=>"000110111",
  14758=>"101110110",
  14759=>"111001000",
  14760=>"100100100",
  14761=>"110010101",
  14762=>"101100100",
  14763=>"100000010",
  14764=>"100000010",
  14765=>"101110010",
  14766=>"000001010",
  14767=>"001110011",
  14768=>"100010101",
  14769=>"110101010",
  14770=>"011101111",
  14771=>"111111111",
  14772=>"100001100",
  14773=>"101101111",
  14774=>"100100111",
  14775=>"111101110",
  14776=>"000010011",
  14777=>"011110010",
  14778=>"010110111",
  14779=>"010010000",
  14780=>"100101010",
  14781=>"000111001",
  14782=>"011101110",
  14783=>"000001100",
  14784=>"000010010",
  14785=>"101011001",
  14786=>"101011000",
  14787=>"011110100",
  14788=>"001101011",
  14789=>"101000000",
  14790=>"110101111",
  14791=>"011000010",
  14792=>"001110101",
  14793=>"000001011",
  14794=>"101011101",
  14795=>"001111101",
  14796=>"001100100",
  14797=>"100111011",
  14798=>"110101010",
  14799=>"000101000",
  14800=>"110000111",
  14801=>"100010100",
  14802=>"010010011",
  14803=>"100111000",
  14804=>"010110010",
  14805=>"010000110",
  14806=>"010111100",
  14807=>"111001010",
  14808=>"100001100",
  14809=>"111111010",
  14810=>"010111000",
  14811=>"010010111",
  14812=>"101111111",
  14813=>"100000000",
  14814=>"010000001",
  14815=>"000111111",
  14816=>"011001101",
  14817=>"101011011",
  14818=>"010000010",
  14819=>"010101000",
  14820=>"010011010",
  14821=>"101001000",
  14822=>"110010010",
  14823=>"001000110",
  14824=>"010000000",
  14825=>"001001111",
  14826=>"100000001",
  14827=>"100000001",
  14828=>"001111101",
  14829=>"110110110",
  14830=>"010010111",
  14831=>"101000000",
  14832=>"101110011",
  14833=>"110110010",
  14834=>"111001000",
  14835=>"010111000",
  14836=>"000111011",
  14837=>"011000010",
  14838=>"011101110",
  14839=>"000101101",
  14840=>"000010100",
  14841=>"111011001",
  14842=>"101010100",
  14843=>"010001010",
  14844=>"101001011",
  14845=>"111110111",
  14846=>"100011010",
  14847=>"001110100",
  14848=>"001001100",
  14849=>"011100101",
  14850=>"110001000",
  14851=>"011100110",
  14852=>"100000101",
  14853=>"101011101",
  14854=>"001001110",
  14855=>"101000101",
  14856=>"101000011",
  14857=>"010100100",
  14858=>"100101100",
  14859=>"101000001",
  14860=>"010110011",
  14861=>"111000000",
  14862=>"011101110",
  14863=>"001110001",
  14864=>"001100100",
  14865=>"111100111",
  14866=>"001110000",
  14867=>"100111011",
  14868=>"001110011",
  14869=>"110100001",
  14870=>"100101101",
  14871=>"111000011",
  14872=>"101010100",
  14873=>"110111000",
  14874=>"101010001",
  14875=>"010001110",
  14876=>"001101001",
  14877=>"001011101",
  14878=>"001111011",
  14879=>"110011000",
  14880=>"000100000",
  14881=>"000001010",
  14882=>"100011000",
  14883=>"101011010",
  14884=>"111001110",
  14885=>"000110001",
  14886=>"100001110",
  14887=>"111011100",
  14888=>"111001001",
  14889=>"000000001",
  14890=>"110100101",
  14891=>"011101010",
  14892=>"010111001",
  14893=>"000011110",
  14894=>"100010000",
  14895=>"010000000",
  14896=>"100111100",
  14897=>"110000000",
  14898=>"101110111",
  14899=>"101111011",
  14900=>"101011101",
  14901=>"101001100",
  14902=>"001101011",
  14903=>"000010100",
  14904=>"011011010",
  14905=>"110011001",
  14906=>"111101001",
  14907=>"111001101",
  14908=>"000100111",
  14909=>"011011011",
  14910=>"011100100",
  14911=>"111000101",
  14912=>"000110000",
  14913=>"001000001",
  14914=>"100010001",
  14915=>"001000011",
  14916=>"100100101",
  14917=>"010100011",
  14918=>"010100100",
  14919=>"011001000",
  14920=>"110111110",
  14921=>"001101011",
  14922=>"011001100",
  14923=>"000110010",
  14924=>"000000100",
  14925=>"000101100",
  14926=>"101001000",
  14927=>"010110101",
  14928=>"011100111",
  14929=>"110000100",
  14930=>"001011011",
  14931=>"101000000",
  14932=>"101000001",
  14933=>"001110001",
  14934=>"100101000",
  14935=>"110000111",
  14936=>"001110101",
  14937=>"110111001",
  14938=>"100001100",
  14939=>"001100101",
  14940=>"100101110",
  14941=>"101001001",
  14942=>"001001001",
  14943=>"011011010",
  14944=>"100010110",
  14945=>"001001100",
  14946=>"010100110",
  14947=>"100101111",
  14948=>"011001010",
  14949=>"011011101",
  14950=>"001000111",
  14951=>"101110001",
  14952=>"000001011",
  14953=>"110101101",
  14954=>"000111101",
  14955=>"101011000",
  14956=>"000100010",
  14957=>"111111110",
  14958=>"110000111",
  14959=>"100011011",
  14960=>"111101011",
  14961=>"011111001",
  14962=>"010011011",
  14963=>"000000101",
  14964=>"001111110",
  14965=>"010100000",
  14966=>"011100001",
  14967=>"001100000",
  14968=>"001111010",
  14969=>"010101101",
  14970=>"110011010",
  14971=>"010111001",
  14972=>"100100010",
  14973=>"000011001",
  14974=>"001001111",
  14975=>"110011111",
  14976=>"100001001",
  14977=>"001001110",
  14978=>"111001001",
  14979=>"101001001",
  14980=>"011100000",
  14981=>"011100010",
  14982=>"001101010",
  14983=>"101001010",
  14984=>"000110001",
  14985=>"100011010",
  14986=>"111100110",
  14987=>"111110001",
  14988=>"101111111",
  14989=>"011110111",
  14990=>"001000000",
  14991=>"000111000",
  14992=>"111001000",
  14993=>"000000111",
  14994=>"001000001",
  14995=>"011001001",
  14996=>"000110101",
  14997=>"000001111",
  14998=>"100101010",
  14999=>"100011110",
  15000=>"000110010",
  15001=>"001100010",
  15002=>"100111000",
  15003=>"101000111",
  15004=>"001000000",
  15005=>"010100000",
  15006=>"001001100",
  15007=>"011100101",
  15008=>"100101011",
  15009=>"110111011",
  15010=>"011010101",
  15011=>"111000100",
  15012=>"010000011",
  15013=>"110101011",
  15014=>"100011000",
  15015=>"101101111",
  15016=>"011100010",
  15017=>"111011001",
  15018=>"010000010",
  15019=>"111011111",
  15020=>"101000111",
  15021=>"101010111",
  15022=>"110000010",
  15023=>"101000101",
  15024=>"010100011",
  15025=>"101001100",
  15026=>"101001100",
  15027=>"100110001",
  15028=>"011000010",
  15029=>"111110110",
  15030=>"001010100",
  15031=>"011111100",
  15032=>"001010011",
  15033=>"000001111",
  15034=>"110011011",
  15035=>"101100110",
  15036=>"001010111",
  15037=>"000101011",
  15038=>"100111100",
  15039=>"101000101",
  15040=>"011100111",
  15041=>"101101111",
  15042=>"110110111",
  15043=>"101111101",
  15044=>"001001111",
  15045=>"011000001",
  15046=>"101100101",
  15047=>"010010010",
  15048=>"010001100",
  15049=>"011001101",
  15050=>"110001011",
  15051=>"111000101",
  15052=>"000101000",
  15053=>"100110100",
  15054=>"110000000",
  15055=>"111011101",
  15056=>"100100101",
  15057=>"011111111",
  15058=>"000011011",
  15059=>"101010110",
  15060=>"100100101",
  15061=>"011011000",
  15062=>"100000010",
  15063=>"001000111",
  15064=>"111111011",
  15065=>"100111000",
  15066=>"001100111",
  15067=>"101100110",
  15068=>"100000110",
  15069=>"101111110",
  15070=>"000000101",
  15071=>"010010001",
  15072=>"110101001",
  15073=>"010000101",
  15074=>"011101110",
  15075=>"100100101",
  15076=>"001111001",
  15077=>"111011011",
  15078=>"111011111",
  15079=>"111110110",
  15080=>"010100111",
  15081=>"111011100",
  15082=>"110011000",
  15083=>"110111010",
  15084=>"011000110",
  15085=>"100011001",
  15086=>"001111101",
  15087=>"000110000",
  15088=>"011100110",
  15089=>"010000110",
  15090=>"111000111",
  15091=>"100011100",
  15092=>"001001111",
  15093=>"101100001",
  15094=>"101101001",
  15095=>"000100001",
  15096=>"010001011",
  15097=>"100010101",
  15098=>"111000110",
  15099=>"100010000",
  15100=>"101100101",
  15101=>"001011101",
  15102=>"000011100",
  15103=>"101100111",
  15104=>"111101101",
  15105=>"000100000",
  15106=>"100011010",
  15107=>"110011001",
  15108=>"010000010",
  15109=>"101111001",
  15110=>"111110100",
  15111=>"111110111",
  15112=>"101001110",
  15113=>"110010001",
  15114=>"100101111",
  15115=>"000101011",
  15116=>"011101110",
  15117=>"101111010",
  15118=>"101000101",
  15119=>"001110101",
  15120=>"100010110",
  15121=>"110110111",
  15122=>"001100001",
  15123=>"101011101",
  15124=>"011100101",
  15125=>"011010111",
  15126=>"001111001",
  15127=>"111010101",
  15128=>"001000110",
  15129=>"100101001",
  15130=>"111110101",
  15131=>"000110111",
  15132=>"000000001",
  15133=>"010110110",
  15134=>"111110111",
  15135=>"000110111",
  15136=>"000001000",
  15137=>"011101000",
  15138=>"111110101",
  15139=>"000000000",
  15140=>"111001100",
  15141=>"111010001",
  15142=>"000100110",
  15143=>"011111111",
  15144=>"011101110",
  15145=>"110100011",
  15146=>"010100110",
  15147=>"000011000",
  15148=>"100000110",
  15149=>"110101011",
  15150=>"111001001",
  15151=>"010110110",
  15152=>"111011000",
  15153=>"110101111",
  15154=>"010001010",
  15155=>"010000001",
  15156=>"010010011",
  15157=>"000010010",
  15158=>"010001010",
  15159=>"101111111",
  15160=>"100110111",
  15161=>"000100101",
  15162=>"010001110",
  15163=>"101100111",
  15164=>"000000110",
  15165=>"001111011",
  15166=>"111101101",
  15167=>"100001100",
  15168=>"000101110",
  15169=>"000011100",
  15170=>"101011100",
  15171=>"001001101",
  15172=>"001101111",
  15173=>"100110000",
  15174=>"100111100",
  15175=>"010001111",
  15176=>"111001111",
  15177=>"100011110",
  15178=>"000010110",
  15179=>"000001111",
  15180=>"101101101",
  15181=>"010001110",
  15182=>"110011000",
  15183=>"100111001",
  15184=>"000111100",
  15185=>"011100111",
  15186=>"010110111",
  15187=>"011011000",
  15188=>"000011001",
  15189=>"010000001",
  15190=>"010000100",
  15191=>"011110001",
  15192=>"000011110",
  15193=>"110100010",
  15194=>"111101111",
  15195=>"101000101",
  15196=>"100110011",
  15197=>"010100100",
  15198=>"001101111",
  15199=>"100000000",
  15200=>"001011110",
  15201=>"100111111",
  15202=>"111011000",
  15203=>"111100100",
  15204=>"000011011",
  15205=>"110100111",
  15206=>"110101101",
  15207=>"010010000",
  15208=>"111001101",
  15209=>"100110100",
  15210=>"001000000",
  15211=>"011010001",
  15212=>"001001011",
  15213=>"110000111",
  15214=>"111101111",
  15215=>"100100101",
  15216=>"010000000",
  15217=>"011110100",
  15218=>"001001010",
  15219=>"000111010",
  15220=>"010100111",
  15221=>"111001000",
  15222=>"001010101",
  15223=>"011101111",
  15224=>"011000110",
  15225=>"111111110",
  15226=>"100010000",
  15227=>"110011110",
  15228=>"011001101",
  15229=>"010001101",
  15230=>"100011010",
  15231=>"011010001",
  15232=>"100111110",
  15233=>"111111111",
  15234=>"000010010",
  15235=>"100000111",
  15236=>"001100011",
  15237=>"011111000",
  15238=>"110100110",
  15239=>"001010010",
  15240=>"100101001",
  15241=>"010001001",
  15242=>"011101001",
  15243=>"111111101",
  15244=>"000000010",
  15245=>"011000100",
  15246=>"111110001",
  15247=>"111100011",
  15248=>"100110011",
  15249=>"001101110",
  15250=>"100100101",
  15251=>"110101110",
  15252=>"001110100",
  15253=>"010011100",
  15254=>"100100111",
  15255=>"111011100",
  15256=>"001100111",
  15257=>"101101011",
  15258=>"110010111",
  15259=>"110110000",
  15260=>"000100101",
  15261=>"111000111",
  15262=>"000100011",
  15263=>"100000001",
  15264=>"110001110",
  15265=>"101100000",
  15266=>"010000011",
  15267=>"010000011",
  15268=>"100011100",
  15269=>"111010000",
  15270=>"000110000",
  15271=>"110011110",
  15272=>"000001111",
  15273=>"101110101",
  15274=>"111011000",
  15275=>"011010101",
  15276=>"111011000",
  15277=>"011100100",
  15278=>"010100101",
  15279=>"010000101",
  15280=>"100111010",
  15281=>"111101001",
  15282=>"011001100",
  15283=>"010001101",
  15284=>"101000101",
  15285=>"001111101",
  15286=>"111111001",
  15287=>"110110010",
  15288=>"000111111",
  15289=>"011001000",
  15290=>"111111100",
  15291=>"001110010",
  15292=>"000100111",
  15293=>"011110000",
  15294=>"100100100",
  15295=>"001100100",
  15296=>"010100101",
  15297=>"010000001",
  15298=>"001011000",
  15299=>"001101110",
  15300=>"111010010",
  15301=>"101100001",
  15302=>"000110000",
  15303=>"110110000",
  15304=>"010110101",
  15305=>"110111100",
  15306=>"011111010",
  15307=>"010100001",
  15308=>"110011110",
  15309=>"001101000",
  15310=>"100000100",
  15311=>"100000010",
  15312=>"010111101",
  15313=>"000100101",
  15314=>"011001110",
  15315=>"100100001",
  15316=>"011000001",
  15317=>"100100011",
  15318=>"101011010",
  15319=>"111111111",
  15320=>"101101111",
  15321=>"111111111",
  15322=>"110010101",
  15323=>"011110000",
  15324=>"000010110",
  15325=>"000010101",
  15326=>"111111000",
  15327=>"011011111",
  15328=>"100110110",
  15329=>"011000111",
  15330=>"100111111",
  15331=>"101100011",
  15332=>"000010011",
  15333=>"111101001",
  15334=>"000111011",
  15335=>"010000101",
  15336=>"011111110",
  15337=>"011011101",
  15338=>"010100000",
  15339=>"001101000",
  15340=>"011001100",
  15341=>"011001101",
  15342=>"001010000",
  15343=>"111111011",
  15344=>"010100010",
  15345=>"100011000",
  15346=>"101011110",
  15347=>"001000011",
  15348=>"010011000",
  15349=>"011100111",
  15350=>"101111110",
  15351=>"001011110",
  15352=>"111010101",
  15353=>"000100010",
  15354=>"011001100",
  15355=>"111100011",
  15356=>"111000100",
  15357=>"011010100",
  15358=>"110100101",
  15359=>"011001011",
  15360=>"001110001",
  15361=>"101111110",
  15362=>"111110000",
  15363=>"100111011",
  15364=>"100011010",
  15365=>"010011011",
  15366=>"110110010",
  15367=>"101111100",
  15368=>"110100001",
  15369=>"000110001",
  15370=>"010001001",
  15371=>"111000101",
  15372=>"001001000",
  15373=>"100111010",
  15374=>"010110111",
  15375=>"111100111",
  15376=>"111010001",
  15377=>"001001100",
  15378=>"101000000",
  15379=>"010100000",
  15380=>"111111000",
  15381=>"010110001",
  15382=>"001011110",
  15383=>"001011101",
  15384=>"111111100",
  15385=>"000011110",
  15386=>"010010000",
  15387=>"010100001",
  15388=>"010000100",
  15389=>"101011000",
  15390=>"101111010",
  15391=>"000001010",
  15392=>"100001010",
  15393=>"111011100",
  15394=>"111111011",
  15395=>"010101011",
  15396=>"000000101",
  15397=>"000001010",
  15398=>"100110001",
  15399=>"110111000",
  15400=>"111100111",
  15401=>"010110001",
  15402=>"000100101",
  15403=>"111101111",
  15404=>"000110111",
  15405=>"011000100",
  15406=>"110101110",
  15407=>"111110010",
  15408=>"001110101",
  15409=>"110011111",
  15410=>"101101011",
  15411=>"100100100",
  15412=>"111000101",
  15413=>"110100110",
  15414=>"000010010",
  15415=>"000010101",
  15416=>"001100101",
  15417=>"011101001",
  15418=>"111100011",
  15419=>"010010000",
  15420=>"101101000",
  15421=>"001010101",
  15422=>"100100100",
  15423=>"111000101",
  15424=>"111011110",
  15425=>"111111011",
  15426=>"110010000",
  15427=>"011010111",
  15428=>"001100001",
  15429=>"000000101",
  15430=>"111001101",
  15431=>"110101110",
  15432=>"000001001",
  15433=>"110001000",
  15434=>"000010000",
  15435=>"001101000",
  15436=>"110100110",
  15437=>"101110011",
  15438=>"000010011",
  15439=>"010010000",
  15440=>"100001000",
  15441=>"000011011",
  15442=>"000000001",
  15443=>"010101011",
  15444=>"100000010",
  15445=>"110110111",
  15446=>"101100101",
  15447=>"001000011",
  15448=>"110110101",
  15449=>"111011000",
  15450=>"101111010",
  15451=>"101110011",
  15452=>"111011000",
  15453=>"101111000",
  15454=>"011001101",
  15455=>"100100110",
  15456=>"010101000",
  15457=>"001011011",
  15458=>"000100001",
  15459=>"010001100",
  15460=>"000100111",
  15461=>"111100111",
  15462=>"001111001",
  15463=>"111011000",
  15464=>"101111101",
  15465=>"111001110",
  15466=>"110010010",
  15467=>"101111100",
  15468=>"111010010",
  15469=>"110010101",
  15470=>"111001101",
  15471=>"010110010",
  15472=>"100111101",
  15473=>"010001110",
  15474=>"100010001",
  15475=>"001111011",
  15476=>"111111110",
  15477=>"000000101",
  15478=>"010001101",
  15479=>"100100111",
  15480=>"111110000",
  15481=>"001100000",
  15482=>"010111001",
  15483=>"101111000",
  15484=>"111111000",
  15485=>"111110111",
  15486=>"011000011",
  15487=>"010101000",
  15488=>"011111011",
  15489=>"010000010",
  15490=>"010000010",
  15491=>"110011001",
  15492=>"100010110",
  15493=>"110100110",
  15494=>"111011010",
  15495=>"011111001",
  15496=>"010010111",
  15497=>"110001111",
  15498=>"011100001",
  15499=>"111101010",
  15500=>"100101100",
  15501=>"101000111",
  15502=>"011010110",
  15503=>"110111001",
  15504=>"010110000",
  15505=>"100100000",
  15506=>"101011010",
  15507=>"010011111",
  15508=>"101101111",
  15509=>"001110110",
  15510=>"001111000",
  15511=>"101001110",
  15512=>"011111100",
  15513=>"011001110",
  15514=>"101111101",
  15515=>"110111010",
  15516=>"011111011",
  15517=>"111001101",
  15518=>"001010010",
  15519=>"001100001",
  15520=>"101010111",
  15521=>"111001111",
  15522=>"010000111",
  15523=>"011100101",
  15524=>"101010011",
  15525=>"110111000",
  15526=>"001001001",
  15527=>"110010110",
  15528=>"111011010",
  15529=>"010101001",
  15530=>"101100101",
  15531=>"011001000",
  15532=>"101001111",
  15533=>"001100001",
  15534=>"000011111",
  15535=>"000110111",
  15536=>"011110111",
  15537=>"101000000",
  15538=>"000000000",
  15539=>"100101101",
  15540=>"010010110",
  15541=>"101011100",
  15542=>"111101101",
  15543=>"011001000",
  15544=>"100001100",
  15545=>"101010111",
  15546=>"011000010",
  15547=>"100010011",
  15548=>"111010111",
  15549=>"001110011",
  15550=>"110010110",
  15551=>"011111111",
  15552=>"111101011",
  15553=>"100010110",
  15554=>"010001001",
  15555=>"010110000",
  15556=>"010110010",
  15557=>"110001010",
  15558=>"001101000",
  15559=>"001110101",
  15560=>"011010000",
  15561=>"100010100",
  15562=>"111111110",
  15563=>"001110011",
  15564=>"100000001",
  15565=>"100101011",
  15566=>"000111111",
  15567=>"100111001",
  15568=>"111010111",
  15569=>"000100001",
  15570=>"111011010",
  15571=>"111000001",
  15572=>"111011100",
  15573=>"110101011",
  15574=>"100001110",
  15575=>"101110001",
  15576=>"010011010",
  15577=>"010110111",
  15578=>"110110110",
  15579=>"111111000",
  15580=>"001111100",
  15581=>"100001101",
  15582=>"010100010",
  15583=>"110011000",
  15584=>"110110100",
  15585=>"100010110",
  15586=>"110111111",
  15587=>"011011101",
  15588=>"000001110",
  15589=>"101001010",
  15590=>"010110101",
  15591=>"000000111",
  15592=>"010101111",
  15593=>"011100110",
  15594=>"010101100",
  15595=>"001100001",
  15596=>"010100000",
  15597=>"111101011",
  15598=>"111110110",
  15599=>"100000001",
  15600=>"111101111",
  15601=>"001100101",
  15602=>"111011110",
  15603=>"000110100",
  15604=>"010010100",
  15605=>"101110101",
  15606=>"010110111",
  15607=>"000011101",
  15608=>"010111011",
  15609=>"011100010",
  15610=>"111110101",
  15611=>"111101010",
  15612=>"111111010",
  15613=>"000101111",
  15614=>"010011001",
  15615=>"111110010",
  15616=>"000010111",
  15617=>"001110100",
  15618=>"101100011",
  15619=>"101101111",
  15620=>"011100011",
  15621=>"111110001",
  15622=>"011101100",
  15623=>"001101101",
  15624=>"111100000",
  15625=>"101101010",
  15626=>"010010011",
  15627=>"110011110",
  15628=>"101111111",
  15629=>"101110010",
  15630=>"000011001",
  15631=>"100010110",
  15632=>"101010000",
  15633=>"110100000",
  15634=>"100100100",
  15635=>"001011001",
  15636=>"010101000",
  15637=>"000111010",
  15638=>"111111111",
  15639=>"111010110",
  15640=>"110100110",
  15641=>"100111010",
  15642=>"110001101",
  15643=>"000011101",
  15644=>"001111101",
  15645=>"000001000",
  15646=>"101011010",
  15647=>"010100011",
  15648=>"110010101",
  15649=>"111101110",
  15650=>"110011011",
  15651=>"101110111",
  15652=>"000000000",
  15653=>"001001011",
  15654=>"010010110",
  15655=>"101100110",
  15656=>"110011000",
  15657=>"111011100",
  15658=>"001101010",
  15659=>"111111011",
  15660=>"111001010",
  15661=>"101011001",
  15662=>"111010001",
  15663=>"101001010",
  15664=>"010111011",
  15665=>"110111110",
  15666=>"110111001",
  15667=>"011010000",
  15668=>"000101110",
  15669=>"100110111",
  15670=>"001000111",
  15671=>"101100010",
  15672=>"011101001",
  15673=>"011100110",
  15674=>"000100110",
  15675=>"100100101",
  15676=>"101000001",
  15677=>"010011010",
  15678=>"010110001",
  15679=>"001010000",
  15680=>"111001101",
  15681=>"111000010",
  15682=>"010010000",
  15683=>"111101110",
  15684=>"000100000",
  15685=>"110001011",
  15686=>"010001100",
  15687=>"000101001",
  15688=>"110101101",
  15689=>"100011110",
  15690=>"010100001",
  15691=>"010001010",
  15692=>"110001110",
  15693=>"111101011",
  15694=>"101110110",
  15695=>"110110011",
  15696=>"100110111",
  15697=>"000110001",
  15698=>"011000111",
  15699=>"111000100",
  15700=>"111000001",
  15701=>"100111001",
  15702=>"101101000",
  15703=>"000100001",
  15704=>"111110101",
  15705=>"011001011",
  15706=>"100111011",
  15707=>"001000111",
  15708=>"101010001",
  15709=>"001011111",
  15710=>"010100101",
  15711=>"001000010",
  15712=>"000001000",
  15713=>"011101001",
  15714=>"000001011",
  15715=>"010101101",
  15716=>"110110110",
  15717=>"010000101",
  15718=>"000110010",
  15719=>"000010000",
  15720=>"001110111",
  15721=>"101100010",
  15722=>"001110011",
  15723=>"110100111",
  15724=>"001101110",
  15725=>"111000111",
  15726=>"100100100",
  15727=>"010000101",
  15728=>"110110111",
  15729=>"111010100",
  15730=>"110000000",
  15731=>"100000111",
  15732=>"001000111",
  15733=>"101101001",
  15734=>"010100010",
  15735=>"010111110",
  15736=>"111111001",
  15737=>"110111100",
  15738=>"110111011",
  15739=>"101010111",
  15740=>"110111101",
  15741=>"100001000",
  15742=>"000100100",
  15743=>"110100001",
  15744=>"010100011",
  15745=>"111010011",
  15746=>"000110011",
  15747=>"010001000",
  15748=>"110101011",
  15749=>"111011100",
  15750=>"001110000",
  15751=>"111000000",
  15752=>"001101000",
  15753=>"000000000",
  15754=>"100000111",
  15755=>"011001000",
  15756=>"100011000",
  15757=>"110011011",
  15758=>"000001000",
  15759=>"100100000",
  15760=>"101001100",
  15761=>"010000010",
  15762=>"011000110",
  15763=>"111010100",
  15764=>"100111000",
  15765=>"101011001",
  15766=>"001001011",
  15767=>"100100100",
  15768=>"100011101",
  15769=>"100001000",
  15770=>"111101111",
  15771=>"011000000",
  15772=>"000011110",
  15773=>"100111111",
  15774=>"000001010",
  15775=>"110101011",
  15776=>"101111111",
  15777=>"100011100",
  15778=>"101011101",
  15779=>"000010110",
  15780=>"101000100",
  15781=>"100110101",
  15782=>"111100001",
  15783=>"101110010",
  15784=>"111001001",
  15785=>"101111111",
  15786=>"111101010",
  15787=>"000011100",
  15788=>"100000010",
  15789=>"001100010",
  15790=>"010001011",
  15791=>"000010101",
  15792=>"101111111",
  15793=>"001001001",
  15794=>"000111111",
  15795=>"000100100",
  15796=>"110101001",
  15797=>"010001111",
  15798=>"111011010",
  15799=>"010100000",
  15800=>"111111111",
  15801=>"011111000",
  15802=>"000011110",
  15803=>"100101010",
  15804=>"000001001",
  15805=>"111011101",
  15806=>"100101110",
  15807=>"001010111",
  15808=>"101011101",
  15809=>"101001111",
  15810=>"101111101",
  15811=>"100010010",
  15812=>"000000110",
  15813=>"110100111",
  15814=>"001101001",
  15815=>"100001100",
  15816=>"000111110",
  15817=>"100111101",
  15818=>"110010111",
  15819=>"011111101",
  15820=>"111111000",
  15821=>"101110110",
  15822=>"000011001",
  15823=>"100110011",
  15824=>"110011000",
  15825=>"110111101",
  15826=>"100110111",
  15827=>"111100010",
  15828=>"000111001",
  15829=>"100100111",
  15830=>"000001100",
  15831=>"010010101",
  15832=>"000101001",
  15833=>"111110101",
  15834=>"011111101",
  15835=>"010100011",
  15836=>"101101011",
  15837=>"001010100",
  15838=>"101000000",
  15839=>"110111100",
  15840=>"011100000",
  15841=>"100010101",
  15842=>"000101010",
  15843=>"100111101",
  15844=>"010010001",
  15845=>"010001011",
  15846=>"111110001",
  15847=>"000000001",
  15848=>"001001000",
  15849=>"111111100",
  15850=>"101110101",
  15851=>"100000011",
  15852=>"010111000",
  15853=>"111000011",
  15854=>"110000011",
  15855=>"000000011",
  15856=>"101101011",
  15857=>"011000000",
  15858=>"110101110",
  15859=>"000110000",
  15860=>"000010100",
  15861=>"011110100",
  15862=>"011101110",
  15863=>"010101001",
  15864=>"010100011",
  15865=>"110010110",
  15866=>"000111010",
  15867=>"000010100",
  15868=>"011011011",
  15869=>"001000100",
  15870=>"110111101",
  15871=>"100001000",
  15872=>"001111101",
  15873=>"000000110",
  15874=>"111101101",
  15875=>"001110101",
  15876=>"011111011",
  15877=>"100111101",
  15878=>"010101000",
  15879=>"111010010",
  15880=>"111100111",
  15881=>"011111101",
  15882=>"001100000",
  15883=>"100110111",
  15884=>"110011010",
  15885=>"100000010",
  15886=>"110011111",
  15887=>"100011000",
  15888=>"000101011",
  15889=>"000011000",
  15890=>"000100011",
  15891=>"110001111",
  15892=>"011001101",
  15893=>"011100011",
  15894=>"110010110",
  15895=>"000010110",
  15896=>"010100010",
  15897=>"100011001",
  15898=>"101100001",
  15899=>"001011101",
  15900=>"000001100",
  15901=>"111110000",
  15902=>"000001110",
  15903=>"111011110",
  15904=>"111111110",
  15905=>"100001110",
  15906=>"001000100",
  15907=>"011000011",
  15908=>"011111111",
  15909=>"110011011",
  15910=>"000111011",
  15911=>"001010000",
  15912=>"000011010",
  15913=>"000000111",
  15914=>"111011011",
  15915=>"101101011",
  15916=>"001101110",
  15917=>"101111010",
  15918=>"011110111",
  15919=>"110010100",
  15920=>"010000000",
  15921=>"000010101",
  15922=>"110101110",
  15923=>"111111111",
  15924=>"011010101",
  15925=>"010110111",
  15926=>"101010110",
  15927=>"011011101",
  15928=>"011001111",
  15929=>"110000001",
  15930=>"001100110",
  15931=>"010111100",
  15932=>"011011011",
  15933=>"010001110",
  15934=>"001000001",
  15935=>"010001001",
  15936=>"110110010",
  15937=>"110000110",
  15938=>"100100010",
  15939=>"001101111",
  15940=>"101001101",
  15941=>"100100001",
  15942=>"001001111",
  15943=>"101111011",
  15944=>"100000100",
  15945=>"010110001",
  15946=>"000101011",
  15947=>"101110100",
  15948=>"111000111",
  15949=>"010010101",
  15950=>"110010000",
  15951=>"000000010",
  15952=>"000011001",
  15953=>"110011110",
  15954=>"011010100",
  15955=>"101010111",
  15956=>"101001011",
  15957=>"101001010",
  15958=>"001100011",
  15959=>"001011110",
  15960=>"110011111",
  15961=>"000100110",
  15962=>"110100001",
  15963=>"001010000",
  15964=>"000010111",
  15965=>"100011011",
  15966=>"100110000",
  15967=>"100001000",
  15968=>"011111101",
  15969=>"001011001",
  15970=>"111110110",
  15971=>"001111101",
  15972=>"100111100",
  15973=>"111011111",
  15974=>"100011100",
  15975=>"010000100",
  15976=>"100110100",
  15977=>"011101000",
  15978=>"101111011",
  15979=>"001100001",
  15980=>"110101000",
  15981=>"001111110",
  15982=>"011100110",
  15983=>"110100110",
  15984=>"110111011",
  15985=>"010111111",
  15986=>"100000111",
  15987=>"110010011",
  15988=>"111111100",
  15989=>"000000101",
  15990=>"011111110",
  15991=>"101111001",
  15992=>"110010010",
  15993=>"100000100",
  15994=>"001001111",
  15995=>"001010110",
  15996=>"100011010",
  15997=>"000010110",
  15998=>"110000000",
  15999=>"110110110",
  16000=>"101100100",
  16001=>"001001001",
  16002=>"101001010",
  16003=>"001000110",
  16004=>"011010100",
  16005=>"111010010",
  16006=>"001011010",
  16007=>"000000000",
  16008=>"100001100",
  16009=>"010110100",
  16010=>"100101100",
  16011=>"011100000",
  16012=>"000110111",
  16013=>"101100100",
  16014=>"111011111",
  16015=>"011001101",
  16016=>"010111110",
  16017=>"000100100",
  16018=>"000001100",
  16019=>"001100100",
  16020=>"100100101",
  16021=>"111001000",
  16022=>"010100111",
  16023=>"011001000",
  16024=>"110010110",
  16025=>"000110101",
  16026=>"000001100",
  16027=>"110101000",
  16028=>"011101100",
  16029=>"000111111",
  16030=>"110100001",
  16031=>"001110010",
  16032=>"111000111",
  16033=>"011000101",
  16034=>"001000110",
  16035=>"010010010",
  16036=>"001010111",
  16037=>"111011000",
  16038=>"001101000",
  16039=>"111011010",
  16040=>"100010000",
  16041=>"100100100",
  16042=>"001010001",
  16043=>"001100100",
  16044=>"000101101",
  16045=>"001100111",
  16046=>"011010110",
  16047=>"001110001",
  16048=>"100100001",
  16049=>"100110010",
  16050=>"111010111",
  16051=>"011101010",
  16052=>"001010100",
  16053=>"010011111",
  16054=>"111110010",
  16055=>"000110110",
  16056=>"111010110",
  16057=>"001001000",
  16058=>"000111110",
  16059=>"101111000",
  16060=>"101101110",
  16061=>"010110001",
  16062=>"101100110",
  16063=>"110101001",
  16064=>"011000000",
  16065=>"111101001",
  16066=>"101110100",
  16067=>"110110010",
  16068=>"101111101",
  16069=>"110000111",
  16070=>"110000111",
  16071=>"111001111",
  16072=>"011000000",
  16073=>"101100010",
  16074=>"010101100",
  16075=>"101111011",
  16076=>"100001100",
  16077=>"000100111",
  16078=>"100100100",
  16079=>"011011110",
  16080=>"100111000",
  16081=>"000010001",
  16082=>"010100001",
  16083=>"010011111",
  16084=>"000010001",
  16085=>"100111100",
  16086=>"000100011",
  16087=>"000111101",
  16088=>"001100111",
  16089=>"111110111",
  16090=>"110011111",
  16091=>"111110100",
  16092=>"101110010",
  16093=>"110000001",
  16094=>"101010011",
  16095=>"000000010",
  16096=>"101001010",
  16097=>"110111101",
  16098=>"110011100",
  16099=>"011010111",
  16100=>"101000110",
  16101=>"001010000",
  16102=>"000000000",
  16103=>"000010101",
  16104=>"011101011",
  16105=>"010110011",
  16106=>"111000000",
  16107=>"100101010",
  16108=>"000111010",
  16109=>"110001001",
  16110=>"010010001",
  16111=>"000011110",
  16112=>"011101110",
  16113=>"111101000",
  16114=>"111111011",
  16115=>"011111110",
  16116=>"010010000",
  16117=>"110111011",
  16118=>"011110101",
  16119=>"011100110",
  16120=>"001010110",
  16121=>"100000111",
  16122=>"100110000",
  16123=>"000010110",
  16124=>"001010000",
  16125=>"110111100",
  16126=>"110111000",
  16127=>"000000000",
  16128=>"001110101",
  16129=>"001011111",
  16130=>"111011000",
  16131=>"010101111",
  16132=>"000100111",
  16133=>"111000000",
  16134=>"010100110",
  16135=>"001010011",
  16136=>"011100000",
  16137=>"000110000",
  16138=>"001011011",
  16139=>"010010011",
  16140=>"001110101",
  16141=>"100010001",
  16142=>"100000111",
  16143=>"111101001",
  16144=>"001000001",
  16145=>"111000101",
  16146=>"000011000",
  16147=>"110010000",
  16148=>"100111100",
  16149=>"110000110",
  16150=>"011110000",
  16151=>"110111001",
  16152=>"111010101",
  16153=>"011010001",
  16154=>"110111010",
  16155=>"100010011",
  16156=>"111011101",
  16157=>"000111011",
  16158=>"011011001",
  16159=>"011100110",
  16160=>"011010010",
  16161=>"111101000",
  16162=>"011111110",
  16163=>"101101001",
  16164=>"010010000",
  16165=>"100011000",
  16166=>"110100101",
  16167=>"001010101",
  16168=>"000101110",
  16169=>"110111110",
  16170=>"100011100",
  16171=>"011100001",
  16172=>"010110111",
  16173=>"101001101",
  16174=>"000000010",
  16175=>"000001100",
  16176=>"110110011",
  16177=>"010011011",
  16178=>"011000100",
  16179=>"010100111",
  16180=>"011100101",
  16181=>"000010000",
  16182=>"101111001",
  16183=>"010001111",
  16184=>"111100010",
  16185=>"000011110",
  16186=>"000000100",
  16187=>"010111000",
  16188=>"110100000",
  16189=>"100111010",
  16190=>"000100100",
  16191=>"111001000",
  16192=>"101011010",
  16193=>"011100011",
  16194=>"111001001",
  16195=>"111011111",
  16196=>"011001011",
  16197=>"111111010",
  16198=>"111010001",
  16199=>"001001111",
  16200=>"100100011",
  16201=>"100010111",
  16202=>"000101011",
  16203=>"011100010",
  16204=>"111010110",
  16205=>"111011110",
  16206=>"100101000",
  16207=>"001011100",
  16208=>"111110000",
  16209=>"010010101",
  16210=>"000110000",
  16211=>"001110111",
  16212=>"101101010",
  16213=>"010011001",
  16214=>"111000001",
  16215=>"111011011",
  16216=>"001000111",
  16217=>"010010110",
  16218=>"101110000",
  16219=>"101011000",
  16220=>"000011011",
  16221=>"010111011",
  16222=>"111101110",
  16223=>"010101010",
  16224=>"110100110",
  16225=>"010110100",
  16226=>"110111110",
  16227=>"001111101",
  16228=>"011111100",
  16229=>"000000101",
  16230=>"010111110",
  16231=>"110010111",
  16232=>"001000110",
  16233=>"011011000",
  16234=>"000001000",
  16235=>"001010001",
  16236=>"001101111",
  16237=>"010111111",
  16238=>"000111101",
  16239=>"101111010",
  16240=>"001000010",
  16241=>"100110000",
  16242=>"001110011",
  16243=>"010101001",
  16244=>"111110101",
  16245=>"010110010",
  16246=>"011101011",
  16247=>"000011000",
  16248=>"101100010",
  16249=>"001101101",
  16250=>"011011111",
  16251=>"011111000",
  16252=>"010000011",
  16253=>"110001011",
  16254=>"000101110",
  16255=>"011100111",
  16256=>"111110010",
  16257=>"100010101",
  16258=>"011101110",
  16259=>"011101000",
  16260=>"000110001",
  16261=>"010001110",
  16262=>"000000010",
  16263=>"100011011",
  16264=>"111001100",
  16265=>"000110100",
  16266=>"100001101",
  16267=>"010100000",
  16268=>"000011100",
  16269=>"010011110",
  16270=>"101000000",
  16271=>"001111001",
  16272=>"101000100",
  16273=>"101010111",
  16274=>"101010111",
  16275=>"110010111",
  16276=>"110000111",
  16277=>"101100101",
  16278=>"000101000",
  16279=>"011110111",
  16280=>"010011101",
  16281=>"100101100",
  16282=>"001110110",
  16283=>"011111111",
  16284=>"011001000",
  16285=>"010001110",
  16286=>"000001000",
  16287=>"111010010",
  16288=>"000010001",
  16289=>"101000000",
  16290=>"101101101",
  16291=>"111100111",
  16292=>"000110000",
  16293=>"000111101",
  16294=>"111010100",
  16295=>"101101011",
  16296=>"001111111",
  16297=>"000010100",
  16298=>"100011111",
  16299=>"110011010",
  16300=>"011100010",
  16301=>"100100000",
  16302=>"000101001",
  16303=>"000011001",
  16304=>"011101110",
  16305=>"000001000",
  16306=>"111011110",
  16307=>"011000110",
  16308=>"100101110",
  16309=>"100110111",
  16310=>"001111011",
  16311=>"000101100",
  16312=>"011110001",
  16313=>"010111001",
  16314=>"011100011",
  16315=>"111101100",
  16316=>"101101111",
  16317=>"001101001",
  16318=>"111001110",
  16319=>"110010100",
  16320=>"010001000",
  16321=>"110101111",
  16322=>"001001000",
  16323=>"000101110",
  16324=>"101111000",
  16325=>"111110100",
  16326=>"101010000",
  16327=>"100001010",
  16328=>"010000001",
  16329=>"011110100",
  16330=>"011110000",
  16331=>"011011100",
  16332=>"100010011",
  16333=>"000010100",
  16334=>"111010000",
  16335=>"110011101",
  16336=>"110011111",
  16337=>"010111010",
  16338=>"111110001",
  16339=>"100011101",
  16340=>"000000101",
  16341=>"000100001",
  16342=>"100000110",
  16343=>"000001110",
  16344=>"000111100",
  16345=>"110101011",
  16346=>"101110010",
  16347=>"111111011",
  16348=>"101000110",
  16349=>"010010101",
  16350=>"101011111",
  16351=>"110010101",
  16352=>"011111100",
  16353=>"100111101",
  16354=>"010110010",
  16355=>"110101111",
  16356=>"111101000",
  16357=>"011101001",
  16358=>"100110101",
  16359=>"110011101",
  16360=>"111011111",
  16361=>"111001101",
  16362=>"000110101",
  16363=>"010011011",
  16364=>"110000011",
  16365=>"101101111",
  16366=>"101011011",
  16367=>"000111000",
  16368=>"011111001",
  16369=>"011010001",
  16370=>"001111111",
  16371=>"111111000",
  16372=>"110100100",
  16373=>"110101111",
  16374=>"110001010",
  16375=>"010010110",
  16376=>"001101111",
  16377=>"111000000",
  16378=>"100001001",
  16379=>"101011111",
  16380=>"101000111",
  16381=>"010010010",
  16382=>"000010110",
  16383=>"111100111",
  16384=>"110010101",
  16385=>"011101111",
  16386=>"011101010",
  16387=>"001111001",
  16388=>"010101110",
  16389=>"100001101",
  16390=>"000010010",
  16391=>"010110110",
  16392=>"100010001",
  16393=>"101000010",
  16394=>"101001001",
  16395=>"110010011",
  16396=>"110000001",
  16397=>"110111110",
  16398=>"000101000",
  16399=>"000011101",
  16400=>"110010110",
  16401=>"100110110",
  16402=>"101011001",
  16403=>"111111001",
  16404=>"000000100",
  16405=>"100010100",
  16406=>"001001110",
  16407=>"100001100",
  16408=>"111111111",
  16409=>"110100000",
  16410=>"111001110",
  16411=>"000111010",
  16412=>"010010011",
  16413=>"011100000",
  16414=>"000000010",
  16415=>"101000100",
  16416=>"101010011",
  16417=>"000100111",
  16418=>"011011100",
  16419=>"011010100",
  16420=>"001111011",
  16421=>"110100100",
  16422=>"000011011",
  16423=>"011010011",
  16424=>"111011111",
  16425=>"000011000",
  16426=>"000101101",
  16427=>"100110001",
  16428=>"011110000",
  16429=>"000110000",
  16430=>"001110000",
  16431=>"010010110",
  16432=>"000011010",
  16433=>"000101000",
  16434=>"111111111",
  16435=>"011001100",
  16436=>"010010100",
  16437=>"011100011",
  16438=>"111000110",
  16439=>"001000010",
  16440=>"001010001",
  16441=>"001001111",
  16442=>"110011001",
  16443=>"000111000",
  16444=>"100011110",
  16445=>"110000111",
  16446=>"000011100",
  16447=>"000000001",
  16448=>"000010100",
  16449=>"100000110",
  16450=>"000101011",
  16451=>"100100010",
  16452=>"111100111",
  16453=>"111101001",
  16454=>"100101100",
  16455=>"000111110",
  16456=>"101101001",
  16457=>"101101010",
  16458=>"110000010",
  16459=>"011010011",
  16460=>"110001111",
  16461=>"101011101",
  16462=>"111110110",
  16463=>"001110000",
  16464=>"100100000",
  16465=>"100010010",
  16466=>"010110101",
  16467=>"001101110",
  16468=>"110110100",
  16469=>"101110111",
  16470=>"010101111",
  16471=>"100110011",
  16472=>"110100001",
  16473=>"101101101",
  16474=>"110011011",
  16475=>"110001110",
  16476=>"100011110",
  16477=>"000010101",
  16478=>"000100000",
  16479=>"001001001",
  16480=>"010000010",
  16481=>"100111110",
  16482=>"011001010",
  16483=>"110010000",
  16484=>"010001000",
  16485=>"011011111",
  16486=>"011011100",
  16487=>"000110000",
  16488=>"101100101",
  16489=>"101101010",
  16490=>"000110001",
  16491=>"010001101",
  16492=>"000010111",
  16493=>"101000111",
  16494=>"110111001",
  16495=>"001001101",
  16496=>"000111010",
  16497=>"000010000",
  16498=>"000100111",
  16499=>"000100000",
  16500=>"000011000",
  16501=>"011110100",
  16502=>"000111010",
  16503=>"010101000",
  16504=>"000010001",
  16505=>"110101110",
  16506=>"111100101",
  16507=>"101110100",
  16508=>"000000100",
  16509=>"011000111",
  16510=>"010101100",
  16511=>"000011101",
  16512=>"011110101",
  16513=>"111101001",
  16514=>"101100000",
  16515=>"101100100",
  16516=>"110010010",
  16517=>"001001000",
  16518=>"110010111",
  16519=>"110010011",
  16520=>"111100001",
  16521=>"010010010",
  16522=>"111100010",
  16523=>"001000101",
  16524=>"010010110",
  16525=>"001001110",
  16526=>"000000010",
  16527=>"111001100",
  16528=>"011010010",
  16529=>"110010001",
  16530=>"000100000",
  16531=>"111100101",
  16532=>"110101000",
  16533=>"010111010",
  16534=>"000101100",
  16535=>"111000101",
  16536=>"000111011",
  16537=>"000010111",
  16538=>"001101010",
  16539=>"110101101",
  16540=>"000001110",
  16541=>"001000011",
  16542=>"101111000",
  16543=>"000111101",
  16544=>"011100110",
  16545=>"111100100",
  16546=>"110110001",
  16547=>"000011000",
  16548=>"010110101",
  16549=>"101100011",
  16550=>"110100111",
  16551=>"000001001",
  16552=>"011111101",
  16553=>"111101110",
  16554=>"000010101",
  16555=>"001101110",
  16556=>"101100110",
  16557=>"011100111",
  16558=>"001001000",
  16559=>"110010101",
  16560=>"111001110",
  16561=>"111001000",
  16562=>"000000101",
  16563=>"010011110",
  16564=>"110101000",
  16565=>"111111100",
  16566=>"100100101",
  16567=>"100110100",
  16568=>"101100010",
  16569=>"000000001",
  16570=>"010010110",
  16571=>"111101101",
  16572=>"000011110",
  16573=>"000110111",
  16574=>"011001100",
  16575=>"000011110",
  16576=>"001001000",
  16577=>"100101101",
  16578=>"110101000",
  16579=>"010101100",
  16580=>"111010100",
  16581=>"001010111",
  16582=>"010111011",
  16583=>"000100001",
  16584=>"110100110",
  16585=>"001011001",
  16586=>"111101001",
  16587=>"010000100",
  16588=>"111111010",
  16589=>"101010011",
  16590=>"010100001",
  16591=>"011001011",
  16592=>"011101000",
  16593=>"100111100",
  16594=>"001000111",
  16595=>"101000110",
  16596=>"110101110",
  16597=>"101010111",
  16598=>"101101000",
  16599=>"011101110",
  16600=>"010010111",
  16601=>"100101001",
  16602=>"011001011",
  16603=>"111000001",
  16604=>"011011001",
  16605=>"011010000",
  16606=>"101100000",
  16607=>"000110100",
  16608=>"111110011",
  16609=>"010110000",
  16610=>"101010101",
  16611=>"011000100",
  16612=>"110100101",
  16613=>"010001000",
  16614=>"000000100",
  16615=>"101110111",
  16616=>"100100011",
  16617=>"100101001",
  16618=>"000110000",
  16619=>"011010111",
  16620=>"110110101",
  16621=>"001010001",
  16622=>"101100100",
  16623=>"111010000",
  16624=>"100011011",
  16625=>"100001110",
  16626=>"110000001",
  16627=>"110110001",
  16628=>"111001111",
  16629=>"111000101",
  16630=>"110001010",
  16631=>"111110001",
  16632=>"000000000",
  16633=>"111010001",
  16634=>"111111100",
  16635=>"000011111",
  16636=>"100110011",
  16637=>"100101000",
  16638=>"100111010",
  16639=>"010100001",
  16640=>"111111100",
  16641=>"001001010",
  16642=>"110111110",
  16643=>"100111000",
  16644=>"111010000",
  16645=>"101101111",
  16646=>"000001101",
  16647=>"001101011",
  16648=>"001010000",
  16649=>"010001110",
  16650=>"100111101",
  16651=>"010100111",
  16652=>"101001001",
  16653=>"000001010",
  16654=>"111111011",
  16655=>"001001010",
  16656=>"001000110",
  16657=>"110011100",
  16658=>"111100011",
  16659=>"000001101",
  16660=>"101011010",
  16661=>"110000000",
  16662=>"001000110",
  16663=>"011011111",
  16664=>"101100101",
  16665=>"110111111",
  16666=>"111010101",
  16667=>"101001111",
  16668=>"010010000",
  16669=>"100101001",
  16670=>"111001100",
  16671=>"110100100",
  16672=>"100011001",
  16673=>"111100111",
  16674=>"110000010",
  16675=>"100100100",
  16676=>"111110101",
  16677=>"000011010",
  16678=>"110110011",
  16679=>"110101011",
  16680=>"111001001",
  16681=>"011000101",
  16682=>"101110010",
  16683=>"100011011",
  16684=>"000110110",
  16685=>"001001000",
  16686=>"100100111",
  16687=>"111110010",
  16688=>"001111000",
  16689=>"000111101",
  16690=>"100100000",
  16691=>"000111001",
  16692=>"001001111",
  16693=>"010011011",
  16694=>"101101000",
  16695=>"111100111",
  16696=>"000000000",
  16697=>"110001110",
  16698=>"100001001",
  16699=>"001110010",
  16700=>"000110000",
  16701=>"110111000",
  16702=>"001111010",
  16703=>"001000100",
  16704=>"000100101",
  16705=>"000000111",
  16706=>"011001010",
  16707=>"110011001",
  16708=>"111100100",
  16709=>"000100010",
  16710=>"010001110",
  16711=>"000001011",
  16712=>"110111010",
  16713=>"011001010",
  16714=>"010101111",
  16715=>"110111000",
  16716=>"111111111",
  16717=>"001000110",
  16718=>"101101100",
  16719=>"101011110",
  16720=>"101101010",
  16721=>"001000010",
  16722=>"011001000",
  16723=>"000100111",
  16724=>"010011001",
  16725=>"011110010",
  16726=>"101010010",
  16727=>"001011001",
  16728=>"000111011",
  16729=>"000100110",
  16730=>"011001011",
  16731=>"001100101",
  16732=>"011100001",
  16733=>"110100101",
  16734=>"111011111",
  16735=>"100111001",
  16736=>"011001001",
  16737=>"110001001",
  16738=>"100111110",
  16739=>"011100101",
  16740=>"011000000",
  16741=>"101001111",
  16742=>"010100010",
  16743=>"110110101",
  16744=>"111001010",
  16745=>"101010100",
  16746=>"111110011",
  16747=>"000010101",
  16748=>"100100011",
  16749=>"000100110",
  16750=>"001011011",
  16751=>"100001011",
  16752=>"100111001",
  16753=>"011000011",
  16754=>"110100110",
  16755=>"010010100",
  16756=>"001011101",
  16757=>"001110001",
  16758=>"000100101",
  16759=>"010000100",
  16760=>"000000100",
  16761=>"010101110",
  16762=>"101111101",
  16763=>"110000001",
  16764=>"001111001",
  16765=>"111011101",
  16766=>"011011010",
  16767=>"101100101",
  16768=>"001111010",
  16769=>"010110000",
  16770=>"010010000",
  16771=>"010100000",
  16772=>"101111100",
  16773=>"011000101",
  16774=>"010010000",
  16775=>"010001010",
  16776=>"110010100",
  16777=>"011110110",
  16778=>"100001111",
  16779=>"111100011",
  16780=>"111011010",
  16781=>"110100000",
  16782=>"100000000",
  16783=>"111000001",
  16784=>"101000111",
  16785=>"111001101",
  16786=>"100011101",
  16787=>"100101011",
  16788=>"000010101",
  16789=>"000011000",
  16790=>"111100100",
  16791=>"000110010",
  16792=>"000000000",
  16793=>"101000100",
  16794=>"010101110",
  16795=>"100100010",
  16796=>"101100001",
  16797=>"001001101",
  16798=>"111111010",
  16799=>"011110000",
  16800=>"101111011",
  16801=>"100010011",
  16802=>"110010111",
  16803=>"011000101",
  16804=>"111000101",
  16805=>"101000100",
  16806=>"101101100",
  16807=>"101110111",
  16808=>"111101110",
  16809=>"100000011",
  16810=>"011010011",
  16811=>"001100010",
  16812=>"001100100",
  16813=>"011110001",
  16814=>"101111100",
  16815=>"111000010",
  16816=>"000100001",
  16817=>"010110101",
  16818=>"010111111",
  16819=>"000100001",
  16820=>"111001110",
  16821=>"111101100",
  16822=>"010011100",
  16823=>"011000011",
  16824=>"100000111",
  16825=>"011001000",
  16826=>"000001100",
  16827=>"000001110",
  16828=>"100011110",
  16829=>"100001011",
  16830=>"000111011",
  16831=>"100001000",
  16832=>"000011100",
  16833=>"000010100",
  16834=>"001000100",
  16835=>"011101011",
  16836=>"100111000",
  16837=>"111101110",
  16838=>"100000100",
  16839=>"101110010",
  16840=>"000010000",
  16841=>"001010000",
  16842=>"101110000",
  16843=>"111001011",
  16844=>"010110100",
  16845=>"110001100",
  16846=>"011011011",
  16847=>"001000001",
  16848=>"001010110",
  16849=>"000010000",
  16850=>"101101000",
  16851=>"001101011",
  16852=>"000101011",
  16853=>"111110110",
  16854=>"100101111",
  16855=>"011001001",
  16856=>"000000101",
  16857=>"010111100",
  16858=>"100110010",
  16859=>"100011110",
  16860=>"110110001",
  16861=>"100010011",
  16862=>"011101110",
  16863=>"110111000",
  16864=>"101011010",
  16865=>"000011100",
  16866=>"100001010",
  16867=>"101000111",
  16868=>"111000001",
  16869=>"011000000",
  16870=>"010110001",
  16871=>"110101011",
  16872=>"000001000",
  16873=>"000110101",
  16874=>"001101100",
  16875=>"010000100",
  16876=>"101110001",
  16877=>"001000010",
  16878=>"111000011",
  16879=>"100101010",
  16880=>"111001100",
  16881=>"010101010",
  16882=>"101110110",
  16883=>"011101000",
  16884=>"111110101",
  16885=>"001000111",
  16886=>"010000001",
  16887=>"000011011",
  16888=>"101101001",
  16889=>"011010111",
  16890=>"001110110",
  16891=>"001101110",
  16892=>"001010001",
  16893=>"111011110",
  16894=>"000010001",
  16895=>"111001111",
  16896=>"011101101",
  16897=>"100000011",
  16898=>"110010110",
  16899=>"001100000",
  16900=>"101011111",
  16901=>"010010000",
  16902=>"110110111",
  16903=>"001011101",
  16904=>"111010101",
  16905=>"100011011",
  16906=>"110010000",
  16907=>"000010010",
  16908=>"100001111",
  16909=>"101000010",
  16910=>"111111000",
  16911=>"100011100",
  16912=>"000011000",
  16913=>"100010101",
  16914=>"010001001",
  16915=>"011100110",
  16916=>"110010010",
  16917=>"001000111",
  16918=>"011111110",
  16919=>"101101101",
  16920=>"000010111",
  16921=>"010111001",
  16922=>"000010001",
  16923=>"001110111",
  16924=>"010110111",
  16925=>"100100110",
  16926=>"001111110",
  16927=>"011111011",
  16928=>"010000111",
  16929=>"011000110",
  16930=>"000010010",
  16931=>"101100111",
  16932=>"100111011",
  16933=>"001001111",
  16934=>"001001101",
  16935=>"101110100",
  16936=>"110110101",
  16937=>"101000110",
  16938=>"011001111",
  16939=>"010001111",
  16940=>"111101110",
  16941=>"101011110",
  16942=>"110011001",
  16943=>"011110111",
  16944=>"110111110",
  16945=>"111111101",
  16946=>"010010110",
  16947=>"011001000",
  16948=>"101010001",
  16949=>"110011011",
  16950=>"011000011",
  16951=>"001001001",
  16952=>"001011000",
  16953=>"011110101",
  16954=>"101011011",
  16955=>"000100100",
  16956=>"000110010",
  16957=>"000001110",
  16958=>"110100101",
  16959=>"111100110",
  16960=>"111100011",
  16961=>"110010000",
  16962=>"110110110",
  16963=>"101001010",
  16964=>"011110111",
  16965=>"100000111",
  16966=>"000100101",
  16967=>"101111100",
  16968=>"100110001",
  16969=>"011101001",
  16970=>"110010101",
  16971=>"111110101",
  16972=>"010111110",
  16973=>"010010010",
  16974=>"110100101",
  16975=>"110111111",
  16976=>"110111101",
  16977=>"111010111",
  16978=>"101101111",
  16979=>"111000000",
  16980=>"001100000",
  16981=>"101000000",
  16982=>"110010010",
  16983=>"001000100",
  16984=>"001100011",
  16985=>"111111010",
  16986=>"001111100",
  16987=>"010000011",
  16988=>"011001101",
  16989=>"000000000",
  16990=>"000000010",
  16991=>"111010011",
  16992=>"110010001",
  16993=>"000000000",
  16994=>"110110111",
  16995=>"101000110",
  16996=>"000001010",
  16997=>"111111110",
  16998=>"000011100",
  16999=>"001000001",
  17000=>"000001001",
  17001=>"100100110",
  17002=>"001101011",
  17003=>"110111001",
  17004=>"000000000",
  17005=>"011100011",
  17006=>"000010000",
  17007=>"110110101",
  17008=>"101011000",
  17009=>"011011011",
  17010=>"100111111",
  17011=>"001000100",
  17012=>"100100000",
  17013=>"010101110",
  17014=>"110001001",
  17015=>"000011101",
  17016=>"010100110",
  17017=>"010111110",
  17018=>"011101001",
  17019=>"100100000",
  17020=>"010101111",
  17021=>"110110110",
  17022=>"011111010",
  17023=>"010000011",
  17024=>"001110100",
  17025=>"011111011",
  17026=>"010010100",
  17027=>"000010001",
  17028=>"000000010",
  17029=>"011111101",
  17030=>"101100111",
  17031=>"111101001",
  17032=>"011001110",
  17033=>"101001111",
  17034=>"111011001",
  17035=>"100100010",
  17036=>"010101001",
  17037=>"111110001",
  17038=>"100100101",
  17039=>"000111100",
  17040=>"000000110",
  17041=>"000001011",
  17042=>"111000111",
  17043=>"100110111",
  17044=>"000001000",
  17045=>"111101001",
  17046=>"111101110",
  17047=>"010101000",
  17048=>"111010100",
  17049=>"111111000",
  17050=>"101001011",
  17051=>"010111111",
  17052=>"010011000",
  17053=>"001001010",
  17054=>"111111101",
  17055=>"101011000",
  17056=>"111110110",
  17057=>"111110000",
  17058=>"001111101",
  17059=>"011000101",
  17060=>"110001111",
  17061=>"101001001",
  17062=>"001111111",
  17063=>"000000010",
  17064=>"000001001",
  17065=>"110100000",
  17066=>"011010111",
  17067=>"000101011",
  17068=>"010010110",
  17069=>"001011110",
  17070=>"011111110",
  17071=>"111101111",
  17072=>"000111010",
  17073=>"110011101",
  17074=>"100010011",
  17075=>"011110001",
  17076=>"000100111",
  17077=>"110000110",
  17078=>"111110011",
  17079=>"100101010",
  17080=>"011100000",
  17081=>"010011011",
  17082=>"110110100",
  17083=>"000001101",
  17084=>"001111100",
  17085=>"010001010",
  17086=>"001011100",
  17087=>"000001011",
  17088=>"111000000",
  17089=>"000001110",
  17090=>"111111000",
  17091=>"000101111",
  17092=>"101110010",
  17093=>"100110001",
  17094=>"010010000",
  17095=>"011101100",
  17096=>"101001111",
  17097=>"111101100",
  17098=>"110110110",
  17099=>"101111000",
  17100=>"001100111",
  17101=>"101011111",
  17102=>"100110000",
  17103=>"010000110",
  17104=>"001101001",
  17105=>"000001001",
  17106=>"110010110",
  17107=>"010011010",
  17108=>"001111010",
  17109=>"011110100",
  17110=>"000001101",
  17111=>"000111100",
  17112=>"001010100",
  17113=>"001001011",
  17114=>"001111101",
  17115=>"101110010",
  17116=>"110001101",
  17117=>"110110011",
  17118=>"001100101",
  17119=>"011011011",
  17120=>"010001001",
  17121=>"000011001",
  17122=>"010110011",
  17123=>"101100100",
  17124=>"000001101",
  17125=>"101101001",
  17126=>"001001111",
  17127=>"000011101",
  17128=>"100000000",
  17129=>"011111100",
  17130=>"010001100",
  17131=>"000010000",
  17132=>"001000101",
  17133=>"000110000",
  17134=>"111000101",
  17135=>"110001000",
  17136=>"110001111",
  17137=>"001111001",
  17138=>"001001101",
  17139=>"010001000",
  17140=>"000000110",
  17141=>"000000010",
  17142=>"101101000",
  17143=>"011011011",
  17144=>"111101101",
  17145=>"011101001",
  17146=>"001001100",
  17147=>"010000010",
  17148=>"011100010",
  17149=>"010110101",
  17150=>"011100000",
  17151=>"000110000",
  17152=>"011100000",
  17153=>"010100000",
  17154=>"100011100",
  17155=>"001111110",
  17156=>"110000110",
  17157=>"111000110",
  17158=>"010101100",
  17159=>"101100110",
  17160=>"000001000",
  17161=>"110100000",
  17162=>"100011110",
  17163=>"111011001",
  17164=>"010100001",
  17165=>"001110011",
  17166=>"011010010",
  17167=>"100110010",
  17168=>"011101111",
  17169=>"111100000",
  17170=>"101100101",
  17171=>"100001111",
  17172=>"101101111",
  17173=>"110101111",
  17174=>"001101010",
  17175=>"111100101",
  17176=>"010010110",
  17177=>"001100101",
  17178=>"101100101",
  17179=>"010101000",
  17180=>"010011010",
  17181=>"111100000",
  17182=>"011100010",
  17183=>"110000100",
  17184=>"010111000",
  17185=>"100111110",
  17186=>"011101011",
  17187=>"010100110",
  17188=>"101010111",
  17189=>"101100111",
  17190=>"001110101",
  17191=>"110001010",
  17192=>"000100010",
  17193=>"101011001",
  17194=>"100111100",
  17195=>"101000000",
  17196=>"110101010",
  17197=>"000001101",
  17198=>"000100111",
  17199=>"000110100",
  17200=>"010100110",
  17201=>"101100110",
  17202=>"000100011",
  17203=>"010101010",
  17204=>"110001011",
  17205=>"000101100",
  17206=>"101111011",
  17207=>"001010001",
  17208=>"000101011",
  17209=>"111110111",
  17210=>"011011001",
  17211=>"111011110",
  17212=>"011101100",
  17213=>"011000101",
  17214=>"100011100",
  17215=>"011111111",
  17216=>"011011001",
  17217=>"011000111",
  17218=>"010011001",
  17219=>"011110100",
  17220=>"100110110",
  17221=>"101100100",
  17222=>"110001111",
  17223=>"011001100",
  17224=>"111011101",
  17225=>"000110110",
  17226=>"110010100",
  17227=>"110100111",
  17228=>"100110011",
  17229=>"101101000",
  17230=>"101110011",
  17231=>"000001011",
  17232=>"111001001",
  17233=>"110001110",
  17234=>"100101011",
  17235=>"011100000",
  17236=>"111100110",
  17237=>"000000011",
  17238=>"001000100",
  17239=>"101101010",
  17240=>"111000100",
  17241=>"010110010",
  17242=>"000101111",
  17243=>"000010000",
  17244=>"011110110",
  17245=>"100001100",
  17246=>"110000000",
  17247=>"000000100",
  17248=>"001111000",
  17249=>"101111111",
  17250=>"000000100",
  17251=>"001011001",
  17252=>"011001100",
  17253=>"000001011",
  17254=>"001111100",
  17255=>"101010010",
  17256=>"010100001",
  17257=>"100001111",
  17258=>"110000001",
  17259=>"011100010",
  17260=>"110011111",
  17261=>"011000010",
  17262=>"111111011",
  17263=>"001110001",
  17264=>"110111000",
  17265=>"111001011",
  17266=>"111100000",
  17267=>"100001101",
  17268=>"001000000",
  17269=>"000000111",
  17270=>"101010011",
  17271=>"101010000",
  17272=>"110001000",
  17273=>"101000001",
  17274=>"101011101",
  17275=>"101110011",
  17276=>"000000000",
  17277=>"010101000",
  17278=>"111000001",
  17279=>"101000000",
  17280=>"001111010",
  17281=>"111000110",
  17282=>"010001010",
  17283=>"000111100",
  17284=>"000000000",
  17285=>"000101100",
  17286=>"000110111",
  17287=>"101000010",
  17288=>"001101110",
  17289=>"111000001",
  17290=>"010101110",
  17291=>"010000000",
  17292=>"100001101",
  17293=>"111110010",
  17294=>"110110100",
  17295=>"001101111",
  17296=>"100101000",
  17297=>"110101100",
  17298=>"101001000",
  17299=>"111000010",
  17300=>"111000011",
  17301=>"110000011",
  17302=>"010011011",
  17303=>"010110010",
  17304=>"110011100",
  17305=>"101001111",
  17306=>"010110000",
  17307=>"011001010",
  17308=>"000001100",
  17309=>"111110010",
  17310=>"011100010",
  17311=>"000000111",
  17312=>"111101001",
  17313=>"100110110",
  17314=>"011000100",
  17315=>"000110100",
  17316=>"010100000",
  17317=>"011111111",
  17318=>"000100100",
  17319=>"010001111",
  17320=>"010000010",
  17321=>"000001100",
  17322=>"000110100",
  17323=>"101001010",
  17324=>"011011101",
  17325=>"010110100",
  17326=>"101011110",
  17327=>"101111100",
  17328=>"110001011",
  17329=>"110110111",
  17330=>"001101101",
  17331=>"001010000",
  17332=>"000011010",
  17333=>"101010011",
  17334=>"000100111",
  17335=>"101000010",
  17336=>"001010110",
  17337=>"001101110",
  17338=>"011111110",
  17339=>"010010011",
  17340=>"111111111",
  17341=>"111111011",
  17342=>"111010010",
  17343=>"001111101",
  17344=>"011100111",
  17345=>"010010111",
  17346=>"011001010",
  17347=>"011110101",
  17348=>"100100000",
  17349=>"001101111",
  17350=>"101010001",
  17351=>"110110100",
  17352=>"000011010",
  17353=>"100100100",
  17354=>"010111100",
  17355=>"011100010",
  17356=>"010010111",
  17357=>"000001100",
  17358=>"000000001",
  17359=>"100101001",
  17360=>"110001011",
  17361=>"000110000",
  17362=>"011101001",
  17363=>"001111101",
  17364=>"010011111",
  17365=>"000101101",
  17366=>"100110100",
  17367=>"000001111",
  17368=>"001010001",
  17369=>"101100111",
  17370=>"000011100",
  17371=>"111110011",
  17372=>"100001011",
  17373=>"010101100",
  17374=>"011011000",
  17375=>"000010101",
  17376=>"001100100",
  17377=>"111101110",
  17378=>"010001010",
  17379=>"101111100",
  17380=>"000000000",
  17381=>"011001001",
  17382=>"010111000",
  17383=>"000111100",
  17384=>"010011111",
  17385=>"001001101",
  17386=>"010010001",
  17387=>"000001000",
  17388=>"001010011",
  17389=>"001100100",
  17390=>"011001000",
  17391=>"111111101",
  17392=>"010110111",
  17393=>"010000100",
  17394=>"100100101",
  17395=>"000001001",
  17396=>"010110110",
  17397=>"010011111",
  17398=>"100010110",
  17399=>"000101011",
  17400=>"111101010",
  17401=>"111101110",
  17402=>"101111010",
  17403=>"010100010",
  17404=>"111111000",
  17405=>"011010010",
  17406=>"011001011",
  17407=>"000100011",
  17408=>"101111111",
  17409=>"000000100",
  17410=>"010100010",
  17411=>"000101110",
  17412=>"111011101",
  17413=>"100000000",
  17414=>"000000010",
  17415=>"010101101",
  17416=>"001011000",
  17417=>"000110101",
  17418=>"101000010",
  17419=>"100110110",
  17420=>"100111111",
  17421=>"001111011",
  17422=>"100001010",
  17423=>"100110100",
  17424=>"000110010",
  17425=>"000110100",
  17426=>"010100010",
  17427=>"000001101",
  17428=>"000111110",
  17429=>"000110100",
  17430=>"001010101",
  17431=>"001100010",
  17432=>"110100000",
  17433=>"001000000",
  17434=>"000101101",
  17435=>"101000111",
  17436=>"100011101",
  17437=>"001111010",
  17438=>"101100000",
  17439=>"010000101",
  17440=>"001000101",
  17441=>"011111101",
  17442=>"000110101",
  17443=>"110111000",
  17444=>"111011100",
  17445=>"100111010",
  17446=>"110001101",
  17447=>"111111111",
  17448=>"011011100",
  17449=>"000001110",
  17450=>"000010011",
  17451=>"001111110",
  17452=>"101001001",
  17453=>"000111000",
  17454=>"101010010",
  17455=>"001110001",
  17456=>"100111010",
  17457=>"110011000",
  17458=>"100111101",
  17459=>"111000101",
  17460=>"011111010",
  17461=>"010101110",
  17462=>"010011101",
  17463=>"101110101",
  17464=>"010011001",
  17465=>"001010110",
  17466=>"111011110",
  17467=>"101000001",
  17468=>"010111000",
  17469=>"010000100",
  17470=>"101100111",
  17471=>"000101101",
  17472=>"111111100",
  17473=>"000010111",
  17474=>"100110100",
  17475=>"100010001",
  17476=>"101110001",
  17477=>"101001110",
  17478=>"110111000",
  17479=>"001001011",
  17480=>"000100000",
  17481=>"010011110",
  17482=>"010101101",
  17483=>"001101001",
  17484=>"010100101",
  17485=>"010100010",
  17486=>"101010001",
  17487=>"100110110",
  17488=>"000100010",
  17489=>"100010111",
  17490=>"001101110",
  17491=>"111111010",
  17492=>"110110111",
  17493=>"010111111",
  17494=>"000100000",
  17495=>"111001010",
  17496=>"011010010",
  17497=>"001110101",
  17498=>"101100100",
  17499=>"111110100",
  17500=>"001110110",
  17501=>"110111010",
  17502=>"110000110",
  17503=>"010000001",
  17504=>"110100001",
  17505=>"101100100",
  17506=>"000011000",
  17507=>"000111111",
  17508=>"001101111",
  17509=>"000011011",
  17510=>"000010100",
  17511=>"101000100",
  17512=>"110100010",
  17513=>"000111110",
  17514=>"101100101",
  17515=>"100001010",
  17516=>"100101101",
  17517=>"010111101",
  17518=>"100101101",
  17519=>"000100001",
  17520=>"111011101",
  17521=>"011011100",
  17522=>"010100001",
  17523=>"101101110",
  17524=>"010101111",
  17525=>"001001100",
  17526=>"100111110",
  17527=>"011000001",
  17528=>"001100001",
  17529=>"001011000",
  17530=>"111001100",
  17531=>"000011011",
  17532=>"000001101",
  17533=>"100001001",
  17534=>"000111111",
  17535=>"100110011",
  17536=>"110010101",
  17537=>"011010101",
  17538=>"011001000",
  17539=>"110100110",
  17540=>"000011000",
  17541=>"011101010",
  17542=>"101010010",
  17543=>"110101000",
  17544=>"101000111",
  17545=>"000010100",
  17546=>"011111011",
  17547=>"111000000",
  17548=>"000101011",
  17549=>"111110111",
  17550=>"000001001",
  17551=>"011111011",
  17552=>"110000101",
  17553=>"100110000",
  17554=>"101100000",
  17555=>"101011110",
  17556=>"101100000",
  17557=>"000101010",
  17558=>"000100110",
  17559=>"010111010",
  17560=>"110101001",
  17561=>"111001010",
  17562=>"010111101",
  17563=>"010011100",
  17564=>"010000100",
  17565=>"000111001",
  17566=>"001100111",
  17567=>"111001101",
  17568=>"100110000",
  17569=>"010101110",
  17570=>"010001010",
  17571=>"100100000",
  17572=>"001001111",
  17573=>"000011111",
  17574=>"100000101",
  17575=>"011011000",
  17576=>"000001000",
  17577=>"010111010",
  17578=>"110001111",
  17579=>"110000101",
  17580=>"011101100",
  17581=>"110101100",
  17582=>"101100100",
  17583=>"111111110",
  17584=>"001010000",
  17585=>"001101010",
  17586=>"111010000",
  17587=>"111100011",
  17588=>"000001011",
  17589=>"001010000",
  17590=>"100000111",
  17591=>"101111000",
  17592=>"100110110",
  17593=>"010010111",
  17594=>"110011100",
  17595=>"101101101",
  17596=>"011010111",
  17597=>"001110101",
  17598=>"011100000",
  17599=>"111100001",
  17600=>"000001010",
  17601=>"010100010",
  17602=>"000011101",
  17603=>"110100000",
  17604=>"000111101",
  17605=>"011101011",
  17606=>"101000100",
  17607=>"101010011",
  17608=>"000101010",
  17609=>"001110111",
  17610=>"101010110",
  17611=>"000101100",
  17612=>"101111101",
  17613=>"100010111",
  17614=>"011010110",
  17615=>"010001000",
  17616=>"001001111",
  17617=>"001000100",
  17618=>"111000111",
  17619=>"011110001",
  17620=>"000000100",
  17621=>"001001001",
  17622=>"111000010",
  17623=>"101110111",
  17624=>"000110101",
  17625=>"010000110",
  17626=>"001001011",
  17627=>"010101000",
  17628=>"011000001",
  17629=>"001111000",
  17630=>"001101001",
  17631=>"001111001",
  17632=>"110001111",
  17633=>"101111110",
  17634=>"111011001",
  17635=>"101100010",
  17636=>"110001000",
  17637=>"101000110",
  17638=>"101000110",
  17639=>"011110001",
  17640=>"100110001",
  17641=>"111001101",
  17642=>"100010011",
  17643=>"010010000",
  17644=>"010111010",
  17645=>"111101100",
  17646=>"000010011",
  17647=>"000001101",
  17648=>"110100000",
  17649=>"011101000",
  17650=>"000010001",
  17651=>"000111100",
  17652=>"010110000",
  17653=>"101010110",
  17654=>"001001010",
  17655=>"101001011",
  17656=>"011110000",
  17657=>"111101000",
  17658=>"101000110",
  17659=>"010000001",
  17660=>"011000010",
  17661=>"001000001",
  17662=>"010110111",
  17663=>"011110000",
  17664=>"111110010",
  17665=>"000100011",
  17666=>"010011100",
  17667=>"001010001",
  17668=>"011001100",
  17669=>"001101110",
  17670=>"011111111",
  17671=>"000000010",
  17672=>"010010001",
  17673=>"101011000",
  17674=>"110100101",
  17675=>"000110010",
  17676=>"010010110",
  17677=>"010111011",
  17678=>"100011011",
  17679=>"000100101",
  17680=>"000010111",
  17681=>"101101111",
  17682=>"111110110",
  17683=>"011111000",
  17684=>"111010000",
  17685=>"101010101",
  17686=>"001100001",
  17687=>"111011110",
  17688=>"110100000",
  17689=>"101001011",
  17690=>"110000110",
  17691=>"000001001",
  17692=>"101100000",
  17693=>"010001000",
  17694=>"110111100",
  17695=>"010111111",
  17696=>"100000011",
  17697=>"000111100",
  17698=>"101101111",
  17699=>"110001110",
  17700=>"111011101",
  17701=>"000110100",
  17702=>"111000101",
  17703=>"001110101",
  17704=>"110100111",
  17705=>"010001110",
  17706=>"100000000",
  17707=>"111100100",
  17708=>"101110010",
  17709=>"001001110",
  17710=>"001111110",
  17711=>"010110010",
  17712=>"011100100",
  17713=>"011101101",
  17714=>"000000100",
  17715=>"011001001",
  17716=>"010000000",
  17717=>"110111000",
  17718=>"111101010",
  17719=>"001100111",
  17720=>"110000001",
  17721=>"001011010",
  17722=>"001001010",
  17723=>"011111111",
  17724=>"000001001",
  17725=>"110100111",
  17726=>"111101110",
  17727=>"000110011",
  17728=>"011010111",
  17729=>"010000110",
  17730=>"101110101",
  17731=>"001001001",
  17732=>"110001101",
  17733=>"101100101",
  17734=>"101100110",
  17735=>"010110011",
  17736=>"111101000",
  17737=>"110011010",
  17738=>"001111110",
  17739=>"011111011",
  17740=>"001011101",
  17741=>"000101011",
  17742=>"010000011",
  17743=>"001001010",
  17744=>"110101010",
  17745=>"000100010",
  17746=>"010000111",
  17747=>"010110100",
  17748=>"010111110",
  17749=>"011001000",
  17750=>"111000100",
  17751=>"011101100",
  17752=>"100000000",
  17753=>"110101100",
  17754=>"001000011",
  17755=>"011101011",
  17756=>"010001001",
  17757=>"010100001",
  17758=>"111001100",
  17759=>"101100111",
  17760=>"101011110",
  17761=>"101100000",
  17762=>"100111110",
  17763=>"101000011",
  17764=>"011010111",
  17765=>"001010111",
  17766=>"011000011",
  17767=>"000000010",
  17768=>"111011001",
  17769=>"011000011",
  17770=>"100111111",
  17771=>"010000000",
  17772=>"010101100",
  17773=>"111011110",
  17774=>"011010101",
  17775=>"101100001",
  17776=>"110110100",
  17777=>"011100000",
  17778=>"110011011",
  17779=>"110010101",
  17780=>"001101011",
  17781=>"100111111",
  17782=>"000001010",
  17783=>"111001000",
  17784=>"010100100",
  17785=>"110000011",
  17786=>"111000100",
  17787=>"110010100",
  17788=>"011101100",
  17789=>"001100111",
  17790=>"000101110",
  17791=>"111000011",
  17792=>"110111111",
  17793=>"101011100",
  17794=>"010000010",
  17795=>"010011011",
  17796=>"010011000",
  17797=>"100010110",
  17798=>"110001000",
  17799=>"101011100",
  17800=>"101000111",
  17801=>"111011111",
  17802=>"110010010",
  17803=>"011000011",
  17804=>"100100000",
  17805=>"010010011",
  17806=>"001001010",
  17807=>"000001011",
  17808=>"100110011",
  17809=>"101101101",
  17810=>"011101000",
  17811=>"111001100",
  17812=>"100101001",
  17813=>"010101011",
  17814=>"010011000",
  17815=>"100001110",
  17816=>"000110100",
  17817=>"010001011",
  17818=>"000100010",
  17819=>"000000111",
  17820=>"010000100",
  17821=>"100011111",
  17822=>"010011001",
  17823=>"110100110",
  17824=>"001001100",
  17825=>"000001111",
  17826=>"001100010",
  17827=>"010010101",
  17828=>"101010001",
  17829=>"010101101",
  17830=>"001111100",
  17831=>"001010110",
  17832=>"100000101",
  17833=>"101101011",
  17834=>"000011100",
  17835=>"010010101",
  17836=>"110110001",
  17837=>"100111011",
  17838=>"111011000",
  17839=>"010010001",
  17840=>"001100110",
  17841=>"101011011",
  17842=>"110111111",
  17843=>"010101111",
  17844=>"111111101",
  17845=>"100110111",
  17846=>"000000101",
  17847=>"011111110",
  17848=>"110000011",
  17849=>"100100011",
  17850=>"001101000",
  17851=>"110010000",
  17852=>"010000001",
  17853=>"101110111",
  17854=>"000111010",
  17855=>"000000100",
  17856=>"011011110",
  17857=>"001111001",
  17858=>"111011000",
  17859=>"101101001",
  17860=>"000101100",
  17861=>"111101000",
  17862=>"011000000",
  17863=>"011110010",
  17864=>"000011000",
  17865=>"110011001",
  17866=>"001000000",
  17867=>"000110000",
  17868=>"001110101",
  17869=>"000001111",
  17870=>"000110010",
  17871=>"000111000",
  17872=>"110111111",
  17873=>"010001001",
  17874=>"101011000",
  17875=>"110001011",
  17876=>"001110011",
  17877=>"001010101",
  17878=>"000011110",
  17879=>"101000000",
  17880=>"101110111",
  17881=>"101011001",
  17882=>"011110011",
  17883=>"111110101",
  17884=>"111101010",
  17885=>"000100110",
  17886=>"101001100",
  17887=>"100100011",
  17888=>"000101101",
  17889=>"011000000",
  17890=>"111111111",
  17891=>"010100100",
  17892=>"001010100",
  17893=>"111010101",
  17894=>"000100110",
  17895=>"011101000",
  17896=>"010011110",
  17897=>"011011000",
  17898=>"100010000",
  17899=>"110110101",
  17900=>"001100000",
  17901=>"011110101",
  17902=>"100011000",
  17903=>"001010100",
  17904=>"110111001",
  17905=>"101100101",
  17906=>"010101000",
  17907=>"011010010",
  17908=>"011101111",
  17909=>"101101110",
  17910=>"000110000",
  17911=>"001100000",
  17912=>"010000101",
  17913=>"110001011",
  17914=>"101110110",
  17915=>"001101100",
  17916=>"010100000",
  17917=>"000010011",
  17918=>"011111011",
  17919=>"110010010",
  17920=>"101111111",
  17921=>"010111111",
  17922=>"010011011",
  17923=>"101111011",
  17924=>"110011001",
  17925=>"000100110",
  17926=>"101100100",
  17927=>"101000000",
  17928=>"011001110",
  17929=>"011011010",
  17930=>"000101000",
  17931=>"110000100",
  17932=>"111111001",
  17933=>"100001111",
  17934=>"100101000",
  17935=>"111000011",
  17936=>"011010110",
  17937=>"010100011",
  17938=>"111001101",
  17939=>"111111111",
  17940=>"000110100",
  17941=>"111110011",
  17942=>"101100000",
  17943=>"110001110",
  17944=>"101100111",
  17945=>"110010101",
  17946=>"011010111",
  17947=>"110010110",
  17948=>"001011010",
  17949=>"011011111",
  17950=>"001101110",
  17951=>"111001001",
  17952=>"110000001",
  17953=>"111000011",
  17954=>"100110101",
  17955=>"000000110",
  17956=>"010100100",
  17957=>"010000001",
  17958=>"101010000",
  17959=>"111110011",
  17960=>"110011010",
  17961=>"101111111",
  17962=>"110000010",
  17963=>"100011001",
  17964=>"001011100",
  17965=>"000100000",
  17966=>"000010001",
  17967=>"000010110",
  17968=>"110010111",
  17969=>"111000011",
  17970=>"011011011",
  17971=>"111001001",
  17972=>"100100101",
  17973=>"110111000",
  17974=>"111100000",
  17975=>"111001110",
  17976=>"000101011",
  17977=>"101100010",
  17978=>"011110100",
  17979=>"100101101",
  17980=>"101111001",
  17981=>"111101100",
  17982=>"011001100",
  17983=>"010010100",
  17984=>"111101001",
  17985=>"011011000",
  17986=>"000000111",
  17987=>"110001110",
  17988=>"100000010",
  17989=>"010010001",
  17990=>"010000010",
  17991=>"010011111",
  17992=>"100100000",
  17993=>"110000011",
  17994=>"001010111",
  17995=>"100001011",
  17996=>"000110010",
  17997=>"010010101",
  17998=>"011100010",
  17999=>"010000000",
  18000=>"001010010",
  18001=>"000001100",
  18002=>"110100001",
  18003=>"001101100",
  18004=>"100011010",
  18005=>"001000101",
  18006=>"101010000",
  18007=>"001101000",
  18008=>"101110100",
  18009=>"010111100",
  18010=>"001110000",
  18011=>"010111101",
  18012=>"011101011",
  18013=>"100010100",
  18014=>"111000111",
  18015=>"111011011",
  18016=>"111011011",
  18017=>"010110010",
  18018=>"101111100",
  18019=>"001001011",
  18020=>"110010000",
  18021=>"011010110",
  18022=>"001111010",
  18023=>"011101010",
  18024=>"010000001",
  18025=>"101010111",
  18026=>"001101000",
  18027=>"001001011",
  18028=>"100011011",
  18029=>"010101111",
  18030=>"001000001",
  18031=>"000000111",
  18032=>"011000111",
  18033=>"000111111",
  18034=>"101101100",
  18035=>"111101101",
  18036=>"011010100",
  18037=>"101100110",
  18038=>"100000000",
  18039=>"111110000",
  18040=>"101100111",
  18041=>"010001011",
  18042=>"010111011",
  18043=>"000101100",
  18044=>"101000111",
  18045=>"011001110",
  18046=>"011001100",
  18047=>"100101011",
  18048=>"101011001",
  18049=>"000110100",
  18050=>"010101000",
  18051=>"111110010",
  18052=>"100011111",
  18053=>"101010001",
  18054=>"100110100",
  18055=>"000000010",
  18056=>"001111111",
  18057=>"001101100",
  18058=>"010101000",
  18059=>"111111110",
  18060=>"001100001",
  18061=>"101101101",
  18062=>"011001101",
  18063=>"010101100",
  18064=>"101001100",
  18065=>"100010000",
  18066=>"001111000",
  18067=>"010111111",
  18068=>"001100010",
  18069=>"010100111",
  18070=>"001101010",
  18071=>"111110111",
  18072=>"110110110",
  18073=>"000110111",
  18074=>"001100000",
  18075=>"111010000",
  18076=>"001001111",
  18077=>"100011000",
  18078=>"000000000",
  18079=>"101101010",
  18080=>"001111000",
  18081=>"100011101",
  18082=>"100010111",
  18083=>"111001101",
  18084=>"001000100",
  18085=>"110111111",
  18086=>"010100000",
  18087=>"000111111",
  18088=>"111001010",
  18089=>"101100100",
  18090=>"011111110",
  18091=>"000101101",
  18092=>"010001000",
  18093=>"101100000",
  18094=>"001110100",
  18095=>"101000001",
  18096=>"011101000",
  18097=>"101111101",
  18098=>"001101010",
  18099=>"011000011",
  18100=>"101110011",
  18101=>"010110101",
  18102=>"001111000",
  18103=>"001110110",
  18104=>"101111000",
  18105=>"001110100",
  18106=>"101101111",
  18107=>"110101101",
  18108=>"000000001",
  18109=>"100010111",
  18110=>"000101110",
  18111=>"110001010",
  18112=>"110111110",
  18113=>"001111001",
  18114=>"011011000",
  18115=>"101101010",
  18116=>"111110111",
  18117=>"101101111",
  18118=>"010101000",
  18119=>"111000100",
  18120=>"100110001",
  18121=>"101011100",
  18122=>"111010111",
  18123=>"011101101",
  18124=>"001000111",
  18125=>"011000111",
  18126=>"001010001",
  18127=>"101011010",
  18128=>"001111100",
  18129=>"101100110",
  18130=>"111010111",
  18131=>"001100101",
  18132=>"110110110",
  18133=>"001001100",
  18134=>"000100111",
  18135=>"110101101",
  18136=>"101000010",
  18137=>"101110010",
  18138=>"000001100",
  18139=>"111011100",
  18140=>"001110001",
  18141=>"011000000",
  18142=>"000010100",
  18143=>"110100111",
  18144=>"110100110",
  18145=>"100110011",
  18146=>"111101000",
  18147=>"011010111",
  18148=>"100011111",
  18149=>"100111110",
  18150=>"010100001",
  18151=>"101001101",
  18152=>"010100100",
  18153=>"111001111",
  18154=>"100100000",
  18155=>"001111001",
  18156=>"111110111",
  18157=>"101000110",
  18158=>"101001101",
  18159=>"001111111",
  18160=>"011001111",
  18161=>"101100000",
  18162=>"100111101",
  18163=>"101011111",
  18164=>"000111010",
  18165=>"000111010",
  18166=>"001011110",
  18167=>"000101011",
  18168=>"110101010",
  18169=>"000100001",
  18170=>"001001110",
  18171=>"100010110",
  18172=>"000110100",
  18173=>"001011101",
  18174=>"111111011",
  18175=>"000101000",
  18176=>"011100001",
  18177=>"001101000",
  18178=>"000100110",
  18179=>"111100110",
  18180=>"100000000",
  18181=>"011010010",
  18182=>"010010011",
  18183=>"100010101",
  18184=>"101010100",
  18185=>"010111010",
  18186=>"001100001",
  18187=>"011110010",
  18188=>"010001111",
  18189=>"000100100",
  18190=>"100010011",
  18191=>"101101111",
  18192=>"101011110",
  18193=>"100011001",
  18194=>"010000001",
  18195=>"100101101",
  18196=>"110010110",
  18197=>"101011010",
  18198=>"100001110",
  18199=>"110000000",
  18200=>"111000110",
  18201=>"101101001",
  18202=>"111100001",
  18203=>"011111101",
  18204=>"100011001",
  18205=>"100101001",
  18206=>"100000111",
  18207=>"001101010",
  18208=>"110111101",
  18209=>"101000000",
  18210=>"110001001",
  18211=>"000100010",
  18212=>"001110101",
  18213=>"110000011",
  18214=>"101000000",
  18215=>"010111111",
  18216=>"101011110",
  18217=>"100111000",
  18218=>"101011111",
  18219=>"000110100",
  18220=>"011111101",
  18221=>"010011110",
  18222=>"001101111",
  18223=>"011001011",
  18224=>"000101010",
  18225=>"110110111",
  18226=>"011110100",
  18227=>"100000001",
  18228=>"001111111",
  18229=>"000100001",
  18230=>"001100100",
  18231=>"011000011",
  18232=>"011001100",
  18233=>"101100110",
  18234=>"110001000",
  18235=>"000000110",
  18236=>"000001011",
  18237=>"011101100",
  18238=>"010111010",
  18239=>"011000110",
  18240=>"110111111",
  18241=>"011100100",
  18242=>"100101010",
  18243=>"101100110",
  18244=>"001010100",
  18245=>"001010011",
  18246=>"010001010",
  18247=>"011000000",
  18248=>"001100101",
  18249=>"110010001",
  18250=>"000001011",
  18251=>"100100100",
  18252=>"101110010",
  18253=>"001111110",
  18254=>"000010111",
  18255=>"010100010",
  18256=>"110000111",
  18257=>"101110101",
  18258=>"011010010",
  18259=>"010110100",
  18260=>"011101111",
  18261=>"111100000",
  18262=>"001111100",
  18263=>"100000101",
  18264=>"110010100",
  18265=>"011111111",
  18266=>"000101011",
  18267=>"101011101",
  18268=>"111010000",
  18269=>"010001111",
  18270=>"001110110",
  18271=>"000001111",
  18272=>"110010000",
  18273=>"010010010",
  18274=>"000111110",
  18275=>"111000001",
  18276=>"110111100",
  18277=>"000111100",
  18278=>"100111100",
  18279=>"001011010",
  18280=>"101000001",
  18281=>"010000010",
  18282=>"000100110",
  18283=>"000110010",
  18284=>"000001000",
  18285=>"110100001",
  18286=>"111011001",
  18287=>"110110110",
  18288=>"101011010",
  18289=>"110011010",
  18290=>"111100101",
  18291=>"001110010",
  18292=>"001011000",
  18293=>"001111010",
  18294=>"100101011",
  18295=>"101101100",
  18296=>"010011011",
  18297=>"100011101",
  18298=>"010011101",
  18299=>"010100001",
  18300=>"111111011",
  18301=>"011101000",
  18302=>"101110111",
  18303=>"110111101",
  18304=>"100010000",
  18305=>"100010010",
  18306=>"111001010",
  18307=>"001000000",
  18308=>"011110011",
  18309=>"000001001",
  18310=>"011110010",
  18311=>"010101100",
  18312=>"111111001",
  18313=>"101111100",
  18314=>"001001011",
  18315=>"110001100",
  18316=>"101111110",
  18317=>"001000000",
  18318=>"100101110",
  18319=>"010100000",
  18320=>"000010100",
  18321=>"011100111",
  18322=>"111100111",
  18323=>"011110010",
  18324=>"110011101",
  18325=>"101010111",
  18326=>"011110010",
  18327=>"110101101",
  18328=>"101000000",
  18329=>"111011001",
  18330=>"100101111",
  18331=>"110000010",
  18332=>"011100001",
  18333=>"010111101",
  18334=>"001010011",
  18335=>"100000011",
  18336=>"100101110",
  18337=>"001101011",
  18338=>"011011000",
  18339=>"100010000",
  18340=>"011110111",
  18341=>"110100001",
  18342=>"111000011",
  18343=>"000001001",
  18344=>"100010101",
  18345=>"101000001",
  18346=>"111000011",
  18347=>"010000110",
  18348=>"100001111",
  18349=>"000010111",
  18350=>"011000101",
  18351=>"110100011",
  18352=>"111101000",
  18353=>"100000110",
  18354=>"100010111",
  18355=>"101010011",
  18356=>"000110111",
  18357=>"100000110",
  18358=>"111101011",
  18359=>"111001010",
  18360=>"100001010",
  18361=>"100101111",
  18362=>"111111010",
  18363=>"000111111",
  18364=>"111011001",
  18365=>"100100010",
  18366=>"001011010",
  18367=>"100100000",
  18368=>"101100000",
  18369=>"100000001",
  18370=>"011110010",
  18371=>"000101010",
  18372=>"010001111",
  18373=>"011110100",
  18374=>"101011101",
  18375=>"000100101",
  18376=>"110110010",
  18377=>"001000000",
  18378=>"111101011",
  18379=>"111001000",
  18380=>"000110110",
  18381=>"111010111",
  18382=>"110000010",
  18383=>"101100001",
  18384=>"111011000",
  18385=>"011011010",
  18386=>"110100111",
  18387=>"100000101",
  18388=>"001111101",
  18389=>"011010101",
  18390=>"110101111",
  18391=>"010111111",
  18392=>"111011100",
  18393=>"100100000",
  18394=>"100101001",
  18395=>"110011011",
  18396=>"101111010",
  18397=>"011111110",
  18398=>"110000011",
  18399=>"000110110",
  18400=>"011001011",
  18401=>"111000011",
  18402=>"011011010",
  18403=>"101001011",
  18404=>"111011110",
  18405=>"101111101",
  18406=>"010111110",
  18407=>"111001000",
  18408=>"110111100",
  18409=>"110000111",
  18410=>"010100111",
  18411=>"011101111",
  18412=>"001110011",
  18413=>"011010100",
  18414=>"101100100",
  18415=>"010000100",
  18416=>"000001011",
  18417=>"101100111",
  18418=>"111101000",
  18419=>"000110111",
  18420=>"100011011",
  18421=>"001000101",
  18422=>"100111000",
  18423=>"001010101",
  18424=>"000011010",
  18425=>"110100101",
  18426=>"100110100",
  18427=>"111111001",
  18428=>"001010001",
  18429=>"101010011",
  18430=>"101101010",
  18431=>"110011100",
  18432=>"001010000",
  18433=>"011100111",
  18434=>"010111011",
  18435=>"111000100",
  18436=>"100010101",
  18437=>"000111000",
  18438=>"010111111",
  18439=>"100100011",
  18440=>"000010011",
  18441=>"100000001",
  18442=>"100011010",
  18443=>"101000001",
  18444=>"110111000",
  18445=>"110100110",
  18446=>"110000010",
  18447=>"010000011",
  18448=>"000001110",
  18449=>"111001010",
  18450=>"111110010",
  18451=>"100111110",
  18452=>"111101010",
  18453=>"111110110",
  18454=>"010111000",
  18455=>"101111100",
  18456=>"011000011",
  18457=>"110110111",
  18458=>"010000000",
  18459=>"110101111",
  18460=>"101010100",
  18461=>"001101010",
  18462=>"110110010",
  18463=>"111100010",
  18464=>"111011010",
  18465=>"110010010",
  18466=>"011111000",
  18467=>"001001110",
  18468=>"111101001",
  18469=>"110101000",
  18470=>"000001001",
  18471=>"100011100",
  18472=>"111010001",
  18473=>"101101010",
  18474=>"000000100",
  18475=>"101110101",
  18476=>"111001101",
  18477=>"100111011",
  18478=>"101111011",
  18479=>"000000100",
  18480=>"111010110",
  18481=>"011110101",
  18482=>"100111111",
  18483=>"010101011",
  18484=>"100110001",
  18485=>"101000101",
  18486=>"110111110",
  18487=>"010010110",
  18488=>"000101111",
  18489=>"101001001",
  18490=>"001100100",
  18491=>"011000101",
  18492=>"010011011",
  18493=>"010101010",
  18494=>"100010001",
  18495=>"111010000",
  18496=>"000111001",
  18497=>"010001110",
  18498=>"011100000",
  18499=>"110111111",
  18500=>"100000101",
  18501=>"111000001",
  18502=>"100001001",
  18503=>"100110000",
  18504=>"010000000",
  18505=>"101001101",
  18506=>"001000101",
  18507=>"001001000",
  18508=>"101111001",
  18509=>"111110111",
  18510=>"101101011",
  18511=>"001010000",
  18512=>"000100100",
  18513=>"011100011",
  18514=>"000011001",
  18515=>"000011100",
  18516=>"100001000",
  18517=>"010110010",
  18518=>"000101110",
  18519=>"101110111",
  18520=>"010101101",
  18521=>"000010011",
  18522=>"101011001",
  18523=>"100110100",
  18524=>"000001000",
  18525=>"000100000",
  18526=>"010110000",
  18527=>"101011110",
  18528=>"100101101",
  18529=>"111011010",
  18530=>"101001100",
  18531=>"011100010",
  18532=>"111010000",
  18533=>"110000100",
  18534=>"101110111",
  18535=>"111011010",
  18536=>"010101110",
  18537=>"001100011",
  18538=>"110110001",
  18539=>"100100001",
  18540=>"000100000",
  18541=>"000001001",
  18542=>"111000101",
  18543=>"101011000",
  18544=>"000010011",
  18545=>"000111101",
  18546=>"110111000",
  18547=>"001001111",
  18548=>"000011010",
  18549=>"100101011",
  18550=>"000010100",
  18551=>"110000101",
  18552=>"010010100",
  18553=>"100001000",
  18554=>"110010010",
  18555=>"011010001",
  18556=>"110011100",
  18557=>"000100111",
  18558=>"111111101",
  18559=>"101001111",
  18560=>"000100010",
  18561=>"001001101",
  18562=>"000001010",
  18563=>"010111101",
  18564=>"000011110",
  18565=>"010101010",
  18566=>"011101111",
  18567=>"100011110",
  18568=>"010101110",
  18569=>"101111101",
  18570=>"110101110",
  18571=>"110101010",
  18572=>"100001011",
  18573=>"110000100",
  18574=>"100001001",
  18575=>"000000110",
  18576=>"101100000",
  18577=>"000110101",
  18578=>"101111100",
  18579=>"011011111",
  18580=>"010010000",
  18581=>"101111000",
  18582=>"101100000",
  18583=>"101101100",
  18584=>"111010110",
  18585=>"000110101",
  18586=>"111101100",
  18587=>"001111111",
  18588=>"100000100",
  18589=>"011110111",
  18590=>"111011101",
  18591=>"000110000",
  18592=>"111111010",
  18593=>"100001000",
  18594=>"000101011",
  18595=>"110011110",
  18596=>"101011011",
  18597=>"100000011",
  18598=>"111010111",
  18599=>"000001000",
  18600=>"100100000",
  18601=>"110010111",
  18602=>"001010010",
  18603=>"000001100",
  18604=>"101011010",
  18605=>"110010111",
  18606=>"001000111",
  18607=>"101100011",
  18608=>"011000111",
  18609=>"111111100",
  18610=>"001000110",
  18611=>"111101011",
  18612=>"000010100",
  18613=>"000001011",
  18614=>"111100101",
  18615=>"110010101",
  18616=>"111001000",
  18617=>"000011111",
  18618=>"001100111",
  18619=>"001001000",
  18620=>"010001101",
  18621=>"010011000",
  18622=>"001000000",
  18623=>"011000101",
  18624=>"111010100",
  18625=>"000000011",
  18626=>"100101110",
  18627=>"010101101",
  18628=>"011101011",
  18629=>"100011110",
  18630=>"011010100",
  18631=>"111000011",
  18632=>"011100011",
  18633=>"101100111",
  18634=>"101011101",
  18635=>"001011100",
  18636=>"101110010",
  18637=>"001001001",
  18638=>"100101000",
  18639=>"000010010",
  18640=>"010000000",
  18641=>"111101010",
  18642=>"101001000",
  18643=>"000101110",
  18644=>"011110101",
  18645=>"100011111",
  18646=>"010110101",
  18647=>"001101101",
  18648=>"001101100",
  18649=>"001100111",
  18650=>"001011110",
  18651=>"101001001",
  18652=>"111110001",
  18653=>"101010111",
  18654=>"110001100",
  18655=>"100001011",
  18656=>"000010011",
  18657=>"011000111",
  18658=>"101110001",
  18659=>"000011100",
  18660=>"000110111",
  18661=>"010000100",
  18662=>"000100010",
  18663=>"110010011",
  18664=>"001001001",
  18665=>"110110000",
  18666=>"111100101",
  18667=>"000011010",
  18668=>"111100101",
  18669=>"100111100",
  18670=>"101111010",
  18671=>"001111110",
  18672=>"100101010",
  18673=>"001000001",
  18674=>"011111111",
  18675=>"011001100",
  18676=>"001101110",
  18677=>"110101010",
  18678=>"000101110",
  18679=>"111111001",
  18680=>"001100010",
  18681=>"010010111",
  18682=>"100001000",
  18683=>"011010100",
  18684=>"000111111",
  18685=>"010111010",
  18686=>"000101111",
  18687=>"001000101",
  18688=>"001101000",
  18689=>"011010111",
  18690=>"110000011",
  18691=>"101110011",
  18692=>"011011001",
  18693=>"100011000",
  18694=>"010001000",
  18695=>"010111101",
  18696=>"110000000",
  18697=>"000111110",
  18698=>"010100011",
  18699=>"110101100",
  18700=>"010010101",
  18701=>"101101001",
  18702=>"101100100",
  18703=>"100101111",
  18704=>"000010111",
  18705=>"100111011",
  18706=>"010000111",
  18707=>"111111100",
  18708=>"110010101",
  18709=>"011010000",
  18710=>"000001111",
  18711=>"000100000",
  18712=>"011010011",
  18713=>"101010100",
  18714=>"111001001",
  18715=>"101010100",
  18716=>"110100100",
  18717=>"110111010",
  18718=>"110011111",
  18719=>"000000100",
  18720=>"001101010",
  18721=>"101011101",
  18722=>"101110111",
  18723=>"011100111",
  18724=>"010110110",
  18725=>"000000101",
  18726=>"001100001",
  18727=>"100001000",
  18728=>"110100111",
  18729=>"011111110",
  18730=>"101101011",
  18731=>"000111110",
  18732=>"010111111",
  18733=>"000000101",
  18734=>"000000001",
  18735=>"001100101",
  18736=>"000110001",
  18737=>"011010001",
  18738=>"101001110",
  18739=>"000101000",
  18740=>"100100000",
  18741=>"000010101",
  18742=>"101101001",
  18743=>"101001111",
  18744=>"101111111",
  18745=>"101000000",
  18746=>"000110111",
  18747=>"100011010",
  18748=>"010101111",
  18749=>"111011101",
  18750=>"111011101",
  18751=>"101100100",
  18752=>"001010001",
  18753=>"110110001",
  18754=>"110110001",
  18755=>"010000110",
  18756=>"010011000",
  18757=>"001001011",
  18758=>"010000100",
  18759=>"101000001",
  18760=>"010100000",
  18761=>"000000011",
  18762=>"001100100",
  18763=>"010001011",
  18764=>"100011011",
  18765=>"100011010",
  18766=>"011110101",
  18767=>"101111100",
  18768=>"110111000",
  18769=>"100011101",
  18770=>"001011101",
  18771=>"010101100",
  18772=>"010100010",
  18773=>"111101000",
  18774=>"001110110",
  18775=>"101110011",
  18776=>"100101011",
  18777=>"110010110",
  18778=>"110001100",
  18779=>"110111111",
  18780=>"111111010",
  18781=>"000001100",
  18782=>"101010001",
  18783=>"100101001",
  18784=>"100001000",
  18785=>"101111001",
  18786=>"100000011",
  18787=>"000101000",
  18788=>"100000110",
  18789=>"000011001",
  18790=>"001011111",
  18791=>"111010100",
  18792=>"010000100",
  18793=>"000111000",
  18794=>"100110000",
  18795=>"010110100",
  18796=>"011111101",
  18797=>"101001101",
  18798=>"001000010",
  18799=>"110101010",
  18800=>"011110111",
  18801=>"010011111",
  18802=>"011001001",
  18803=>"000101001",
  18804=>"110101100",
  18805=>"101010110",
  18806=>"000111000",
  18807=>"010100100",
  18808=>"110001001",
  18809=>"000101000",
  18810=>"111110001",
  18811=>"010110000",
  18812=>"001100101",
  18813=>"000011010",
  18814=>"100110101",
  18815=>"101110110",
  18816=>"101001111",
  18817=>"100011000",
  18818=>"110011011",
  18819=>"000100001",
  18820=>"010110010",
  18821=>"100010000",
  18822=>"101001101",
  18823=>"000100000",
  18824=>"110111010",
  18825=>"111111000",
  18826=>"000010001",
  18827=>"110001110",
  18828=>"111111001",
  18829=>"001000011",
  18830=>"110111001",
  18831=>"111001000",
  18832=>"010111010",
  18833=>"000010010",
  18834=>"010111110",
  18835=>"000101011",
  18836=>"101111110",
  18837=>"011011000",
  18838=>"010000000",
  18839=>"000010110",
  18840=>"000000011",
  18841=>"000010010",
  18842=>"111001011",
  18843=>"110111000",
  18844=>"111011011",
  18845=>"100110111",
  18846=>"000110101",
  18847=>"110100011",
  18848=>"011010111",
  18849=>"001101001",
  18850=>"010001110",
  18851=>"101101110",
  18852=>"110010101",
  18853=>"001101110",
  18854=>"101010101",
  18855=>"001110101",
  18856=>"010100001",
  18857=>"000001110",
  18858=>"000010001",
  18859=>"001001000",
  18860=>"111111000",
  18861=>"101011101",
  18862=>"101101100",
  18863=>"111100010",
  18864=>"000001010",
  18865=>"001011000",
  18866=>"101010110",
  18867=>"001000011",
  18868=>"100000110",
  18869=>"111011101",
  18870=>"010001010",
  18871=>"110110011",
  18872=>"010110111",
  18873=>"001011100",
  18874=>"001011001",
  18875=>"011010010",
  18876=>"000001001",
  18877=>"001001010",
  18878=>"101010110",
  18879=>"000100111",
  18880=>"000000011",
  18881=>"101001010",
  18882=>"110010011",
  18883=>"000111010",
  18884=>"111011001",
  18885=>"000001101",
  18886=>"100111110",
  18887=>"110110000",
  18888=>"100111111",
  18889=>"110011000",
  18890=>"101001010",
  18891=>"111111100",
  18892=>"000011100",
  18893=>"001001000",
  18894=>"001011101",
  18895=>"101000011",
  18896=>"000101011",
  18897=>"000000010",
  18898=>"001101110",
  18899=>"110100011",
  18900=>"101111001",
  18901=>"000011110",
  18902=>"111111101",
  18903=>"001100000",
  18904=>"101010111",
  18905=>"111100100",
  18906=>"001000001",
  18907=>"010100010",
  18908=>"110110010",
  18909=>"001111100",
  18910=>"000001000",
  18911=>"110100011",
  18912=>"110101000",
  18913=>"010001101",
  18914=>"100111011",
  18915=>"001000001",
  18916=>"111010010",
  18917=>"111111111",
  18918=>"101101000",
  18919=>"111010100",
  18920=>"001100000",
  18921=>"000010111",
  18922=>"110111010",
  18923=>"000110111",
  18924=>"100010000",
  18925=>"111001010",
  18926=>"101111011",
  18927=>"111011101",
  18928=>"011000000",
  18929=>"110111110",
  18930=>"010100010",
  18931=>"101110000",
  18932=>"001101001",
  18933=>"110101000",
  18934=>"111100001",
  18935=>"001110111",
  18936=>"010000001",
  18937=>"111110001",
  18938=>"001010001",
  18939=>"000101010",
  18940=>"001010001",
  18941=>"011010100",
  18942=>"000110001",
  18943=>"000111010",
  18944=>"001010010",
  18945=>"110001000",
  18946=>"100100110",
  18947=>"101100010",
  18948=>"100000010",
  18949=>"110001000",
  18950=>"111000000",
  18951=>"010110011",
  18952=>"101100001",
  18953=>"111101100",
  18954=>"111010110",
  18955=>"011101101",
  18956=>"100011111",
  18957=>"000000001",
  18958=>"110100000",
  18959=>"011000000",
  18960=>"101110001",
  18961=>"111111111",
  18962=>"010101101",
  18963=>"110110100",
  18964=>"001000010",
  18965=>"001001101",
  18966=>"010010011",
  18967=>"100001111",
  18968=>"000101110",
  18969=>"000010010",
  18970=>"011010011",
  18971=>"011010111",
  18972=>"111100001",
  18973=>"100000011",
  18974=>"011000010",
  18975=>"001101101",
  18976=>"000001000",
  18977=>"110101010",
  18978=>"111010110",
  18979=>"101000000",
  18980=>"010110000",
  18981=>"111011111",
  18982=>"010101110",
  18983=>"100010111",
  18984=>"110010010",
  18985=>"111111010",
  18986=>"001010011",
  18987=>"111000011",
  18988=>"110110110",
  18989=>"101111111",
  18990=>"110001010",
  18991=>"100011111",
  18992=>"101110101",
  18993=>"010110010",
  18994=>"000110100",
  18995=>"011001101",
  18996=>"101011111",
  18997=>"111001111",
  18998=>"111000101",
  18999=>"100001011",
  19000=>"000101000",
  19001=>"010111010",
  19002=>"101101000",
  19003=>"111010010",
  19004=>"001011101",
  19005=>"010110100",
  19006=>"111110110",
  19007=>"111010101",
  19008=>"110010100",
  19009=>"101110000",
  19010=>"110011011",
  19011=>"001011110",
  19012=>"000000111",
  19013=>"100001100",
  19014=>"000000010",
  19015=>"010111101",
  19016=>"011111100",
  19017=>"110101110",
  19018=>"010101111",
  19019=>"011111010",
  19020=>"011101100",
  19021=>"010110001",
  19022=>"011110110",
  19023=>"001101111",
  19024=>"010001100",
  19025=>"101000100",
  19026=>"000010011",
  19027=>"101101111",
  19028=>"111000111",
  19029=>"000111110",
  19030=>"001010100",
  19031=>"000011000",
  19032=>"111010111",
  19033=>"111101101",
  19034=>"101010111",
  19035=>"010001000",
  19036=>"110110110",
  19037=>"100001000",
  19038=>"010011000",
  19039=>"001000101",
  19040=>"001111001",
  19041=>"100000000",
  19042=>"100001111",
  19043=>"000011101",
  19044=>"011001001",
  19045=>"011110001",
  19046=>"100100001",
  19047=>"110001110",
  19048=>"011010011",
  19049=>"001101000",
  19050=>"011011111",
  19051=>"100011011",
  19052=>"100001100",
  19053=>"101111101",
  19054=>"111101011",
  19055=>"100101100",
  19056=>"101011111",
  19057=>"001101000",
  19058=>"000100001",
  19059=>"111011011",
  19060=>"001010011",
  19061=>"111001010",
  19062=>"100010101",
  19063=>"111100111",
  19064=>"110010110",
  19065=>"100010000",
  19066=>"100111010",
  19067=>"101010100",
  19068=>"001100010",
  19069=>"000010100",
  19070=>"110101110",
  19071=>"110110111",
  19072=>"011011101",
  19073=>"001110011",
  19074=>"100111010",
  19075=>"000011101",
  19076=>"100011100",
  19077=>"000110010",
  19078=>"110000000",
  19079=>"110011011",
  19080=>"110101101",
  19081=>"000011000",
  19082=>"011011011",
  19083=>"101011010",
  19084=>"100001011",
  19085=>"001000101",
  19086=>"100010010",
  19087=>"001001000",
  19088=>"110110001",
  19089=>"001100011",
  19090=>"101000000",
  19091=>"011010011",
  19092=>"100000000",
  19093=>"001101000",
  19094=>"101100011",
  19095=>"011001001",
  19096=>"110111101",
  19097=>"110100011",
  19098=>"101001111",
  19099=>"010001100",
  19100=>"011100111",
  19101=>"000000101",
  19102=>"001010101",
  19103=>"111111111",
  19104=>"011101010",
  19105=>"100011100",
  19106=>"001110110",
  19107=>"000100000",
  19108=>"001000001",
  19109=>"010000001",
  19110=>"100001110",
  19111=>"000100000",
  19112=>"111111111",
  19113=>"010000110",
  19114=>"110001101",
  19115=>"100101111",
  19116=>"010100001",
  19117=>"100011011",
  19118=>"110001010",
  19119=>"010011111",
  19120=>"110000110",
  19121=>"001000110",
  19122=>"010000011",
  19123=>"001000011",
  19124=>"101111100",
  19125=>"011111000",
  19126=>"011000100",
  19127=>"011001100",
  19128=>"001100100",
  19129=>"100100010",
  19130=>"101110111",
  19131=>"001010101",
  19132=>"101011110",
  19133=>"110000101",
  19134=>"110001000",
  19135=>"000001000",
  19136=>"011111110",
  19137=>"100100011",
  19138=>"000000101",
  19139=>"001001101",
  19140=>"010111011",
  19141=>"011011111",
  19142=>"010001110",
  19143=>"100010101",
  19144=>"000010000",
  19145=>"001001111",
  19146=>"111100001",
  19147=>"100010111",
  19148=>"001011000",
  19149=>"001111011",
  19150=>"000010000",
  19151=>"100000000",
  19152=>"011111101",
  19153=>"000110000",
  19154=>"101101111",
  19155=>"111100110",
  19156=>"111010100",
  19157=>"010001111",
  19158=>"111000100",
  19159=>"010101110",
  19160=>"001000111",
  19161=>"010100010",
  19162=>"111010111",
  19163=>"000100111",
  19164=>"000111010",
  19165=>"110111011",
  19166=>"100001100",
  19167=>"010011101",
  19168=>"000100101",
  19169=>"100100011",
  19170=>"001010110",
  19171=>"000111000",
  19172=>"010101101",
  19173=>"000101111",
  19174=>"111101000",
  19175=>"010011010",
  19176=>"111111010",
  19177=>"101100111",
  19178=>"100001011",
  19179=>"100101001",
  19180=>"100100100",
  19181=>"000000001",
  19182=>"011000010",
  19183=>"100010011",
  19184=>"110101001",
  19185=>"011101101",
  19186=>"011111111",
  19187=>"111011111",
  19188=>"000101101",
  19189=>"110000111",
  19190=>"100111001",
  19191=>"110010000",
  19192=>"000000000",
  19193=>"100101110",
  19194=>"011100001",
  19195=>"000010001",
  19196=>"110001011",
  19197=>"100110111",
  19198=>"101111011",
  19199=>"111000001",
  19200=>"101111111",
  19201=>"100101100",
  19202=>"000111011",
  19203=>"001000110",
  19204=>"100001000",
  19205=>"010111110",
  19206=>"010100101",
  19207=>"010110101",
  19208=>"101100010",
  19209=>"001111111",
  19210=>"110010000",
  19211=>"100010010",
  19212=>"110011001",
  19213=>"110110101",
  19214=>"100001111",
  19215=>"100000000",
  19216=>"011100001",
  19217=>"011010101",
  19218=>"011101110",
  19219=>"011100011",
  19220=>"110000001",
  19221=>"111011010",
  19222=>"011011000",
  19223=>"001011101",
  19224=>"110110110",
  19225=>"011000001",
  19226=>"011000011",
  19227=>"101011111",
  19228=>"111101001",
  19229=>"110001111",
  19230=>"110111101",
  19231=>"000001101",
  19232=>"000000101",
  19233=>"000100000",
  19234=>"110011000",
  19235=>"010000100",
  19236=>"011010010",
  19237=>"111110110",
  19238=>"001000111",
  19239=>"111111110",
  19240=>"100000001",
  19241=>"101001110",
  19242=>"010101101",
  19243=>"001101011",
  19244=>"010111110",
  19245=>"000101010",
  19246=>"000111001",
  19247=>"100111111",
  19248=>"010101100",
  19249=>"101111001",
  19250=>"100100100",
  19251=>"111001110",
  19252=>"010001110",
  19253=>"111111110",
  19254=>"010010001",
  19255=>"101000000",
  19256=>"000100011",
  19257=>"001010000",
  19258=>"100111011",
  19259=>"011110100",
  19260=>"110101110",
  19261=>"100100100",
  19262=>"111111111",
  19263=>"000000011",
  19264=>"100001010",
  19265=>"111100110",
  19266=>"001110111",
  19267=>"011111010",
  19268=>"100111010",
  19269=>"100000011",
  19270=>"111101010",
  19271=>"010010000",
  19272=>"011111011",
  19273=>"111001100",
  19274=>"001111100",
  19275=>"111101111",
  19276=>"000011001",
  19277=>"011001110",
  19278=>"011101100",
  19279=>"100101111",
  19280=>"111111010",
  19281=>"010101100",
  19282=>"100111010",
  19283=>"001101111",
  19284=>"100100101",
  19285=>"111001011",
  19286=>"000101101",
  19287=>"001111000",
  19288=>"000001100",
  19289=>"101110100",
  19290=>"101011101",
  19291=>"001100000",
  19292=>"000001010",
  19293=>"010101000",
  19294=>"101001011",
  19295=>"000000110",
  19296=>"001110001",
  19297=>"000000110",
  19298=>"100100110",
  19299=>"111000100",
  19300=>"001000011",
  19301=>"111101010",
  19302=>"110111110",
  19303=>"111001000",
  19304=>"101110011",
  19305=>"011010111",
  19306=>"000111101",
  19307=>"001110001",
  19308=>"110010100",
  19309=>"000110011",
  19310=>"100111111",
  19311=>"111111010",
  19312=>"111100010",
  19313=>"111111111",
  19314=>"000101010",
  19315=>"011110000",
  19316=>"010100000",
  19317=>"011100110",
  19318=>"110110000",
  19319=>"101001110",
  19320=>"111010011",
  19321=>"010111101",
  19322=>"101000000",
  19323=>"010111001",
  19324=>"001000100",
  19325=>"101110111",
  19326=>"111011001",
  19327=>"111001011",
  19328=>"101011101",
  19329=>"000101111",
  19330=>"000001010",
  19331=>"000110010",
  19332=>"001110000",
  19333=>"010111001",
  19334=>"011001011",
  19335=>"101010101",
  19336=>"101010001",
  19337=>"110110000",
  19338=>"000011101",
  19339=>"110011100",
  19340=>"001000111",
  19341=>"100011010",
  19342=>"000011001",
  19343=>"001001100",
  19344=>"010011110",
  19345=>"010100010",
  19346=>"101011110",
  19347=>"110110000",
  19348=>"011010111",
  19349=>"111011110",
  19350=>"101100011",
  19351=>"001100100",
  19352=>"001100100",
  19353=>"001100110",
  19354=>"000100100",
  19355=>"110010010",
  19356=>"101110100",
  19357=>"110000111",
  19358=>"101000001",
  19359=>"111101110",
  19360=>"100000000",
  19361=>"010011010",
  19362=>"111111111",
  19363=>"101100001",
  19364=>"001001000",
  19365=>"100011011",
  19366=>"000000000",
  19367=>"101110010",
  19368=>"001000100",
  19369=>"111111111",
  19370=>"011100111",
  19371=>"101011001",
  19372=>"010100110",
  19373=>"111100101",
  19374=>"010010001",
  19375=>"001111101",
  19376=>"000100000",
  19377=>"100010011",
  19378=>"101000000",
  19379=>"101000010",
  19380=>"100111111",
  19381=>"011011000",
  19382=>"000100001",
  19383=>"101110001",
  19384=>"101001100",
  19385=>"100111010",
  19386=>"100010011",
  19387=>"001001000",
  19388=>"100100001",
  19389=>"101110000",
  19390=>"011000000",
  19391=>"010000100",
  19392=>"011001101",
  19393=>"100111101",
  19394=>"110011101",
  19395=>"010110010",
  19396=>"010111010",
  19397=>"111110011",
  19398=>"011010000",
  19399=>"000000010",
  19400=>"111111010",
  19401=>"011110111",
  19402=>"001010101",
  19403=>"101100111",
  19404=>"110000101",
  19405=>"111111000",
  19406=>"111111001",
  19407=>"101011101",
  19408=>"110001101",
  19409=>"111011110",
  19410=>"011001011",
  19411=>"101111100",
  19412=>"100000001",
  19413=>"100010100",
  19414=>"100101110",
  19415=>"011100011",
  19416=>"011011011",
  19417=>"001100000",
  19418=>"010101111",
  19419=>"100011110",
  19420=>"110001001",
  19421=>"000001010",
  19422=>"010010111",
  19423=>"010010001",
  19424=>"110111110",
  19425=>"101110111",
  19426=>"101111110",
  19427=>"010111100",
  19428=>"000110111",
  19429=>"101101111",
  19430=>"011011110",
  19431=>"011101001",
  19432=>"000001011",
  19433=>"000000010",
  19434=>"011000010",
  19435=>"001010000",
  19436=>"010101000",
  19437=>"110011001",
  19438=>"111111111",
  19439=>"001101001",
  19440=>"100110100",
  19441=>"110010101",
  19442=>"011101100",
  19443=>"000111111",
  19444=>"110101011",
  19445=>"000001100",
  19446=>"100000100",
  19447=>"011101000",
  19448=>"011110101",
  19449=>"100100101",
  19450=>"111001101",
  19451=>"100101111",
  19452=>"010110100",
  19453=>"000100000",
  19454=>"100110111",
  19455=>"001000011",
  19456=>"110110000",
  19457=>"001011101",
  19458=>"110000111",
  19459=>"110110100",
  19460=>"000101111",
  19461=>"110010000",
  19462=>"111111101",
  19463=>"100101011",
  19464=>"101100100",
  19465=>"010011011",
  19466=>"011001111",
  19467=>"100101111",
  19468=>"011011101",
  19469=>"000010101",
  19470=>"001011101",
  19471=>"001011110",
  19472=>"011000101",
  19473=>"000010110",
  19474=>"111111000",
  19475=>"110101001",
  19476=>"010000001",
  19477=>"101010100",
  19478=>"110110100",
  19479=>"001001011",
  19480=>"100100101",
  19481=>"100010101",
  19482=>"111001110",
  19483=>"000000001",
  19484=>"110110111",
  19485=>"001101110",
  19486=>"101010001",
  19487=>"111101010",
  19488=>"110011011",
  19489=>"100011011",
  19490=>"000011000",
  19491=>"010001111",
  19492=>"101101001",
  19493=>"101111001",
  19494=>"001000010",
  19495=>"011000100",
  19496=>"100001110",
  19497=>"000101011",
  19498=>"010000011",
  19499=>"011001101",
  19500=>"001101000",
  19501=>"000000111",
  19502=>"011110000",
  19503=>"011011111",
  19504=>"110111010",
  19505=>"101111011",
  19506=>"111011101",
  19507=>"110111011",
  19508=>"110111100",
  19509=>"111101100",
  19510=>"001110110",
  19511=>"111111111",
  19512=>"001011011",
  19513=>"000000001",
  19514=>"001001011",
  19515=>"000101110",
  19516=>"110100110",
  19517=>"111111101",
  19518=>"001101100",
  19519=>"111011000",
  19520=>"010111011",
  19521=>"101110011",
  19522=>"111100000",
  19523=>"000000100",
  19524=>"001100010",
  19525=>"111110111",
  19526=>"001000010",
  19527=>"101111101",
  19528=>"111000100",
  19529=>"001111111",
  19530=>"111000111",
  19531=>"001000101",
  19532=>"100000101",
  19533=>"110110110",
  19534=>"010110111",
  19535=>"011111100",
  19536=>"000000001",
  19537=>"111001111",
  19538=>"000110011",
  19539=>"010101001",
  19540=>"011101011",
  19541=>"101101110",
  19542=>"101110101",
  19543=>"000010101",
  19544=>"111111111",
  19545=>"101111100",
  19546=>"001110011",
  19547=>"010111101",
  19548=>"000100000",
  19549=>"000111110",
  19550=>"101111101",
  19551=>"110001110",
  19552=>"001101001",
  19553=>"001000011",
  19554=>"111101100",
  19555=>"000000011",
  19556=>"100110111",
  19557=>"100010011",
  19558=>"100010000",
  19559=>"000100111",
  19560=>"101000111",
  19561=>"011111111",
  19562=>"101001101",
  19563=>"010111110",
  19564=>"111110000",
  19565=>"111011101",
  19566=>"100000100",
  19567=>"110001000",
  19568=>"110000000",
  19569=>"000010110",
  19570=>"000000011",
  19571=>"000101011",
  19572=>"100010101",
  19573=>"001100010",
  19574=>"111101100",
  19575=>"001000110",
  19576=>"010011101",
  19577=>"111100111",
  19578=>"101100110",
  19579=>"101100000",
  19580=>"001001101",
  19581=>"110110011",
  19582=>"000000000",
  19583=>"100011011",
  19584=>"100101011",
  19585=>"010000011",
  19586=>"111110000",
  19587=>"000001001",
  19588=>"000100011",
  19589=>"100000100",
  19590=>"110110011",
  19591=>"100100100",
  19592=>"000110001",
  19593=>"101100110",
  19594=>"110010000",
  19595=>"110111111",
  19596=>"001110100",
  19597=>"010101101",
  19598=>"110000100",
  19599=>"011111111",
  19600=>"110001011",
  19601=>"000100000",
  19602=>"010010010",
  19603=>"010110011",
  19604=>"000011111",
  19605=>"001111010",
  19606=>"000000001",
  19607=>"001000101",
  19608=>"100010011",
  19609=>"011101011",
  19610=>"101110111",
  19611=>"111110100",
  19612=>"000011011",
  19613=>"110101110",
  19614=>"000110011",
  19615=>"100001011",
  19616=>"011000101",
  19617=>"101101011",
  19618=>"101001101",
  19619=>"111100001",
  19620=>"000010000",
  19621=>"010101001",
  19622=>"000011101",
  19623=>"100010001",
  19624=>"100011101",
  19625=>"111011010",
  19626=>"110000110",
  19627=>"100111101",
  19628=>"110101001",
  19629=>"111110011",
  19630=>"100100010",
  19631=>"110110110",
  19632=>"001010110",
  19633=>"010111011",
  19634=>"111101000",
  19635=>"000010000",
  19636=>"001101000",
  19637=>"100111110",
  19638=>"010100010",
  19639=>"010000011",
  19640=>"011110110",
  19641=>"001111110",
  19642=>"011001101",
  19643=>"011011110",
  19644=>"001011000",
  19645=>"101101111",
  19646=>"110001101",
  19647=>"110101100",
  19648=>"100000011",
  19649=>"111011001",
  19650=>"001111001",
  19651=>"101110110",
  19652=>"110001000",
  19653=>"111010011",
  19654=>"110000000",
  19655=>"011111100",
  19656=>"011010000",
  19657=>"001100101",
  19658=>"010111101",
  19659=>"011001100",
  19660=>"001100000",
  19661=>"101110110",
  19662=>"100001010",
  19663=>"110000011",
  19664=>"100000011",
  19665=>"001000111",
  19666=>"010110001",
  19667=>"010001001",
  19668=>"111010010",
  19669=>"001101001",
  19670=>"101011100",
  19671=>"111000110",
  19672=>"011000010",
  19673=>"000100100",
  19674=>"000011101",
  19675=>"001000010",
  19676=>"010001111",
  19677=>"010011101",
  19678=>"001010110",
  19679=>"011101111",
  19680=>"001010100",
  19681=>"011000011",
  19682=>"000110110",
  19683=>"011011001",
  19684=>"101010011",
  19685=>"000011101",
  19686=>"111110010",
  19687=>"011111010",
  19688=>"110110001",
  19689=>"111100010",
  19690=>"011100111",
  19691=>"000010001",
  19692=>"110001000",
  19693=>"100010110",
  19694=>"100000010",
  19695=>"001010001",
  19696=>"001110010",
  19697=>"110010001",
  19698=>"101011001",
  19699=>"111111001",
  19700=>"111100101",
  19701=>"010011110",
  19702=>"110101010",
  19703=>"001010111",
  19704=>"000111110",
  19705=>"110111000",
  19706=>"010110100",
  19707=>"011110110",
  19708=>"110101101",
  19709=>"101010010",
  19710=>"100100111",
  19711=>"111100101",
  19712=>"110010011",
  19713=>"101110010",
  19714=>"000000110",
  19715=>"110010100",
  19716=>"100110110",
  19717=>"111110000",
  19718=>"010010111",
  19719=>"011010101",
  19720=>"010000000",
  19721=>"010011000",
  19722=>"111010011",
  19723=>"010110001",
  19724=>"000101111",
  19725=>"100000010",
  19726=>"010011010",
  19727=>"000011001",
  19728=>"011001010",
  19729=>"110101000",
  19730=>"010010100",
  19731=>"001110011",
  19732=>"000010000",
  19733=>"000001101",
  19734=>"001011101",
  19735=>"000001110",
  19736=>"001101110",
  19737=>"111001010",
  19738=>"110011101",
  19739=>"001111111",
  19740=>"111001110",
  19741=>"010000110",
  19742=>"011000101",
  19743=>"011110011",
  19744=>"000010001",
  19745=>"001101101",
  19746=>"001101100",
  19747=>"010010000",
  19748=>"111001000",
  19749=>"110110111",
  19750=>"011100100",
  19751=>"000100011",
  19752=>"011011110",
  19753=>"000110110",
  19754=>"010001101",
  19755=>"100000010",
  19756=>"101000100",
  19757=>"001001100",
  19758=>"000000000",
  19759=>"000101001",
  19760=>"100110111",
  19761=>"101101111",
  19762=>"111100011",
  19763=>"000101100",
  19764=>"011100000",
  19765=>"101011011",
  19766=>"101000100",
  19767=>"101100111",
  19768=>"001001011",
  19769=>"010000101",
  19770=>"000110011",
  19771=>"100111001",
  19772=>"100010011",
  19773=>"011111011",
  19774=>"000101011",
  19775=>"101110100",
  19776=>"111111011",
  19777=>"010111011",
  19778=>"011110110",
  19779=>"101100111",
  19780=>"001100010",
  19781=>"111011111",
  19782=>"010110001",
  19783=>"000001101",
  19784=>"000000110",
  19785=>"101011000",
  19786=>"011110001",
  19787=>"100001100",
  19788=>"001010001",
  19789=>"010111111",
  19790=>"110010000",
  19791=>"101110110",
  19792=>"111111000",
  19793=>"111111101",
  19794=>"000110111",
  19795=>"101010111",
  19796=>"101001000",
  19797=>"101111111",
  19798=>"000100100",
  19799=>"011011101",
  19800=>"000100011",
  19801=>"000101001",
  19802=>"110100100",
  19803=>"100100110",
  19804=>"010001000",
  19805=>"000010000",
  19806=>"100101111",
  19807=>"010100000",
  19808=>"111111011",
  19809=>"100010010",
  19810=>"010110011",
  19811=>"000000101",
  19812=>"001101001",
  19813=>"000100001",
  19814=>"111110001",
  19815=>"011000101",
  19816=>"100110100",
  19817=>"101101001",
  19818=>"111011011",
  19819=>"111000101",
  19820=>"110011011",
  19821=>"101010000",
  19822=>"100111010",
  19823=>"100110110",
  19824=>"100101110",
  19825=>"110010000",
  19826=>"011110111",
  19827=>"111101101",
  19828=>"000001100",
  19829=>"011011001",
  19830=>"000011011",
  19831=>"110011110",
  19832=>"110111111",
  19833=>"100000110",
  19834=>"111011001",
  19835=>"001100111",
  19836=>"111001010",
  19837=>"110000011",
  19838=>"111100110",
  19839=>"011110101",
  19840=>"000100111",
  19841=>"011100101",
  19842=>"110010011",
  19843=>"100011110",
  19844=>"010011010",
  19845=>"100000100",
  19846=>"111100010",
  19847=>"110010001",
  19848=>"000001101",
  19849=>"111110011",
  19850=>"111010000",
  19851=>"000010101",
  19852=>"011101100",
  19853=>"010010110",
  19854=>"010000000",
  19855=>"010100010",
  19856=>"011110001",
  19857=>"000000111",
  19858=>"001101101",
  19859=>"011011101",
  19860=>"000111001",
  19861=>"011101100",
  19862=>"011011001",
  19863=>"101100001",
  19864=>"010111100",
  19865=>"000100111",
  19866=>"100000100",
  19867=>"011110111",
  19868=>"101011000",
  19869=>"101111100",
  19870=>"100001110",
  19871=>"111111111",
  19872=>"001011101",
  19873=>"110110100",
  19874=>"100001111",
  19875=>"000100110",
  19876=>"110110100",
  19877=>"101011001",
  19878=>"010101000",
  19879=>"111100000",
  19880=>"110110111",
  19881=>"011101111",
  19882=>"001111010",
  19883=>"000010011",
  19884=>"001011111",
  19885=>"111001011",
  19886=>"000111001",
  19887=>"001011110",
  19888=>"111000011",
  19889=>"011101101",
  19890=>"000001111",
  19891=>"000110101",
  19892=>"000110111",
  19893=>"001000000",
  19894=>"000110000",
  19895=>"111000111",
  19896=>"110010011",
  19897=>"000100100",
  19898=>"000100000",
  19899=>"010101000",
  19900=>"011010111",
  19901=>"110111001",
  19902=>"110011110",
  19903=>"011101101",
  19904=>"110111111",
  19905=>"000010001",
  19906=>"001010011",
  19907=>"111001010",
  19908=>"000010000",
  19909=>"100001010",
  19910=>"111000011",
  19911=>"101000101",
  19912=>"101010111",
  19913=>"000100101",
  19914=>"100000101",
  19915=>"111111101",
  19916=>"000111001",
  19917=>"011110000",
  19918=>"000000110",
  19919=>"111110111",
  19920=>"100000001",
  19921=>"000010010",
  19922=>"010001001",
  19923=>"001011000",
  19924=>"110101110",
  19925=>"110101010",
  19926=>"011101101",
  19927=>"010001110",
  19928=>"011100100",
  19929=>"111111110",
  19930=>"001011010",
  19931=>"000011100",
  19932=>"001000001",
  19933=>"010000000",
  19934=>"011000100",
  19935=>"001101110",
  19936=>"110010011",
  19937=>"111111000",
  19938=>"110100111",
  19939=>"011011011",
  19940=>"110011100",
  19941=>"011010111",
  19942=>"000101100",
  19943=>"111010111",
  19944=>"000110001",
  19945=>"011111101",
  19946=>"011100110",
  19947=>"011000101",
  19948=>"110100000",
  19949=>"100010000",
  19950=>"100111111",
  19951=>"101101111",
  19952=>"100011110",
  19953=>"111001000",
  19954=>"010101001",
  19955=>"011011011",
  19956=>"100011100",
  19957=>"100001100",
  19958=>"010011110",
  19959=>"010110011",
  19960=>"100101011",
  19961=>"101111011",
  19962=>"000100100",
  19963=>"000101000",
  19964=>"001100100",
  19965=>"001101010",
  19966=>"011100100",
  19967=>"011111100",
  19968=>"100011101",
  19969=>"101000110",
  19970=>"101011100",
  19971=>"101111110",
  19972=>"011000100",
  19973=>"001010001",
  19974=>"110010100",
  19975=>"101000011",
  19976=>"011110110",
  19977=>"110100101",
  19978=>"001001001",
  19979=>"000111000",
  19980=>"100110111",
  19981=>"000111101",
  19982=>"100001100",
  19983=>"010011000",
  19984=>"100111101",
  19985=>"101010001",
  19986=>"111001100",
  19987=>"000101101",
  19988=>"011000110",
  19989=>"100000000",
  19990=>"110001100",
  19991=>"000110111",
  19992=>"011111011",
  19993=>"000011100",
  19994=>"010001110",
  19995=>"110011111",
  19996=>"010001011",
  19997=>"001000110",
  19998=>"100101001",
  19999=>"100010101",
  20000=>"111001110",
  20001=>"010000100",
  20002=>"000000100",
  20003=>"101001001",
  20004=>"001100101",
  20005=>"001101111",
  20006=>"010101111",
  20007=>"010000110",
  20008=>"001101000",
  20009=>"110111100",
  20010=>"111101101",
  20011=>"011110000",
  20012=>"110010001",
  20013=>"000000000",
  20014=>"001001111",
  20015=>"110010111",
  20016=>"110110000",
  20017=>"110011111",
  20018=>"110110010",
  20019=>"010111110",
  20020=>"000010011",
  20021=>"111101010",
  20022=>"100100111",
  20023=>"110011100",
  20024=>"100101100",
  20025=>"001000110",
  20026=>"110111011",
  20027=>"101100001",
  20028=>"011000010",
  20029=>"010010001",
  20030=>"000111111",
  20031=>"010011010",
  20032=>"001101000",
  20033=>"010011111",
  20034=>"010010100",
  20035=>"000000000",
  20036=>"111100001",
  20037=>"111000100",
  20038=>"110000010",
  20039=>"010110100",
  20040=>"000010110",
  20041=>"011011110",
  20042=>"010000101",
  20043=>"110011100",
  20044=>"110101111",
  20045=>"110100001",
  20046=>"100100111",
  20047=>"011011011",
  20048=>"001110111",
  20049=>"101111100",
  20050=>"110110101",
  20051=>"001000001",
  20052=>"001001011",
  20053=>"000001101",
  20054=>"101010101",
  20055=>"101110100",
  20056=>"000001010",
  20057=>"001011110",
  20058=>"010111111",
  20059=>"101011000",
  20060=>"001100001",
  20061=>"001001111",
  20062=>"101011111",
  20063=>"010111101",
  20064=>"011111110",
  20065=>"001010011",
  20066=>"111101000",
  20067=>"101101100",
  20068=>"111110100",
  20069=>"100101100",
  20070=>"100110111",
  20071=>"000000010",
  20072=>"000001000",
  20073=>"100110110",
  20074=>"011010100",
  20075=>"110011111",
  20076=>"000111100",
  20077=>"100111110",
  20078=>"111100100",
  20079=>"101101111",
  20080=>"001100001",
  20081=>"010000100",
  20082=>"101010110",
  20083=>"100011010",
  20084=>"110010110",
  20085=>"001101111",
  20086=>"110001010",
  20087=>"000010101",
  20088=>"101001110",
  20089=>"101011100",
  20090=>"111011010",
  20091=>"000000101",
  20092=>"000111000",
  20093=>"001000100",
  20094=>"111101001",
  20095=>"100001101",
  20096=>"100011111",
  20097=>"110011101",
  20098=>"111011100",
  20099=>"001010111",
  20100=>"101101110",
  20101=>"001000010",
  20102=>"000011110",
  20103=>"111100110",
  20104=>"100101111",
  20105=>"011010111",
  20106=>"011010101",
  20107=>"110000000",
  20108=>"111001010",
  20109=>"000011011",
  20110=>"111000001",
  20111=>"111011000",
  20112=>"010101011",
  20113=>"010001000",
  20114=>"111111110",
  20115=>"001001100",
  20116=>"001011000",
  20117=>"001101101",
  20118=>"011101010",
  20119=>"001011011",
  20120=>"101111100",
  20121=>"110110000",
  20122=>"011110001",
  20123=>"001100001",
  20124=>"001101111",
  20125=>"100110100",
  20126=>"110111101",
  20127=>"111000111",
  20128=>"111001000",
  20129=>"001010111",
  20130=>"001000000",
  20131=>"110011100",
  20132=>"000110000",
  20133=>"010001110",
  20134=>"100111101",
  20135=>"000000000",
  20136=>"010111110",
  20137=>"101100011",
  20138=>"010110001",
  20139=>"101000101",
  20140=>"101110111",
  20141=>"110101001",
  20142=>"001010000",
  20143=>"011001111",
  20144=>"001100111",
  20145=>"010000001",
  20146=>"001111011",
  20147=>"010110000",
  20148=>"101011001",
  20149=>"000111110",
  20150=>"100000000",
  20151=>"010111011",
  20152=>"101100110",
  20153=>"110111010",
  20154=>"011011100",
  20155=>"110110100",
  20156=>"100001111",
  20157=>"110011101",
  20158=>"001000011",
  20159=>"111110101",
  20160=>"101100100",
  20161=>"110000011",
  20162=>"001011010",
  20163=>"010111000",
  20164=>"011011100",
  20165=>"000110000",
  20166=>"100101001",
  20167=>"101111111",
  20168=>"101001001",
  20169=>"111101000",
  20170=>"000100011",
  20171=>"101001100",
  20172=>"100011110",
  20173=>"111101110",
  20174=>"000000110",
  20175=>"000110110",
  20176=>"110110000",
  20177=>"100000000",
  20178=>"000010111",
  20179=>"001001110",
  20180=>"011010001",
  20181=>"100001100",
  20182=>"110101111",
  20183=>"000110111",
  20184=>"001100111",
  20185=>"001101101",
  20186=>"011000100",
  20187=>"110100101",
  20188=>"000110111",
  20189=>"111010000",
  20190=>"100110111",
  20191=>"100001001",
  20192=>"000111001",
  20193=>"000110011",
  20194=>"111101100",
  20195=>"000011011",
  20196=>"010000010",
  20197=>"011001101",
  20198=>"110000100",
  20199=>"011010010",
  20200=>"100100100",
  20201=>"101010010",
  20202=>"110111101",
  20203=>"011001110",
  20204=>"001111110",
  20205=>"100101001",
  20206=>"011111110",
  20207=>"001111010",
  20208=>"100011011",
  20209=>"001100001",
  20210=>"010011101",
  20211=>"000001101",
  20212=>"010110001",
  20213=>"111001111",
  20214=>"101010100",
  20215=>"011110011",
  20216=>"100111000",
  20217=>"101000001",
  20218=>"111101000",
  20219=>"100000100",
  20220=>"101100111",
  20221=>"111101101",
  20222=>"001110001",
  20223=>"100100100",
  20224=>"011011110",
  20225=>"000011011",
  20226=>"010100111",
  20227=>"001101010",
  20228=>"010001100",
  20229=>"100110111",
  20230=>"000111110",
  20231=>"101101011",
  20232=>"110010100",
  20233=>"101101001",
  20234=>"001011110",
  20235=>"011111110",
  20236=>"001000001",
  20237=>"000011100",
  20238=>"010011011",
  20239=>"110000111",
  20240=>"101111111",
  20241=>"001010110",
  20242=>"011110010",
  20243=>"110100111",
  20244=>"110010011",
  20245=>"001110000",
  20246=>"111010011",
  20247=>"000100000",
  20248=>"111011010",
  20249=>"101010010",
  20250=>"010000001",
  20251=>"101110100",
  20252=>"001011001",
  20253=>"000010011",
  20254=>"111101100",
  20255=>"100000011",
  20256=>"111000100",
  20257=>"010111011",
  20258=>"101000101",
  20259=>"001001111",
  20260=>"001001101",
  20261=>"000100110",
  20262=>"101111000",
  20263=>"001011000",
  20264=>"110011111",
  20265=>"101001110",
  20266=>"101110101",
  20267=>"100100010",
  20268=>"001000101",
  20269=>"001111010",
  20270=>"101101010",
  20271=>"000000001",
  20272=>"000010111",
  20273=>"100001101",
  20274=>"100010010",
  20275=>"111000111",
  20276=>"111101111",
  20277=>"011010111",
  20278=>"100000111",
  20279=>"101000111",
  20280=>"101000111",
  20281=>"110101010",
  20282=>"101010000",
  20283=>"111011010",
  20284=>"111110000",
  20285=>"000010000",
  20286=>"100010101",
  20287=>"100010110",
  20288=>"010111100",
  20289=>"011001001",
  20290=>"101001000",
  20291=>"101101111",
  20292=>"110101000",
  20293=>"011000000",
  20294=>"000101111",
  20295=>"011000000",
  20296=>"011111011",
  20297=>"000011100",
  20298=>"001011110",
  20299=>"000101010",
  20300=>"010001110",
  20301=>"001010011",
  20302=>"001001000",
  20303=>"111010010",
  20304=>"101010101",
  20305=>"100111110",
  20306=>"000011001",
  20307=>"000001101",
  20308=>"011010001",
  20309=>"011001011",
  20310=>"011100000",
  20311=>"010000000",
  20312=>"111010001",
  20313=>"000010010",
  20314=>"010110011",
  20315=>"011000000",
  20316=>"110111010",
  20317=>"000100100",
  20318=>"101111101",
  20319=>"001000110",
  20320=>"010010000",
  20321=>"111011101",
  20322=>"011101111",
  20323=>"001010010",
  20324=>"111000101",
  20325=>"100011101",
  20326=>"100101000",
  20327=>"011101001",
  20328=>"001001010",
  20329=>"101101101",
  20330=>"000111111",
  20331=>"010001111",
  20332=>"010011011",
  20333=>"100111110",
  20334=>"001001100",
  20335=>"011101010",
  20336=>"110100110",
  20337=>"010100000",
  20338=>"111101111",
  20339=>"000111101",
  20340=>"000100010",
  20341=>"000110110",
  20342=>"100110111",
  20343=>"100000111",
  20344=>"100101010",
  20345=>"001101111",
  20346=>"110111100",
  20347=>"000111011",
  20348=>"100001100",
  20349=>"111001001",
  20350=>"100000100",
  20351=>"001001101",
  20352=>"010110010",
  20353=>"000010011",
  20354=>"011010000",
  20355=>"011100000",
  20356=>"001001111",
  20357=>"011100100",
  20358=>"000011100",
  20359=>"101111000",
  20360=>"100001100",
  20361=>"100000111",
  20362=>"111100011",
  20363=>"100000111",
  20364=>"000100101",
  20365=>"110001011",
  20366=>"010010001",
  20367=>"100110100",
  20368=>"010110101",
  20369=>"111111111",
  20370=>"100110011",
  20371=>"101111101",
  20372=>"100001110",
  20373=>"001101000",
  20374=>"001001000",
  20375=>"111001111",
  20376=>"001111000",
  20377=>"010000101",
  20378=>"101110011",
  20379=>"111110001",
  20380=>"010111101",
  20381=>"010100100",
  20382=>"000011011",
  20383=>"000010101",
  20384=>"000000011",
  20385=>"111000111",
  20386=>"000110100",
  20387=>"111101101",
  20388=>"011000011",
  20389=>"001010111",
  20390=>"010001001",
  20391=>"100001010",
  20392=>"100011001",
  20393=>"001001110",
  20394=>"010100101",
  20395=>"111001111",
  20396=>"011101111",
  20397=>"000000101",
  20398=>"011110010",
  20399=>"001101100",
  20400=>"100111001",
  20401=>"010110111",
  20402=>"111101111",
  20403=>"011100011",
  20404=>"111100100",
  20405=>"101101011",
  20406=>"011101011",
  20407=>"010000111",
  20408=>"011100011",
  20409=>"000100110",
  20410=>"000111011",
  20411=>"110100010",
  20412=>"100000101",
  20413=>"110100110",
  20414=>"101000010",
  20415=>"110000001",
  20416=>"101111101",
  20417=>"001001010",
  20418=>"101001000",
  20419=>"111001010",
  20420=>"011110110",
  20421=>"101110010",
  20422=>"000011000",
  20423=>"110011111",
  20424=>"000000010",
  20425=>"101101001",
  20426=>"011111111",
  20427=>"110011101",
  20428=>"010100011",
  20429=>"000100110",
  20430=>"010011111",
  20431=>"101010100",
  20432=>"110011111",
  20433=>"001000001",
  20434=>"111010100",
  20435=>"010000011",
  20436=>"100100111",
  20437=>"100110001",
  20438=>"101100100",
  20439=>"101100111",
  20440=>"000101011",
  20441=>"001110101",
  20442=>"001001011",
  20443=>"011001001",
  20444=>"101000000",
  20445=>"000111000",
  20446=>"000010100",
  20447=>"001000011",
  20448=>"010111110",
  20449=>"010111111",
  20450=>"110110101",
  20451=>"100010111",
  20452=>"011000110",
  20453=>"000010000",
  20454=>"001010011",
  20455=>"000000110",
  20456=>"001001010",
  20457=>"111010110",
  20458=>"011101100",
  20459=>"100101101",
  20460=>"000000001",
  20461=>"110110100",
  20462=>"010011101",
  20463=>"010000111",
  20464=>"000011110",
  20465=>"001011100",
  20466=>"011010000",
  20467=>"110000100",
  20468=>"011100000",
  20469=>"000011101",
  20470=>"000111101",
  20471=>"010001011",
  20472=>"000000110",
  20473=>"110000010",
  20474=>"010011110",
  20475=>"101110111",
  20476=>"010000010",
  20477=>"000011111",
  20478=>"010101110",
  20479=>"110011110",
  20480=>"100000010",
  20481=>"011001110",
  20482=>"000100111",
  20483=>"101110101",
  20484=>"000011110",
  20485=>"111000010",
  20486=>"011000000",
  20487=>"001110010",
  20488=>"010111011",
  20489=>"001111101",
  20490=>"111010111",
  20491=>"100000011",
  20492=>"111100111",
  20493=>"010101111",
  20494=>"100100001",
  20495=>"011011001",
  20496=>"000000010",
  20497=>"001000110",
  20498=>"010101000",
  20499=>"111011101",
  20500=>"011110111",
  20501=>"100100011",
  20502=>"000111101",
  20503=>"111011101",
  20504=>"010001101",
  20505=>"001111001",
  20506=>"010001000",
  20507=>"011110011",
  20508=>"111010111",
  20509=>"110110010",
  20510=>"101000111",
  20511=>"101111011",
  20512=>"010011111",
  20513=>"111001101",
  20514=>"101101011",
  20515=>"010100011",
  20516=>"100101000",
  20517=>"111101011",
  20518=>"101011101",
  20519=>"100001110",
  20520=>"110010101",
  20521=>"111011110",
  20522=>"000111011",
  20523=>"111101111",
  20524=>"001110011",
  20525=>"110011111",
  20526=>"000001010",
  20527=>"111011100",
  20528=>"000101001",
  20529=>"111001101",
  20530=>"011000101",
  20531=>"001110100",
  20532=>"000000100",
  20533=>"001000010",
  20534=>"101011000",
  20535=>"010001101",
  20536=>"110100001",
  20537=>"101110101",
  20538=>"001111101",
  20539=>"111001000",
  20540=>"000011010",
  20541=>"001100110",
  20542=>"110000000",
  20543=>"100000010",
  20544=>"101001001",
  20545=>"000001010",
  20546=>"000110011",
  20547=>"101101000",
  20548=>"010100101",
  20549=>"101001001",
  20550=>"101111100",
  20551=>"101110011",
  20552=>"011001100",
  20553=>"110111000",
  20554=>"100011111",
  20555=>"100010010",
  20556=>"110100010",
  20557=>"110110010",
  20558=>"010110101",
  20559=>"001111011",
  20560=>"111011001",
  20561=>"111111011",
  20562=>"001011111",
  20563=>"001011000",
  20564=>"011100111",
  20565=>"101100111",
  20566=>"111101000",
  20567=>"110111011",
  20568=>"111101100",
  20569=>"111010000",
  20570=>"111001100",
  20571=>"010000000",
  20572=>"111001110",
  20573=>"010100010",
  20574=>"011011100",
  20575=>"000110001",
  20576=>"000000000",
  20577=>"011100111",
  20578=>"101100000",
  20579=>"010010101",
  20580=>"101011101",
  20581=>"000100101",
  20582=>"011000000",
  20583=>"010111110",
  20584=>"011110011",
  20585=>"110110011",
  20586=>"101111011",
  20587=>"001100000",
  20588=>"100111000",
  20589=>"011101100",
  20590=>"011110000",
  20591=>"111010011",
  20592=>"000011000",
  20593=>"010100101",
  20594=>"111111111",
  20595=>"100100100",
  20596=>"101111001",
  20597=>"111000100",
  20598=>"011110001",
  20599=>"110010001",
  20600=>"000111100",
  20601=>"010000011",
  20602=>"001111100",
  20603=>"001010000",
  20604=>"100000011",
  20605=>"111101010",
  20606=>"011100100",
  20607=>"000000000",
  20608=>"111001110",
  20609=>"110001010",
  20610=>"100011111",
  20611=>"110000100",
  20612=>"110110100",
  20613=>"111100100",
  20614=>"111111110",
  20615=>"011101100",
  20616=>"111100110",
  20617=>"111100010",
  20618=>"110001110",
  20619=>"011000000",
  20620=>"101111110",
  20621=>"000010000",
  20622=>"011111011",
  20623=>"111100110",
  20624=>"001001011",
  20625=>"001101000",
  20626=>"010101011",
  20627=>"001000010",
  20628=>"000100001",
  20629=>"111010010",
  20630=>"110100011",
  20631=>"010110111",
  20632=>"011011000",
  20633=>"110111101",
  20634=>"000000101",
  20635=>"011100110",
  20636=>"011101101",
  20637=>"101000101",
  20638=>"010100101",
  20639=>"110000000",
  20640=>"110111100",
  20641=>"100001100",
  20642=>"110011110",
  20643=>"000100010",
  20644=>"011011001",
  20645=>"111011000",
  20646=>"000111111",
  20647=>"101100111",
  20648=>"001110100",
  20649=>"100110000",
  20650=>"111101110",
  20651=>"000010011",
  20652=>"010101101",
  20653=>"001011000",
  20654=>"101000100",
  20655=>"111111101",
  20656=>"011010000",
  20657=>"100001100",
  20658=>"010010011",
  20659=>"011110110",
  20660=>"111011110",
  20661=>"010000010",
  20662=>"011111010",
  20663=>"000100000",
  20664=>"001001111",
  20665=>"000000000",
  20666=>"101000011",
  20667=>"111101111",
  20668=>"000010000",
  20669=>"111101101",
  20670=>"010110001",
  20671=>"110101111",
  20672=>"101011101",
  20673=>"010110011",
  20674=>"001010000",
  20675=>"011111010",
  20676=>"111111010",
  20677=>"100111011",
  20678=>"000101101",
  20679=>"001100100",
  20680=>"000100011",
  20681=>"010011010",
  20682=>"000000000",
  20683=>"101110010",
  20684=>"011100100",
  20685=>"111100111",
  20686=>"010100100",
  20687=>"001111011",
  20688=>"101001111",
  20689=>"011010110",
  20690=>"001110000",
  20691=>"100000001",
  20692=>"101100110",
  20693=>"111010001",
  20694=>"010011011",
  20695=>"101000110",
  20696=>"000000101",
  20697=>"000010011",
  20698=>"101111001",
  20699=>"001100000",
  20700=>"011010101",
  20701=>"101101000",
  20702=>"111101001",
  20703=>"000011011",
  20704=>"111010100",
  20705=>"100000100",
  20706=>"000011100",
  20707=>"110011110",
  20708=>"000001100",
  20709=>"110000110",
  20710=>"000011000",
  20711=>"100111010",
  20712=>"111111111",
  20713=>"000000110",
  20714=>"000011011",
  20715=>"011010101",
  20716=>"101011010",
  20717=>"101101111",
  20718=>"101011110",
  20719=>"111100111",
  20720=>"011010011",
  20721=>"101111110",
  20722=>"101100100",
  20723=>"100110011",
  20724=>"111011100",
  20725=>"011001111",
  20726=>"000011110",
  20727=>"000010001",
  20728=>"010001010",
  20729=>"000010100",
  20730=>"010010111",
  20731=>"101111110",
  20732=>"000101101",
  20733=>"011101110",
  20734=>"100111000",
  20735=>"000000000",
  20736=>"011110000",
  20737=>"100100010",
  20738=>"001111100",
  20739=>"111111000",
  20740=>"110000001",
  20741=>"101010011",
  20742=>"101001000",
  20743=>"010000010",
  20744=>"001000100",
  20745=>"111100110",
  20746=>"111100001",
  20747=>"111101100",
  20748=>"101100101",
  20749=>"110100000",
  20750=>"111100000",
  20751=>"011000000",
  20752=>"000110001",
  20753=>"001110000",
  20754=>"110000110",
  20755=>"111011110",
  20756=>"011101011",
  20757=>"100001000",
  20758=>"101100001",
  20759=>"100000010",
  20760=>"100101110",
  20761=>"111101000",
  20762=>"000001100",
  20763=>"011010100",
  20764=>"010001000",
  20765=>"010111011",
  20766=>"111110101",
  20767=>"011111100",
  20768=>"111011101",
  20769=>"001010110",
  20770=>"110111101",
  20771=>"001101011",
  20772=>"100100110",
  20773=>"001010000",
  20774=>"011101110",
  20775=>"001101110",
  20776=>"010001011",
  20777=>"100000110",
  20778=>"100100100",
  20779=>"100100010",
  20780=>"001001000",
  20781=>"001000100",
  20782=>"000000100",
  20783=>"010001000",
  20784=>"001011010",
  20785=>"111001001",
  20786=>"111011101",
  20787=>"000010010",
  20788=>"101011001",
  20789=>"000000010",
  20790=>"001010001",
  20791=>"101101101",
  20792=>"000000100",
  20793=>"011100100",
  20794=>"111000010",
  20795=>"100111000",
  20796=>"010101011",
  20797=>"000001111",
  20798=>"011111110",
  20799=>"111011101",
  20800=>"111100110",
  20801=>"000010111",
  20802=>"100011101",
  20803=>"010101010",
  20804=>"111100011",
  20805=>"000011001",
  20806=>"011000001",
  20807=>"001011011",
  20808=>"001001111",
  20809=>"011111001",
  20810=>"101100110",
  20811=>"010010010",
  20812=>"011110100",
  20813=>"110011001",
  20814=>"111110101",
  20815=>"111010010",
  20816=>"000110101",
  20817=>"000001101",
  20818=>"111110000",
  20819=>"001000111",
  20820=>"011110111",
  20821=>"101101100",
  20822=>"100001110",
  20823=>"100101100",
  20824=>"001010011",
  20825=>"000101101",
  20826=>"011011000",
  20827=>"010000010",
  20828=>"010000100",
  20829=>"111011111",
  20830=>"111011100",
  20831=>"101010010",
  20832=>"111010010",
  20833=>"011111101",
  20834=>"000000100",
  20835=>"011100100",
  20836=>"100101000",
  20837=>"010101100",
  20838=>"101010111",
  20839=>"011010001",
  20840=>"001001001",
  20841=>"110011011",
  20842=>"111010101",
  20843=>"010110101",
  20844=>"101100011",
  20845=>"100001100",
  20846=>"000100001",
  20847=>"110001100",
  20848=>"000000100",
  20849=>"100010111",
  20850=>"110110011",
  20851=>"101100001",
  20852=>"100110110",
  20853=>"010100001",
  20854=>"100111000",
  20855=>"000000010",
  20856=>"100101000",
  20857=>"110001000",
  20858=>"010010111",
  20859=>"011000000",
  20860=>"111110001",
  20861=>"111011100",
  20862=>"111010000",
  20863=>"010101001",
  20864=>"111011111",
  20865=>"010100010",
  20866=>"110100001",
  20867=>"101000001",
  20868=>"001010101",
  20869=>"010010101",
  20870=>"010111100",
  20871=>"011111111",
  20872=>"000001110",
  20873=>"101000101",
  20874=>"111111011",
  20875=>"011100111",
  20876=>"110111010",
  20877=>"010100001",
  20878=>"011111101",
  20879=>"010100110",
  20880=>"001000101",
  20881=>"110001000",
  20882=>"111101010",
  20883=>"010000010",
  20884=>"011011001",
  20885=>"011111100",
  20886=>"000000010",
  20887=>"001001100",
  20888=>"111111111",
  20889=>"010101111",
  20890=>"110111111",
  20891=>"000111001",
  20892=>"100111100",
  20893=>"000010111",
  20894=>"000011111",
  20895=>"001110000",
  20896=>"100011100",
  20897=>"110100110",
  20898=>"101001101",
  20899=>"000001111",
  20900=>"001101011",
  20901=>"110000101",
  20902=>"110000001",
  20903=>"100010010",
  20904=>"110001101",
  20905=>"110110100",
  20906=>"111100011",
  20907=>"000111100",
  20908=>"111100111",
  20909=>"000000111",
  20910=>"111001100",
  20911=>"101110011",
  20912=>"111011011",
  20913=>"111110011",
  20914=>"001101001",
  20915=>"010101000",
  20916=>"111011100",
  20917=>"011011111",
  20918=>"110011110",
  20919=>"010110101",
  20920=>"001001100",
  20921=>"001000100",
  20922=>"001001000",
  20923=>"011111110",
  20924=>"001000000",
  20925=>"111101110",
  20926=>"010101110",
  20927=>"110101100",
  20928=>"111001010",
  20929=>"101011111",
  20930=>"001011011",
  20931=>"000100010",
  20932=>"010010010",
  20933=>"001000010",
  20934=>"101101110",
  20935=>"101111100",
  20936=>"011110111",
  20937=>"110110101",
  20938=>"111100111",
  20939=>"001011010",
  20940=>"000110011",
  20941=>"011001111",
  20942=>"110111101",
  20943=>"001010100",
  20944=>"110001001",
  20945=>"001000110",
  20946=>"110010000",
  20947=>"010000010",
  20948=>"111111011",
  20949=>"111101110",
  20950=>"011001100",
  20951=>"111011100",
  20952=>"010000011",
  20953=>"110010100",
  20954=>"101110100",
  20955=>"110111001",
  20956=>"001111010",
  20957=>"111100100",
  20958=>"001000100",
  20959=>"000000101",
  20960=>"001111010",
  20961=>"111010010",
  20962=>"100110000",
  20963=>"101110001",
  20964=>"011000100",
  20965=>"000001010",
  20966=>"101011000",
  20967=>"000001100",
  20968=>"110111111",
  20969=>"001011100",
  20970=>"100010111",
  20971=>"111100111",
  20972=>"111111011",
  20973=>"111011100",
  20974=>"110001100",
  20975=>"010011100",
  20976=>"010101111",
  20977=>"001010111",
  20978=>"010111101",
  20979=>"000000110",
  20980=>"111001010",
  20981=>"000100110",
  20982=>"110111111",
  20983=>"001001100",
  20984=>"100001111",
  20985=>"111100010",
  20986=>"101100010",
  20987=>"000101110",
  20988=>"111001101",
  20989=>"001100111",
  20990=>"110111010",
  20991=>"001111001",
  20992=>"001000000",
  20993=>"010100000",
  20994=>"110010110",
  20995=>"010100111",
  20996=>"011111111",
  20997=>"010111110",
  20998=>"001111100",
  20999=>"111001000",
  21000=>"110011000",
  21001=>"111111101",
  21002=>"010011010",
  21003=>"010100100",
  21004=>"101010000",
  21005=>"000010000",
  21006=>"000010100",
  21007=>"100111100",
  21008=>"100100011",
  21009=>"111000110",
  21010=>"011001101",
  21011=>"001101000",
  21012=>"010011010",
  21013=>"101110110",
  21014=>"000010001",
  21015=>"011011011",
  21016=>"010111000",
  21017=>"000110110",
  21018=>"111100110",
  21019=>"101011100",
  21020=>"001110111",
  21021=>"001010011",
  21022=>"000000011",
  21023=>"001110011",
  21024=>"101001111",
  21025=>"010101100",
  21026=>"111010000",
  21027=>"010000101",
  21028=>"111011111",
  21029=>"001100111",
  21030=>"110111001",
  21031=>"010000001",
  21032=>"101001111",
  21033=>"001001000",
  21034=>"000010011",
  21035=>"010000101",
  21036=>"000101001",
  21037=>"110110010",
  21038=>"001100010",
  21039=>"011101010",
  21040=>"101111110",
  21041=>"001111010",
  21042=>"010111111",
  21043=>"101111111",
  21044=>"011111000",
  21045=>"001010111",
  21046=>"000010100",
  21047=>"100101011",
  21048=>"100101110",
  21049=>"110010100",
  21050=>"111111111",
  21051=>"111001101",
  21052=>"010110110",
  21053=>"000010011",
  21054=>"110001010",
  21055=>"100110001",
  21056=>"001011101",
  21057=>"001000101",
  21058=>"100101001",
  21059=>"111110110",
  21060=>"100111101",
  21061=>"010111010",
  21062=>"010111110",
  21063=>"010010110",
  21064=>"000100101",
  21065=>"110100010",
  21066=>"010111101",
  21067=>"010010111",
  21068=>"101100101",
  21069=>"111010101",
  21070=>"111111100",
  21071=>"111010100",
  21072=>"010111000",
  21073=>"001001111",
  21074=>"111111110",
  21075=>"010100000",
  21076=>"001111110",
  21077=>"011101110",
  21078=>"100011110",
  21079=>"000011000",
  21080=>"011011101",
  21081=>"111100111",
  21082=>"111111101",
  21083=>"001000100",
  21084=>"011000100",
  21085=>"001111101",
  21086=>"100111100",
  21087=>"010100101",
  21088=>"000000001",
  21089=>"110110111",
  21090=>"011001011",
  21091=>"111110100",
  21092=>"011001011",
  21093=>"100000110",
  21094=>"000101111",
  21095=>"010111011",
  21096=>"101111100",
  21097=>"011000000",
  21098=>"110000010",
  21099=>"001010011",
  21100=>"010110000",
  21101=>"010100100",
  21102=>"110110111",
  21103=>"011010111",
  21104=>"111101011",
  21105=>"010110110",
  21106=>"110111011",
  21107=>"000011111",
  21108=>"011001110",
  21109=>"001000010",
  21110=>"100100100",
  21111=>"001010100",
  21112=>"111110000",
  21113=>"010100111",
  21114=>"101111110",
  21115=>"111001001",
  21116=>"111111000",
  21117=>"100111010",
  21118=>"110000100",
  21119=>"010010110",
  21120=>"100000100",
  21121=>"011111110",
  21122=>"001010100",
  21123=>"010010101",
  21124=>"110101010",
  21125=>"110111101",
  21126=>"101001000",
  21127=>"101100100",
  21128=>"000101101",
  21129=>"001101010",
  21130=>"100000111",
  21131=>"110000001",
  21132=>"010101000",
  21133=>"111110010",
  21134=>"000000101",
  21135=>"011111100",
  21136=>"110100100",
  21137=>"100011001",
  21138=>"010010111",
  21139=>"110100000",
  21140=>"000111001",
  21141=>"111101100",
  21142=>"000011000",
  21143=>"011110010",
  21144=>"111110100",
  21145=>"010100100",
  21146=>"101010000",
  21147=>"000100001",
  21148=>"000010010",
  21149=>"110100010",
  21150=>"100001000",
  21151=>"000001011",
  21152=>"000011000",
  21153=>"011011110",
  21154=>"101101110",
  21155=>"111001110",
  21156=>"101111111",
  21157=>"000100011",
  21158=>"110110010",
  21159=>"010000011",
  21160=>"001010100",
  21161=>"000101000",
  21162=>"000111101",
  21163=>"011100100",
  21164=>"111000011",
  21165=>"101010001",
  21166=>"011111111",
  21167=>"111001011",
  21168=>"011010111",
  21169=>"001101100",
  21170=>"110101110",
  21171=>"111001010",
  21172=>"010110011",
  21173=>"110100101",
  21174=>"110101110",
  21175=>"010111001",
  21176=>"011110001",
  21177=>"001110100",
  21178=>"111001010",
  21179=>"001000100",
  21180=>"001111111",
  21181=>"000011001",
  21182=>"000111110",
  21183=>"010111011",
  21184=>"100000010",
  21185=>"001111011",
  21186=>"010010100",
  21187=>"010011100",
  21188=>"110010100",
  21189=>"111010110",
  21190=>"101010100",
  21191=>"000101110",
  21192=>"111111011",
  21193=>"100000100",
  21194=>"011001100",
  21195=>"001101111",
  21196=>"001010010",
  21197=>"011110001",
  21198=>"011001000",
  21199=>"011000010",
  21200=>"110111011",
  21201=>"101001000",
  21202=>"000010000",
  21203=>"000000010",
  21204=>"000110100",
  21205=>"101100111",
  21206=>"010110101",
  21207=>"111011101",
  21208=>"111001011",
  21209=>"011000010",
  21210=>"110001010",
  21211=>"111111010",
  21212=>"010000010",
  21213=>"000011100",
  21214=>"111000011",
  21215=>"000100111",
  21216=>"010010101",
  21217=>"001110010",
  21218=>"000100010",
  21219=>"111111100",
  21220=>"011101100",
  21221=>"100010011",
  21222=>"110001101",
  21223=>"101000110",
  21224=>"111111011",
  21225=>"101011010",
  21226=>"010100001",
  21227=>"110011100",
  21228=>"001010011",
  21229=>"100111000",
  21230=>"100000001",
  21231=>"010100100",
  21232=>"101001100",
  21233=>"000111001",
  21234=>"000011100",
  21235=>"101111000",
  21236=>"110111001",
  21237=>"101010001",
  21238=>"010110000",
  21239=>"010011000",
  21240=>"010100000",
  21241=>"010000011",
  21242=>"110100101",
  21243=>"010111110",
  21244=>"011000001",
  21245=>"111111111",
  21246=>"001101101",
  21247=>"010011000",
  21248=>"111011000",
  21249=>"101000101",
  21250=>"011111111",
  21251=>"001101111",
  21252=>"000101110",
  21253=>"000100111",
  21254=>"000001000",
  21255=>"110000010",
  21256=>"001001001",
  21257=>"101110111",
  21258=>"011000010",
  21259=>"110101010",
  21260=>"001011000",
  21261=>"000111000",
  21262=>"111000001",
  21263=>"011001010",
  21264=>"001000101",
  21265=>"100111100",
  21266=>"100110001",
  21267=>"001111000",
  21268=>"011000111",
  21269=>"100100010",
  21270=>"001000100",
  21271=>"001101110",
  21272=>"101110110",
  21273=>"111110001",
  21274=>"011000000",
  21275=>"110010111",
  21276=>"100011111",
  21277=>"011101101",
  21278=>"000111111",
  21279=>"010110010",
  21280=>"011110111",
  21281=>"000010000",
  21282=>"100000001",
  21283=>"000100001",
  21284=>"100010110",
  21285=>"000111111",
  21286=>"101110110",
  21287=>"001111000",
  21288=>"110111001",
  21289=>"000010100",
  21290=>"101001101",
  21291=>"101101010",
  21292=>"101010111",
  21293=>"010010010",
  21294=>"111101000",
  21295=>"010100101",
  21296=>"101101110",
  21297=>"010010001",
  21298=>"010011011",
  21299=>"011001000",
  21300=>"010011111",
  21301=>"011011011",
  21302=>"110000010",
  21303=>"010010000",
  21304=>"001000010",
  21305=>"111111010",
  21306=>"001101011",
  21307=>"100011010",
  21308=>"000100101",
  21309=>"001101011",
  21310=>"001011001",
  21311=>"100011111",
  21312=>"001001100",
  21313=>"111111011",
  21314=>"111011111",
  21315=>"111011110",
  21316=>"100100100",
  21317=>"011000110",
  21318=>"010001011",
  21319=>"110111101",
  21320=>"110001100",
  21321=>"111100001",
  21322=>"010101010",
  21323=>"010011011",
  21324=>"011101011",
  21325=>"000101010",
  21326=>"001001101",
  21327=>"111010110",
  21328=>"010000000",
  21329=>"000000111",
  21330=>"011000110",
  21331=>"001100100",
  21332=>"011011110",
  21333=>"011100000",
  21334=>"001000001",
  21335=>"010101111",
  21336=>"000100110",
  21337=>"001001010",
  21338=>"011001001",
  21339=>"100000100",
  21340=>"100000101",
  21341=>"111101101",
  21342=>"001111100",
  21343=>"111110111",
  21344=>"100111011",
  21345=>"110010010",
  21346=>"000010000",
  21347=>"110101111",
  21348=>"101111101",
  21349=>"110011111",
  21350=>"100000011",
  21351=>"111101110",
  21352=>"111000101",
  21353=>"110111101",
  21354=>"101000010",
  21355=>"101000000",
  21356=>"001001111",
  21357=>"011000110",
  21358=>"111110111",
  21359=>"000111011",
  21360=>"010111000",
  21361=>"000110111",
  21362=>"010110101",
  21363=>"011010100",
  21364=>"111110110",
  21365=>"101000110",
  21366=>"100111110",
  21367=>"100011011",
  21368=>"100101110",
  21369=>"001101000",
  21370=>"010111011",
  21371=>"110111110",
  21372=>"101110001",
  21373=>"011001100",
  21374=>"001011110",
  21375=>"001101111",
  21376=>"101100011",
  21377=>"011011000",
  21378=>"110101111",
  21379=>"100001111",
  21380=>"101011001",
  21381=>"100110111",
  21382=>"000010000",
  21383=>"010011100",
  21384=>"111100111",
  21385=>"110011101",
  21386=>"111001110",
  21387=>"101000101",
  21388=>"100111001",
  21389=>"111101001",
  21390=>"110011100",
  21391=>"010110111",
  21392=>"111101000",
  21393=>"111101100",
  21394=>"001011000",
  21395=>"101111000",
  21396=>"011111001",
  21397=>"010011100",
  21398=>"010000000",
  21399=>"010101000",
  21400=>"011000110",
  21401=>"101101001",
  21402=>"110000000",
  21403=>"001000101",
  21404=>"011001011",
  21405=>"000111101",
  21406=>"110010101",
  21407=>"100000000",
  21408=>"100110101",
  21409=>"100101101",
  21410=>"010111001",
  21411=>"000001001",
  21412=>"111110111",
  21413=>"001111111",
  21414=>"011011000",
  21415=>"010100111",
  21416=>"010110010",
  21417=>"000000011",
  21418=>"101101101",
  21419=>"101100110",
  21420=>"110000011",
  21421=>"000111110",
  21422=>"111011101",
  21423=>"010010001",
  21424=>"101000101",
  21425=>"100100010",
  21426=>"101010110",
  21427=>"010001111",
  21428=>"000000111",
  21429=>"110001100",
  21430=>"011111011",
  21431=>"111110110",
  21432=>"001101101",
  21433=>"110100011",
  21434=>"110100001",
  21435=>"011111001",
  21436=>"010100010",
  21437=>"100001000",
  21438=>"000000111",
  21439=>"100011010",
  21440=>"011011001",
  21441=>"000111011",
  21442=>"000000011",
  21443=>"000100010",
  21444=>"101111001",
  21445=>"000111110",
  21446=>"001000110",
  21447=>"000000100",
  21448=>"001010100",
  21449=>"011011010",
  21450=>"001111100",
  21451=>"011000110",
  21452=>"001000011",
  21453=>"001000000",
  21454=>"100011011",
  21455=>"110110100",
  21456=>"111011010",
  21457=>"000111010",
  21458=>"011100000",
  21459=>"111100010",
  21460=>"000000110",
  21461=>"110100101",
  21462=>"100010111",
  21463=>"011000101",
  21464=>"010011111",
  21465=>"001000001",
  21466=>"001111101",
  21467=>"000000101",
  21468=>"000111111",
  21469=>"110101100",
  21470=>"100110110",
  21471=>"101100001",
  21472=>"100110010",
  21473=>"100101011",
  21474=>"000100001",
  21475=>"110010010",
  21476=>"111100100",
  21477=>"001011110",
  21478=>"011100100",
  21479=>"011000011",
  21480=>"000000110",
  21481=>"011011000",
  21482=>"111111011",
  21483=>"111101111",
  21484=>"001011000",
  21485=>"110101110",
  21486=>"001001110",
  21487=>"000010100",
  21488=>"100101000",
  21489=>"111000000",
  21490=>"110001000",
  21491=>"111011111",
  21492=>"011111011",
  21493=>"111011111",
  21494=>"110011110",
  21495=>"100110001",
  21496=>"101001000",
  21497=>"101001100",
  21498=>"000110000",
  21499=>"110001101",
  21500=>"010100011",
  21501=>"110010010",
  21502=>"001010000",
  21503=>"101100111",
  21504=>"011110110",
  21505=>"011110110",
  21506=>"110011010",
  21507=>"111011111",
  21508=>"011011010",
  21509=>"101101111",
  21510=>"011110100",
  21511=>"001100100",
  21512=>"010011000",
  21513=>"001111000",
  21514=>"111101011",
  21515=>"100110110",
  21516=>"000001010",
  21517=>"001101011",
  21518=>"101010010",
  21519=>"110100010",
  21520=>"100001111",
  21521=>"110001011",
  21522=>"100101100",
  21523=>"111110010",
  21524=>"110001111",
  21525=>"010101010",
  21526=>"001010011",
  21527=>"010010010",
  21528=>"101110011",
  21529=>"000011101",
  21530=>"110010101",
  21531=>"111001101",
  21532=>"000011111",
  21533=>"000111000",
  21534=>"111110011",
  21535=>"001110101",
  21536=>"100111111",
  21537=>"111100010",
  21538=>"101000010",
  21539=>"110011111",
  21540=>"011101010",
  21541=>"100100110",
  21542=>"000011101",
  21543=>"110011101",
  21544=>"111100101",
  21545=>"000001100",
  21546=>"101010110",
  21547=>"011010001",
  21548=>"100000010",
  21549=>"001101111",
  21550=>"010000011",
  21551=>"011001000",
  21552=>"100101111",
  21553=>"110011100",
  21554=>"101001110",
  21555=>"101001010",
  21556=>"011000110",
  21557=>"110001000",
  21558=>"100001001",
  21559=>"111010111",
  21560=>"001100000",
  21561=>"111111111",
  21562=>"000010011",
  21563=>"111110010",
  21564=>"011000101",
  21565=>"111100111",
  21566=>"111100000",
  21567=>"010110000",
  21568=>"100010101",
  21569=>"000110011",
  21570=>"011000010",
  21571=>"100110000",
  21572=>"011011111",
  21573=>"110000100",
  21574=>"000011110",
  21575=>"011000100",
  21576=>"101011101",
  21577=>"011000100",
  21578=>"011101001",
  21579=>"000101000",
  21580=>"001100111",
  21581=>"111001101",
  21582=>"110100000",
  21583=>"111010010",
  21584=>"100000000",
  21585=>"101110011",
  21586=>"110001011",
  21587=>"010111010",
  21588=>"111001101",
  21589=>"010111100",
  21590=>"110000110",
  21591=>"001110010",
  21592=>"010101000",
  21593=>"101010000",
  21594=>"010100000",
  21595=>"010011110",
  21596=>"100100011",
  21597=>"010000011",
  21598=>"100101101",
  21599=>"011111100",
  21600=>"100110110",
  21601=>"011110010",
  21602=>"001101100",
  21603=>"010110101",
  21604=>"101001000",
  21605=>"001001000",
  21606=>"110100001",
  21607=>"101000100",
  21608=>"101001110",
  21609=>"110110011",
  21610=>"010100100",
  21611=>"100001011",
  21612=>"001001100",
  21613=>"010011010",
  21614=>"011010101",
  21615=>"101000011",
  21616=>"101000010",
  21617=>"000011001",
  21618=>"011101110",
  21619=>"101111100",
  21620=>"101010000",
  21621=>"000100111",
  21622=>"000000010",
  21623=>"100001101",
  21624=>"001010110",
  21625=>"100001011",
  21626=>"111111011",
  21627=>"010111100",
  21628=>"100100101",
  21629=>"000000100",
  21630=>"101101101",
  21631=>"110111101",
  21632=>"010100001",
  21633=>"001111100",
  21634=>"001100000",
  21635=>"100100100",
  21636=>"001101111",
  21637=>"100110010",
  21638=>"011110101",
  21639=>"101000100",
  21640=>"001011011",
  21641=>"000011101",
  21642=>"001011000",
  21643=>"111111111",
  21644=>"100010110",
  21645=>"110010100",
  21646=>"111000101",
  21647=>"011110001",
  21648=>"111100110",
  21649=>"011100001",
  21650=>"111001001",
  21651=>"001001100",
  21652=>"000010111",
  21653=>"111001000",
  21654=>"110000000",
  21655=>"001101101",
  21656=>"000010000",
  21657=>"000000010",
  21658=>"001011110",
  21659=>"111001000",
  21660=>"000011000",
  21661=>"101101100",
  21662=>"100111001",
  21663=>"101000000",
  21664=>"101111100",
  21665=>"100001000",
  21666=>"110000001",
  21667=>"100000100",
  21668=>"011101010",
  21669=>"100010101",
  21670=>"011110010",
  21671=>"101111000",
  21672=>"011011111",
  21673=>"000111110",
  21674=>"010001100",
  21675=>"111111010",
  21676=>"011011010",
  21677=>"001100111",
  21678=>"011100111",
  21679=>"001011111",
  21680=>"100001100",
  21681=>"100011000",
  21682=>"100001110",
  21683=>"001101100",
  21684=>"101101100",
  21685=>"111100101",
  21686=>"000011000",
  21687=>"001111001",
  21688=>"010100100",
  21689=>"000010000",
  21690=>"000011110",
  21691=>"101100000",
  21692=>"010100010",
  21693=>"100101001",
  21694=>"000011001",
  21695=>"100111000",
  21696=>"111110000",
  21697=>"011011101",
  21698=>"001000011",
  21699=>"011001000",
  21700=>"011011011",
  21701=>"000001011",
  21702=>"101101110",
  21703=>"111110001",
  21704=>"001111000",
  21705=>"010011011",
  21706=>"110001000",
  21707=>"111011101",
  21708=>"110100000",
  21709=>"110000101",
  21710=>"011110111",
  21711=>"011001001",
  21712=>"000101100",
  21713=>"110100011",
  21714=>"111011111",
  21715=>"001000010",
  21716=>"011010101",
  21717=>"011101110",
  21718=>"001110101",
  21719=>"100110101",
  21720=>"010011110",
  21721=>"001100000",
  21722=>"111010101",
  21723=>"110111011",
  21724=>"101010011",
  21725=>"001111010",
  21726=>"001100001",
  21727=>"100101000",
  21728=>"001101101",
  21729=>"000110111",
  21730=>"111101101",
  21731=>"000110010",
  21732=>"011100011",
  21733=>"010011100",
  21734=>"100010101",
  21735=>"111000101",
  21736=>"000110011",
  21737=>"110011110",
  21738=>"101001000",
  21739=>"100000100",
  21740=>"001001000",
  21741=>"000011001",
  21742=>"010011010",
  21743=>"010011010",
  21744=>"000101111",
  21745=>"000000011",
  21746=>"000010101",
  21747=>"001001010",
  21748=>"110010111",
  21749=>"101001110",
  21750=>"101111000",
  21751=>"000001000",
  21752=>"100011101",
  21753=>"011111100",
  21754=>"111111101",
  21755=>"111011011",
  21756=>"111100100",
  21757=>"010000101",
  21758=>"100111010",
  21759=>"001110111",
  21760=>"101001000",
  21761=>"100000100",
  21762=>"001111001",
  21763=>"010010010",
  21764=>"100000011",
  21765=>"101110001",
  21766=>"000011100",
  21767=>"101100000",
  21768=>"011001011",
  21769=>"000010010",
  21770=>"010111111",
  21771=>"111111010",
  21772=>"011101000",
  21773=>"010010011",
  21774=>"100010011",
  21775=>"100000101",
  21776=>"001011111",
  21777=>"000001111",
  21778=>"100101100",
  21779=>"110001010",
  21780=>"110011110",
  21781=>"110110000",
  21782=>"000001000",
  21783=>"001001100",
  21784=>"000111110",
  21785=>"111000000",
  21786=>"010001011",
  21787=>"000010100",
  21788=>"011111101",
  21789=>"110100010",
  21790=>"010000000",
  21791=>"001000000",
  21792=>"011100001",
  21793=>"011000100",
  21794=>"110010111",
  21795=>"010110011",
  21796=>"111010100",
  21797=>"011010110",
  21798=>"011001001",
  21799=>"110010100",
  21800=>"000000011",
  21801=>"110110000",
  21802=>"001101010",
  21803=>"001001100",
  21804=>"110001000",
  21805=>"011100101",
  21806=>"001110100",
  21807=>"000011010",
  21808=>"000110000",
  21809=>"001111111",
  21810=>"011001101",
  21811=>"111111111",
  21812=>"000000101",
  21813=>"100110010",
  21814=>"011000110",
  21815=>"110010101",
  21816=>"000100001",
  21817=>"001101111",
  21818=>"010110111",
  21819=>"100010110",
  21820=>"101001010",
  21821=>"110111100",
  21822=>"000011000",
  21823=>"011101101",
  21824=>"111110100",
  21825=>"000100100",
  21826=>"100111110",
  21827=>"101010001",
  21828=>"000010111",
  21829=>"000010010",
  21830=>"011000010",
  21831=>"111000011",
  21832=>"100001011",
  21833=>"100000001",
  21834=>"001111101",
  21835=>"000001110",
  21836=>"010010111",
  21837=>"100100010",
  21838=>"010100010",
  21839=>"111101101",
  21840=>"110110101",
  21841=>"010110010",
  21842=>"000101101",
  21843=>"010111010",
  21844=>"101011000",
  21845=>"010110111",
  21846=>"101111101",
  21847=>"010101101",
  21848=>"001000000",
  21849=>"110000001",
  21850=>"010001101",
  21851=>"001110111",
  21852=>"011111100",
  21853=>"110100100",
  21854=>"111011110",
  21855=>"011111110",
  21856=>"110110000",
  21857=>"010000000",
  21858=>"101111101",
  21859=>"010011100",
  21860=>"101111011",
  21861=>"010011011",
  21862=>"100000001",
  21863=>"001110010",
  21864=>"111101000",
  21865=>"110001100",
  21866=>"111011011",
  21867=>"100010011",
  21868=>"001101111",
  21869=>"111111101",
  21870=>"010010110",
  21871=>"011100111",
  21872=>"000100101",
  21873=>"011101110",
  21874=>"010010101",
  21875=>"010111011",
  21876=>"001011101",
  21877=>"101100001",
  21878=>"000000110",
  21879=>"001111110",
  21880=>"001001101",
  21881=>"100110110",
  21882=>"100001101",
  21883=>"110001101",
  21884=>"011010001",
  21885=>"100001000",
  21886=>"100110000",
  21887=>"111111110",
  21888=>"111001101",
  21889=>"101111101",
  21890=>"001101010",
  21891=>"110011111",
  21892=>"011001111",
  21893=>"110011000",
  21894=>"001000111",
  21895=>"000110110",
  21896=>"011000010",
  21897=>"100001110",
  21898=>"000011111",
  21899=>"100011000",
  21900=>"101100101",
  21901=>"101111001",
  21902=>"000111000",
  21903=>"100011101",
  21904=>"000111001",
  21905=>"001111001",
  21906=>"110010011",
  21907=>"010000001",
  21908=>"111010011",
  21909=>"110110110",
  21910=>"011101000",
  21911=>"010101111",
  21912=>"010110111",
  21913=>"100101101",
  21914=>"101110011",
  21915=>"100111001",
  21916=>"000010111",
  21917=>"010110011",
  21918=>"010011000",
  21919=>"000110110",
  21920=>"010010011",
  21921=>"010001111",
  21922=>"101100101",
  21923=>"100000011",
  21924=>"001110001",
  21925=>"011100010",
  21926=>"110011110",
  21927=>"011000101",
  21928=>"001001100",
  21929=>"000001011",
  21930=>"000010010",
  21931=>"001101100",
  21932=>"110101111",
  21933=>"001000101",
  21934=>"100000100",
  21935=>"001001100",
  21936=>"111110010",
  21937=>"011110010",
  21938=>"111001000",
  21939=>"010000010",
  21940=>"101100001",
  21941=>"101010101",
  21942=>"001111010",
  21943=>"000010001",
  21944=>"111110010",
  21945=>"100111000",
  21946=>"000010000",
  21947=>"000100111",
  21948=>"001000111",
  21949=>"100001101",
  21950=>"001010111",
  21951=>"110011111",
  21952=>"110101101",
  21953=>"100001100",
  21954=>"010101110",
  21955=>"110000100",
  21956=>"000100010",
  21957=>"110000000",
  21958=>"101000001",
  21959=>"011110111",
  21960=>"011001111",
  21961=>"110110110",
  21962=>"100000000",
  21963=>"111011010",
  21964=>"101010111",
  21965=>"101011110",
  21966=>"111110111",
  21967=>"010111001",
  21968=>"101011111",
  21969=>"000001100",
  21970=>"000110001",
  21971=>"111000110",
  21972=>"100001001",
  21973=>"100001000",
  21974=>"001001011",
  21975=>"000010010",
  21976=>"111110010",
  21977=>"100001000",
  21978=>"100111110",
  21979=>"000110001",
  21980=>"111001000",
  21981=>"000100111",
  21982=>"101011001",
  21983=>"010011010",
  21984=>"000011111",
  21985=>"111111011",
  21986=>"101001010",
  21987=>"101001011",
  21988=>"101100110",
  21989=>"111010001",
  21990=>"011101001",
  21991=>"000011001",
  21992=>"001111000",
  21993=>"100000001",
  21994=>"100100010",
  21995=>"011101101",
  21996=>"011100010",
  21997=>"110011101",
  21998=>"001001101",
  21999=>"011100001",
  22000=>"011101011",
  22001=>"110111111",
  22002=>"001101101",
  22003=>"000001100",
  22004=>"001000101",
  22005=>"001000101",
  22006=>"000001000",
  22007=>"101100101",
  22008=>"100100010",
  22009=>"101011100",
  22010=>"110001011",
  22011=>"110000101",
  22012=>"010010110",
  22013=>"000000010",
  22014=>"110101111",
  22015=>"000011010",
  22016=>"100011000",
  22017=>"011100101",
  22018=>"100100111",
  22019=>"110111010",
  22020=>"100111110",
  22021=>"000101100",
  22022=>"001111010",
  22023=>"010110010",
  22024=>"101010100",
  22025=>"001001101",
  22026=>"001101100",
  22027=>"000000100",
  22028=>"001001101",
  22029=>"101010000",
  22030=>"010110000",
  22031=>"001001011",
  22032=>"100100100",
  22033=>"111000000",
  22034=>"000011110",
  22035=>"111001001",
  22036=>"010000010",
  22037=>"101011111",
  22038=>"100111010",
  22039=>"010101010",
  22040=>"000011000",
  22041=>"110001111",
  22042=>"010100111",
  22043=>"100000110",
  22044=>"111110000",
  22045=>"110010100",
  22046=>"000110011",
  22047=>"111011110",
  22048=>"110000000",
  22049=>"110110110",
  22050=>"110111011",
  22051=>"100000100",
  22052=>"110101011",
  22053=>"100000100",
  22054=>"101000000",
  22055=>"001010111",
  22056=>"000011001",
  22057=>"101110100",
  22058=>"001111111",
  22059=>"010100011",
  22060=>"001111011",
  22061=>"000001110",
  22062=>"101011110",
  22063=>"000100000",
  22064=>"010001101",
  22065=>"001010000",
  22066=>"001101000",
  22067=>"100111000",
  22068=>"110111000",
  22069=>"000011100",
  22070=>"110101001",
  22071=>"101000011",
  22072=>"101001000",
  22073=>"001010110",
  22074=>"110011011",
  22075=>"001000010",
  22076=>"111111101",
  22077=>"100010100",
  22078=>"100000111",
  22079=>"110001101",
  22080=>"010010100",
  22081=>"010000111",
  22082=>"100010111",
  22083=>"000000001",
  22084=>"001101010",
  22085=>"000001110",
  22086=>"000011010",
  22087=>"001011010",
  22088=>"011000110",
  22089=>"010101111",
  22090=>"110100010",
  22091=>"000000101",
  22092=>"010110111",
  22093=>"001011010",
  22094=>"101001101",
  22095=>"110100010",
  22096=>"011101101",
  22097=>"100111101",
  22098=>"111011101",
  22099=>"100100000",
  22100=>"010101001",
  22101=>"010010000",
  22102=>"001011111",
  22103=>"101101001",
  22104=>"011110100",
  22105=>"011101001",
  22106=>"010100001",
  22107=>"011011110",
  22108=>"001100111",
  22109=>"001100011",
  22110=>"000011011",
  22111=>"100011111",
  22112=>"001011101",
  22113=>"001010001",
  22114=>"000111001",
  22115=>"110101101",
  22116=>"101110110",
  22117=>"100111100",
  22118=>"000000000",
  22119=>"000000001",
  22120=>"000111100",
  22121=>"001010110",
  22122=>"101010100",
  22123=>"001001001",
  22124=>"010001010",
  22125=>"000010111",
  22126=>"100111111",
  22127=>"101011000",
  22128=>"101101000",
  22129=>"011010011",
  22130=>"101111101",
  22131=>"001001001",
  22132=>"100000111",
  22133=>"010001100",
  22134=>"111110010",
  22135=>"100000001",
  22136=>"100011110",
  22137=>"010110001",
  22138=>"001110101",
  22139=>"001110001",
  22140=>"101000000",
  22141=>"110010010",
  22142=>"011011010",
  22143=>"011011010",
  22144=>"110101110",
  22145=>"000111111",
  22146=>"010101110",
  22147=>"000000011",
  22148=>"111001111",
  22149=>"111010000",
  22150=>"011010110",
  22151=>"101011001",
  22152=>"011100101",
  22153=>"000000101",
  22154=>"001001001",
  22155=>"111110101",
  22156=>"001000111",
  22157=>"100111111",
  22158=>"000001110",
  22159=>"011110100",
  22160=>"101000111",
  22161=>"101001101",
  22162=>"111011111",
  22163=>"101000110",
  22164=>"000000110",
  22165=>"101000000",
  22166=>"001100011",
  22167=>"000100100",
  22168=>"111100010",
  22169=>"101000110",
  22170=>"101111100",
  22171=>"111000010",
  22172=>"001100100",
  22173=>"101000111",
  22174=>"000010001",
  22175=>"000111100",
  22176=>"100101101",
  22177=>"110010100",
  22178=>"000111001",
  22179=>"000011111",
  22180=>"010111111",
  22181=>"011110010",
  22182=>"001101111",
  22183=>"100100110",
  22184=>"010000010",
  22185=>"001000000",
  22186=>"111111000",
  22187=>"000110001",
  22188=>"001010001",
  22189=>"001010111",
  22190=>"010110100",
  22191=>"100000011",
  22192=>"111000010",
  22193=>"000010101",
  22194=>"101010011",
  22195=>"101101101",
  22196=>"111101011",
  22197=>"001101100",
  22198=>"011001111",
  22199=>"110011111",
  22200=>"100010111",
  22201=>"111101101",
  22202=>"101010101",
  22203=>"100001101",
  22204=>"000110100",
  22205=>"000001011",
  22206=>"000011101",
  22207=>"111000100",
  22208=>"000111011",
  22209=>"000111111",
  22210=>"001011100",
  22211=>"100100001",
  22212=>"101100100",
  22213=>"000010010",
  22214=>"111011010",
  22215=>"010111000",
  22216=>"101011001",
  22217=>"100000101",
  22218=>"010010100",
  22219=>"010101011",
  22220=>"010010011",
  22221=>"100011111",
  22222=>"111111010",
  22223=>"001001000",
  22224=>"110011000",
  22225=>"010111001",
  22226=>"010000001",
  22227=>"010100111",
  22228=>"011100111",
  22229=>"100010110",
  22230=>"000101110",
  22231=>"101011010",
  22232=>"100101010",
  22233=>"011010100",
  22234=>"100101111",
  22235=>"000011010",
  22236=>"101000011",
  22237=>"000011101",
  22238=>"000001111",
  22239=>"100100101",
  22240=>"011110000",
  22241=>"111001011",
  22242=>"111000100",
  22243=>"111110011",
  22244=>"101111000",
  22245=>"100111100",
  22246=>"100000100",
  22247=>"111101001",
  22248=>"001000110",
  22249=>"000001100",
  22250=>"110111100",
  22251=>"110111000",
  22252=>"110100010",
  22253=>"101101000",
  22254=>"101000110",
  22255=>"000000011",
  22256=>"111110111",
  22257=>"010111101",
  22258=>"001100110",
  22259=>"000001011",
  22260=>"110010110",
  22261=>"000001110",
  22262=>"010111101",
  22263=>"111001110",
  22264=>"100100100",
  22265=>"100111001",
  22266=>"011000000",
  22267=>"111011000",
  22268=>"010101100",
  22269=>"000100111",
  22270=>"110000101",
  22271=>"101001100",
  22272=>"010101000",
  22273=>"000100000",
  22274=>"000111100",
  22275=>"000010000",
  22276=>"000011110",
  22277=>"110011010",
  22278=>"000101100",
  22279=>"011010010",
  22280=>"011001001",
  22281=>"000001111",
  22282=>"011111101",
  22283=>"000011000",
  22284=>"011101100",
  22285=>"110100101",
  22286=>"010111011",
  22287=>"001000001",
  22288=>"101001001",
  22289=>"001010000",
  22290=>"110010000",
  22291=>"101000101",
  22292=>"101001100",
  22293=>"111100111",
  22294=>"111000110",
  22295=>"000111101",
  22296=>"010110010",
  22297=>"001010011",
  22298=>"110111011",
  22299=>"101001111",
  22300=>"100100010",
  22301=>"000111111",
  22302=>"010001100",
  22303=>"010010101",
  22304=>"001011111",
  22305=>"100000000",
  22306=>"101011110",
  22307=>"110001011",
  22308=>"100000110",
  22309=>"111010101",
  22310=>"001001111",
  22311=>"110011101",
  22312=>"110001010",
  22313=>"000000110",
  22314=>"111101001",
  22315=>"111011100",
  22316=>"001110011",
  22317=>"111011110",
  22318=>"010110010",
  22319=>"110111110",
  22320=>"000110110",
  22321=>"100110111",
  22322=>"110101000",
  22323=>"110010011",
  22324=>"101001100",
  22325=>"011000101",
  22326=>"001101101",
  22327=>"100101010",
  22328=>"100010110",
  22329=>"011111000",
  22330=>"000100111",
  22331=>"000000000",
  22332=>"000111010",
  22333=>"011100000",
  22334=>"010110001",
  22335=>"010111101",
  22336=>"001101101",
  22337=>"111110110",
  22338=>"011000110",
  22339=>"011010000",
  22340=>"111010010",
  22341=>"000111010",
  22342=>"100100110",
  22343=>"101011110",
  22344=>"001101110",
  22345=>"100110011",
  22346=>"011101110",
  22347=>"000010101",
  22348=>"111001101",
  22349=>"110111000",
  22350=>"111010000",
  22351=>"111110001",
  22352=>"110111010",
  22353=>"001001101",
  22354=>"011111000",
  22355=>"110111100",
  22356=>"100000000",
  22357=>"111111010",
  22358=>"101010111",
  22359=>"001101010",
  22360=>"010111100",
  22361=>"010110010",
  22362=>"111101000",
  22363=>"001111101",
  22364=>"111101110",
  22365=>"010011001",
  22366=>"011001110",
  22367=>"011101101",
  22368=>"000100111",
  22369=>"110010100",
  22370=>"010011010",
  22371=>"100111100",
  22372=>"000001011",
  22373=>"011110001",
  22374=>"000011110",
  22375=>"101101110",
  22376=>"000010011",
  22377=>"011001101",
  22378=>"000011000",
  22379=>"100001000",
  22380=>"100010010",
  22381=>"001101011",
  22382=>"010111001",
  22383=>"110001111",
  22384=>"110011110",
  22385=>"101011100",
  22386=>"110101100",
  22387=>"011100000",
  22388=>"100111101",
  22389=>"111001111",
  22390=>"101111001",
  22391=>"111000001",
  22392=>"101011100",
  22393=>"111000110",
  22394=>"001010000",
  22395=>"100110111",
  22396=>"001001010",
  22397=>"101010110",
  22398=>"000110110",
  22399=>"101111101",
  22400=>"111101100",
  22401=>"101110101",
  22402=>"000011110",
  22403=>"010100010",
  22404=>"000001110",
  22405=>"000010111",
  22406=>"000000001",
  22407=>"000011001",
  22408=>"001110010",
  22409=>"111001011",
  22410=>"000001101",
  22411=>"000000100",
  22412=>"010001011",
  22413=>"101111110",
  22414=>"100111000",
  22415=>"101010011",
  22416=>"010010100",
  22417=>"100101011",
  22418=>"010001010",
  22419=>"101011111",
  22420=>"011000000",
  22421=>"010011010",
  22422=>"101110101",
  22423=>"101010011",
  22424=>"010100101",
  22425=>"100100110",
  22426=>"010100001",
  22427=>"100110001",
  22428=>"001100101",
  22429=>"110110010",
  22430=>"000001110",
  22431=>"011100110",
  22432=>"110000010",
  22433=>"010000010",
  22434=>"000111101",
  22435=>"011110001",
  22436=>"000100111",
  22437=>"011101111",
  22438=>"001011111",
  22439=>"000011100",
  22440=>"110111001",
  22441=>"011111101",
  22442=>"111001000",
  22443=>"111010001",
  22444=>"101000100",
  22445=>"110001101",
  22446=>"110110010",
  22447=>"110001111",
  22448=>"111101011",
  22449=>"010101010",
  22450=>"110111110",
  22451=>"001000001",
  22452=>"111110111",
  22453=>"010101111",
  22454=>"010100111",
  22455=>"000000011",
  22456=>"010100000",
  22457=>"000110001",
  22458=>"000001111",
  22459=>"111000101",
  22460=>"101001101",
  22461=>"100000101",
  22462=>"111101111",
  22463=>"001110110",
  22464=>"100001110",
  22465=>"000110011",
  22466=>"110110010",
  22467=>"110010111",
  22468=>"000111010",
  22469=>"010111001",
  22470=>"111001110",
  22471=>"000111001",
  22472=>"000000101",
  22473=>"010000011",
  22474=>"100001100",
  22475=>"000111000",
  22476=>"000001010",
  22477=>"110011101",
  22478=>"000100001",
  22479=>"010110111",
  22480=>"110100110",
  22481=>"010001010",
  22482=>"000001011",
  22483=>"010001000",
  22484=>"100111111",
  22485=>"111001111",
  22486=>"011101111",
  22487=>"010111101",
  22488=>"000000110",
  22489=>"011001000",
  22490=>"010101010",
  22491=>"100001010",
  22492=>"111001110",
  22493=>"101010110",
  22494=>"110100110",
  22495=>"001111010",
  22496=>"000000100",
  22497=>"011000101",
  22498=>"100111110",
  22499=>"010101101",
  22500=>"001000010",
  22501=>"100001110",
  22502=>"010110100",
  22503=>"100111001",
  22504=>"000001111",
  22505=>"001011000",
  22506=>"111000011",
  22507=>"100100001",
  22508=>"000100110",
  22509=>"000111000",
  22510=>"110111110",
  22511=>"111001100",
  22512=>"111001001",
  22513=>"010110001",
  22514=>"100100000",
  22515=>"010010010",
  22516=>"001001010",
  22517=>"001010010",
  22518=>"100011000",
  22519=>"111011101",
  22520=>"001101111",
  22521=>"001100101",
  22522=>"110101011",
  22523=>"111010011",
  22524=>"111110010",
  22525=>"001100010",
  22526=>"111100011",
  22527=>"111110001",
  22528=>"000011010",
  22529=>"110111100",
  22530=>"110110001",
  22531=>"001010000",
  22532=>"011111110",
  22533=>"101001110",
  22534=>"000011010",
  22535=>"001100100",
  22536=>"000110001",
  22537=>"000011000",
  22538=>"101000101",
  22539=>"111101111",
  22540=>"101100010",
  22541=>"000001000",
  22542=>"001111111",
  22543=>"000011010",
  22544=>"001101010",
  22545=>"110001111",
  22546=>"110011100",
  22547=>"101111100",
  22548=>"111101001",
  22549=>"111010001",
  22550=>"100011110",
  22551=>"000100110",
  22552=>"111111101",
  22553=>"000000111",
  22554=>"000001111",
  22555=>"111010011",
  22556=>"100111000",
  22557=>"111001101",
  22558=>"011000110",
  22559=>"111110101",
  22560=>"000000000",
  22561=>"010100101",
  22562=>"010001000",
  22563=>"011000010",
  22564=>"111011111",
  22565=>"101011010",
  22566=>"000100011",
  22567=>"000101001",
  22568=>"111001000",
  22569=>"110110111",
  22570=>"000111101",
  22571=>"101010101",
  22572=>"101001100",
  22573=>"001010100",
  22574=>"010101111",
  22575=>"011100111",
  22576=>"011110111",
  22577=>"101101000",
  22578=>"101101101",
  22579=>"011101011",
  22580=>"100010011",
  22581=>"100000011",
  22582=>"101101001",
  22583=>"010111101",
  22584=>"001011011",
  22585=>"010001000",
  22586=>"100000000",
  22587=>"100111011",
  22588=>"111101100",
  22589=>"101000100",
  22590=>"110111100",
  22591=>"110101010",
  22592=>"110001101",
  22593=>"110000000",
  22594=>"001101011",
  22595=>"000000111",
  22596=>"101001101",
  22597=>"011000000",
  22598=>"101111000",
  22599=>"111010000",
  22600=>"101001011",
  22601=>"110010101",
  22602=>"110101101",
  22603=>"101001011",
  22604=>"000000101",
  22605=>"100111110",
  22606=>"100011001",
  22607=>"000111100",
  22608=>"011101001",
  22609=>"001011100",
  22610=>"111011011",
  22611=>"001100001",
  22612=>"001110010",
  22613=>"111000101",
  22614=>"110010010",
  22615=>"011110100",
  22616=>"111100010",
  22617=>"111100011",
  22618=>"000110010",
  22619=>"001000101",
  22620=>"000110011",
  22621=>"110011111",
  22622=>"000011100",
  22623=>"000011110",
  22624=>"001000010",
  22625=>"010000101",
  22626=>"101101101",
  22627=>"011001000",
  22628=>"111011001",
  22629=>"010000011",
  22630=>"011111111",
  22631=>"011100101",
  22632=>"010011010",
  22633=>"111110011",
  22634=>"110001110",
  22635=>"101110111",
  22636=>"101000111",
  22637=>"101111011",
  22638=>"111000100",
  22639=>"111001000",
  22640=>"111000000",
  22641=>"000001111",
  22642=>"111100011",
  22643=>"011101000",
  22644=>"110010111",
  22645=>"110101111",
  22646=>"100101100",
  22647=>"111000010",
  22648=>"001011011",
  22649=>"101001111",
  22650=>"110011110",
  22651=>"110110110",
  22652=>"000011000",
  22653=>"100110101",
  22654=>"101100000",
  22655=>"001011000",
  22656=>"101001010",
  22657=>"110111011",
  22658=>"110110001",
  22659=>"001100100",
  22660=>"100110101",
  22661=>"000001001",
  22662=>"111110010",
  22663=>"010100011",
  22664=>"010101111",
  22665=>"000011000",
  22666=>"110001001",
  22667=>"101100101",
  22668=>"010000000",
  22669=>"110000100",
  22670=>"111001110",
  22671=>"100010101",
  22672=>"111001111",
  22673=>"001110001",
  22674=>"010011101",
  22675=>"111011111",
  22676=>"111011011",
  22677=>"101001000",
  22678=>"001011000",
  22679=>"110111011",
  22680=>"100110111",
  22681=>"101100000",
  22682=>"010111100",
  22683=>"100001100",
  22684=>"111001000",
  22685=>"001010000",
  22686=>"100011000",
  22687=>"110010000",
  22688=>"101000111",
  22689=>"000011111",
  22690=>"001001011",
  22691=>"111101010",
  22692=>"011010110",
  22693=>"010111101",
  22694=>"000100010",
  22695=>"000011011",
  22696=>"111111111",
  22697=>"011000000",
  22698=>"110111011",
  22699=>"011101010",
  22700=>"001101101",
  22701=>"011000000",
  22702=>"110111111",
  22703=>"011101000",
  22704=>"011010001",
  22705=>"010111110",
  22706=>"101111001",
  22707=>"001111001",
  22708=>"111101100",
  22709=>"001010111",
  22710=>"101100111",
  22711=>"100010010",
  22712=>"100000100",
  22713=>"111101101",
  22714=>"110000110",
  22715=>"111000110",
  22716=>"001000000",
  22717=>"010100111",
  22718=>"000101110",
  22719=>"101100111",
  22720=>"011011001",
  22721=>"101001000",
  22722=>"111001100",
  22723=>"100000100",
  22724=>"110100001",
  22725=>"100101111",
  22726=>"101000110",
  22727=>"001101101",
  22728=>"000001001",
  22729=>"010101111",
  22730=>"110011100",
  22731=>"000001011",
  22732=>"110100110",
  22733=>"001001101",
  22734=>"011001100",
  22735=>"011001001",
  22736=>"011100100",
  22737=>"000110100",
  22738=>"001100111",
  22739=>"011101111",
  22740=>"100111011",
  22741=>"101111100",
  22742=>"011010111",
  22743=>"101100101",
  22744=>"000111100",
  22745=>"001001000",
  22746=>"101000011",
  22747=>"101010111",
  22748=>"100011001",
  22749=>"000110100",
  22750=>"010110000",
  22751=>"110000000",
  22752=>"010100000",
  22753=>"001110000",
  22754=>"111011110",
  22755=>"011010100",
  22756=>"011101000",
  22757=>"101110111",
  22758=>"011000000",
  22759=>"110011100",
  22760=>"110000100",
  22761=>"011101111",
  22762=>"001110111",
  22763=>"011011111",
  22764=>"100000000",
  22765=>"000100101",
  22766=>"111001110",
  22767=>"000001001",
  22768=>"000100101",
  22769=>"010001101",
  22770=>"010101101",
  22771=>"111011010",
  22772=>"110110111",
  22773=>"110111000",
  22774=>"100101001",
  22775=>"010100001",
  22776=>"001111100",
  22777=>"100101010",
  22778=>"000000101",
  22779=>"100100001",
  22780=>"000001111",
  22781=>"000111010",
  22782=>"000010001",
  22783=>"100110100",
  22784=>"000010000",
  22785=>"001011000",
  22786=>"011101110",
  22787=>"000011101",
  22788=>"111011101",
  22789=>"111110010",
  22790=>"011111001",
  22791=>"101011111",
  22792=>"111000111",
  22793=>"001000001",
  22794=>"100001010",
  22795=>"101000100",
  22796=>"100110111",
  22797=>"101110101",
  22798=>"001110111",
  22799=>"100101100",
  22800=>"010010000",
  22801=>"000110100",
  22802=>"111010101",
  22803=>"010000001",
  22804=>"100110100",
  22805=>"010111010",
  22806=>"111110101",
  22807=>"111100100",
  22808=>"000011101",
  22809=>"000101011",
  22810=>"001101110",
  22811=>"011001110",
  22812=>"000111000",
  22813=>"001100101",
  22814=>"101100101",
  22815=>"011101010",
  22816=>"111010111",
  22817=>"010100010",
  22818=>"101011101",
  22819=>"001101101",
  22820=>"000001001",
  22821=>"001100111",
  22822=>"001010110",
  22823=>"001111110",
  22824=>"100101101",
  22825=>"101000010",
  22826=>"001110001",
  22827=>"011001110",
  22828=>"001000110",
  22829=>"100101000",
  22830=>"100000010",
  22831=>"000111101",
  22832=>"010011010",
  22833=>"111100011",
  22834=>"001000010",
  22835=>"000010010",
  22836=>"001011100",
  22837=>"110110011",
  22838=>"110111101",
  22839=>"001001000",
  22840=>"001001100",
  22841=>"101001110",
  22842=>"110010011",
  22843=>"010101100",
  22844=>"010111101",
  22845=>"111011100",
  22846=>"110100101",
  22847=>"110101010",
  22848=>"110100101",
  22849=>"010100000",
  22850=>"101110111",
  22851=>"011110010",
  22852=>"110110111",
  22853=>"100000110",
  22854=>"101011110",
  22855=>"110001001",
  22856=>"111111111",
  22857=>"000011001",
  22858=>"100010101",
  22859=>"011001111",
  22860=>"110001110",
  22861=>"111011101",
  22862=>"111100000",
  22863=>"010100100",
  22864=>"001100000",
  22865=>"100111011",
  22866=>"110100010",
  22867=>"001001100",
  22868=>"001000000",
  22869=>"000011111",
  22870=>"110110101",
  22871=>"100101110",
  22872=>"000111000",
  22873=>"011001001",
  22874=>"111001010",
  22875=>"000001001",
  22876=>"111001000",
  22877=>"110000011",
  22878=>"011110000",
  22879=>"111100111",
  22880=>"110101010",
  22881=>"010001011",
  22882=>"011111000",
  22883=>"001011100",
  22884=>"001111001",
  22885=>"101100110",
  22886=>"011101010",
  22887=>"001001000",
  22888=>"101101111",
  22889=>"000001011",
  22890=>"101000100",
  22891=>"100000100",
  22892=>"011000000",
  22893=>"110111001",
  22894=>"100111110",
  22895=>"110010000",
  22896=>"001010111",
  22897=>"110000000",
  22898=>"000001101",
  22899=>"000110010",
  22900=>"001110101",
  22901=>"011111100",
  22902=>"100000011",
  22903=>"011101001",
  22904=>"101001011",
  22905=>"011001100",
  22906=>"101110111",
  22907=>"011011000",
  22908=>"110001111",
  22909=>"101100111",
  22910=>"100011001",
  22911=>"001010010",
  22912=>"010111111",
  22913=>"111111001",
  22914=>"111011111",
  22915=>"000100100",
  22916=>"011111100",
  22917=>"011000101",
  22918=>"111111101",
  22919=>"011000100",
  22920=>"000110111",
  22921=>"110000111",
  22922=>"011011101",
  22923=>"001100000",
  22924=>"000011000",
  22925=>"101110111",
  22926=>"000100111",
  22927=>"010100110",
  22928=>"101111000",
  22929=>"000000001",
  22930=>"101100001",
  22931=>"010100010",
  22932=>"011001100",
  22933=>"010010101",
  22934=>"101110011",
  22935=>"010111101",
  22936=>"010000101",
  22937=>"010010010",
  22938=>"111101111",
  22939=>"111011101",
  22940=>"111111001",
  22941=>"101000010",
  22942=>"101010001",
  22943=>"110001001",
  22944=>"111110000",
  22945=>"000000010",
  22946=>"110001000",
  22947=>"000100101",
  22948=>"100010000",
  22949=>"110101001",
  22950=>"001110100",
  22951=>"011011011",
  22952=>"000101011",
  22953=>"100101111",
  22954=>"111011111",
  22955=>"100111111",
  22956=>"111001101",
  22957=>"011101111",
  22958=>"100001110",
  22959=>"111100111",
  22960=>"111000001",
  22961=>"110000111",
  22962=>"100101010",
  22963=>"001000110",
  22964=>"111111110",
  22965=>"001101011",
  22966=>"001000010",
  22967=>"001101111",
  22968=>"001011101",
  22969=>"000101010",
  22970=>"001100000",
  22971=>"011010111",
  22972=>"011000101",
  22973=>"010110110",
  22974=>"101101001",
  22975=>"001110111",
  22976=>"001100000",
  22977=>"011000100",
  22978=>"101010111",
  22979=>"000110101",
  22980=>"000101111",
  22981=>"111000011",
  22982=>"011111110",
  22983=>"011011000",
  22984=>"000111000",
  22985=>"101101010",
  22986=>"010100000",
  22987=>"001110000",
  22988=>"110011011",
  22989=>"111111011",
  22990=>"001010110",
  22991=>"011010011",
  22992=>"010001101",
  22993=>"000000001",
  22994=>"001100101",
  22995=>"001100001",
  22996=>"001110001",
  22997=>"001111000",
  22998=>"111001101",
  22999=>"000000010",
  23000=>"110100001",
  23001=>"001101001",
  23002=>"101100010",
  23003=>"110000010",
  23004=>"100001101",
  23005=>"000001001",
  23006=>"000010001",
  23007=>"110111000",
  23008=>"111111010",
  23009=>"111111000",
  23010=>"011000101",
  23011=>"110110000",
  23012=>"010010100",
  23013=>"000010101",
  23014=>"010000001",
  23015=>"111010000",
  23016=>"010010111",
  23017=>"010110001",
  23018=>"001000100",
  23019=>"010000111",
  23020=>"011110010",
  23021=>"000111001",
  23022=>"100000010",
  23023=>"000001011",
  23024=>"011111000",
  23025=>"110110011",
  23026=>"100111000",
  23027=>"000101011",
  23028=>"110110010",
  23029=>"001101001",
  23030=>"000101001",
  23031=>"001101010",
  23032=>"001000001",
  23033=>"011111010",
  23034=>"110111011",
  23035=>"111001111",
  23036=>"011001101",
  23037=>"100100010",
  23038=>"011111111",
  23039=>"111000000",
  23040=>"101110110",
  23041=>"001001001",
  23042=>"011010001",
  23043=>"000000010",
  23044=>"010110010",
  23045=>"000000100",
  23046=>"101011111",
  23047=>"001000011",
  23048=>"101011110",
  23049=>"111001110",
  23050=>"010011101",
  23051=>"011100100",
  23052=>"110011000",
  23053=>"111010101",
  23054=>"000001000",
  23055=>"011111100",
  23056=>"111100110",
  23057=>"100110000",
  23058=>"100010110",
  23059=>"011100011",
  23060=>"000101000",
  23061=>"101101101",
  23062=>"110001111",
  23063=>"000100001",
  23064=>"100011111",
  23065=>"100100011",
  23066=>"100010101",
  23067=>"000100100",
  23068=>"001001000",
  23069=>"000111000",
  23070=>"001000000",
  23071=>"111100101",
  23072=>"101101011",
  23073=>"110000111",
  23074=>"101010111",
  23075=>"101010000",
  23076=>"010110110",
  23077=>"010100111",
  23078=>"001101011",
  23079=>"101101111",
  23080=>"011010011",
  23081=>"000000111",
  23082=>"000011011",
  23083=>"001010110",
  23084=>"100010001",
  23085=>"100111000",
  23086=>"100101110",
  23087=>"100000010",
  23088=>"101100011",
  23089=>"101101110",
  23090=>"010001001",
  23091=>"110001111",
  23092=>"011011001",
  23093=>"011110111",
  23094=>"011011011",
  23095=>"001111010",
  23096=>"110111100",
  23097=>"101001010",
  23098=>"100100010",
  23099=>"101000110",
  23100=>"010100011",
  23101=>"011001101",
  23102=>"011011010",
  23103=>"000011100",
  23104=>"011011100",
  23105=>"110101000",
  23106=>"000011000",
  23107=>"010001101",
  23108=>"011010111",
  23109=>"011100111",
  23110=>"000000100",
  23111=>"001100110",
  23112=>"001111101",
  23113=>"101101100",
  23114=>"000010111",
  23115=>"001001011",
  23116=>"000000011",
  23117=>"011011101",
  23118=>"100100011",
  23119=>"111110110",
  23120=>"100100101",
  23121=>"010010001",
  23122=>"100000001",
  23123=>"001001111",
  23124=>"101111010",
  23125=>"001010101",
  23126=>"100100010",
  23127=>"010110110",
  23128=>"001111011",
  23129=>"011101100",
  23130=>"010011011",
  23131=>"111100100",
  23132=>"110111011",
  23133=>"011110100",
  23134=>"110000000",
  23135=>"111011101",
  23136=>"101111100",
  23137=>"001110100",
  23138=>"101001000",
  23139=>"000011110",
  23140=>"001101010",
  23141=>"101101100",
  23142=>"011011110",
  23143=>"111011110",
  23144=>"110010111",
  23145=>"100100011",
  23146=>"111111111",
  23147=>"110111011",
  23148=>"010001100",
  23149=>"110111111",
  23150=>"001101100",
  23151=>"100011000",
  23152=>"110000001",
  23153=>"011110010",
  23154=>"010000010",
  23155=>"110111010",
  23156=>"000000100",
  23157=>"101010111",
  23158=>"101110010",
  23159=>"111011110",
  23160=>"110101110",
  23161=>"000001100",
  23162=>"000001000",
  23163=>"000000100",
  23164=>"110000101",
  23165=>"000110100",
  23166=>"101000110",
  23167=>"111100101",
  23168=>"110001010",
  23169=>"110011101",
  23170=>"101000111",
  23171=>"111110110",
  23172=>"001011110",
  23173=>"110100001",
  23174=>"001111011",
  23175=>"101101010",
  23176=>"100001100",
  23177=>"011001111",
  23178=>"100101111",
  23179=>"111010000",
  23180=>"010000000",
  23181=>"000000010",
  23182=>"111101101",
  23183=>"101111111",
  23184=>"010101100",
  23185=>"001000101",
  23186=>"001011111",
  23187=>"100011110",
  23188=>"110111100",
  23189=>"111001001",
  23190=>"000111100",
  23191=>"111001000",
  23192=>"001110010",
  23193=>"001111000",
  23194=>"001100101",
  23195=>"001110100",
  23196=>"010100011",
  23197=>"111000100",
  23198=>"010001000",
  23199=>"001001111",
  23200=>"101001011",
  23201=>"001011111",
  23202=>"000110011",
  23203=>"000111010",
  23204=>"101000001",
  23205=>"100101110",
  23206=>"100000100",
  23207=>"000110000",
  23208=>"100010100",
  23209=>"110010111",
  23210=>"010010001",
  23211=>"011000011",
  23212=>"001001010",
  23213=>"110111000",
  23214=>"011000000",
  23215=>"000101110",
  23216=>"000101101",
  23217=>"001100010",
  23218=>"110000001",
  23219=>"111101011",
  23220=>"110000001",
  23221=>"101101101",
  23222=>"001111011",
  23223=>"110110100",
  23224=>"010111111",
  23225=>"011010110",
  23226=>"101011110",
  23227=>"001110010",
  23228=>"001100111",
  23229=>"000010000",
  23230=>"111000111",
  23231=>"100101001",
  23232=>"000000100",
  23233=>"101100101",
  23234=>"101011011",
  23235=>"110110110",
  23236=>"001101010",
  23237=>"100010111",
  23238=>"010001010",
  23239=>"110010111",
  23240=>"100101011",
  23241=>"011101001",
  23242=>"100010100",
  23243=>"011110000",
  23244=>"000111111",
  23245=>"001001100",
  23246=>"111110111",
  23247=>"110001101",
  23248=>"100110011",
  23249=>"111001100",
  23250=>"100101110",
  23251=>"000000110",
  23252=>"110001000",
  23253=>"101001111",
  23254=>"111100100",
  23255=>"111110111",
  23256=>"000000010",
  23257=>"000010101",
  23258=>"100110101",
  23259=>"110101111",
  23260=>"110001000",
  23261=>"011000000",
  23262=>"010010001",
  23263=>"110010110",
  23264=>"010001000",
  23265=>"111110010",
  23266=>"111000010",
  23267=>"001101110",
  23268=>"100010001",
  23269=>"011000001",
  23270=>"001110111",
  23271=>"001001101",
  23272=>"111101011",
  23273=>"111100010",
  23274=>"000001110",
  23275=>"110010100",
  23276=>"001000000",
  23277=>"010100101",
  23278=>"111100000",
  23279=>"001110000",
  23280=>"101000110",
  23281=>"110000000",
  23282=>"001010101",
  23283=>"101000101",
  23284=>"000001010",
  23285=>"111000001",
  23286=>"001000000",
  23287=>"001100000",
  23288=>"010101011",
  23289=>"001001000",
  23290=>"011111001",
  23291=>"110101100",
  23292=>"101111010",
  23293=>"111100011",
  23294=>"001111011",
  23295=>"010001000",
  23296=>"100000100",
  23297=>"100110010",
  23298=>"001100010",
  23299=>"010011000",
  23300=>"110011011",
  23301=>"100001000",
  23302=>"111111000",
  23303=>"111110010",
  23304=>"011110001",
  23305=>"101100100",
  23306=>"100001101",
  23307=>"001001011",
  23308=>"001000100",
  23309=>"010011011",
  23310=>"011011001",
  23311=>"011100110",
  23312=>"000100111",
  23313=>"000101011",
  23314=>"110101110",
  23315=>"101110001",
  23316=>"000100000",
  23317=>"000100100",
  23318=>"111010000",
  23319=>"011111010",
  23320=>"111110110",
  23321=>"001001010",
  23322=>"010100011",
  23323=>"000111001",
  23324=>"011110111",
  23325=>"110100010",
  23326=>"100000111",
  23327=>"100001000",
  23328=>"111011111",
  23329=>"101111100",
  23330=>"011110111",
  23331=>"101011000",
  23332=>"101101000",
  23333=>"000000010",
  23334=>"011100111",
  23335=>"101101110",
  23336=>"000101001",
  23337=>"101100100",
  23338=>"110100010",
  23339=>"111010110",
  23340=>"001110010",
  23341=>"111010010",
  23342=>"000111011",
  23343=>"101111111",
  23344=>"100110110",
  23345=>"101000101",
  23346=>"001000011",
  23347=>"000100100",
  23348=>"110100011",
  23349=>"111011101",
  23350=>"100110100",
  23351=>"000001000",
  23352=>"110101000",
  23353=>"111010101",
  23354=>"010010101",
  23355=>"110011000",
  23356=>"110010000",
  23357=>"010101001",
  23358=>"001011010",
  23359=>"001111010",
  23360=>"010010110",
  23361=>"111001000",
  23362=>"010100100",
  23363=>"001001011",
  23364=>"011000110",
  23365=>"001111001",
  23366=>"111111110",
  23367=>"110101101",
  23368=>"001001000",
  23369=>"010000001",
  23370=>"010000010",
  23371=>"011001100",
  23372=>"101110001",
  23373=>"001011110",
  23374=>"000110100",
  23375=>"111010110",
  23376=>"100111110",
  23377=>"100101100",
  23378=>"010000100",
  23379=>"101101010",
  23380=>"101111100",
  23381=>"100101000",
  23382=>"100100101",
  23383=>"000100111",
  23384=>"110101001",
  23385=>"010001111",
  23386=>"000111011",
  23387=>"001010011",
  23388=>"111110010",
  23389=>"100101111",
  23390=>"111000111",
  23391=>"010110110",
  23392=>"010111010",
  23393=>"101010001",
  23394=>"010010110",
  23395=>"010101101",
  23396=>"000101101",
  23397=>"101010101",
  23398=>"001000010",
  23399=>"010001000",
  23400=>"000001000",
  23401=>"101001110",
  23402=>"100011000",
  23403=>"010001100",
  23404=>"001111111",
  23405=>"000101110",
  23406=>"101001001",
  23407=>"110100010",
  23408=>"101010101",
  23409=>"101011011",
  23410=>"100101101",
  23411=>"001000011",
  23412=>"101000011",
  23413=>"011011000",
  23414=>"000011001",
  23415=>"001000010",
  23416=>"011100010",
  23417=>"100111101",
  23418=>"101110011",
  23419=>"011110011",
  23420=>"000110011",
  23421=>"001100001",
  23422=>"111110110",
  23423=>"011100100",
  23424=>"111010011",
  23425=>"000011001",
  23426=>"000101000",
  23427=>"110001011",
  23428=>"101011101",
  23429=>"101011001",
  23430=>"010011111",
  23431=>"001001110",
  23432=>"000011100",
  23433=>"100111111",
  23434=>"000010010",
  23435=>"110011111",
  23436=>"111100001",
  23437=>"110100111",
  23438=>"011010000",
  23439=>"100111010",
  23440=>"011101011",
  23441=>"111100010",
  23442=>"000010110",
  23443=>"111010101",
  23444=>"010000110",
  23445=>"001011101",
  23446=>"011010111",
  23447=>"111010101",
  23448=>"111011100",
  23449=>"011101100",
  23450=>"000001111",
  23451=>"101001101",
  23452=>"000110000",
  23453=>"000000100",
  23454=>"010000011",
  23455=>"101111111",
  23456=>"101100000",
  23457=>"001000001",
  23458=>"111011101",
  23459=>"111001000",
  23460=>"000100001",
  23461=>"110100101",
  23462=>"001011100",
  23463=>"111010010",
  23464=>"001000110",
  23465=>"101011001",
  23466=>"001100000",
  23467=>"001011000",
  23468=>"011010000",
  23469=>"110010100",
  23470=>"111111001",
  23471=>"000000011",
  23472=>"100110001",
  23473=>"110101010",
  23474=>"000000011",
  23475=>"001011011",
  23476=>"011001001",
  23477=>"011111100",
  23478=>"101011011",
  23479=>"000110100",
  23480=>"011001111",
  23481=>"111101110",
  23482=>"010010111",
  23483=>"100001111",
  23484=>"001001111",
  23485=>"100101101",
  23486=>"000100101",
  23487=>"100111010",
  23488=>"111010111",
  23489=>"110010110",
  23490=>"000101000",
  23491=>"101000110",
  23492=>"111000010",
  23493=>"001001001",
  23494=>"100100001",
  23495=>"001010011",
  23496=>"111000010",
  23497=>"110101111",
  23498=>"011000111",
  23499=>"110000010",
  23500=>"010111000",
  23501=>"110010011",
  23502=>"000001110",
  23503=>"101000001",
  23504=>"010011101",
  23505=>"011100101",
  23506=>"010100001",
  23507=>"010011000",
  23508=>"110100000",
  23509=>"110010101",
  23510=>"110100100",
  23511=>"110100010",
  23512=>"000010111",
  23513=>"110110101",
  23514=>"011000000",
  23515=>"000110010",
  23516=>"111101101",
  23517=>"001101001",
  23518=>"010100001",
  23519=>"001000010",
  23520=>"010100010",
  23521=>"001011010",
  23522=>"010001110",
  23523=>"000000110",
  23524=>"100000101",
  23525=>"101110111",
  23526=>"110001011",
  23527=>"101111101",
  23528=>"000000101",
  23529=>"100000101",
  23530=>"111111011",
  23531=>"001011111",
  23532=>"100101011",
  23533=>"101100111",
  23534=>"110001010",
  23535=>"100001110",
  23536=>"111000001",
  23537=>"000011000",
  23538=>"000011101",
  23539=>"110000000",
  23540=>"011001101",
  23541=>"101011000",
  23542=>"001110111",
  23543=>"111001011",
  23544=>"100101000",
  23545=>"111011100",
  23546=>"000001000",
  23547=>"011101000",
  23548=>"100001111",
  23549=>"011110100",
  23550=>"111110011",
  23551=>"011010111",
  23552=>"110110111",
  23553=>"101100110",
  23554=>"101110110",
  23555=>"101111011",
  23556=>"100101101",
  23557=>"010001000",
  23558=>"111111100",
  23559=>"110010001",
  23560=>"111011100",
  23561=>"000001011",
  23562=>"111000001",
  23563=>"110101010",
  23564=>"100000010",
  23565=>"111011011",
  23566=>"010001000",
  23567=>"100111010",
  23568=>"101001111",
  23569=>"010000001",
  23570=>"111010011",
  23571=>"111101101",
  23572=>"101011011",
  23573=>"110011110",
  23574=>"001100101",
  23575=>"011100101",
  23576=>"110000111",
  23577=>"011110000",
  23578=>"110010011",
  23579=>"010100011",
  23580=>"000111101",
  23581=>"101100000",
  23582=>"000011111",
  23583=>"110100101",
  23584=>"110011011",
  23585=>"110101101",
  23586=>"010110000",
  23587=>"001000000",
  23588=>"000000110",
  23589=>"001011111",
  23590=>"000011011",
  23591=>"101000010",
  23592=>"100111110",
  23593=>"110110101",
  23594=>"001011100",
  23595=>"101101001",
  23596=>"101000011",
  23597=>"101110011",
  23598=>"010100001",
  23599=>"000111011",
  23600=>"001001011",
  23601=>"000001010",
  23602=>"100101001",
  23603=>"000111000",
  23604=>"110010000",
  23605=>"010100001",
  23606=>"101000110",
  23607=>"110001001",
  23608=>"011111011",
  23609=>"100011001",
  23610=>"100110101",
  23611=>"101001000",
  23612=>"100100111",
  23613=>"010000010",
  23614=>"111111111",
  23615=>"010011000",
  23616=>"010000001",
  23617=>"101011100",
  23618=>"110111001",
  23619=>"001011101",
  23620=>"111010011",
  23621=>"001001001",
  23622=>"001010110",
  23623=>"000000000",
  23624=>"010111101",
  23625=>"010100000",
  23626=>"010001101",
  23627=>"011010100",
  23628=>"010010000",
  23629=>"110111100",
  23630=>"101101010",
  23631=>"001100010",
  23632=>"011010010",
  23633=>"001101100",
  23634=>"000000010",
  23635=>"101001011",
  23636=>"100011100",
  23637=>"110000010",
  23638=>"110100101",
  23639=>"100000000",
  23640=>"000110000",
  23641=>"001000001",
  23642=>"101010010",
  23643=>"111111001",
  23644=>"011010100",
  23645=>"010000010",
  23646=>"100010110",
  23647=>"101001000",
  23648=>"001001110",
  23649=>"001001001",
  23650=>"000000111",
  23651=>"011110101",
  23652=>"101101100",
  23653=>"100001110",
  23654=>"001011011",
  23655=>"000101010",
  23656=>"011011110",
  23657=>"111111100",
  23658=>"101001100",
  23659=>"111111001",
  23660=>"000011111",
  23661=>"101100001",
  23662=>"111100110",
  23663=>"100000011",
  23664=>"100011001",
  23665=>"010100100",
  23666=>"110010111",
  23667=>"000110000",
  23668=>"101010000",
  23669=>"101111100",
  23670=>"000010011",
  23671=>"110001111",
  23672=>"000100110",
  23673=>"010101001",
  23674=>"110110111",
  23675=>"100101010",
  23676=>"001101110",
  23677=>"101111111",
  23678=>"100011111",
  23679=>"011100111",
  23680=>"110110011",
  23681=>"110111101",
  23682=>"101110001",
  23683=>"111001011",
  23684=>"011111000",
  23685=>"001111001",
  23686=>"010000100",
  23687=>"010000001",
  23688=>"011110111",
  23689=>"000000000",
  23690=>"100111000",
  23691=>"010001011",
  23692=>"000010111",
  23693=>"001010010",
  23694=>"010011110",
  23695=>"000100011",
  23696=>"000111011",
  23697=>"110100001",
  23698=>"010101100",
  23699=>"001000100",
  23700=>"001001011",
  23701=>"100010101",
  23702=>"000111010",
  23703=>"100111000",
  23704=>"000000110",
  23705=>"011100111",
  23706=>"000011101",
  23707=>"101011000",
  23708=>"000101100",
  23709=>"011011101",
  23710=>"000010001",
  23711=>"000000010",
  23712=>"010010100",
  23713=>"101111101",
  23714=>"011111110",
  23715=>"001001000",
  23716=>"100000010",
  23717=>"111110011",
  23718=>"011010010",
  23719=>"101110100",
  23720=>"000001000",
  23721=>"010011010",
  23722=>"110101101",
  23723=>"011110000",
  23724=>"111010100",
  23725=>"011101010",
  23726=>"101010111",
  23727=>"010001111",
  23728=>"001011011",
  23729=>"000001011",
  23730=>"000001010",
  23731=>"000111110",
  23732=>"000001001",
  23733=>"011011110",
  23734=>"101000011",
  23735=>"011100100",
  23736=>"001000100",
  23737=>"101100101",
  23738=>"010011010",
  23739=>"000011101",
  23740=>"111100100",
  23741=>"101000001",
  23742=>"001001000",
  23743=>"000100101",
  23744=>"100100000",
  23745=>"111001010",
  23746=>"100001000",
  23747=>"111111111",
  23748=>"111101011",
  23749=>"011101010",
  23750=>"101000111",
  23751=>"000111110",
  23752=>"000011111",
  23753=>"100010010",
  23754=>"100000010",
  23755=>"110111100",
  23756=>"101001000",
  23757=>"111000010",
  23758=>"000100110",
  23759=>"011000000",
  23760=>"100100101",
  23761=>"101110000",
  23762=>"111011101",
  23763=>"110001000",
  23764=>"000011110",
  23765=>"110101111",
  23766=>"001000000",
  23767=>"011001000",
  23768=>"000010111",
  23769=>"100110011",
  23770=>"100001100",
  23771=>"011001010",
  23772=>"000100010",
  23773=>"000011001",
  23774=>"010101000",
  23775=>"111000000",
  23776=>"100001111",
  23777=>"000100111",
  23778=>"100101000",
  23779=>"000100011",
  23780=>"101001000",
  23781=>"100010010",
  23782=>"001011110",
  23783=>"011110001",
  23784=>"001011101",
  23785=>"100011101",
  23786=>"100001001",
  23787=>"001000111",
  23788=>"111000100",
  23789=>"101011001",
  23790=>"001110110",
  23791=>"100000011",
  23792=>"110101100",
  23793=>"010001000",
  23794=>"110111001",
  23795=>"010101101",
  23796=>"010011011",
  23797=>"101001000",
  23798=>"110110100",
  23799=>"100000001",
  23800=>"001111101",
  23801=>"000100001",
  23802=>"001111010",
  23803=>"001001001",
  23804=>"110101010",
  23805=>"100011100",
  23806=>"101010011",
  23807=>"010101011",
  23808=>"111101001",
  23809=>"101100100",
  23810=>"111010111",
  23811=>"001101001",
  23812=>"111100000",
  23813=>"111010000",
  23814=>"111100111",
  23815=>"001110110",
  23816=>"101010110",
  23817=>"010010000",
  23818=>"111010110",
  23819=>"110011001",
  23820=>"001110111",
  23821=>"110101111",
  23822=>"111100000",
  23823=>"101010101",
  23824=>"001010011",
  23825=>"110111000",
  23826=>"001111111",
  23827=>"111110010",
  23828=>"111110011",
  23829=>"000000100",
  23830=>"101000010",
  23831=>"000010010",
  23832=>"111101110",
  23833=>"111101000",
  23834=>"110010001",
  23835=>"101101001",
  23836=>"001110000",
  23837=>"011001010",
  23838=>"100111011",
  23839=>"101111000",
  23840=>"011110001",
  23841=>"100100010",
  23842=>"000001010",
  23843=>"011000011",
  23844=>"001110011",
  23845=>"010111111",
  23846=>"000110000",
  23847=>"000000000",
  23848=>"001110000",
  23849=>"100111101",
  23850=>"110010001",
  23851=>"101011110",
  23852=>"110111111",
  23853=>"101100100",
  23854=>"110010011",
  23855=>"111101010",
  23856=>"111000010",
  23857=>"100010001",
  23858=>"111100010",
  23859=>"110000010",
  23860=>"000010110",
  23861=>"000001111",
  23862=>"000010100",
  23863=>"100101111",
  23864=>"010000111",
  23865=>"110110100",
  23866=>"111001101",
  23867=>"000000111",
  23868=>"001110001",
  23869=>"111110011",
  23870=>"001111000",
  23871=>"011111001",
  23872=>"000000110",
  23873=>"000111101",
  23874=>"101110100",
  23875=>"101110010",
  23876=>"000001101",
  23877=>"010100001",
  23878=>"001000110",
  23879=>"000001110",
  23880=>"011010000",
  23881=>"100010100",
  23882=>"000101010",
  23883=>"101110011",
  23884=>"110001111",
  23885=>"101001100",
  23886=>"001010110",
  23887=>"000100000",
  23888=>"100100001",
  23889=>"010010010",
  23890=>"010110111",
  23891=>"011110100",
  23892=>"011000000",
  23893=>"010110110",
  23894=>"001111100",
  23895=>"101001101",
  23896=>"000000110",
  23897=>"100100100",
  23898=>"011111111",
  23899=>"100110010",
  23900=>"011000101",
  23901=>"001010100",
  23902=>"111000111",
  23903=>"000000000",
  23904=>"000110110",
  23905=>"011001011",
  23906=>"010010001",
  23907=>"101010111",
  23908=>"101011101",
  23909=>"001011010",
  23910=>"101000010",
  23911=>"000101000",
  23912=>"101111010",
  23913=>"000101110",
  23914=>"011001000",
  23915=>"111001100",
  23916=>"000100001",
  23917=>"110011101",
  23918=>"111100000",
  23919=>"001010111",
  23920=>"111111110",
  23921=>"010101000",
  23922=>"011010101",
  23923=>"110001111",
  23924=>"000001111",
  23925=>"001011000",
  23926=>"010100011",
  23927=>"000110000",
  23928=>"010101010",
  23929=>"111110011",
  23930=>"010011101",
  23931=>"011111101",
  23932=>"111000110",
  23933=>"100110000",
  23934=>"011100111",
  23935=>"110001001",
  23936=>"010011101",
  23937=>"001001100",
  23938=>"101110001",
  23939=>"001011111",
  23940=>"111100101",
  23941=>"000000001",
  23942=>"101010001",
  23943=>"101001011",
  23944=>"001011000",
  23945=>"010100100",
  23946=>"100101011",
  23947=>"101011101",
  23948=>"100101000",
  23949=>"011010100",
  23950=>"001100101",
  23951=>"000000000",
  23952=>"000100000",
  23953=>"000010000",
  23954=>"010001001",
  23955=>"001001110",
  23956=>"111110000",
  23957=>"000111010",
  23958=>"100010101",
  23959=>"100111111",
  23960=>"101010001",
  23961=>"000111001",
  23962=>"110010110",
  23963=>"010000010",
  23964=>"101101011",
  23965=>"001011011",
  23966=>"001111100",
  23967=>"100010011",
  23968=>"101000000",
  23969=>"001110100",
  23970=>"111010011",
  23971=>"101011110",
  23972=>"101101111",
  23973=>"100001100",
  23974=>"010100001",
  23975=>"101111010",
  23976=>"000111100",
  23977=>"100000000",
  23978=>"010001000",
  23979=>"101101101",
  23980=>"100110000",
  23981=>"000011100",
  23982=>"000101101",
  23983=>"110110100",
  23984=>"100101111",
  23985=>"111010010",
  23986=>"101110101",
  23987=>"001001010",
  23988=>"111001000",
  23989=>"110110011",
  23990=>"110111011",
  23991=>"001000011",
  23992=>"100000000",
  23993=>"010010000",
  23994=>"000000011",
  23995=>"010010011",
  23996=>"000100111",
  23997=>"000100111",
  23998=>"011111000",
  23999=>"101011110",
  24000=>"000011011",
  24001=>"101011100",
  24002=>"001001011",
  24003=>"000000101",
  24004=>"100100111",
  24005=>"110111101",
  24006=>"000010011",
  24007=>"101001101",
  24008=>"111100100",
  24009=>"110101100",
  24010=>"101010000",
  24011=>"011110001",
  24012=>"111100100",
  24013=>"000101011",
  24014=>"101100001",
  24015=>"111001110",
  24016=>"001111000",
  24017=>"111010110",
  24018=>"011000110",
  24019=>"001010000",
  24020=>"011000011",
  24021=>"000010111",
  24022=>"100011100",
  24023=>"001000101",
  24024=>"011010011",
  24025=>"110001011",
  24026=>"111111000",
  24027=>"111000001",
  24028=>"111000111",
  24029=>"100001001",
  24030=>"011011001",
  24031=>"111011100",
  24032=>"101001100",
  24033=>"110010000",
  24034=>"100100110",
  24035=>"001000110",
  24036=>"101101010",
  24037=>"111110001",
  24038=>"111000000",
  24039=>"001010010",
  24040=>"110111111",
  24041=>"111111100",
  24042=>"100011101",
  24043=>"001011110",
  24044=>"001100100",
  24045=>"100100000",
  24046=>"000000110",
  24047=>"000001101",
  24048=>"000001001",
  24049=>"100111011",
  24050=>"101001010",
  24051=>"000001001",
  24052=>"111110010",
  24053=>"011010011",
  24054=>"101000110",
  24055=>"111111101",
  24056=>"000010001",
  24057=>"000101110",
  24058=>"000000110",
  24059=>"000111011",
  24060=>"000000101",
  24061=>"101101010",
  24062=>"111110010",
  24063=>"001010111",
  24064=>"101110000",
  24065=>"110101000",
  24066=>"101110110",
  24067=>"110010000",
  24068=>"000110001",
  24069=>"111100001",
  24070=>"101101110",
  24071=>"011001111",
  24072=>"011110100",
  24073=>"111100110",
  24074=>"011001001",
  24075=>"001111000",
  24076=>"001010111",
  24077=>"100000000",
  24078=>"101100001",
  24079=>"110100100",
  24080=>"101100000",
  24081=>"000000001",
  24082=>"011000000",
  24083=>"000101001",
  24084=>"100001011",
  24085=>"100011111",
  24086=>"010011100",
  24087=>"000001100",
  24088=>"010000001",
  24089=>"110110101",
  24090=>"001110101",
  24091=>"010000100",
  24092=>"100100110",
  24093=>"110111100",
  24094=>"101111001",
  24095=>"010101011",
  24096=>"011100001",
  24097=>"111110001",
  24098=>"101111010",
  24099=>"110101110",
  24100=>"111111110",
  24101=>"100011111",
  24102=>"111110111",
  24103=>"000100010",
  24104=>"101111000",
  24105=>"000010100",
  24106=>"101000101",
  24107=>"000001101",
  24108=>"010010101",
  24109=>"110000011",
  24110=>"010101001",
  24111=>"000011011",
  24112=>"001000001",
  24113=>"101101101",
  24114=>"011110001",
  24115=>"100001011",
  24116=>"111011000",
  24117=>"111111111",
  24118=>"111011100",
  24119=>"001111110",
  24120=>"110010100",
  24121=>"110001011",
  24122=>"001110011",
  24123=>"110011111",
  24124=>"111101011",
  24125=>"010110001",
  24126=>"110100101",
  24127=>"111000001",
  24128=>"101100000",
  24129=>"111100111",
  24130=>"011011101",
  24131=>"000110000",
  24132=>"010101010",
  24133=>"111011100",
  24134=>"110001100",
  24135=>"010011001",
  24136=>"001001100",
  24137=>"000110010",
  24138=>"001100011",
  24139=>"101100101",
  24140=>"001110011",
  24141=>"100001100",
  24142=>"001111110",
  24143=>"000100110",
  24144=>"000101001",
  24145=>"000010110",
  24146=>"001001110",
  24147=>"111110010",
  24148=>"101000110",
  24149=>"001010001",
  24150=>"100100100",
  24151=>"001011110",
  24152=>"000001011",
  24153=>"010011111",
  24154=>"001011111",
  24155=>"101000010",
  24156=>"110101100",
  24157=>"000101000",
  24158=>"100101101",
  24159=>"000010110",
  24160=>"011011110",
  24161=>"000110110",
  24162=>"001100001",
  24163=>"000110001",
  24164=>"011000100",
  24165=>"001100000",
  24166=>"011110010",
  24167=>"100110011",
  24168=>"101111000",
  24169=>"000111111",
  24170=>"001001111",
  24171=>"010101010",
  24172=>"110001001",
  24173=>"110111101",
  24174=>"111011010",
  24175=>"101001001",
  24176=>"011101001",
  24177=>"101101001",
  24178=>"101101100",
  24179=>"010001101",
  24180=>"000001111",
  24181=>"100111010",
  24182=>"011001001",
  24183=>"001010100",
  24184=>"000010000",
  24185=>"110111110",
  24186=>"001011001",
  24187=>"011111101",
  24188=>"000011110",
  24189=>"000010010",
  24190=>"010000110",
  24191=>"110110100",
  24192=>"011100110",
  24193=>"100100001",
  24194=>"001001011",
  24195=>"011011011",
  24196=>"111001110",
  24197=>"101100000",
  24198=>"100011001",
  24199=>"000001010",
  24200=>"000100000",
  24201=>"000101100",
  24202=>"111001111",
  24203=>"111100110",
  24204=>"101011101",
  24205=>"000111110",
  24206=>"011101111",
  24207=>"111011110",
  24208=>"100100001",
  24209=>"111011111",
  24210=>"000000101",
  24211=>"000110101",
  24212=>"101101001",
  24213=>"100011111",
  24214=>"010100001",
  24215=>"010011000",
  24216=>"101011100",
  24217=>"000000001",
  24218=>"101111110",
  24219=>"010010010",
  24220=>"111000111",
  24221=>"111000111",
  24222=>"001000111",
  24223=>"001101100",
  24224=>"111100111",
  24225=>"100110001",
  24226=>"111101111",
  24227=>"010000101",
  24228=>"011110000",
  24229=>"010001110",
  24230=>"111101110",
  24231=>"000010111",
  24232=>"010011000",
  24233=>"010001011",
  24234=>"100100100",
  24235=>"001100010",
  24236=>"111100000",
  24237=>"110001001",
  24238=>"101100101",
  24239=>"000000101",
  24240=>"100111100",
  24241=>"110111111",
  24242=>"000100100",
  24243=>"001101111",
  24244=>"001111011",
  24245=>"100101111",
  24246=>"010111001",
  24247=>"011001011",
  24248=>"111100100",
  24249=>"110100101",
  24250=>"110100000",
  24251=>"000111100",
  24252=>"101011101",
  24253=>"101101011",
  24254=>"010000110",
  24255=>"000101011",
  24256=>"000001001",
  24257=>"100100110",
  24258=>"000111010",
  24259=>"100111110",
  24260=>"010010111",
  24261=>"100000110",
  24262=>"100000010",
  24263=>"010000001",
  24264=>"110111001",
  24265=>"111101101",
  24266=>"010010110",
  24267=>"100111101",
  24268=>"101100001",
  24269=>"010101010",
  24270=>"100010001",
  24271=>"010110101",
  24272=>"111111011",
  24273=>"101010011",
  24274=>"000101101",
  24275=>"010011111",
  24276=>"010011010",
  24277=>"010010000",
  24278=>"000110110",
  24279=>"001011101",
  24280=>"000001001",
  24281=>"100100000",
  24282=>"011000011",
  24283=>"010110100",
  24284=>"010110010",
  24285=>"111101010",
  24286=>"010001111",
  24287=>"110001100",
  24288=>"000000000",
  24289=>"110000011",
  24290=>"101110111",
  24291=>"111011011",
  24292=>"100101010",
  24293=>"011011101",
  24294=>"111000001",
  24295=>"101100101",
  24296=>"101100101",
  24297=>"100100001",
  24298=>"111111001",
  24299=>"011001100",
  24300=>"011011001",
  24301=>"000101110",
  24302=>"000110101",
  24303=>"100100001",
  24304=>"101000100",
  24305=>"000001100",
  24306=>"110111100",
  24307=>"011101100",
  24308=>"101001010",
  24309=>"101101000",
  24310=>"001001101",
  24311=>"110110111",
  24312=>"100111010",
  24313=>"000001101",
  24314=>"000010011",
  24315=>"111100000",
  24316=>"111100010",
  24317=>"100111111",
  24318=>"100100110",
  24319=>"111110111",
  24320=>"011000001",
  24321=>"010111000",
  24322=>"001111011",
  24323=>"010011110",
  24324=>"011111000",
  24325=>"011011101",
  24326=>"101010110",
  24327=>"111010110",
  24328=>"001101100",
  24329=>"001010000",
  24330=>"110100100",
  24331=>"001101100",
  24332=>"010100100",
  24333=>"100000010",
  24334=>"111111110",
  24335=>"101100100",
  24336=>"011000100",
  24337=>"101010000",
  24338=>"011011000",
  24339=>"100101100",
  24340=>"111011000",
  24341=>"001011000",
  24342=>"101111001",
  24343=>"101110100",
  24344=>"100011100",
  24345=>"100001000",
  24346=>"011101001",
  24347=>"010111111",
  24348=>"101100001",
  24349=>"101010110",
  24350=>"100101010",
  24351=>"011110110",
  24352=>"110111011",
  24353=>"000000101",
  24354=>"111110000",
  24355=>"111111100",
  24356=>"011000000",
  24357=>"101010111",
  24358=>"110100101",
  24359=>"010000000",
  24360=>"011001100",
  24361=>"001101100",
  24362=>"010100011",
  24363=>"110101101",
  24364=>"100001001",
  24365=>"101000000",
  24366=>"110100100",
  24367=>"111101010",
  24368=>"100000111",
  24369=>"011101101",
  24370=>"000011010",
  24371=>"100011100",
  24372=>"111001011",
  24373=>"110110100",
  24374=>"001101011",
  24375=>"100110110",
  24376=>"111001111",
  24377=>"111110110",
  24378=>"010010110",
  24379=>"101111100",
  24380=>"000000000",
  24381=>"010101110",
  24382=>"001011000",
  24383=>"000000100",
  24384=>"000100100",
  24385=>"110010101",
  24386=>"110001111",
  24387=>"100111000",
  24388=>"101010000",
  24389=>"001110001",
  24390=>"010001001",
  24391=>"110000100",
  24392=>"111111011",
  24393=>"111111101",
  24394=>"101001001",
  24395=>"000001100",
  24396=>"011101111",
  24397=>"101010010",
  24398=>"001111110",
  24399=>"100111111",
  24400=>"100010000",
  24401=>"110110001",
  24402=>"110101101",
  24403=>"011011001",
  24404=>"010000101",
  24405=>"111000110",
  24406=>"111010100",
  24407=>"100001110",
  24408=>"100110000",
  24409=>"110111011",
  24410=>"001100111",
  24411=>"101001011",
  24412=>"101011010",
  24413=>"011100101",
  24414=>"100001001",
  24415=>"110000100",
  24416=>"111101110",
  24417=>"100000010",
  24418=>"010010111",
  24419=>"110100100",
  24420=>"111101101",
  24421=>"110000110",
  24422=>"111111000",
  24423=>"101100100",
  24424=>"011011110",
  24425=>"011001010",
  24426=>"001001100",
  24427=>"111000000",
  24428=>"110101100",
  24429=>"101100111",
  24430=>"001101001",
  24431=>"010110110",
  24432=>"000000001",
  24433=>"111010000",
  24434=>"110111110",
  24435=>"100111001",
  24436=>"111110000",
  24437=>"101010000",
  24438=>"101110010",
  24439=>"011011010",
  24440=>"110110110",
  24441=>"110111100",
  24442=>"110000101",
  24443=>"000110111",
  24444=>"100100000",
  24445=>"101000110",
  24446=>"101101111",
  24447=>"101100101",
  24448=>"110110011",
  24449=>"101111010",
  24450=>"010111101",
  24451=>"110110111",
  24452=>"100010000",
  24453=>"111111010",
  24454=>"000100000",
  24455=>"101100011",
  24456=>"110001101",
  24457=>"001100110",
  24458=>"001011001",
  24459=>"111011111",
  24460=>"010000010",
  24461=>"010000001",
  24462=>"011000111",
  24463=>"101001011",
  24464=>"101111000",
  24465=>"101101100",
  24466=>"011011100",
  24467=>"110111001",
  24468=>"111011000",
  24469=>"000000001",
  24470=>"001110110",
  24471=>"000010110",
  24472=>"100101011",
  24473=>"010000011",
  24474=>"111101001",
  24475=>"101111011",
  24476=>"100111111",
  24477=>"101110010",
  24478=>"101101011",
  24479=>"100001010",
  24480=>"000000010",
  24481=>"111111000",
  24482=>"001100001",
  24483=>"110101110",
  24484=>"001011000",
  24485=>"000001001",
  24486=>"010100101",
  24487=>"110111110",
  24488=>"011111110",
  24489=>"010001010",
  24490=>"011111100",
  24491=>"011101011",
  24492=>"011001001",
  24493=>"001001100",
  24494=>"101010000",
  24495=>"100000110",
  24496=>"011101000",
  24497=>"011011111",
  24498=>"110001010",
  24499=>"010000000",
  24500=>"111010110",
  24501=>"001000001",
  24502=>"001110100",
  24503=>"101100111",
  24504=>"101000101",
  24505=>"010110111",
  24506=>"100011111",
  24507=>"101010010",
  24508=>"010101101",
  24509=>"010010010",
  24510=>"101100111",
  24511=>"111011001",
  24512=>"010111010",
  24513=>"101100100",
  24514=>"110101111",
  24515=>"110111111",
  24516=>"000011010",
  24517=>"000100001",
  24518=>"110000000",
  24519=>"010010100",
  24520=>"111100011",
  24521=>"101011101",
  24522=>"111111000",
  24523=>"001110110",
  24524=>"110110010",
  24525=>"000110110",
  24526=>"110000110",
  24527=>"000101111",
  24528=>"001101101",
  24529=>"000010001",
  24530=>"010000111",
  24531=>"111101110",
  24532=>"001010101",
  24533=>"011111100",
  24534=>"011111001",
  24535=>"001000000",
  24536=>"010000010",
  24537=>"010111011",
  24538=>"000011100",
  24539=>"011001101",
  24540=>"010001001",
  24541=>"011111011",
  24542=>"011111001",
  24543=>"100000110",
  24544=>"111110011",
  24545=>"101000001",
  24546=>"100100111",
  24547=>"110001011",
  24548=>"100101010",
  24549=>"000000010",
  24550=>"000001011",
  24551=>"110001110",
  24552=>"100110111",
  24553=>"000111000",
  24554=>"111111100",
  24555=>"100110001",
  24556=>"111010011",
  24557=>"100001111",
  24558=>"011000101",
  24559=>"010001100",
  24560=>"101100011",
  24561=>"101110111",
  24562=>"110010111",
  24563=>"011010111",
  24564=>"000000110",
  24565=>"000001010",
  24566=>"100001011",
  24567=>"010001000",
  24568=>"010101101",
  24569=>"100110001",
  24570=>"011111111",
  24571=>"111010000",
  24572=>"000001111",
  24573=>"011010110",
  24574=>"001101010",
  24575=>"001000010",
  24576=>"001010010",
  24577=>"111110011",
  24578=>"010110111",
  24579=>"001101010",
  24580=>"011000110",
  24581=>"000100111",
  24582=>"010110010",
  24583=>"111011100",
  24584=>"111101010",
  24585=>"000111001",
  24586=>"010101101",
  24587=>"111110111",
  24588=>"000101100",
  24589=>"101011110",
  24590=>"011111111",
  24591=>"001101010",
  24592=>"111101101",
  24593=>"010011101",
  24594=>"000010011",
  24595=>"011110001",
  24596=>"010111111",
  24597=>"010001100",
  24598=>"010000011",
  24599=>"100001001",
  24600=>"111000001",
  24601=>"101001011",
  24602=>"001011100",
  24603=>"111000010",
  24604=>"101101010",
  24605=>"010100010",
  24606=>"000010110",
  24607=>"000000010",
  24608=>"001000101",
  24609=>"000010000",
  24610=>"100000001",
  24611=>"000111111",
  24612=>"001111010",
  24613=>"101010001",
  24614=>"001110010",
  24615=>"000101100",
  24616=>"110110010",
  24617=>"111101101",
  24618=>"110011010",
  24619=>"001100100",
  24620=>"001111011",
  24621=>"101101000",
  24622=>"111001110",
  24623=>"111111111",
  24624=>"000000001",
  24625=>"101101001",
  24626=>"010100000",
  24627=>"011111100",
  24628=>"000100110",
  24629=>"001111001",
  24630=>"001111101",
  24631=>"001000000",
  24632=>"110011100",
  24633=>"010000001",
  24634=>"111011000",
  24635=>"110100011",
  24636=>"001001011",
  24637=>"010101111",
  24638=>"101111011",
  24639=>"010111111",
  24640=>"111100101",
  24641=>"111001000",
  24642=>"101001001",
  24643=>"011101111",
  24644=>"110110000",
  24645=>"001101110",
  24646=>"100001000",
  24647=>"110111101",
  24648=>"111100010",
  24649=>"011101111",
  24650=>"111101101",
  24651=>"000001101",
  24652=>"111010001",
  24653=>"010000110",
  24654=>"011011011",
  24655=>"010010110",
  24656=>"000111010",
  24657=>"001110000",
  24658=>"010111100",
  24659=>"111100001",
  24660=>"010011111",
  24661=>"000001011",
  24662=>"011011010",
  24663=>"111110100",
  24664=>"101001110",
  24665=>"000001111",
  24666=>"000111111",
  24667=>"111101111",
  24668=>"111101111",
  24669=>"111001000",
  24670=>"010101100",
  24671=>"100011011",
  24672=>"010010011",
  24673=>"100011110",
  24674=>"001110100",
  24675=>"101011111",
  24676=>"010011010",
  24677=>"000100110",
  24678=>"110101111",
  24679=>"111101100",
  24680=>"000111111",
  24681=>"001001100",
  24682=>"111111110",
  24683=>"110101011",
  24684=>"111110100",
  24685=>"111001000",
  24686=>"101011001",
  24687=>"100001000",
  24688=>"110010110",
  24689=>"101101010",
  24690=>"011010011",
  24691=>"100011110",
  24692=>"110000011",
  24693=>"010100101",
  24694=>"001100001",
  24695=>"001001111",
  24696=>"100011011",
  24697=>"101111100",
  24698=>"000001011",
  24699=>"001001011",
  24700=>"000001100",
  24701=>"110101010",
  24702=>"011100001",
  24703=>"000011001",
  24704=>"010000101",
  24705=>"010010010",
  24706=>"101110110",
  24707=>"100010101",
  24708=>"010101000",
  24709=>"110111110",
  24710=>"010000110",
  24711=>"110111011",
  24712=>"100000101",
  24713=>"111000010",
  24714=>"100100000",
  24715=>"111100011",
  24716=>"001101001",
  24717=>"000100001",
  24718=>"000001011",
  24719=>"010101111",
  24720=>"000001100",
  24721=>"111111110",
  24722=>"001111011",
  24723=>"000000010",
  24724=>"101000111",
  24725=>"100111110",
  24726=>"101001110",
  24727=>"111110000",
  24728=>"100011111",
  24729=>"101111001",
  24730=>"001011000",
  24731=>"011111110",
  24732=>"110111001",
  24733=>"111111101",
  24734=>"000101000",
  24735=>"110010101",
  24736=>"010101001",
  24737=>"011011000",
  24738=>"010010110",
  24739=>"100110100",
  24740=>"111000001",
  24741=>"001000111",
  24742=>"011010110",
  24743=>"111001011",
  24744=>"010001010",
  24745=>"110011100",
  24746=>"001001110",
  24747=>"011000001",
  24748=>"011100000",
  24749=>"001101101",
  24750=>"010101000",
  24751=>"111001110",
  24752=>"100000000",
  24753=>"000110010",
  24754=>"000011100",
  24755=>"110110010",
  24756=>"001100001",
  24757=>"101010010",
  24758=>"010011100",
  24759=>"100110000",
  24760=>"110101010",
  24761=>"100111101",
  24762=>"111000001",
  24763=>"111101011",
  24764=>"101011010",
  24765=>"011100100",
  24766=>"110101000",
  24767=>"101000001",
  24768=>"000001000",
  24769=>"011111111",
  24770=>"100101111",
  24771=>"111100111",
  24772=>"110110000",
  24773=>"101110110",
  24774=>"000110100",
  24775=>"001110000",
  24776=>"100100100",
  24777=>"011001101",
  24778=>"001001000",
  24779=>"011100100",
  24780=>"010010100",
  24781=>"101011001",
  24782=>"111000011",
  24783=>"001111100",
  24784=>"111111011",
  24785=>"010011001",
  24786=>"100001111",
  24787=>"001101010",
  24788=>"000100001",
  24789=>"101111010",
  24790=>"111101010",
  24791=>"101001001",
  24792=>"000000011",
  24793=>"011010100",
  24794=>"100101101",
  24795=>"001011001",
  24796=>"001010101",
  24797=>"010110000",
  24798=>"111011001",
  24799=>"101111011",
  24800=>"111111110",
  24801=>"011110100",
  24802=>"100001110",
  24803=>"110011111",
  24804=>"000101010",
  24805=>"110000110",
  24806=>"000011011",
  24807=>"010000001",
  24808=>"111110010",
  24809=>"101111001",
  24810=>"111001010",
  24811=>"110100001",
  24812=>"101110001",
  24813=>"111001111",
  24814=>"010011101",
  24815=>"010010111",
  24816=>"000110111",
  24817=>"010100010",
  24818=>"100110111",
  24819=>"010011100",
  24820=>"100101100",
  24821=>"011000001",
  24822=>"111000100",
  24823=>"111101010",
  24824=>"010011111",
  24825=>"000000110",
  24826=>"010001100",
  24827=>"100101001",
  24828=>"101100100",
  24829=>"111000000",
  24830=>"000011111",
  24831=>"010110000",
  24832=>"000000000",
  24833=>"011111001",
  24834=>"010001011",
  24835=>"001100111",
  24836=>"011111011",
  24837=>"001100111",
  24838=>"111001010",
  24839=>"111000010",
  24840=>"101001101",
  24841=>"100010000",
  24842=>"010000110",
  24843=>"010100110",
  24844=>"011101011",
  24845=>"000001110",
  24846=>"111010001",
  24847=>"101000100",
  24848=>"101000011",
  24849=>"110010010",
  24850=>"101111000",
  24851=>"010101011",
  24852=>"111011110",
  24853=>"100100110",
  24854=>"010100101",
  24855=>"010000011",
  24856=>"111111111",
  24857=>"011100001",
  24858=>"111000110",
  24859=>"111101011",
  24860=>"100000000",
  24861=>"001000111",
  24862=>"100001010",
  24863=>"111000101",
  24864=>"001111001",
  24865=>"110011101",
  24866=>"101101110",
  24867=>"011110101",
  24868=>"111001111",
  24869=>"011000000",
  24870=>"110010111",
  24871=>"110101110",
  24872=>"101011111",
  24873=>"111011110",
  24874=>"110010110",
  24875=>"110000101",
  24876=>"001001000",
  24877=>"010000110",
  24878=>"101000001",
  24879=>"000010110",
  24880=>"011100011",
  24881=>"011011100",
  24882=>"110111110",
  24883=>"011111010",
  24884=>"110011100",
  24885=>"101100001",
  24886=>"101010100",
  24887=>"101110100",
  24888=>"100010111",
  24889=>"011010011",
  24890=>"001000010",
  24891=>"110000000",
  24892=>"011111100",
  24893=>"101110001",
  24894=>"111100101",
  24895=>"010000001",
  24896=>"100110110",
  24897=>"001110110",
  24898=>"010011000",
  24899=>"101011011",
  24900=>"000110100",
  24901=>"011100101",
  24902=>"110000110",
  24903=>"001110001",
  24904=>"101001001",
  24905=>"000001001",
  24906=>"101000000",
  24907=>"000000011",
  24908=>"010000010",
  24909=>"100110100",
  24910=>"001100010",
  24911=>"110110101",
  24912=>"110100000",
  24913=>"110100011",
  24914=>"111110000",
  24915=>"000111011",
  24916=>"100100001",
  24917=>"110000101",
  24918=>"000000110",
  24919=>"001000010",
  24920=>"110000011",
  24921=>"111001000",
  24922=>"001110100",
  24923=>"000000100",
  24924=>"000110110",
  24925=>"001011001",
  24926=>"010000010",
  24927=>"101010111",
  24928=>"101111011",
  24929=>"001101011",
  24930=>"000101001",
  24931=>"010000100",
  24932=>"110010001",
  24933=>"111110001",
  24934=>"011011010",
  24935=>"110010011",
  24936=>"100001011",
  24937=>"101000010",
  24938=>"110011000",
  24939=>"101011000",
  24940=>"010100001",
  24941=>"101101100",
  24942=>"111111011",
  24943=>"101101101",
  24944=>"010001100",
  24945=>"000010101",
  24946=>"000001100",
  24947=>"100111110",
  24948=>"000100110",
  24949=>"001110010",
  24950=>"111101000",
  24951=>"001011001",
  24952=>"110100011",
  24953=>"010111011",
  24954=>"011101011",
  24955=>"011101011",
  24956=>"001000010",
  24957=>"001011101",
  24958=>"100000100",
  24959=>"000110011",
  24960=>"110101100",
  24961=>"000001100",
  24962=>"110001000",
  24963=>"100001111",
  24964=>"000011101",
  24965=>"010010110",
  24966=>"000101101",
  24967=>"101101011",
  24968=>"011101011",
  24969=>"000011100",
  24970=>"101001011",
  24971=>"101101001",
  24972=>"000100011",
  24973=>"001010010",
  24974=>"010100110",
  24975=>"000100101",
  24976=>"000111111",
  24977=>"101000000",
  24978=>"000000101",
  24979=>"000001000",
  24980=>"000010101",
  24981=>"101000100",
  24982=>"011000011",
  24983=>"111001001",
  24984=>"111010101",
  24985=>"010001100",
  24986=>"101001001",
  24987=>"100111011",
  24988=>"110011110",
  24989=>"000101001",
  24990=>"111000000",
  24991=>"011011010",
  24992=>"001010100",
  24993=>"010101110",
  24994=>"001010110",
  24995=>"001110110",
  24996=>"101101101",
  24997=>"101111010",
  24998=>"000010001",
  24999=>"001101110",
  25000=>"001011100",
  25001=>"101100011",
  25002=>"100000100",
  25003=>"111110101",
  25004=>"011101000",
  25005=>"001010111",
  25006=>"001011010",
  25007=>"101010101",
  25008=>"110000000",
  25009=>"001000000",
  25010=>"000110111",
  25011=>"110111110",
  25012=>"011011010",
  25013=>"101000001",
  25014=>"111011100",
  25015=>"100110101",
  25016=>"111111111",
  25017=>"111001010",
  25018=>"101011111",
  25019=>"101110100",
  25020=>"000011001",
  25021=>"110110000",
  25022=>"011101010",
  25023=>"111001001",
  25024=>"100110010",
  25025=>"100110011",
  25026=>"100011011",
  25027=>"101100010",
  25028=>"001010101",
  25029=>"110000011",
  25030=>"011011011",
  25031=>"011101110",
  25032=>"101010111",
  25033=>"101101110",
  25034=>"011011101",
  25035=>"010101010",
  25036=>"001111010",
  25037=>"101000010",
  25038=>"101011101",
  25039=>"111011111",
  25040=>"100001000",
  25041=>"011100110",
  25042=>"010011110",
  25043=>"010100011",
  25044=>"110001000",
  25045=>"000101110",
  25046=>"110001000",
  25047=>"111101110",
  25048=>"110110101",
  25049=>"001111111",
  25050=>"001110101",
  25051=>"001011100",
  25052=>"010000101",
  25053=>"001011101",
  25054=>"010100111",
  25055=>"111010010",
  25056=>"011001100",
  25057=>"101001001",
  25058=>"011010000",
  25059=>"010100010",
  25060=>"010000001",
  25061=>"111101000",
  25062=>"000000000",
  25063=>"010010101",
  25064=>"101100010",
  25065=>"001011110",
  25066=>"111010010",
  25067=>"111010100",
  25068=>"011111001",
  25069=>"011011010",
  25070=>"100011100",
  25071=>"000101001",
  25072=>"111011000",
  25073=>"110000100",
  25074=>"000001111",
  25075=>"010001101",
  25076=>"110111011",
  25077=>"010111000",
  25078=>"110000100",
  25079=>"100001010",
  25080=>"000001101",
  25081=>"101010101",
  25082=>"111000010",
  25083=>"010110111",
  25084=>"111011111",
  25085=>"010111010",
  25086=>"100001001",
  25087=>"101010011",
  25088=>"000100110",
  25089=>"100000100",
  25090=>"100000000",
  25091=>"001100101",
  25092=>"100001001",
  25093=>"101100111",
  25094=>"011100100",
  25095=>"011011011",
  25096=>"010100111",
  25097=>"010000010",
  25098=>"010110001",
  25099=>"001000001",
  25100=>"101100110",
  25101=>"110101011",
  25102=>"001000011",
  25103=>"011111100",
  25104=>"011101101",
  25105=>"111000011",
  25106=>"010101110",
  25107=>"101100111",
  25108=>"011001011",
  25109=>"010111001",
  25110=>"101000100",
  25111=>"011100001",
  25112=>"000111010",
  25113=>"111110001",
  25114=>"000101110",
  25115=>"100001000",
  25116=>"000111111",
  25117=>"011011110",
  25118=>"001111100",
  25119=>"110110100",
  25120=>"111001011",
  25121=>"000111000",
  25122=>"011011100",
  25123=>"110111100",
  25124=>"110000111",
  25125=>"010011110",
  25126=>"000110111",
  25127=>"100011000",
  25128=>"001000011",
  25129=>"001010000",
  25130=>"101111111",
  25131=>"100100001",
  25132=>"110111011",
  25133=>"001000010",
  25134=>"111110100",
  25135=>"001000100",
  25136=>"110010001",
  25137=>"000011011",
  25138=>"000000001",
  25139=>"100111110",
  25140=>"010100000",
  25141=>"001110111",
  25142=>"101111110",
  25143=>"010010110",
  25144=>"010001010",
  25145=>"001000101",
  25146=>"101010111",
  25147=>"111011101",
  25148=>"010001000",
  25149=>"000011100",
  25150=>"110111011",
  25151=>"100111111",
  25152=>"001101001",
  25153=>"111111000",
  25154=>"011111111",
  25155=>"010100101",
  25156=>"010001000",
  25157=>"001100101",
  25158=>"110000010",
  25159=>"111001100",
  25160=>"110011101",
  25161=>"101011101",
  25162=>"101000111",
  25163=>"111111010",
  25164=>"100001001",
  25165=>"011010010",
  25166=>"110111100",
  25167=>"000100110",
  25168=>"001011100",
  25169=>"000100111",
  25170=>"001110100",
  25171=>"011100011",
  25172=>"011000111",
  25173=>"111100111",
  25174=>"110100111",
  25175=>"010010000",
  25176=>"000000111",
  25177=>"001000011",
  25178=>"010101011",
  25179=>"010100111",
  25180=>"011110010",
  25181=>"011011110",
  25182=>"011001011",
  25183=>"011111101",
  25184=>"110101100",
  25185=>"111101011",
  25186=>"110111010",
  25187=>"101111111",
  25188=>"110010101",
  25189=>"101000010",
  25190=>"011001011",
  25191=>"110000100",
  25192=>"001011010",
  25193=>"101011011",
  25194=>"101111101",
  25195=>"000101010",
  25196=>"000001000",
  25197=>"111100011",
  25198=>"110100101",
  25199=>"001100010",
  25200=>"111110111",
  25201=>"110010110",
  25202=>"011001010",
  25203=>"011111100",
  25204=>"111011110",
  25205=>"111111110",
  25206=>"100100101",
  25207=>"000100011",
  25208=>"111000001",
  25209=>"111001000",
  25210=>"111000101",
  25211=>"011100011",
  25212=>"011000001",
  25213=>"000010110",
  25214=>"000000101",
  25215=>"011001110",
  25216=>"111111101",
  25217=>"110010111",
  25218=>"010000101",
  25219=>"000011011",
  25220=>"001111010",
  25221=>"000100010",
  25222=>"011110101",
  25223=>"010110110",
  25224=>"101010010",
  25225=>"111100110",
  25226=>"011000101",
  25227=>"010001111",
  25228=>"110000010",
  25229=>"101110000",
  25230=>"110111111",
  25231=>"111111100",
  25232=>"000110011",
  25233=>"011111110",
  25234=>"110000011",
  25235=>"010001001",
  25236=>"000010011",
  25237=>"111000111",
  25238=>"111101101",
  25239=>"111000011",
  25240=>"111010101",
  25241=>"010100000",
  25242=>"111000010",
  25243=>"001011101",
  25244=>"111101111",
  25245=>"000100011",
  25246=>"010001000",
  25247=>"100100010",
  25248=>"110101111",
  25249=>"101111101",
  25250=>"000100011",
  25251=>"101101001",
  25252=>"111111001",
  25253=>"101110111",
  25254=>"100110001",
  25255=>"011000101",
  25256=>"101100110",
  25257=>"111100011",
  25258=>"000011110",
  25259=>"011101110",
  25260=>"110111110",
  25261=>"110001100",
  25262=>"000001010",
  25263=>"100011011",
  25264=>"010110101",
  25265=>"010000010",
  25266=>"010010010",
  25267=>"110011101",
  25268=>"101110110",
  25269=>"100011111",
  25270=>"101101111",
  25271=>"001101011",
  25272=>"001101110",
  25273=>"101001111",
  25274=>"010000010",
  25275=>"110001000",
  25276=>"101010100",
  25277=>"011001111",
  25278=>"011100111",
  25279=>"110010010",
  25280=>"010000010",
  25281=>"101110010",
  25282=>"010010000",
  25283=>"000101111",
  25284=>"000101010",
  25285=>"110101000",
  25286=>"010101111",
  25287=>"011001110",
  25288=>"110101100",
  25289=>"001110001",
  25290=>"110000000",
  25291=>"011001000",
  25292=>"010101011",
  25293=>"111001111",
  25294=>"100010111",
  25295=>"101011101",
  25296=>"011000001",
  25297=>"111111010",
  25298=>"010001100",
  25299=>"101010110",
  25300=>"100010011",
  25301=>"110101000",
  25302=>"101111010",
  25303=>"010010100",
  25304=>"100010110",
  25305=>"111111100",
  25306=>"000111001",
  25307=>"010111001",
  25308=>"001011010",
  25309=>"100001011",
  25310=>"001110010",
  25311=>"010011000",
  25312=>"100001101",
  25313=>"111011110",
  25314=>"110101011",
  25315=>"111110010",
  25316=>"100111001",
  25317=>"110000110",
  25318=>"011111000",
  25319=>"111100010",
  25320=>"111110101",
  25321=>"111001001",
  25322=>"000001110",
  25323=>"010110000",
  25324=>"000010111",
  25325=>"011000001",
  25326=>"011110100",
  25327=>"011011001",
  25328=>"100010011",
  25329=>"001011101",
  25330=>"011011011",
  25331=>"111000110",
  25332=>"110101110",
  25333=>"101000100",
  25334=>"001001111",
  25335=>"101101110",
  25336=>"111111101",
  25337=>"010001000",
  25338=>"101110010",
  25339=>"000101111",
  25340=>"000000011",
  25341=>"010001011",
  25342=>"100011001",
  25343=>"111000101",
  25344=>"111010110",
  25345=>"111101100",
  25346=>"111111111",
  25347=>"111100110",
  25348=>"001000010",
  25349=>"011110101",
  25350=>"010110010",
  25351=>"100111100",
  25352=>"110110111",
  25353=>"000000110",
  25354=>"001100100",
  25355=>"110011001",
  25356=>"010010000",
  25357=>"010001011",
  25358=>"011000001",
  25359=>"010110101",
  25360=>"100011010",
  25361=>"101000001",
  25362=>"100101011",
  25363=>"011010011",
  25364=>"000000011",
  25365=>"000000001",
  25366=>"001010111",
  25367=>"001110000",
  25368=>"110010111",
  25369=>"111001101",
  25370=>"100101010",
  25371=>"000110001",
  25372=>"100110010",
  25373=>"000101010",
  25374=>"000010110",
  25375=>"110101011",
  25376=>"010100011",
  25377=>"010111111",
  25378=>"111100101",
  25379=>"000101101",
  25380=>"000110011",
  25381=>"101110010",
  25382=>"101011000",
  25383=>"100011110",
  25384=>"010110100",
  25385=>"101110011",
  25386=>"101010001",
  25387=>"000001000",
  25388=>"110111101",
  25389=>"100010010",
  25390=>"001101111",
  25391=>"000111111",
  25392=>"101111001",
  25393=>"001011110",
  25394=>"110001000",
  25395=>"011100000",
  25396=>"001100001",
  25397=>"001100010",
  25398=>"100000000",
  25399=>"011111000",
  25400=>"010000111",
  25401=>"101010111",
  25402=>"111000111",
  25403=>"110111011",
  25404=>"111101001",
  25405=>"011000100",
  25406=>"010100000",
  25407=>"011001111",
  25408=>"100111111",
  25409=>"001011110",
  25410=>"111110100",
  25411=>"000010001",
  25412=>"001110111",
  25413=>"001000110",
  25414=>"100010010",
  25415=>"101101010",
  25416=>"110110000",
  25417=>"000101101",
  25418=>"111101011",
  25419=>"101000010",
  25420=>"110100000",
  25421=>"001100101",
  25422=>"101100010",
  25423=>"111100000",
  25424=>"001100000",
  25425=>"000111101",
  25426=>"110100000",
  25427=>"001101110",
  25428=>"101111001",
  25429=>"111100101",
  25430=>"101011110",
  25431=>"110101110",
  25432=>"111001011",
  25433=>"010011111",
  25434=>"110011110",
  25435=>"000000100",
  25436=>"001010101",
  25437=>"110111111",
  25438=>"001100000",
  25439=>"101010010",
  25440=>"000111000",
  25441=>"000111111",
  25442=>"110000101",
  25443=>"011001001",
  25444=>"011111100",
  25445=>"011101100",
  25446=>"001011111",
  25447=>"010101010",
  25448=>"011100111",
  25449=>"110101001",
  25450=>"011110001",
  25451=>"010110010",
  25452=>"100110101",
  25453=>"011010110",
  25454=>"010100000",
  25455=>"011100111",
  25456=>"110011001",
  25457=>"010100011",
  25458=>"000101000",
  25459=>"110011001",
  25460=>"001001100",
  25461=>"110100101",
  25462=>"011100100",
  25463=>"100100100",
  25464=>"110110101",
  25465=>"010110100",
  25466=>"001100110",
  25467=>"011001111",
  25468=>"111011101",
  25469=>"100110101",
  25470=>"001110110",
  25471=>"110011011",
  25472=>"110010001",
  25473=>"110010111",
  25474=>"111001000",
  25475=>"011101100",
  25476=>"010001011",
  25477=>"101100000",
  25478=>"101100101",
  25479=>"000101010",
  25480=>"001110000",
  25481=>"100011110",
  25482=>"110010011",
  25483=>"010010010",
  25484=>"000000101",
  25485=>"101110010",
  25486=>"011011101",
  25487=>"100000000",
  25488=>"011001101",
  25489=>"000110011",
  25490=>"011110101",
  25491=>"001111010",
  25492=>"110100010",
  25493=>"001001110",
  25494=>"001101001",
  25495=>"000000100",
  25496=>"001011010",
  25497=>"111000001",
  25498=>"110001100",
  25499=>"100100111",
  25500=>"111110001",
  25501=>"100100100",
  25502=>"001011011",
  25503=>"000000110",
  25504=>"100110100",
  25505=>"101111001",
  25506=>"010011111",
  25507=>"011001011",
  25508=>"111101100",
  25509=>"010010011",
  25510=>"001000111",
  25511=>"110101100",
  25512=>"010011111",
  25513=>"101110111",
  25514=>"110110100",
  25515=>"000101111",
  25516=>"101000010",
  25517=>"011111000",
  25518=>"010010100",
  25519=>"100111101",
  25520=>"111110101",
  25521=>"110011101",
  25522=>"011011001",
  25523=>"110011111",
  25524=>"010001010",
  25525=>"000010010",
  25526=>"001011100",
  25527=>"000001011",
  25528=>"011111110",
  25529=>"000100011",
  25530=>"110000011",
  25531=>"100100011",
  25532=>"111001010",
  25533=>"000011000",
  25534=>"111100111",
  25535=>"101010011",
  25536=>"000111111",
  25537=>"111101110",
  25538=>"101011001",
  25539=>"101011000",
  25540=>"001101010",
  25541=>"001010111",
  25542=>"101111111",
  25543=>"001100100",
  25544=>"000000000",
  25545=>"000100101",
  25546=>"111100001",
  25547=>"001110100",
  25548=>"011010010",
  25549=>"011010000",
  25550=>"001000000",
  25551=>"010001011",
  25552=>"010000010",
  25553=>"101011110",
  25554=>"111110001",
  25555=>"001000011",
  25556=>"010000100",
  25557=>"100110010",
  25558=>"100001010",
  25559=>"111111000",
  25560=>"101111010",
  25561=>"000000001",
  25562=>"010110001",
  25563=>"000001001",
  25564=>"100000100",
  25565=>"111001100",
  25566=>"111110000",
  25567=>"111001001",
  25568=>"111111000",
  25569=>"000001011",
  25570=>"000111111",
  25571=>"001001010",
  25572=>"101101011",
  25573=>"011001010",
  25574=>"010100101",
  25575=>"000000101",
  25576=>"111111101",
  25577=>"011110011",
  25578=>"111000100",
  25579=>"010110101",
  25580=>"010101001",
  25581=>"101010100",
  25582=>"100000111",
  25583=>"010100011",
  25584=>"001111111",
  25585=>"000110111",
  25586=>"000001001",
  25587=>"111010111",
  25588=>"001000001",
  25589=>"110100101",
  25590=>"111100110",
  25591=>"111111100",
  25592=>"110100100",
  25593=>"010011100",
  25594=>"001010010",
  25595=>"000110010",
  25596=>"000000111",
  25597=>"110001100",
  25598=>"010000110",
  25599=>"111001011",
  25600=>"110101001",
  25601=>"110001111",
  25602=>"001001001",
  25603=>"010111101",
  25604=>"110010100",
  25605=>"011011000",
  25606=>"101100010",
  25607=>"010000011",
  25608=>"110101111",
  25609=>"100111000",
  25610=>"001010000",
  25611=>"001010100",
  25612=>"001010011",
  25613=>"010001001",
  25614=>"101110101",
  25615=>"110000011",
  25616=>"010010001",
  25617=>"001100100",
  25618=>"011010000",
  25619=>"001010110",
  25620=>"110100101",
  25621=>"111111011",
  25622=>"001001110",
  25623=>"111001010",
  25624=>"010101101",
  25625=>"011111110",
  25626=>"011100000",
  25627=>"100101101",
  25628=>"110101010",
  25629=>"010010010",
  25630=>"111101010",
  25631=>"010100000",
  25632=>"100011101",
  25633=>"111111111",
  25634=>"111111000",
  25635=>"000001000",
  25636=>"010110000",
  25637=>"010001101",
  25638=>"100100010",
  25639=>"011010111",
  25640=>"000101000",
  25641=>"110010000",
  25642=>"010101001",
  25643=>"111101101",
  25644=>"110100110",
  25645=>"011110101",
  25646=>"001001001",
  25647=>"101100100",
  25648=>"110100110",
  25649=>"000100110",
  25650=>"111111010",
  25651=>"110110010",
  25652=>"100000010",
  25653=>"010000010",
  25654=>"111000101",
  25655=>"110100101",
  25656=>"011001001",
  25657=>"111011110",
  25658=>"000011011",
  25659=>"001110010",
  25660=>"000001100",
  25661=>"000100111",
  25662=>"100101011",
  25663=>"100011010",
  25664=>"010000011",
  25665=>"000011000",
  25666=>"111010001",
  25667=>"000010011",
  25668=>"001110000",
  25669=>"111110000",
  25670=>"100000001",
  25671=>"111010110",
  25672=>"011000000",
  25673=>"011001010",
  25674=>"110111100",
  25675=>"110000010",
  25676=>"111001101",
  25677=>"111110010",
  25678=>"100110010",
  25679=>"011100000",
  25680=>"001011110",
  25681=>"101101001",
  25682=>"011000011",
  25683=>"100011011",
  25684=>"111001000",
  25685=>"100011011",
  25686=>"101110011",
  25687=>"100100001",
  25688=>"100111111",
  25689=>"111011110",
  25690=>"100100010",
  25691=>"110010100",
  25692=>"011101000",
  25693=>"101000010",
  25694=>"111001101",
  25695=>"001011011",
  25696=>"110000101",
  25697=>"010001010",
  25698=>"011111110",
  25699=>"010010111",
  25700=>"110011000",
  25701=>"011000001",
  25702=>"001111011",
  25703=>"111000010",
  25704=>"010011100",
  25705=>"010011100",
  25706=>"110010100",
  25707=>"000000110",
  25708=>"100101000",
  25709=>"010001001",
  25710=>"111100100",
  25711=>"101010010",
  25712=>"011100011",
  25713=>"001101111",
  25714=>"111100001",
  25715=>"011110011",
  25716=>"101000100",
  25717=>"011110101",
  25718=>"000101111",
  25719=>"100110000",
  25720=>"111101101",
  25721=>"000101101",
  25722=>"111011101",
  25723=>"111011101",
  25724=>"111001110",
  25725=>"010110111",
  25726=>"000011000",
  25727=>"100010000",
  25728=>"010000101",
  25729=>"110101101",
  25730=>"101101011",
  25731=>"001111110",
  25732=>"111101100",
  25733=>"011000100",
  25734=>"110110000",
  25735=>"001100011",
  25736=>"111100000",
  25737=>"000101110",
  25738=>"001110100",
  25739=>"101111101",
  25740=>"100111111",
  25741=>"001000111",
  25742=>"000001010",
  25743=>"110101110",
  25744=>"001011010",
  25745=>"111010100",
  25746=>"000101011",
  25747=>"111011101",
  25748=>"101101111",
  25749=>"001010011",
  25750=>"100111010",
  25751=>"110111111",
  25752=>"000001011",
  25753=>"001111111",
  25754=>"110100000",
  25755=>"000100001",
  25756=>"000010101",
  25757=>"000111000",
  25758=>"100110110",
  25759=>"001000001",
  25760=>"010010101",
  25761=>"001001110",
  25762=>"011000111",
  25763=>"011111111",
  25764=>"100000010",
  25765=>"001010001",
  25766=>"101101110",
  25767=>"010001010",
  25768=>"001110010",
  25769=>"100010100",
  25770=>"111001000",
  25771=>"000011000",
  25772=>"110101000",
  25773=>"101111010",
  25774=>"001101011",
  25775=>"011110100",
  25776=>"100001100",
  25777=>"110100011",
  25778=>"000100011",
  25779=>"011101000",
  25780=>"101001001",
  25781=>"111111111",
  25782=>"110001100",
  25783=>"101110101",
  25784=>"000001100",
  25785=>"001001110",
  25786=>"100010110",
  25787=>"100001001",
  25788=>"000101111",
  25789=>"000100010",
  25790=>"010001010",
  25791=>"101100100",
  25792=>"000010011",
  25793=>"100000000",
  25794=>"110110001",
  25795=>"101011101",
  25796=>"100100111",
  25797=>"001111001",
  25798=>"001100100",
  25799=>"100010000",
  25800=>"100011010",
  25801=>"100101101",
  25802=>"101011010",
  25803=>"110010000",
  25804=>"000010111",
  25805=>"110110110",
  25806=>"011101111",
  25807=>"111011001",
  25808=>"110010001",
  25809=>"100110000",
  25810=>"000001001",
  25811=>"110101001",
  25812=>"011100001",
  25813=>"010110110",
  25814=>"110111111",
  25815=>"000111100",
  25816=>"000000100",
  25817=>"101001111",
  25818=>"110011110",
  25819=>"100101100",
  25820=>"101101100",
  25821=>"011000110",
  25822=>"000111011",
  25823=>"100001111",
  25824=>"110110010",
  25825=>"110011111",
  25826=>"000010010",
  25827=>"010100011",
  25828=>"011101011",
  25829=>"001101111",
  25830=>"000101000",
  25831=>"000111010",
  25832=>"011101111",
  25833=>"110000010",
  25834=>"010001010",
  25835=>"100101000",
  25836=>"010111111",
  25837=>"101010000",
  25838=>"010000111",
  25839=>"010000001",
  25840=>"001001110",
  25841=>"001100111",
  25842=>"001011001",
  25843=>"010100011",
  25844=>"000011010",
  25845=>"111111110",
  25846=>"010001101",
  25847=>"111000111",
  25848=>"101111111",
  25849=>"100111110",
  25850=>"000101010",
  25851=>"110000110",
  25852=>"111101100",
  25853=>"100010110",
  25854=>"001011011",
  25855=>"011010100",
  25856=>"111110110",
  25857=>"000101100",
  25858=>"100111000",
  25859=>"000110010",
  25860=>"101111010",
  25861=>"110111111",
  25862=>"011001101",
  25863=>"010000001",
  25864=>"011010101",
  25865=>"000100111",
  25866=>"110011000",
  25867=>"010110110",
  25868=>"100010100",
  25869=>"001000010",
  25870=>"001101111",
  25871=>"001011101",
  25872=>"101110101",
  25873=>"000001011",
  25874=>"111010000",
  25875=>"000101101",
  25876=>"101101000",
  25877=>"100110100",
  25878=>"110011010",
  25879=>"000100111",
  25880=>"010111010",
  25881=>"001000000",
  25882=>"011010110",
  25883=>"000110001",
  25884=>"011110001",
  25885=>"010011001",
  25886=>"110100011",
  25887=>"110001111",
  25888=>"010100110",
  25889=>"110110010",
  25890=>"110011100",
  25891=>"001001111",
  25892=>"010000001",
  25893=>"100101111",
  25894=>"001101001",
  25895=>"111101100",
  25896=>"010001100",
  25897=>"011011101",
  25898=>"111111101",
  25899=>"000001110",
  25900=>"111110111",
  25901=>"011111010",
  25902=>"000001000",
  25903=>"000000110",
  25904=>"100000100",
  25905=>"011110001",
  25906=>"100010101",
  25907=>"011010100",
  25908=>"101100000",
  25909=>"101001000",
  25910=>"010010100",
  25911=>"101001000",
  25912=>"110000010",
  25913=>"101111011",
  25914=>"111111101",
  25915=>"000000111",
  25916=>"001111100",
  25917=>"111000101",
  25918=>"011000001",
  25919=>"110000001",
  25920=>"100011010",
  25921=>"000001000",
  25922=>"101111111",
  25923=>"010010011",
  25924=>"011010111",
  25925=>"101111010",
  25926=>"101100101",
  25927=>"110010011",
  25928=>"000011001",
  25929=>"110000111",
  25930=>"101010101",
  25931=>"001110011",
  25932=>"000001001",
  25933=>"000001110",
  25934=>"111111110",
  25935=>"100110110",
  25936=>"011011101",
  25937=>"001111011",
  25938=>"100011000",
  25939=>"011011101",
  25940=>"010110100",
  25941=>"111010110",
  25942=>"011110110",
  25943=>"110011010",
  25944=>"000111000",
  25945=>"011001010",
  25946=>"110011010",
  25947=>"000011001",
  25948=>"110100110",
  25949=>"110001111",
  25950=>"001101100",
  25951=>"001100000",
  25952=>"010100010",
  25953=>"011111110",
  25954=>"001101111",
  25955=>"000110101",
  25956=>"000001000",
  25957=>"000011101",
  25958=>"001001000",
  25959=>"001001100",
  25960=>"111011010",
  25961=>"011111110",
  25962=>"000110100",
  25963=>"011100110",
  25964=>"000101111",
  25965=>"111101001",
  25966=>"001101000",
  25967=>"010100000",
  25968=>"011101010",
  25969=>"100000001",
  25970=>"011001001",
  25971=>"011011101",
  25972=>"101101110",
  25973=>"000100110",
  25974=>"010000110",
  25975=>"000011110",
  25976=>"100100000",
  25977=>"111101100",
  25978=>"100011101",
  25979=>"000111110",
  25980=>"110010110",
  25981=>"111111011",
  25982=>"000010000",
  25983=>"001011010",
  25984=>"011000000",
  25985=>"100011101",
  25986=>"110110111",
  25987=>"001111000",
  25988=>"110000110",
  25989=>"110010001",
  25990=>"001010001",
  25991=>"110011000",
  25992=>"001010010",
  25993=>"111111100",
  25994=>"100100100",
  25995=>"100110101",
  25996=>"111010001",
  25997=>"001110011",
  25998=>"110010010",
  25999=>"100100000",
  26000=>"111101111",
  26001=>"100100111",
  26002=>"100101111",
  26003=>"000011001",
  26004=>"100111110",
  26005=>"011111101",
  26006=>"011101101",
  26007=>"111001011",
  26008=>"000011011",
  26009=>"100001001",
  26010=>"000011110",
  26011=>"010011101",
  26012=>"100000111",
  26013=>"001001010",
  26014=>"001001101",
  26015=>"011000010",
  26016=>"110010010",
  26017=>"011010000",
  26018=>"000010011",
  26019=>"000010100",
  26020=>"000001001",
  26021=>"000100010",
  26022=>"010100010",
  26023=>"100101010",
  26024=>"110101111",
  26025=>"000000010",
  26026=>"111100000",
  26027=>"000100000",
  26028=>"111001111",
  26029=>"011100001",
  26030=>"100101001",
  26031=>"101011100",
  26032=>"001001110",
  26033=>"000011001",
  26034=>"011000100",
  26035=>"110100101",
  26036=>"100110011",
  26037=>"100101100",
  26038=>"101111010",
  26039=>"101010001",
  26040=>"110100110",
  26041=>"101101011",
  26042=>"001000101",
  26043=>"001000001",
  26044=>"101010010",
  26045=>"010100000",
  26046=>"110001110",
  26047=>"010010000",
  26048=>"001001011",
  26049=>"100101000",
  26050=>"100010000",
  26051=>"100110111",
  26052=>"111001001",
  26053=>"001000101",
  26054=>"011001001",
  26055=>"110011000",
  26056=>"110010000",
  26057=>"000000100",
  26058=>"111001010",
  26059=>"010101001",
  26060=>"010100001",
  26061=>"111111111",
  26062=>"100110000",
  26063=>"010000110",
  26064=>"100110111",
  26065=>"000011111",
  26066=>"100101011",
  26067=>"101101110",
  26068=>"111110111",
  26069=>"001001110",
  26070=>"000010000",
  26071=>"100011011",
  26072=>"000011111",
  26073=>"111110101",
  26074=>"001110000",
  26075=>"000001111",
  26076=>"111001001",
  26077=>"000100100",
  26078=>"101101000",
  26079=>"011100110",
  26080=>"110010101",
  26081=>"001110011",
  26082=>"001001110",
  26083=>"111001010",
  26084=>"100000000",
  26085=>"100000010",
  26086=>"000101000",
  26087=>"010011000",
  26088=>"010111000",
  26089=>"010110100",
  26090=>"111000011",
  26091=>"101100011",
  26092=>"111101010",
  26093=>"010001000",
  26094=>"110000001",
  26095=>"101000010",
  26096=>"110100101",
  26097=>"111011001",
  26098=>"100110100",
  26099=>"101010111",
  26100=>"101001000",
  26101=>"100001000",
  26102=>"111011111",
  26103=>"100001000",
  26104=>"010000010",
  26105=>"101011000",
  26106=>"110011100",
  26107=>"101000111",
  26108=>"111011001",
  26109=>"110110011",
  26110=>"101101100",
  26111=>"111101001",
  26112=>"010001000",
  26113=>"000001001",
  26114=>"111011011",
  26115=>"000110110",
  26116=>"100010000",
  26117=>"101100100",
  26118=>"000000001",
  26119=>"101100001",
  26120=>"101001000",
  26121=>"111001100",
  26122=>"111011001",
  26123=>"010001111",
  26124=>"110101011",
  26125=>"100010101",
  26126=>"100101001",
  26127=>"100100100",
  26128=>"101100100",
  26129=>"100100111",
  26130=>"111000000",
  26131=>"100111101",
  26132=>"000001011",
  26133=>"111010010",
  26134=>"000100000",
  26135=>"111111010",
  26136=>"000111110",
  26137=>"110100001",
  26138=>"101100000",
  26139=>"000100100",
  26140=>"111101110",
  26141=>"110000111",
  26142=>"001010101",
  26143=>"000011011",
  26144=>"110000000",
  26145=>"111001011",
  26146=>"010100000",
  26147=>"101111011",
  26148=>"110110100",
  26149=>"001110110",
  26150=>"010011000",
  26151=>"110000011",
  26152=>"001110011",
  26153=>"111010100",
  26154=>"000101110",
  26155=>"101010000",
  26156=>"101110100",
  26157=>"110110010",
  26158=>"010000011",
  26159=>"000010011",
  26160=>"000011000",
  26161=>"010101101",
  26162=>"101110100",
  26163=>"011011001",
  26164=>"110000110",
  26165=>"000001011",
  26166=>"011010111",
  26167=>"110110100",
  26168=>"011100100",
  26169=>"110011110",
  26170=>"000101011",
  26171=>"001000010",
  26172=>"111100111",
  26173=>"110111110",
  26174=>"111000000",
  26175=>"000100011",
  26176=>"111101101",
  26177=>"100100010",
  26178=>"011000000",
  26179=>"110111100",
  26180=>"000100010",
  26181=>"101011111",
  26182=>"100001101",
  26183=>"010000000",
  26184=>"110001000",
  26185=>"101111110",
  26186=>"000100010",
  26187=>"011100010",
  26188=>"111111111",
  26189=>"010100011",
  26190=>"011000011",
  26191=>"000000010",
  26192=>"000111011",
  26193=>"110010001",
  26194=>"111001010",
  26195=>"110001010",
  26196=>"110001100",
  26197=>"101101110",
  26198=>"100100000",
  26199=>"000011011",
  26200=>"100011011",
  26201=>"010000010",
  26202=>"110110110",
  26203=>"001000100",
  26204=>"101001011",
  26205=>"011000111",
  26206=>"010100111",
  26207=>"101011100",
  26208=>"101000111",
  26209=>"001001001",
  26210=>"110001101",
  26211=>"100111100",
  26212=>"011100101",
  26213=>"001000001",
  26214=>"100001100",
  26215=>"001000011",
  26216=>"111011111",
  26217=>"000101001",
  26218=>"110001011",
  26219=>"100110110",
  26220=>"010010010",
  26221=>"001010000",
  26222=>"010100010",
  26223=>"101101101",
  26224=>"111010110",
  26225=>"111010010",
  26226=>"010000010",
  26227=>"001000000",
  26228=>"000110000",
  26229=>"101011110",
  26230=>"111111111",
  26231=>"110000010",
  26232=>"000010100",
  26233=>"111101110",
  26234=>"000001011",
  26235=>"010010100",
  26236=>"000101110",
  26237=>"000110011",
  26238=>"011001011",
  26239=>"111101010",
  26240=>"100010000",
  26241=>"101001001",
  26242=>"110000100",
  26243=>"001000000",
  26244=>"010101010",
  26245=>"100001100",
  26246=>"101111100",
  26247=>"111111101",
  26248=>"100000111",
  26249=>"000000010",
  26250=>"110101000",
  26251=>"100110000",
  26252=>"100000000",
  26253=>"100010110",
  26254=>"001101100",
  26255=>"100111101",
  26256=>"010100011",
  26257=>"000110011",
  26258=>"001101111",
  26259=>"010101101",
  26260=>"000100101",
  26261=>"101010100",
  26262=>"100100000",
  26263=>"100101100",
  26264=>"111110000",
  26265=>"000011010",
  26266=>"110011100",
  26267=>"001101010",
  26268=>"100100010",
  26269=>"110100101",
  26270=>"010100000",
  26271=>"100000111",
  26272=>"001110010",
  26273=>"001011000",
  26274=>"110111111",
  26275=>"011101011",
  26276=>"101000011",
  26277=>"000010111",
  26278=>"001110000",
  26279=>"010110101",
  26280=>"101011111",
  26281=>"110110011",
  26282=>"010000000",
  26283=>"111100011",
  26284=>"110011101",
  26285=>"110100110",
  26286=>"010111010",
  26287=>"110011101",
  26288=>"110000000",
  26289=>"111110010",
  26290=>"000010001",
  26291=>"100011011",
  26292=>"011111010",
  26293=>"110011001",
  26294=>"011000000",
  26295=>"000010000",
  26296=>"001011111",
  26297=>"000110110",
  26298=>"000001111",
  26299=>"010100010",
  26300=>"000110011",
  26301=>"001110101",
  26302=>"000001010",
  26303=>"110111100",
  26304=>"001010101",
  26305=>"010110010",
  26306=>"100011010",
  26307=>"000011010",
  26308=>"011010010",
  26309=>"010100000",
  26310=>"000011100",
  26311=>"000011001",
  26312=>"010100100",
  26313=>"101011011",
  26314=>"101010000",
  26315=>"100110010",
  26316=>"011101101",
  26317=>"000001000",
  26318=>"111110101",
  26319=>"100000010",
  26320=>"111010011",
  26321=>"110001100",
  26322=>"010111110",
  26323=>"100111000",
  26324=>"010011010",
  26325=>"000100101",
  26326=>"010001001",
  26327=>"001110111",
  26328=>"110111010",
  26329=>"000011000",
  26330=>"111001110",
  26331=>"110010101",
  26332=>"001001011",
  26333=>"111110110",
  26334=>"000111100",
  26335=>"110111110",
  26336=>"001110100",
  26337=>"101010011",
  26338=>"000001100",
  26339=>"011001001",
  26340=>"110100000",
  26341=>"111110101",
  26342=>"111010101",
  26343=>"111111100",
  26344=>"011010100",
  26345=>"111010010",
  26346=>"110010001",
  26347=>"111110010",
  26348=>"110111000",
  26349=>"000001100",
  26350=>"001101000",
  26351=>"010110101",
  26352=>"000010000",
  26353=>"001110101",
  26354=>"001001101",
  26355=>"111111010",
  26356=>"011110011",
  26357=>"101001011",
  26358=>"110101110",
  26359=>"111010110",
  26360=>"001111000",
  26361=>"101111100",
  26362=>"110011101",
  26363=>"000001110",
  26364=>"111101001",
  26365=>"111111111",
  26366=>"010000111",
  26367=>"011001100",
  26368=>"110000011",
  26369=>"101111001",
  26370=>"011111000",
  26371=>"000110110",
  26372=>"111110111",
  26373=>"011000010",
  26374=>"000011110",
  26375=>"100101101",
  26376=>"110100100",
  26377=>"100101011",
  26378=>"101010010",
  26379=>"000101010",
  26380=>"010110011",
  26381=>"110110110",
  26382=>"110011011",
  26383=>"011010000",
  26384=>"101011010",
  26385=>"000000000",
  26386=>"001000100",
  26387=>"000111101",
  26388=>"000110101",
  26389=>"110100101",
  26390=>"001000101",
  26391=>"011000111",
  26392=>"000100101",
  26393=>"001100011",
  26394=>"001001001",
  26395=>"010001110",
  26396=>"111011001",
  26397=>"011110001",
  26398=>"001000010",
  26399=>"011000111",
  26400=>"100000011",
  26401=>"100001100",
  26402=>"101001111",
  26403=>"010001111",
  26404=>"000001000",
  26405=>"111111101",
  26406=>"100000101",
  26407=>"110001011",
  26408=>"001011110",
  26409=>"010000101",
  26410=>"110000110",
  26411=>"001000000",
  26412=>"100001100",
  26413=>"000011110",
  26414=>"111111110",
  26415=>"110000010",
  26416=>"110100101",
  26417=>"010010100",
  26418=>"101001100",
  26419=>"000001101",
  26420=>"010110111",
  26421=>"110010011",
  26422=>"101110101",
  26423=>"010001010",
  26424=>"000101001",
  26425=>"110000000",
  26426=>"000110100",
  26427=>"111011111",
  26428=>"010101001",
  26429=>"000110010",
  26430=>"000101000",
  26431=>"100110111",
  26432=>"111110110",
  26433=>"011101100",
  26434=>"010011000",
  26435=>"011110110",
  26436=>"001111001",
  26437=>"011000111",
  26438=>"110000100",
  26439=>"111101010",
  26440=>"110100111",
  26441=>"001000001",
  26442=>"101101010",
  26443=>"011011110",
  26444=>"100010010",
  26445=>"010000000",
  26446=>"100000100",
  26447=>"101000010",
  26448=>"011011110",
  26449=>"010011111",
  26450=>"010001010",
  26451=>"101100110",
  26452=>"011100000",
  26453=>"111110010",
  26454=>"100010101",
  26455=>"011000011",
  26456=>"111111100",
  26457=>"101101101",
  26458=>"101101011",
  26459=>"001000001",
  26460=>"111100111",
  26461=>"101000001",
  26462=>"000111011",
  26463=>"001000011",
  26464=>"110001010",
  26465=>"000000110",
  26466=>"101001011",
  26467=>"100011010",
  26468=>"011000110",
  26469=>"000000011",
  26470=>"101010011",
  26471=>"101001010",
  26472=>"001001000",
  26473=>"100100000",
  26474=>"101000110",
  26475=>"111001000",
  26476=>"011000000",
  26477=>"110100000",
  26478=>"100011111",
  26479=>"111100001",
  26480=>"011110010",
  26481=>"011110110",
  26482=>"111001111",
  26483=>"010100111",
  26484=>"110000011",
  26485=>"000001101",
  26486=>"101001001",
  26487=>"110010100",
  26488=>"100101100",
  26489=>"000010100",
  26490=>"010100111",
  26491=>"011110110",
  26492=>"000001101",
  26493=>"110100101",
  26494=>"010011010",
  26495=>"000001011",
  26496=>"010010110",
  26497=>"000010010",
  26498=>"010010101",
  26499=>"111010000",
  26500=>"100011011",
  26501=>"100100110",
  26502=>"010100101",
  26503=>"110111110",
  26504=>"101011100",
  26505=>"111000001",
  26506=>"011011101",
  26507=>"011000101",
  26508=>"100001110",
  26509=>"100000000",
  26510=>"110010001",
  26511=>"001111000",
  26512=>"111001010",
  26513=>"010100010",
  26514=>"010010110",
  26515=>"100100100",
  26516=>"110100001",
  26517=>"000110100",
  26518=>"010010000",
  26519=>"000111000",
  26520=>"011110000",
  26521=>"000000001",
  26522=>"100010001",
  26523=>"010111011",
  26524=>"010001110",
  26525=>"110010110",
  26526=>"001110011",
  26527=>"100110110",
  26528=>"100111000",
  26529=>"100001101",
  26530=>"000101001",
  26531=>"010000101",
  26532=>"000000010",
  26533=>"011101100",
  26534=>"110100111",
  26535=>"110011011",
  26536=>"110001101",
  26537=>"110010010",
  26538=>"110111110",
  26539=>"111001010",
  26540=>"100100000",
  26541=>"111100111",
  26542=>"111000000",
  26543=>"011010001",
  26544=>"101011001",
  26545=>"001100111",
  26546=>"011100000",
  26547=>"110001011",
  26548=>"100001101",
  26549=>"101001111",
  26550=>"001011100",
  26551=>"101010101",
  26552=>"001010110",
  26553=>"010110000",
  26554=>"010001001",
  26555=>"111001001",
  26556=>"110111111",
  26557=>"001111111",
  26558=>"000001011",
  26559=>"010111001",
  26560=>"110100000",
  26561=>"110111010",
  26562=>"101111110",
  26563=>"010010100",
  26564=>"011011101",
  26565=>"001100100",
  26566=>"011011110",
  26567=>"111110100",
  26568=>"010000011",
  26569=>"101100010",
  26570=>"100001001",
  26571=>"011000011",
  26572=>"010101000",
  26573=>"100101111",
  26574=>"111001110",
  26575=>"101001000",
  26576=>"100000011",
  26577=>"110010000",
  26578=>"000000101",
  26579=>"111000000",
  26580=>"110000101",
  26581=>"111001100",
  26582=>"001001000",
  26583=>"010111111",
  26584=>"110000011",
  26585=>"110111101",
  26586=>"100010011",
  26587=>"010110101",
  26588=>"110000000",
  26589=>"100110010",
  26590=>"010001010",
  26591=>"000010010",
  26592=>"101010111",
  26593=>"111001111",
  26594=>"111100001",
  26595=>"111010001",
  26596=>"011000111",
  26597=>"000000011",
  26598=>"000010101",
  26599=>"101111110",
  26600=>"110001100",
  26601=>"101101101",
  26602=>"111000001",
  26603=>"101100010",
  26604=>"011111101",
  26605=>"111000000",
  26606=>"011001100",
  26607=>"110111010",
  26608=>"000010000",
  26609=>"101011010",
  26610=>"011100100",
  26611=>"011010100",
  26612=>"110000010",
  26613=>"000000011",
  26614=>"110101111",
  26615=>"000001000",
  26616=>"100010001",
  26617=>"111110111",
  26618=>"100001000",
  26619=>"011101011",
  26620=>"100000100",
  26621=>"001110000",
  26622=>"010100111",
  26623=>"010000011",
  26624=>"100100000",
  26625=>"111000110",
  26626=>"110100011",
  26627=>"110100101",
  26628=>"111010111",
  26629=>"001100000",
  26630=>"101110000",
  26631=>"011011111",
  26632=>"010111010",
  26633=>"010101100",
  26634=>"100000011",
  26635=>"110000010",
  26636=>"001001010",
  26637=>"110100010",
  26638=>"010111011",
  26639=>"001101000",
  26640=>"111100011",
  26641=>"101001010",
  26642=>"010010100",
  26643=>"101101101",
  26644=>"101101101",
  26645=>"001110010",
  26646=>"010101110",
  26647=>"001101110",
  26648=>"011100001",
  26649=>"100110010",
  26650=>"001000100",
  26651=>"110111110",
  26652=>"100010111",
  26653=>"110110101",
  26654=>"010111111",
  26655=>"011000110",
  26656=>"101111011",
  26657=>"101011010",
  26658=>"011101110",
  26659=>"101110100",
  26660=>"101000101",
  26661=>"011100001",
  26662=>"110100101",
  26663=>"100111111",
  26664=>"110110000",
  26665=>"111100101",
  26666=>"110000000",
  26667=>"111111001",
  26668=>"010111001",
  26669=>"110001111",
  26670=>"011110110",
  26671=>"011100110",
  26672=>"111010001",
  26673=>"001111000",
  26674=>"110111000",
  26675=>"110100000",
  26676=>"111100011",
  26677=>"101101110",
  26678=>"000000000",
  26679=>"111011001",
  26680=>"111010010",
  26681=>"111101110",
  26682=>"001000011",
  26683=>"110100100",
  26684=>"000010000",
  26685=>"000101110",
  26686=>"111111100",
  26687=>"111000111",
  26688=>"100011010",
  26689=>"100001111",
  26690=>"011100111",
  26691=>"100101111",
  26692=>"110110111",
  26693=>"100011000",
  26694=>"100110100",
  26695=>"001010001",
  26696=>"101111110",
  26697=>"101011001",
  26698=>"111110111",
  26699=>"000000111",
  26700=>"011101111",
  26701=>"011001000",
  26702=>"010010010",
  26703=>"000011011",
  26704=>"011100111",
  26705=>"000011001",
  26706=>"111000010",
  26707=>"100101000",
  26708=>"111111110",
  26709=>"101111010",
  26710=>"001111110",
  26711=>"100110111",
  26712=>"001111001",
  26713=>"011011011",
  26714=>"010000100",
  26715=>"011100110",
  26716=>"101111111",
  26717=>"111110111",
  26718=>"000110110",
  26719=>"100011101",
  26720=>"000010100",
  26721=>"001110100",
  26722=>"111010010",
  26723=>"100101000",
  26724=>"000000001",
  26725=>"000111101",
  26726=>"110111010",
  26727=>"101000111",
  26728=>"101101101",
  26729=>"110011100",
  26730=>"111111000",
  26731=>"100000111",
  26732=>"101101101",
  26733=>"001111101",
  26734=>"110101101",
  26735=>"000100111",
  26736=>"000110101",
  26737=>"100111101",
  26738=>"000000011",
  26739=>"110011011",
  26740=>"110101100",
  26741=>"000011011",
  26742=>"011110000",
  26743=>"100111001",
  26744=>"100100000",
  26745=>"111111111",
  26746=>"011011001",
  26747=>"100100000",
  26748=>"101100110",
  26749=>"001101011",
  26750=>"011110011",
  26751=>"111110110",
  26752=>"010101110",
  26753=>"101001001",
  26754=>"101101010",
  26755=>"000000100",
  26756=>"110110111",
  26757=>"111001111",
  26758=>"011011110",
  26759=>"011111110",
  26760=>"101010101",
  26761=>"100101010",
  26762=>"010011000",
  26763=>"111110111",
  26764=>"101001000",
  26765=>"010111100",
  26766=>"001100001",
  26767=>"001000010",
  26768=>"011001001",
  26769=>"000001111",
  26770=>"001010101",
  26771=>"000100000",
  26772=>"001101100",
  26773=>"000011111",
  26774=>"001101010",
  26775=>"011011100",
  26776=>"101101010",
  26777=>"101010010",
  26778=>"010011000",
  26779=>"001011111",
  26780=>"110111100",
  26781=>"100000000",
  26782=>"010000000",
  26783=>"001101100",
  26784=>"010100011",
  26785=>"001000110",
  26786=>"001011111",
  26787=>"000110011",
  26788=>"000100011",
  26789=>"110011000",
  26790=>"011100000",
  26791=>"011010000",
  26792=>"111010101",
  26793=>"010111001",
  26794=>"110111110",
  26795=>"100000010",
  26796=>"111010111",
  26797=>"000011011",
  26798=>"111111011",
  26799=>"100011101",
  26800=>"100100000",
  26801=>"100110111",
  26802=>"001011101",
  26803=>"111011111",
  26804=>"010110100",
  26805=>"100000010",
  26806=>"110101111",
  26807=>"000001010",
  26808=>"110100100",
  26809=>"111111111",
  26810=>"010110110",
  26811=>"100111010",
  26812=>"110100101",
  26813=>"111000010",
  26814=>"010100100",
  26815=>"110010110",
  26816=>"101110010",
  26817=>"110100011",
  26818=>"110111110",
  26819=>"001010100",
  26820=>"001101001",
  26821=>"111111110",
  26822=>"011001011",
  26823=>"110101110",
  26824=>"000111110",
  26825=>"001000100",
  26826=>"110101111",
  26827=>"101111100",
  26828=>"010111100",
  26829=>"000011000",
  26830=>"000010001",
  26831=>"110100110",
  26832=>"110100100",
  26833=>"111000101",
  26834=>"101101011",
  26835=>"011101101",
  26836=>"000001000",
  26837=>"010011001",
  26838=>"011111100",
  26839=>"100000111",
  26840=>"101111010",
  26841=>"111110010",
  26842=>"011011100",
  26843=>"110010001",
  26844=>"110000100",
  26845=>"011011100",
  26846=>"110100110",
  26847=>"001010101",
  26848=>"001111110",
  26849=>"010011010",
  26850=>"111111111",
  26851=>"111011100",
  26852=>"001001011",
  26853=>"001000100",
  26854=>"110001000",
  26855=>"001011100",
  26856=>"111111011",
  26857=>"111111111",
  26858=>"100011110",
  26859=>"010111001",
  26860=>"100010001",
  26861=>"001100100",
  26862=>"110101010",
  26863=>"100111111",
  26864=>"000101111",
  26865=>"110001001",
  26866=>"101001111",
  26867=>"010110011",
  26868=>"101110111",
  26869=>"010010100",
  26870=>"110001000",
  26871=>"101001111",
  26872=>"000010001",
  26873=>"000111101",
  26874=>"001100100",
  26875=>"101110110",
  26876=>"111101101",
  26877=>"001010010",
  26878=>"001101110",
  26879=>"011101111",
  26880=>"110000011",
  26881=>"000111001",
  26882=>"100001001",
  26883=>"101111101",
  26884=>"101010000",
  26885=>"110111111",
  26886=>"110110100",
  26887=>"001010101",
  26888=>"010011100",
  26889=>"110001011",
  26890=>"000100100",
  26891=>"010000110",
  26892=>"111000000",
  26893=>"000110110",
  26894=>"001011100",
  26895=>"001001101",
  26896=>"011010010",
  26897=>"111001111",
  26898=>"101100100",
  26899=>"101001011",
  26900=>"011001011",
  26901=>"111101100",
  26902=>"111001101",
  26903=>"110010001",
  26904=>"100001011",
  26905=>"100101000",
  26906=>"100010110",
  26907=>"100001100",
  26908=>"000000000",
  26909=>"011101011",
  26910=>"010011101",
  26911=>"111100110",
  26912=>"001111000",
  26913=>"000111000",
  26914=>"110000000",
  26915=>"110110111",
  26916=>"011010111",
  26917=>"011001111",
  26918=>"001111101",
  26919=>"101010000",
  26920=>"011110101",
  26921=>"001101011",
  26922=>"100111110",
  26923=>"000001101",
  26924=>"011000000",
  26925=>"010010001",
  26926=>"111101111",
  26927=>"110001000",
  26928=>"011110101",
  26929=>"101101011",
  26930=>"111111011",
  26931=>"011001110",
  26932=>"000001010",
  26933=>"010111011",
  26934=>"110010001",
  26935=>"100001101",
  26936=>"101111111",
  26937=>"111010100",
  26938=>"000101111",
  26939=>"100101101",
  26940=>"000100011",
  26941=>"000100001",
  26942=>"000100010",
  26943=>"101000000",
  26944=>"001000000",
  26945=>"100001100",
  26946=>"011100111",
  26947=>"101010000",
  26948=>"000100011",
  26949=>"000010000",
  26950=>"000000000",
  26951=>"100110101",
  26952=>"111010101",
  26953=>"100110111",
  26954=>"111110010",
  26955=>"100110001",
  26956=>"011010001",
  26957=>"111011010",
  26958=>"111101010",
  26959=>"101111110",
  26960=>"101111000",
  26961=>"111111100",
  26962=>"010000110",
  26963=>"001111011",
  26964=>"100100111",
  26965=>"100100110",
  26966=>"000010110",
  26967=>"111100000",
  26968=>"010000011",
  26969=>"111111110",
  26970=>"001101101",
  26971=>"101011110",
  26972=>"011100111",
  26973=>"110001000",
  26974=>"110111110",
  26975=>"111111001",
  26976=>"111011100",
  26977=>"100000011",
  26978=>"101110000",
  26979=>"101111101",
  26980=>"111100110",
  26981=>"100100000",
  26982=>"000100000",
  26983=>"111110101",
  26984=>"001101111",
  26985=>"101100000",
  26986=>"110000111",
  26987=>"111111011",
  26988=>"110110111",
  26989=>"100011011",
  26990=>"001101000",
  26991=>"000101001",
  26992=>"001011000",
  26993=>"000011110",
  26994=>"100001001",
  26995=>"000010110",
  26996=>"100001000",
  26997=>"010001011",
  26998=>"111100111",
  26999=>"101011010",
  27000=>"101000110",
  27001=>"001111111",
  27002=>"010111010",
  27003=>"010111000",
  27004=>"111010010",
  27005=>"011010001",
  27006=>"001000101",
  27007=>"111100100",
  27008=>"100100111",
  27009=>"001111100",
  27010=>"011100001",
  27011=>"111010101",
  27012=>"101100000",
  27013=>"010110011",
  27014=>"011011000",
  27015=>"011001101",
  27016=>"101111011",
  27017=>"001011110",
  27018=>"101100000",
  27019=>"011000101",
  27020=>"100111110",
  27021=>"110000101",
  27022=>"011111110",
  27023=>"110001100",
  27024=>"011111101",
  27025=>"010101001",
  27026=>"110000110",
  27027=>"001010101",
  27028=>"111001010",
  27029=>"010111000",
  27030=>"000100010",
  27031=>"110100010",
  27032=>"100010001",
  27033=>"011101110",
  27034=>"000001110",
  27035=>"110010010",
  27036=>"100100000",
  27037=>"011010000",
  27038=>"111111100",
  27039=>"010000111",
  27040=>"101000100",
  27041=>"001010010",
  27042=>"101011000",
  27043=>"101001101",
  27044=>"000100000",
  27045=>"101001101",
  27046=>"101111011",
  27047=>"110110010",
  27048=>"010011110",
  27049=>"100010010",
  27050=>"111110000",
  27051=>"000111011",
  27052=>"111010010",
  27053=>"111110111",
  27054=>"011001100",
  27055=>"010000101",
  27056=>"000100010",
  27057=>"110011101",
  27058=>"110101000",
  27059=>"010100000",
  27060=>"111100101",
  27061=>"101111011",
  27062=>"111011110",
  27063=>"010100100",
  27064=>"101110111",
  27065=>"111110010",
  27066=>"111111010",
  27067=>"100001101",
  27068=>"010110001",
  27069=>"110001101",
  27070=>"011100100",
  27071=>"101000000",
  27072=>"110010010",
  27073=>"011011101",
  27074=>"100010101",
  27075=>"011000110",
  27076=>"101000110",
  27077=>"011000110",
  27078=>"000100000",
  27079=>"000110101",
  27080=>"100001010",
  27081=>"111110111",
  27082=>"000111100",
  27083=>"101001010",
  27084=>"010101111",
  27085=>"110111100",
  27086=>"110011100",
  27087=>"010111110",
  27088=>"101010001",
  27089=>"001011110",
  27090=>"010100110",
  27091=>"010000010",
  27092=>"001010010",
  27093=>"010011010",
  27094=>"001111101",
  27095=>"111101111",
  27096=>"011011001",
  27097=>"100110101",
  27098=>"001010011",
  27099=>"001101000",
  27100=>"111101111",
  27101=>"101011010",
  27102=>"001110101",
  27103=>"100101010",
  27104=>"001110010",
  27105=>"011000001",
  27106=>"001111111",
  27107=>"100101100",
  27108=>"010010101",
  27109=>"010110010",
  27110=>"010000100",
  27111=>"001100100",
  27112=>"000101101",
  27113=>"111110101",
  27114=>"010000010",
  27115=>"011010101",
  27116=>"111000110",
  27117=>"010100110",
  27118=>"110001111",
  27119=>"011100110",
  27120=>"100100010",
  27121=>"011011010",
  27122=>"011010101",
  27123=>"110100010",
  27124=>"010000011",
  27125=>"001010010",
  27126=>"101000001",
  27127=>"001010000",
  27128=>"101110011",
  27129=>"111101010",
  27130=>"000011110",
  27131=>"001010001",
  27132=>"001001110",
  27133=>"001101111",
  27134=>"010110000",
  27135=>"000111111",
  27136=>"101111100",
  27137=>"100011111",
  27138=>"101011000",
  27139=>"010000111",
  27140=>"100110101",
  27141=>"010111101",
  27142=>"111110110",
  27143=>"001111001",
  27144=>"010010100",
  27145=>"110001111",
  27146=>"110011110",
  27147=>"100000011",
  27148=>"110110100",
  27149=>"100110101",
  27150=>"001111000",
  27151=>"110111000",
  27152=>"010001111",
  27153=>"111111001",
  27154=>"111111111",
  27155=>"111110011",
  27156=>"100011010",
  27157=>"001100111",
  27158=>"110111011",
  27159=>"010100110",
  27160=>"111111110",
  27161=>"100011111",
  27162=>"010100010",
  27163=>"011101100",
  27164=>"111111111",
  27165=>"001000001",
  27166=>"001000011",
  27167=>"110001110",
  27168=>"010100101",
  27169=>"010011101",
  27170=>"001010110",
  27171=>"000111100",
  27172=>"011101101",
  27173=>"011001101",
  27174=>"110101101",
  27175=>"100001000",
  27176=>"000110110",
  27177=>"101001110",
  27178=>"110010101",
  27179=>"001000111",
  27180=>"111000100",
  27181=>"100111101",
  27182=>"011111100",
  27183=>"100111111",
  27184=>"010100100",
  27185=>"110001011",
  27186=>"011001101",
  27187=>"011101000",
  27188=>"101110101",
  27189=>"100001010",
  27190=>"001100100",
  27191=>"000010100",
  27192=>"000111000",
  27193=>"001101100",
  27194=>"010000010",
  27195=>"111110000",
  27196=>"010011000",
  27197=>"000001101",
  27198=>"011110011",
  27199=>"001000111",
  27200=>"001001010",
  27201=>"100110000",
  27202=>"011010101",
  27203=>"110000011",
  27204=>"010001110",
  27205=>"111000001",
  27206=>"010111001",
  27207=>"001000011",
  27208=>"110010100",
  27209=>"001100100",
  27210=>"100110011",
  27211=>"100000110",
  27212=>"000010101",
  27213=>"001101111",
  27214=>"001011000",
  27215=>"111100101",
  27216=>"010111000",
  27217=>"000000110",
  27218=>"110100100",
  27219=>"111100010",
  27220=>"000011110",
  27221=>"111001000",
  27222=>"101100110",
  27223=>"100111110",
  27224=>"000101101",
  27225=>"011000000",
  27226=>"110010111",
  27227=>"101011001",
  27228=>"010101111",
  27229=>"100011101",
  27230=>"111101101",
  27231=>"111011101",
  27232=>"000011001",
  27233=>"011110101",
  27234=>"000111110",
  27235=>"100110010",
  27236=>"010101100",
  27237=>"101000001",
  27238=>"001110101",
  27239=>"111111011",
  27240=>"011010101",
  27241=>"111011100",
  27242=>"101110111",
  27243=>"000100111",
  27244=>"100011111",
  27245=>"110110000",
  27246=>"100000101",
  27247=>"010100110",
  27248=>"110111110",
  27249=>"111000001",
  27250=>"100011000",
  27251=>"000101111",
  27252=>"100100010",
  27253=>"101011111",
  27254=>"000111100",
  27255=>"001010011",
  27256=>"010110001",
  27257=>"011001010",
  27258=>"001010111",
  27259=>"010100111",
  27260=>"100100100",
  27261=>"011110111",
  27262=>"110110111",
  27263=>"000000011",
  27264=>"001001001",
  27265=>"001010100",
  27266=>"101100110",
  27267=>"011110110",
  27268=>"011101101",
  27269=>"110011000",
  27270=>"001111110",
  27271=>"111011110",
  27272=>"101100000",
  27273=>"001110111",
  27274=>"010100101",
  27275=>"001101011",
  27276=>"100100110",
  27277=>"100011111",
  27278=>"100110000",
  27279=>"010101111",
  27280=>"011000111",
  27281=>"001010001",
  27282=>"000101010",
  27283=>"110101101",
  27284=>"110000100",
  27285=>"101101000",
  27286=>"000001011",
  27287=>"100000100",
  27288=>"001100110",
  27289=>"010111111",
  27290=>"101110000",
  27291=>"000101011",
  27292=>"001101010",
  27293=>"110000111",
  27294=>"010100111",
  27295=>"111000010",
  27296=>"100011010",
  27297=>"110111110",
  27298=>"001101000",
  27299=>"110100111",
  27300=>"110100100",
  27301=>"110010100",
  27302=>"111101101",
  27303=>"100111010",
  27304=>"110101101",
  27305=>"001100111",
  27306=>"011001111",
  27307=>"000011110",
  27308=>"001010000",
  27309=>"000100011",
  27310=>"011011000",
  27311=>"110100110",
  27312=>"001001001",
  27313=>"110101101",
  27314=>"110000000",
  27315=>"101000111",
  27316=>"111010111",
  27317=>"011000111",
  27318=>"100000101",
  27319=>"110011011",
  27320=>"001110101",
  27321=>"011111000",
  27322=>"000110101",
  27323=>"101011011",
  27324=>"001111110",
  27325=>"110101111",
  27326=>"111110011",
  27327=>"111110011",
  27328=>"100111101",
  27329=>"001011111",
  27330=>"010110100",
  27331=>"100010100",
  27332=>"101110011",
  27333=>"110110110",
  27334=>"000011000",
  27335=>"101111010",
  27336=>"000011101",
  27337=>"000010010",
  27338=>"101001111",
  27339=>"010100010",
  27340=>"101010111",
  27341=>"001001001",
  27342=>"000110100",
  27343=>"001100111",
  27344=>"100001111",
  27345=>"000000011",
  27346=>"000110001",
  27347=>"010101000",
  27348=>"100000110",
  27349=>"101010100",
  27350=>"011000100",
  27351=>"111100011",
  27352=>"000000000",
  27353=>"100000100",
  27354=>"010101100",
  27355=>"100100110",
  27356=>"110110011",
  27357=>"100111000",
  27358=>"001001101",
  27359=>"010011001",
  27360=>"111010111",
  27361=>"110100111",
  27362=>"101100010",
  27363=>"110100111",
  27364=>"110100101",
  27365=>"011000101",
  27366=>"011010110",
  27367=>"000001110",
  27368=>"000111011",
  27369=>"110011111",
  27370=>"111011101",
  27371=>"111111111",
  27372=>"010111110",
  27373=>"010100000",
  27374=>"000011100",
  27375=>"101000010",
  27376=>"000101001",
  27377=>"010010001",
  27378=>"010100001",
  27379=>"101100101",
  27380=>"000000010",
  27381=>"110011011",
  27382=>"010000011",
  27383=>"010000100",
  27384=>"111100101",
  27385=>"011000011",
  27386=>"111100101",
  27387=>"100101101",
  27388=>"110000010",
  27389=>"010111000",
  27390=>"101001010",
  27391=>"010000000",
  27392=>"000111101",
  27393=>"110100000",
  27394=>"101011101",
  27395=>"111100110",
  27396=>"000000010",
  27397=>"000101100",
  27398=>"000110100",
  27399=>"010001101",
  27400=>"101011001",
  27401=>"000000101",
  27402=>"010001101",
  27403=>"110110010",
  27404=>"110111101",
  27405=>"110101001",
  27406=>"100101110",
  27407=>"001001111",
  27408=>"000001000",
  27409=>"001000010",
  27410=>"010100010",
  27411=>"000010001",
  27412=>"001011101",
  27413=>"101011101",
  27414=>"110011010",
  27415=>"101000001",
  27416=>"011000011",
  27417=>"100000110",
  27418=>"011101011",
  27419=>"001001011",
  27420=>"101110100",
  27421=>"011000111",
  27422=>"001111101",
  27423=>"100000100",
  27424=>"110100100",
  27425=>"000000001",
  27426=>"111110111",
  27427=>"001101100",
  27428=>"010001001",
  27429=>"001001010",
  27430=>"110111111",
  27431=>"011011101",
  27432=>"110001110",
  27433=>"100100111",
  27434=>"000111000",
  27435=>"010101001",
  27436=>"101101101",
  27437=>"111000001",
  27438=>"111011110",
  27439=>"011011101",
  27440=>"000001111",
  27441=>"110111111",
  27442=>"101110101",
  27443=>"010000101",
  27444=>"000001010",
  27445=>"110001101",
  27446=>"010000011",
  27447=>"110000011",
  27448=>"000010010",
  27449=>"111000001",
  27450=>"110100110",
  27451=>"001101010",
  27452=>"010010001",
  27453=>"001000111",
  27454=>"011011111",
  27455=>"110000110",
  27456=>"001110100",
  27457=>"000001100",
  27458=>"100100001",
  27459=>"010110011",
  27460=>"001100110",
  27461=>"010101011",
  27462=>"011101111",
  27463=>"101111100",
  27464=>"100111001",
  27465=>"111111000",
  27466=>"010010101",
  27467=>"100110100",
  27468=>"101100011",
  27469=>"010000001",
  27470=>"010000100",
  27471=>"000001111",
  27472=>"100100100",
  27473=>"111111101",
  27474=>"011011110",
  27475=>"010011101",
  27476=>"000011111",
  27477=>"111011010",
  27478=>"010100111",
  27479=>"111111101",
  27480=>"100011010",
  27481=>"110010000",
  27482=>"100001110",
  27483=>"101000011",
  27484=>"111010110",
  27485=>"101010010",
  27486=>"111100001",
  27487=>"100110100",
  27488=>"011110011",
  27489=>"011110101",
  27490=>"111111011",
  27491=>"010001010",
  27492=>"100110000",
  27493=>"110010011",
  27494=>"001010001",
  27495=>"111100111",
  27496=>"100100010",
  27497=>"101101100",
  27498=>"001100111",
  27499=>"001001101",
  27500=>"101001001",
  27501=>"110110111",
  27502=>"010111101",
  27503=>"011010101",
  27504=>"001010010",
  27505=>"101010100",
  27506=>"000010010",
  27507=>"100011110",
  27508=>"010111111",
  27509=>"110011101",
  27510=>"000111110",
  27511=>"110000111",
  27512=>"101000110",
  27513=>"001101011",
  27514=>"011100111",
  27515=>"011000101",
  27516=>"010000110",
  27517=>"110011010",
  27518=>"111010110",
  27519=>"011111101",
  27520=>"100010000",
  27521=>"001010010",
  27522=>"111111111",
  27523=>"001101000",
  27524=>"110111100",
  27525=>"000000000",
  27526=>"101010110",
  27527=>"110001101",
  27528=>"101110010",
  27529=>"010111100",
  27530=>"101111000",
  27531=>"010101100",
  27532=>"110000001",
  27533=>"101111011",
  27534=>"011001110",
  27535=>"101100011",
  27536=>"000100111",
  27537=>"101111011",
  27538=>"000011100",
  27539=>"001110110",
  27540=>"000100110",
  27541=>"000101000",
  27542=>"011000010",
  27543=>"011010010",
  27544=>"011111100",
  27545=>"110110010",
  27546=>"010100110",
  27547=>"101000010",
  27548=>"000011000",
  27549=>"111101001",
  27550=>"010010001",
  27551=>"100111010",
  27552=>"101011011",
  27553=>"110101001",
  27554=>"111100011",
  27555=>"101010000",
  27556=>"001101011",
  27557=>"101111101",
  27558=>"100100110",
  27559=>"100001101",
  27560=>"001000001",
  27561=>"111111111",
  27562=>"000101010",
  27563=>"011001000",
  27564=>"000001011",
  27565=>"000011010",
  27566=>"101100010",
  27567=>"110100000",
  27568=>"001000101",
  27569=>"101101000",
  27570=>"011101011",
  27571=>"011000010",
  27572=>"011001111",
  27573=>"101111101",
  27574=>"000010000",
  27575=>"100011111",
  27576=>"011110110",
  27577=>"011101011",
  27578=>"101000001",
  27579=>"011110110",
  27580=>"111010110",
  27581=>"010010010",
  27582=>"011110010",
  27583=>"011000000",
  27584=>"111101010",
  27585=>"011111101",
  27586=>"011001000",
  27587=>"111100011",
  27588=>"110111101",
  27589=>"110010100",
  27590=>"001110000",
  27591=>"100100100",
  27592=>"110000110",
  27593=>"101111001",
  27594=>"011010101",
  27595=>"101100111",
  27596=>"110001110",
  27597=>"100010100",
  27598=>"111001110",
  27599=>"000001011",
  27600=>"101001100",
  27601=>"010001111",
  27602=>"111000000",
  27603=>"110000101",
  27604=>"101100110",
  27605=>"111111010",
  27606=>"100010001",
  27607=>"111111110",
  27608=>"110111101",
  27609=>"010000110",
  27610=>"001101001",
  27611=>"001110001",
  27612=>"010111100",
  27613=>"010110010",
  27614=>"001000100",
  27615=>"110101111",
  27616=>"111111101",
  27617=>"100001110",
  27618=>"001010100",
  27619=>"010110101",
  27620=>"011110011",
  27621=>"111111001",
  27622=>"011100001",
  27623=>"011001100",
  27624=>"111111100",
  27625=>"110110111",
  27626=>"100110010",
  27627=>"100011011",
  27628=>"000110010",
  27629=>"000100101",
  27630=>"110011110",
  27631=>"010001101",
  27632=>"100111111",
  27633=>"100101010",
  27634=>"001000011",
  27635=>"000101010",
  27636=>"010101000",
  27637=>"101001000",
  27638=>"100101101",
  27639=>"011001100",
  27640=>"010011111",
  27641=>"100110001",
  27642=>"100111101",
  27643=>"110000011",
  27644=>"100011011",
  27645=>"010001010",
  27646=>"110111110",
  27647=>"101010100",
  27648=>"101100101",
  27649=>"001011101",
  27650=>"000110100",
  27651=>"101110110",
  27652=>"001011000",
  27653=>"111001111",
  27654=>"101010110",
  27655=>"111110001",
  27656=>"000110000",
  27657=>"011111110",
  27658=>"110100110",
  27659=>"100100010",
  27660=>"010000011",
  27661=>"111100000",
  27662=>"011101000",
  27663=>"101111111",
  27664=>"111110101",
  27665=>"011000000",
  27666=>"100000000",
  27667=>"011001111",
  27668=>"011111001",
  27669=>"110111011",
  27670=>"011110011",
  27671=>"111010001",
  27672=>"100100111",
  27673=>"101010000",
  27674=>"001000010",
  27675=>"011010000",
  27676=>"111100000",
  27677=>"101100111",
  27678=>"000010110",
  27679=>"101000000",
  27680=>"101100000",
  27681=>"011010000",
  27682=>"101000110",
  27683=>"011010000",
  27684=>"000110110",
  27685=>"000001111",
  27686=>"100010100",
  27687=>"100111000",
  27688=>"011011100",
  27689=>"010001011",
  27690=>"111110101",
  27691=>"000110001",
  27692=>"011001100",
  27693=>"010100111",
  27694=>"111100100",
  27695=>"010110000",
  27696=>"001101111",
  27697=>"101010011",
  27698=>"101111000",
  27699=>"000110011",
  27700=>"100101111",
  27701=>"100001000",
  27702=>"110111000",
  27703=>"010000100",
  27704=>"000000101",
  27705=>"110110000",
  27706=>"111000110",
  27707=>"110000001",
  27708=>"111100100",
  27709=>"011010110",
  27710=>"010001100",
  27711=>"111100111",
  27712=>"010111010",
  27713=>"000111111",
  27714=>"110110000",
  27715=>"000011001",
  27716=>"001000100",
  27717=>"001010010",
  27718=>"001111000",
  27719=>"000010111",
  27720=>"100010110",
  27721=>"101110000",
  27722=>"010001100",
  27723=>"110111110",
  27724=>"110100101",
  27725=>"001101111",
  27726=>"101001011",
  27727=>"011100101",
  27728=>"010001110",
  27729=>"110001001",
  27730=>"011010100",
  27731=>"000010111",
  27732=>"110001001",
  27733=>"101001111",
  27734=>"101010111",
  27735=>"001100100",
  27736=>"000010001",
  27737=>"111000111",
  27738=>"001011101",
  27739=>"100000000",
  27740=>"000100100",
  27741=>"000100001",
  27742=>"010010011",
  27743=>"010001011",
  27744=>"111011111",
  27745=>"000100011",
  27746=>"011100111",
  27747=>"001010110",
  27748=>"001001100",
  27749=>"011110101",
  27750=>"000111100",
  27751=>"111100101",
  27752=>"001000100",
  27753=>"011001100",
  27754=>"010110010",
  27755=>"101010010",
  27756=>"110110000",
  27757=>"110010000",
  27758=>"110000011",
  27759=>"001010110",
  27760=>"110110110",
  27761=>"100000001",
  27762=>"000111111",
  27763=>"010000110",
  27764=>"100101011",
  27765=>"001000101",
  27766=>"110110101",
  27767=>"001010110",
  27768=>"011101000",
  27769=>"110001111",
  27770=>"000110111",
  27771=>"110110100",
  27772=>"100100101",
  27773=>"100100011",
  27774=>"111110111",
  27775=>"111010000",
  27776=>"101101111",
  27777=>"101010000",
  27778=>"011011110",
  27779=>"010010100",
  27780=>"101010100",
  27781=>"100010010",
  27782=>"110011100",
  27783=>"100110110",
  27784=>"010010110",
  27785=>"100011011",
  27786=>"100000000",
  27787=>"100100011",
  27788=>"001101101",
  27789=>"101100101",
  27790=>"011000000",
  27791=>"101110010",
  27792=>"111001100",
  27793=>"000110101",
  27794=>"111011011",
  27795=>"000010001",
  27796=>"011010111",
  27797=>"001111011",
  27798=>"011000000",
  27799=>"100000010",
  27800=>"001101100",
  27801=>"011010010",
  27802=>"111101000",
  27803=>"110011010",
  27804=>"010100000",
  27805=>"000011010",
  27806=>"001011111",
  27807=>"010011010",
  27808=>"010101001",
  27809=>"011011000",
  27810=>"110010101",
  27811=>"000010111",
  27812=>"110001000",
  27813=>"111100101",
  27814=>"010110100",
  27815=>"101011000",
  27816=>"100101111",
  27817=>"100111101",
  27818=>"000010000",
  27819=>"110101101",
  27820=>"011001101",
  27821=>"110000101",
  27822=>"110011000",
  27823=>"000111110",
  27824=>"000010000",
  27825=>"010011011",
  27826=>"000001100",
  27827=>"011100100",
  27828=>"100000011",
  27829=>"001100010",
  27830=>"101111111",
  27831=>"101000001",
  27832=>"000000001",
  27833=>"010011001",
  27834=>"010010000",
  27835=>"111000111",
  27836=>"100010111",
  27837=>"111011011",
  27838=>"101010000",
  27839=>"011100001",
  27840=>"000100111",
  27841=>"001000001",
  27842=>"000111111",
  27843=>"100111101",
  27844=>"001111010",
  27845=>"001011011",
  27846=>"010100000",
  27847=>"111001010",
  27848=>"000010101",
  27849=>"111010011",
  27850=>"111001011",
  27851=>"111000000",
  27852=>"100110010",
  27853=>"100001100",
  27854=>"100000010",
  27855=>"111101110",
  27856=>"100010011",
  27857=>"010000101",
  27858=>"100110000",
  27859=>"010010010",
  27860=>"100101000",
  27861=>"001010111",
  27862=>"101101011",
  27863=>"000101111",
  27864=>"000001101",
  27865=>"101111010",
  27866=>"011110010",
  27867=>"101001100",
  27868=>"001101011",
  27869=>"000110010",
  27870=>"000001001",
  27871=>"111100110",
  27872=>"000101110",
  27873=>"010011101",
  27874=>"010100111",
  27875=>"110001010",
  27876=>"110011100",
  27877=>"011110111",
  27878=>"111011010",
  27879=>"000101101",
  27880=>"110101001",
  27881=>"001000111",
  27882=>"000000000",
  27883=>"011010001",
  27884=>"001010011",
  27885=>"010111100",
  27886=>"010001111",
  27887=>"111000010",
  27888=>"110111110",
  27889=>"001000010",
  27890=>"010110010",
  27891=>"101010000",
  27892=>"111110110",
  27893=>"001010000",
  27894=>"111010011",
  27895=>"111100000",
  27896=>"010101001",
  27897=>"110101111",
  27898=>"110101100",
  27899=>"010000101",
  27900=>"011000001",
  27901=>"110110110",
  27902=>"000110110",
  27903=>"000101011",
  27904=>"010010111",
  27905=>"010100010",
  27906=>"011001101",
  27907=>"010110010",
  27908=>"000010111",
  27909=>"011010100",
  27910=>"101000110",
  27911=>"100010110",
  27912=>"010110010",
  27913=>"010111000",
  27914=>"111111110",
  27915=>"010111111",
  27916=>"000000100",
  27917=>"000011010",
  27918=>"000001100",
  27919=>"110001101",
  27920=>"011000010",
  27921=>"000101110",
  27922=>"110001011",
  27923=>"100000110",
  27924=>"100000111",
  27925=>"101110000",
  27926=>"101110001",
  27927=>"011111101",
  27928=>"011101111",
  27929=>"001001101",
  27930=>"000101000",
  27931=>"001100001",
  27932=>"101100001",
  27933=>"001010001",
  27934=>"010110001",
  27935=>"101101001",
  27936=>"111010001",
  27937=>"000011000",
  27938=>"110001110",
  27939=>"010001001",
  27940=>"110101100",
  27941=>"010001110",
  27942=>"011111000",
  27943=>"000010010",
  27944=>"101100011",
  27945=>"110110010",
  27946=>"011001101",
  27947=>"110110000",
  27948=>"111010001",
  27949=>"110010000",
  27950=>"001000000",
  27951=>"101010100",
  27952=>"111101001",
  27953=>"101111000",
  27954=>"010100000",
  27955=>"000100110",
  27956=>"101011100",
  27957=>"111110100",
  27958=>"110000100",
  27959=>"110011010",
  27960=>"010100010",
  27961=>"001100100",
  27962=>"001110101",
  27963=>"011000010",
  27964=>"011100000",
  27965=>"111011101",
  27966=>"111111001",
  27967=>"110000000",
  27968=>"011111010",
  27969=>"010110110",
  27970=>"011010111",
  27971=>"001100001",
  27972=>"101010001",
  27973=>"100110011",
  27974=>"001111010",
  27975=>"000001010",
  27976=>"001011011",
  27977=>"010000110",
  27978=>"100101111",
  27979=>"110100000",
  27980=>"011101110",
  27981=>"010000001",
  27982=>"000110100",
  27983=>"011001000",
  27984=>"011101101",
  27985=>"111011111",
  27986=>"101001101",
  27987=>"111110111",
  27988=>"110011111",
  27989=>"100011001",
  27990=>"110110100",
  27991=>"000100111",
  27992=>"110011111",
  27993=>"011011010",
  27994=>"111111100",
  27995=>"100001010",
  27996=>"110110000",
  27997=>"011011100",
  27998=>"100001111",
  27999=>"011110000",
  28000=>"010011001",
  28001=>"010110000",
  28002=>"000010110",
  28003=>"000100101",
  28004=>"101001011",
  28005=>"111110010",
  28006=>"010010101",
  28007=>"100110000",
  28008=>"100001010",
  28009=>"110001101",
  28010=>"000110010",
  28011=>"000110000",
  28012=>"110001000",
  28013=>"101111111",
  28014=>"000011000",
  28015=>"001101100",
  28016=>"100000001",
  28017=>"010100010",
  28018=>"101011010",
  28019=>"100001000",
  28020=>"010000010",
  28021=>"111110111",
  28022=>"010001100",
  28023=>"000110000",
  28024=>"010001011",
  28025=>"001000001",
  28026=>"000011111",
  28027=>"101000010",
  28028=>"000001010",
  28029=>"101100011",
  28030=>"000101100",
  28031=>"000110010",
  28032=>"100100101",
  28033=>"100001100",
  28034=>"001100111",
  28035=>"010101101",
  28036=>"101110101",
  28037=>"111011110",
  28038=>"011011000",
  28039=>"011001010",
  28040=>"111110011",
  28041=>"011001000",
  28042=>"000011111",
  28043=>"001001101",
  28044=>"000111000",
  28045=>"111011110",
  28046=>"110100111",
  28047=>"001101111",
  28048=>"111010100",
  28049=>"001001000",
  28050=>"111100010",
  28051=>"011100110",
  28052=>"010011100",
  28053=>"101101011",
  28054=>"000000101",
  28055=>"010110110",
  28056=>"111011101",
  28057=>"100110101",
  28058=>"100011101",
  28059=>"011001100",
  28060=>"101010100",
  28061=>"010010010",
  28062=>"000011011",
  28063=>"101000111",
  28064=>"011011000",
  28065=>"111000000",
  28066=>"010111001",
  28067=>"001000000",
  28068=>"110111110",
  28069=>"000101011",
  28070=>"001111010",
  28071=>"011111111",
  28072=>"001001010",
  28073=>"001010101",
  28074=>"110100110",
  28075=>"011010001",
  28076=>"111111101",
  28077=>"011111011",
  28078=>"110111011",
  28079=>"010111011",
  28080=>"100010000",
  28081=>"011111110",
  28082=>"110111110",
  28083=>"010111000",
  28084=>"000010000",
  28085=>"100001100",
  28086=>"001101000",
  28087=>"110111011",
  28088=>"011010100",
  28089=>"001101101",
  28090=>"101010110",
  28091=>"011110001",
  28092=>"110001111",
  28093=>"101000101",
  28094=>"110000110",
  28095=>"010000000",
  28096=>"100101101",
  28097=>"100010101",
  28098=>"011000101",
  28099=>"101000010",
  28100=>"011001101",
  28101=>"011111001",
  28102=>"011110101",
  28103=>"010011011",
  28104=>"000111001",
  28105=>"001111111",
  28106=>"110011101",
  28107=>"100111100",
  28108=>"110010001",
  28109=>"111010110",
  28110=>"000001100",
  28111=>"111110100",
  28112=>"011011100",
  28113=>"010001000",
  28114=>"011011100",
  28115=>"011000010",
  28116=>"110011101",
  28117=>"000110101",
  28118=>"000010100",
  28119=>"101110110",
  28120=>"100101011",
  28121=>"110101000",
  28122=>"011011001",
  28123=>"010110101",
  28124=>"100100001",
  28125=>"100100110",
  28126=>"011101101",
  28127=>"000111111",
  28128=>"011100100",
  28129=>"001101010",
  28130=>"110100110",
  28131=>"001011000",
  28132=>"010110001",
  28133=>"011000010",
  28134=>"010101101",
  28135=>"001010100",
  28136=>"011111001",
  28137=>"111010101",
  28138=>"101000010",
  28139=>"011100010",
  28140=>"000101111",
  28141=>"000110000",
  28142=>"010000110",
  28143=>"100001001",
  28144=>"011111111",
  28145=>"101001001",
  28146=>"100101001",
  28147=>"111111001",
  28148=>"010110111",
  28149=>"000010010",
  28150=>"000000011",
  28151=>"101001000",
  28152=>"100011011",
  28153=>"101101001",
  28154=>"110001011",
  28155=>"110110101",
  28156=>"000100111",
  28157=>"111010001",
  28158=>"101101010",
  28159=>"000001001",
  28160=>"101000010",
  28161=>"100010011",
  28162=>"110000101",
  28163=>"101110101",
  28164=>"110000010",
  28165=>"110001010",
  28166=>"001101101",
  28167=>"111110011",
  28168=>"100100101",
  28169=>"111011011",
  28170=>"100101111",
  28171=>"010100111",
  28172=>"001100010",
  28173=>"111000101",
  28174=>"000110111",
  28175=>"100111111",
  28176=>"010000111",
  28177=>"101100000",
  28178=>"010010010",
  28179=>"101100000",
  28180=>"000100111",
  28181=>"001111111",
  28182=>"000100001",
  28183=>"100111011",
  28184=>"011010101",
  28185=>"001000111",
  28186=>"000011011",
  28187=>"110101100",
  28188=>"101111100",
  28189=>"110001100",
  28190=>"110011100",
  28191=>"000101111",
  28192=>"111100111",
  28193=>"111101110",
  28194=>"000011111",
  28195=>"000010011",
  28196=>"111011000",
  28197=>"110100010",
  28198=>"101100000",
  28199=>"001010110",
  28200=>"111111101",
  28201=>"000101110",
  28202=>"101011100",
  28203=>"010000101",
  28204=>"011100111",
  28205=>"100000000",
  28206=>"101000101",
  28207=>"010010111",
  28208=>"110001010",
  28209=>"110010101",
  28210=>"111001001",
  28211=>"100010101",
  28212=>"100110111",
  28213=>"011100101",
  28214=>"100110000",
  28215=>"000100101",
  28216=>"111110100",
  28217=>"000010000",
  28218=>"110111101",
  28219=>"101101000",
  28220=>"010100100",
  28221=>"010001111",
  28222=>"000001001",
  28223=>"101111010",
  28224=>"001000100",
  28225=>"100011110",
  28226=>"100011000",
  28227=>"001010000",
  28228=>"100010111",
  28229=>"111011101",
  28230=>"001110110",
  28231=>"000101111",
  28232=>"100111111",
  28233=>"000101101",
  28234=>"000001001",
  28235=>"010011110",
  28236=>"100110110",
  28237=>"010010000",
  28238=>"110010011",
  28239=>"001101111",
  28240=>"111110111",
  28241=>"000011111",
  28242=>"110101101",
  28243=>"000001101",
  28244=>"110101110",
  28245=>"000001000",
  28246=>"010010100",
  28247=>"010010110",
  28248=>"000100111",
  28249=>"101110100",
  28250=>"000010010",
  28251=>"101011000",
  28252=>"110011001",
  28253=>"000100011",
  28254=>"111100000",
  28255=>"111100011",
  28256=>"010100100",
  28257=>"100100100",
  28258=>"011001000",
  28259=>"001110110",
  28260=>"011111100",
  28261=>"101000111",
  28262=>"111011110",
  28263=>"100011100",
  28264=>"111011100",
  28265=>"100101000",
  28266=>"111000011",
  28267=>"011111010",
  28268=>"010000100",
  28269=>"100000101",
  28270=>"001011000",
  28271=>"110001000",
  28272=>"001111011",
  28273=>"011000100",
  28274=>"000100000",
  28275=>"110011100",
  28276=>"010001100",
  28277=>"000001001",
  28278=>"110110010",
  28279=>"010110010",
  28280=>"110010010",
  28281=>"001010111",
  28282=>"111110110",
  28283=>"100101001",
  28284=>"111001111",
  28285=>"010111010",
  28286=>"010000000",
  28287=>"010110010",
  28288=>"111110100",
  28289=>"111111000",
  28290=>"010110011",
  28291=>"101000100",
  28292=>"000110010",
  28293=>"110000001",
  28294=>"110001011",
  28295=>"111011000",
  28296=>"000100011",
  28297=>"011011010",
  28298=>"111100110",
  28299=>"011110101",
  28300=>"001001100",
  28301=>"000000001",
  28302=>"001001110",
  28303=>"100011000",
  28304=>"010100011",
  28305=>"111101011",
  28306=>"010001111",
  28307=>"000101101",
  28308=>"000000011",
  28309=>"000101110",
  28310=>"111001110",
  28311=>"100001111",
  28312=>"001100011",
  28313=>"100000010",
  28314=>"001001011",
  28315=>"011111111",
  28316=>"111110111",
  28317=>"110010101",
  28318=>"010011101",
  28319=>"000000011",
  28320=>"001101101",
  28321=>"000110111",
  28322=>"110000111",
  28323=>"110100000",
  28324=>"101011000",
  28325=>"001110011",
  28326=>"000100010",
  28327=>"101000111",
  28328=>"001010010",
  28329=>"110011110",
  28330=>"101010010",
  28331=>"001110100",
  28332=>"111011100",
  28333=>"000000000",
  28334=>"010101001",
  28335=>"100100001",
  28336=>"011100011",
  28337=>"010000010",
  28338=>"000110101",
  28339=>"111100011",
  28340=>"011001010",
  28341=>"100110001",
  28342=>"100101001",
  28343=>"000100101",
  28344=>"101110111",
  28345=>"100100111",
  28346=>"111100010",
  28347=>"000000110",
  28348=>"001100100",
  28349=>"001010111",
  28350=>"010001101",
  28351=>"011010000",
  28352=>"000001111",
  28353=>"000111100",
  28354=>"001000101",
  28355=>"010010111",
  28356=>"010011010",
  28357=>"000000001",
  28358=>"101010011",
  28359=>"011101101",
  28360=>"010010000",
  28361=>"001110111",
  28362=>"111010011",
  28363=>"101111111",
  28364=>"101101100",
  28365=>"111111101",
  28366=>"000101110",
  28367=>"000110011",
  28368=>"110000010",
  28369=>"111110110",
  28370=>"000110100",
  28371=>"000101000",
  28372=>"010011101",
  28373=>"111011010",
  28374=>"000001101",
  28375=>"000010111",
  28376=>"110011010",
  28377=>"000100011",
  28378=>"110001010",
  28379=>"110101100",
  28380=>"100111110",
  28381=>"111011000",
  28382=>"110010000",
  28383=>"111010011",
  28384=>"100110111",
  28385=>"001111010",
  28386=>"000110001",
  28387=>"000001111",
  28388=>"101011001",
  28389=>"111010101",
  28390=>"011000100",
  28391=>"110011000",
  28392=>"101101111",
  28393=>"100101100",
  28394=>"111001010",
  28395=>"111011110",
  28396=>"101100010",
  28397=>"011001010",
  28398=>"110011111",
  28399=>"010101001",
  28400=>"101100111",
  28401=>"110100101",
  28402=>"110000110",
  28403=>"000001001",
  28404=>"010001111",
  28405=>"110101101",
  28406=>"000111000",
  28407=>"100000110",
  28408=>"000011001",
  28409=>"000110000",
  28410=>"100101010",
  28411=>"101110100",
  28412=>"111011011",
  28413=>"110110111",
  28414=>"100011101",
  28415=>"001010111",
  28416=>"100001001",
  28417=>"101011111",
  28418=>"011010110",
  28419=>"011101100",
  28420=>"111111011",
  28421=>"010110011",
  28422=>"001010111",
  28423=>"100101010",
  28424=>"110010010",
  28425=>"110101001",
  28426=>"110001001",
  28427=>"100010001",
  28428=>"111010000",
  28429=>"001100111",
  28430=>"011010010",
  28431=>"000101101",
  28432=>"101000111",
  28433=>"011101110",
  28434=>"110001001",
  28435=>"101010000",
  28436=>"110000001",
  28437=>"110011011",
  28438=>"000000010",
  28439=>"010100000",
  28440=>"100110100",
  28441=>"001010110",
  28442=>"111001011",
  28443=>"110101000",
  28444=>"011010001",
  28445=>"111111111",
  28446=>"000010010",
  28447=>"111000110",
  28448=>"100100101",
  28449=>"001101001",
  28450=>"010000100",
  28451=>"110110001",
  28452=>"000000001",
  28453=>"010110000",
  28454=>"110010011",
  28455=>"110100010",
  28456=>"101100101",
  28457=>"101000000",
  28458=>"101011010",
  28459=>"110000111",
  28460=>"111111011",
  28461=>"000110110",
  28462=>"011100101",
  28463=>"000010001",
  28464=>"000000001",
  28465=>"011000001",
  28466=>"010000110",
  28467=>"101010111",
  28468=>"001110100",
  28469=>"000110100",
  28470=>"001010000",
  28471=>"001101000",
  28472=>"010001110",
  28473=>"111101100",
  28474=>"101110111",
  28475=>"000010100",
  28476=>"010110010",
  28477=>"000101111",
  28478=>"010001000",
  28479=>"000100110",
  28480=>"100100000",
  28481=>"111010010",
  28482=>"001001100",
  28483=>"101010011",
  28484=>"000110110",
  28485=>"101100111",
  28486=>"011000001",
  28487=>"111000010",
  28488=>"101000010",
  28489=>"111010101",
  28490=>"010100101",
  28491=>"011010000",
  28492=>"001000010",
  28493=>"101011000",
  28494=>"001110101",
  28495=>"111111101",
  28496=>"010111110",
  28497=>"001000100",
  28498=>"110111101",
  28499=>"110001010",
  28500=>"000111010",
  28501=>"111000001",
  28502=>"000001001",
  28503=>"011101011",
  28504=>"101101001",
  28505=>"110101111",
  28506=>"010001011",
  28507=>"110001101",
  28508=>"111101011",
  28509=>"000111111",
  28510=>"111111000",
  28511=>"111010010",
  28512=>"001101100",
  28513=>"111001100",
  28514=>"001100011",
  28515=>"001001010",
  28516=>"110000000",
  28517=>"001111110",
  28518=>"111111010",
  28519=>"110111100",
  28520=>"001110000",
  28521=>"011010001",
  28522=>"101001001",
  28523=>"100101101",
  28524=>"100010101",
  28525=>"001010101",
  28526=>"101001000",
  28527=>"010111010",
  28528=>"010111111",
  28529=>"010001111",
  28530=>"101010001",
  28531=>"001000101",
  28532=>"010100001",
  28533=>"100101000",
  28534=>"110010001",
  28535=>"000001000",
  28536=>"011111001",
  28537=>"000110010",
  28538=>"111111111",
  28539=>"111111010",
  28540=>"000001001",
  28541=>"110001010",
  28542=>"110010000",
  28543=>"000001100",
  28544=>"101011101",
  28545=>"001101010",
  28546=>"011000001",
  28547=>"111000111",
  28548=>"001000000",
  28549=>"101011101",
  28550=>"100101001",
  28551=>"010011011",
  28552=>"001000101",
  28553=>"010010011",
  28554=>"111101000",
  28555=>"110010010",
  28556=>"011000001",
  28557=>"101001101",
  28558=>"110101101",
  28559=>"000010101",
  28560=>"011110010",
  28561=>"011110011",
  28562=>"000000110",
  28563=>"110011100",
  28564=>"010110111",
  28565=>"000100011",
  28566=>"101010110",
  28567=>"011111011",
  28568=>"001000111",
  28569=>"101001000",
  28570=>"011010111",
  28571=>"011110000",
  28572=>"100100011",
  28573=>"001101001",
  28574=>"110001011",
  28575=>"000101011",
  28576=>"101001000",
  28577=>"110000010",
  28578=>"000010001",
  28579=>"100000000",
  28580=>"110111010",
  28581=>"111101100",
  28582=>"111100010",
  28583=>"011010101",
  28584=>"011100110",
  28585=>"010101001",
  28586=>"101000111",
  28587=>"111010100",
  28588=>"000000010",
  28589=>"000000101",
  28590=>"000111101",
  28591=>"000101111",
  28592=>"111111011",
  28593=>"111011011",
  28594=>"000101010",
  28595=>"111100101",
  28596=>"111100000",
  28597=>"010010111",
  28598=>"011111110",
  28599=>"000001111",
  28600=>"000111111",
  28601=>"010110100",
  28602=>"011000111",
  28603=>"000100101",
  28604=>"111110001",
  28605=>"000110011",
  28606=>"000001000",
  28607=>"000010111",
  28608=>"100111111",
  28609=>"110000100",
  28610=>"001011000",
  28611=>"111110010",
  28612=>"111000111",
  28613=>"000001010",
  28614=>"111100110",
  28615=>"011010000",
  28616=>"101100111",
  28617=>"110010101",
  28618=>"001001000",
  28619=>"110101100",
  28620=>"101011110",
  28621=>"011111001",
  28622=>"100000111",
  28623=>"101100101",
  28624=>"100111101",
  28625=>"111001101",
  28626=>"111010000",
  28627=>"001010111",
  28628=>"110001111",
  28629=>"111101110",
  28630=>"111101101",
  28631=>"111100101",
  28632=>"011000100",
  28633=>"111101001",
  28634=>"101111111",
  28635=>"111011011",
  28636=>"011111111",
  28637=>"000010110",
  28638=>"110011011",
  28639=>"110000000",
  28640=>"000011110",
  28641=>"110101100",
  28642=>"110010100",
  28643=>"000010101",
  28644=>"111001000",
  28645=>"110100110",
  28646=>"000111101",
  28647=>"101100100",
  28648=>"100010000",
  28649=>"111111101",
  28650=>"011011110",
  28651=>"011100111",
  28652=>"000110101",
  28653=>"101011111",
  28654=>"101010000",
  28655=>"011001110",
  28656=>"100011110",
  28657=>"010011001",
  28658=>"100100110",
  28659=>"110101110",
  28660=>"000011100",
  28661=>"001111011",
  28662=>"011100110",
  28663=>"000001011",
  28664=>"001110111",
  28665=>"111000100",
  28666=>"100010111",
  28667=>"001111110",
  28668=>"001100111",
  28669=>"100000101",
  28670=>"011000100",
  28671=>"111100010",
  28672=>"101001110",
  28673=>"100100101",
  28674=>"111000101",
  28675=>"011110001",
  28676=>"010010110",
  28677=>"001000101",
  28678=>"001010001",
  28679=>"111111100",
  28680=>"101001000",
  28681=>"000011000",
  28682=>"101111101",
  28683=>"000001100",
  28684=>"111000001",
  28685=>"001110011",
  28686=>"001000010",
  28687=>"101100001",
  28688=>"101110100",
  28689=>"111011110",
  28690=>"001010111",
  28691=>"001000101",
  28692=>"110001000",
  28693=>"000000110",
  28694=>"110111101",
  28695=>"000001000",
  28696=>"010111100",
  28697=>"011010001",
  28698=>"111110100",
  28699=>"111111011",
  28700=>"111111111",
  28701=>"111011011",
  28702=>"011000010",
  28703=>"111111011",
  28704=>"101111010",
  28705=>"101110001",
  28706=>"010100001",
  28707=>"111000000",
  28708=>"001101000",
  28709=>"110001111",
  28710=>"000001101",
  28711=>"011011111",
  28712=>"000000100",
  28713=>"111010001",
  28714=>"010111000",
  28715=>"010100010",
  28716=>"100011011",
  28717=>"101100100",
  28718=>"010110110",
  28719=>"011100100",
  28720=>"111010100",
  28721=>"101000001",
  28722=>"010101010",
  28723=>"111101010",
  28724=>"111111110",
  28725=>"110011100",
  28726=>"111101111",
  28727=>"111101101",
  28728=>"000001011",
  28729=>"000001101",
  28730=>"000111110",
  28731=>"000100101",
  28732=>"010110111",
  28733=>"011001011",
  28734=>"010001110",
  28735=>"111100101",
  28736=>"111010100",
  28737=>"111101000",
  28738=>"111110101",
  28739=>"010001110",
  28740=>"000000111",
  28741=>"011100100",
  28742=>"010101100",
  28743=>"111110100",
  28744=>"000001100",
  28745=>"011011111",
  28746=>"110101111",
  28747=>"101010010",
  28748=>"010110101",
  28749=>"101110110",
  28750=>"100100110",
  28751=>"100111001",
  28752=>"000000111",
  28753=>"111000000",
  28754=>"110011111",
  28755=>"010010111",
  28756=>"100101010",
  28757=>"101011101",
  28758=>"011101110",
  28759=>"011111111",
  28760=>"101011111",
  28761=>"101101101",
  28762=>"110101011",
  28763=>"011010011",
  28764=>"001110001",
  28765=>"111000100",
  28766=>"010011110",
  28767=>"100110101",
  28768=>"111000101",
  28769=>"011101100",
  28770=>"000111111",
  28771=>"101100000",
  28772=>"101100101",
  28773=>"010110101",
  28774=>"000101101",
  28775=>"000111010",
  28776=>"111010001",
  28777=>"010000100",
  28778=>"111000111",
  28779=>"011001010",
  28780=>"101010001",
  28781=>"110010110",
  28782=>"100110010",
  28783=>"001111001",
  28784=>"111100000",
  28785=>"001100111",
  28786=>"101010100",
  28787=>"110110010",
  28788=>"000000111",
  28789=>"000001000",
  28790=>"101001001",
  28791=>"111111110",
  28792=>"111101101",
  28793=>"100100100",
  28794=>"011011100",
  28795=>"010110000",
  28796=>"010111110",
  28797=>"000010001",
  28798=>"000011100",
  28799=>"010110110",
  28800=>"011110000",
  28801=>"100110100",
  28802=>"111111010",
  28803=>"111100000",
  28804=>"110010111",
  28805=>"010001100",
  28806=>"100001111",
  28807=>"000101011",
  28808=>"000010111",
  28809=>"101100100",
  28810=>"001011100",
  28811=>"110101110",
  28812=>"111010111",
  28813=>"100110101",
  28814=>"010001110",
  28815=>"010000101",
  28816=>"111111011",
  28817=>"101111101",
  28818=>"101100110",
  28819=>"101110011",
  28820=>"001111100",
  28821=>"101001110",
  28822=>"011100011",
  28823=>"011011110",
  28824=>"001010100",
  28825=>"000101101",
  28826=>"100111011",
  28827=>"010100000",
  28828=>"101011100",
  28829=>"100100110",
  28830=>"001000011",
  28831=>"100010100",
  28832=>"010010101",
  28833=>"010001010",
  28834=>"101100000",
  28835=>"000001101",
  28836=>"111001110",
  28837=>"110110000",
  28838=>"111101010",
  28839=>"000111111",
  28840=>"110001011",
  28841=>"001101111",
  28842=>"000100110",
  28843=>"010100000",
  28844=>"010111101",
  28845=>"000100001",
  28846=>"000100001",
  28847=>"100101011",
  28848=>"011101000",
  28849=>"100110001",
  28850=>"011000101",
  28851=>"001100101",
  28852=>"011010101",
  28853=>"000110110",
  28854=>"000110110",
  28855=>"101101101",
  28856=>"111010101",
  28857=>"101001111",
  28858=>"010000101",
  28859=>"001000010",
  28860=>"001100000",
  28861=>"010001000",
  28862=>"100101001",
  28863=>"000011010",
  28864=>"111100100",
  28865=>"011011000",
  28866=>"011101001",
  28867=>"111011100",
  28868=>"011011000",
  28869=>"010001000",
  28870=>"111111111",
  28871=>"101101000",
  28872=>"011010101",
  28873=>"001110011",
  28874=>"100010010",
  28875=>"100110010",
  28876=>"000111100",
  28877=>"101000110",
  28878=>"001100011",
  28879=>"110110100",
  28880=>"101101000",
  28881=>"111011100",
  28882=>"001101000",
  28883=>"100010010",
  28884=>"000001000",
  28885=>"000000101",
  28886=>"110100100",
  28887=>"001001011",
  28888=>"101100010",
  28889=>"000111000",
  28890=>"000000011",
  28891=>"001001011",
  28892=>"000111101",
  28893=>"101010101",
  28894=>"110010000",
  28895=>"101101011",
  28896=>"110010101",
  28897=>"011100111",
  28898=>"010110011",
  28899=>"111011011",
  28900=>"111111010",
  28901=>"001011110",
  28902=>"111111110",
  28903=>"011110010",
  28904=>"011010100",
  28905=>"001101010",
  28906=>"001000000",
  28907=>"001101111",
  28908=>"001100011",
  28909=>"001111110",
  28910=>"010101111",
  28911=>"001000110",
  28912=>"000110111",
  28913=>"110000010",
  28914=>"111110010",
  28915=>"011100001",
  28916=>"101000000",
  28917=>"010010000",
  28918=>"000010011",
  28919=>"101001010",
  28920=>"111011000",
  28921=>"101011110",
  28922=>"001101100",
  28923=>"001001101",
  28924=>"011101010",
  28925=>"001110101",
  28926=>"011000100",
  28927=>"111000101",
  28928=>"000011000",
  28929=>"011100101",
  28930=>"101101100",
  28931=>"010111000",
  28932=>"100110110",
  28933=>"001000010",
  28934=>"011001111",
  28935=>"010111001",
  28936=>"100101110",
  28937=>"000101100",
  28938=>"111000110",
  28939=>"110001011",
  28940=>"011011111",
  28941=>"010000100",
  28942=>"011001000",
  28943=>"010000101",
  28944=>"111111101",
  28945=>"111100111",
  28946=>"110100100",
  28947=>"001000010",
  28948=>"000100101",
  28949=>"010111111",
  28950=>"101000010",
  28951=>"101110010",
  28952=>"100100101",
  28953=>"110101010",
  28954=>"110111010",
  28955=>"011100100",
  28956=>"001110011",
  28957=>"111001010",
  28958=>"001000111",
  28959=>"010110010",
  28960=>"001111100",
  28961=>"101111000",
  28962=>"110100100",
  28963=>"010010010",
  28964=>"000000000",
  28965=>"010010100",
  28966=>"000000011",
  28967=>"010010000",
  28968=>"101100000",
  28969=>"011111000",
  28970=>"101011111",
  28971=>"111101111",
  28972=>"100010100",
  28973=>"100100101",
  28974=>"011111010",
  28975=>"001100101",
  28976=>"101000000",
  28977=>"110000110",
  28978=>"111101101",
  28979=>"100100011",
  28980=>"011000101",
  28981=>"101001100",
  28982=>"011110111",
  28983=>"001110000",
  28984=>"111111110",
  28985=>"000110111",
  28986=>"000011011",
  28987=>"001010000",
  28988=>"100111100",
  28989=>"101100111",
  28990=>"100000010",
  28991=>"111000001",
  28992=>"110011111",
  28993=>"110101010",
  28994=>"110000001",
  28995=>"011011011",
  28996=>"100100001",
  28997=>"100100011",
  28998=>"110000001",
  28999=>"110001000",
  29000=>"000010111",
  29001=>"110100110",
  29002=>"110010100",
  29003=>"011011000",
  29004=>"010001110",
  29005=>"111111000",
  29006=>"001111001",
  29007=>"011100101",
  29008=>"110000100",
  29009=>"101001010",
  29010=>"010011110",
  29011=>"111100000",
  29012=>"000100001",
  29013=>"110101101",
  29014=>"111100001",
  29015=>"000101111",
  29016=>"000111100",
  29017=>"110101101",
  29018=>"101010100",
  29019=>"110100101",
  29020=>"100110111",
  29021=>"100101110",
  29022=>"100110000",
  29023=>"011011101",
  29024=>"010101011",
  29025=>"100111110",
  29026=>"110000101",
  29027=>"000011111",
  29028=>"111011110",
  29029=>"111001001",
  29030=>"010000111",
  29031=>"111100010",
  29032=>"110011110",
  29033=>"001011111",
  29034=>"000100000",
  29035=>"111111110",
  29036=>"110100000",
  29037=>"001100101",
  29038=>"000010101",
  29039=>"001100010",
  29040=>"111101011",
  29041=>"100011010",
  29042=>"100011110",
  29043=>"011101011",
  29044=>"010000011",
  29045=>"111100001",
  29046=>"110110010",
  29047=>"101000111",
  29048=>"111000110",
  29049=>"001100000",
  29050=>"110101110",
  29051=>"111100011",
  29052=>"001111110",
  29053=>"010000101",
  29054=>"110100111",
  29055=>"100101010",
  29056=>"101011110",
  29057=>"110101011",
  29058=>"001101010",
  29059=>"111010110",
  29060=>"101001011",
  29061=>"010101101",
  29062=>"100100100",
  29063=>"001010011",
  29064=>"000010100",
  29065=>"101111011",
  29066=>"000010010",
  29067=>"001000111",
  29068=>"101011110",
  29069=>"011000001",
  29070=>"000100100",
  29071=>"110110011",
  29072=>"101001111",
  29073=>"001010111",
  29074=>"101000001",
  29075=>"110101000",
  29076=>"100110111",
  29077=>"110111010",
  29078=>"001110001",
  29079=>"110001000",
  29080=>"110010001",
  29081=>"101011000",
  29082=>"101101101",
  29083=>"001111000",
  29084=>"000100001",
  29085=>"010110111",
  29086=>"100001011",
  29087=>"100100111",
  29088=>"000010001",
  29089=>"101000110",
  29090=>"010110110",
  29091=>"000010010",
  29092=>"011001011",
  29093=>"101111100",
  29094=>"111000101",
  29095=>"001000001",
  29096=>"111110001",
  29097=>"001001011",
  29098=>"101000011",
  29099=>"110001001",
  29100=>"000100111",
  29101=>"010001011",
  29102=>"111100111",
  29103=>"110010011",
  29104=>"000000111",
  29105=>"000000111",
  29106=>"010010100",
  29107=>"111001001",
  29108=>"101011000",
  29109=>"101000100",
  29110=>"100100111",
  29111=>"000000100",
  29112=>"110111111",
  29113=>"110111101",
  29114=>"010110111",
  29115=>"111101100",
  29116=>"010010111",
  29117=>"010111111",
  29118=>"011100111",
  29119=>"011101011",
  29120=>"001010000",
  29121=>"001000101",
  29122=>"010100110",
  29123=>"110111010",
  29124=>"001110111",
  29125=>"000110111",
  29126=>"110001011",
  29127=>"100000110",
  29128=>"111110001",
  29129=>"010000111",
  29130=>"010010111",
  29131=>"111000110",
  29132=>"001100001",
  29133=>"110000100",
  29134=>"110011011",
  29135=>"111101010",
  29136=>"000000110",
  29137=>"011110111",
  29138=>"111101101",
  29139=>"101101010",
  29140=>"101110110",
  29141=>"101010111",
  29142=>"001011100",
  29143=>"110100010",
  29144=>"111101110",
  29145=>"000110011",
  29146=>"010110010",
  29147=>"000011100",
  29148=>"100110101",
  29149=>"111000010",
  29150=>"001111101",
  29151=>"110101110",
  29152=>"110100000",
  29153=>"110110101",
  29154=>"111001111",
  29155=>"011000101",
  29156=>"010010011",
  29157=>"101001011",
  29158=>"001011101",
  29159=>"000001010",
  29160=>"001010000",
  29161=>"111110101",
  29162=>"110101101",
  29163=>"101010010",
  29164=>"101100000",
  29165=>"100010000",
  29166=>"100101111",
  29167=>"111100000",
  29168=>"111111000",
  29169=>"001000110",
  29170=>"011001100",
  29171=>"110000111",
  29172=>"100011101",
  29173=>"001000001",
  29174=>"101100000",
  29175=>"010010001",
  29176=>"010110000",
  29177=>"001101000",
  29178=>"000100110",
  29179=>"000000010",
  29180=>"000101100",
  29181=>"110111000",
  29182=>"011001100",
  29183=>"101101010",
  29184=>"100000010",
  29185=>"100110100",
  29186=>"010000001",
  29187=>"001000100",
  29188=>"010010100",
  29189=>"000000111",
  29190=>"001100110",
  29191=>"011010101",
  29192=>"001000001",
  29193=>"101011110",
  29194=>"000100011",
  29195=>"001100110",
  29196=>"111110110",
  29197=>"001101111",
  29198=>"000101101",
  29199=>"010010000",
  29200=>"011100111",
  29201=>"011001100",
  29202=>"000001010",
  29203=>"000100100",
  29204=>"111001000",
  29205=>"001011011",
  29206=>"101011100",
  29207=>"100100110",
  29208=>"001000001",
  29209=>"011011111",
  29210=>"101110000",
  29211=>"001001011",
  29212=>"000001111",
  29213=>"010011011",
  29214=>"001000110",
  29215=>"010011001",
  29216=>"011111011",
  29217=>"101100111",
  29218=>"111001101",
  29219=>"011110010",
  29220=>"110000101",
  29221=>"001110100",
  29222=>"111110111",
  29223=>"110000001",
  29224=>"010001000",
  29225=>"101010100",
  29226=>"111011010",
  29227=>"011000101",
  29228=>"011111000",
  29229=>"111111000",
  29230=>"100101010",
  29231=>"000000100",
  29232=>"000110111",
  29233=>"000100101",
  29234=>"101110011",
  29235=>"111110110",
  29236=>"101100101",
  29237=>"111110111",
  29238=>"111100010",
  29239=>"101101110",
  29240=>"100000000",
  29241=>"011011101",
  29242=>"100010100",
  29243=>"100110001",
  29244=>"111111010",
  29245=>"100001001",
  29246=>"000010001",
  29247=>"000110000",
  29248=>"011010101",
  29249=>"001110011",
  29250=>"011011001",
  29251=>"100111001",
  29252=>"001010110",
  29253=>"011111000",
  29254=>"001000001",
  29255=>"011100010",
  29256=>"000111111",
  29257=>"010100001",
  29258=>"000010111",
  29259=>"000110111",
  29260=>"101110110",
  29261=>"110101111",
  29262=>"001000011",
  29263=>"000111001",
  29264=>"111101001",
  29265=>"100001110",
  29266=>"001101010",
  29267=>"000111110",
  29268=>"010011001",
  29269=>"111111111",
  29270=>"111010111",
  29271=>"000001111",
  29272=>"001010110",
  29273=>"101000001",
  29274=>"010000010",
  29275=>"000011101",
  29276=>"101111011",
  29277=>"110000010",
  29278=>"011010100",
  29279=>"010000110",
  29280=>"101111101",
  29281=>"011011111",
  29282=>"011001001",
  29283=>"110101110",
  29284=>"011110101",
  29285=>"110011100",
  29286=>"101000010",
  29287=>"110010110",
  29288=>"101111111",
  29289=>"001111111",
  29290=>"101000111",
  29291=>"100100011",
  29292=>"000100110",
  29293=>"010010111",
  29294=>"111100101",
  29295=>"000111000",
  29296=>"011101100",
  29297=>"011111111",
  29298=>"111010011",
  29299=>"111101110",
  29300=>"011010001",
  29301=>"110110100",
  29302=>"100001000",
  29303=>"010001010",
  29304=>"100011111",
  29305=>"111000010",
  29306=>"000000010",
  29307=>"110111010",
  29308=>"111001110",
  29309=>"111011000",
  29310=>"101011010",
  29311=>"110010110",
  29312=>"000001001",
  29313=>"010111011",
  29314=>"101001101",
  29315=>"100000001",
  29316=>"000111010",
  29317=>"110000100",
  29318=>"101001000",
  29319=>"110011011",
  29320=>"011111010",
  29321=>"011010110",
  29322=>"111100110",
  29323=>"101011010",
  29324=>"110000001",
  29325=>"010101100",
  29326=>"100011111",
  29327=>"100011000",
  29328=>"101010001",
  29329=>"111011011",
  29330=>"111101001",
  29331=>"111001100",
  29332=>"111100101",
  29333=>"111000101",
  29334=>"000101001",
  29335=>"010111000",
  29336=>"111110001",
  29337=>"011001001",
  29338=>"111101010",
  29339=>"100000010",
  29340=>"010001101",
  29341=>"000000001",
  29342=>"100100000",
  29343=>"011101101",
  29344=>"010101011",
  29345=>"110111000",
  29346=>"101110101",
  29347=>"011001010",
  29348=>"001001000",
  29349=>"011101101",
  29350=>"001101100",
  29351=>"101100010",
  29352=>"110001111",
  29353=>"000010101",
  29354=>"110100110",
  29355=>"010001000",
  29356=>"100101110",
  29357=>"101101011",
  29358=>"011010000",
  29359=>"011001000",
  29360=>"111110101",
  29361=>"100100111",
  29362=>"110000100",
  29363=>"111001101",
  29364=>"010110001",
  29365=>"010010011",
  29366=>"011110110",
  29367=>"010011000",
  29368=>"001011110",
  29369=>"001111000",
  29370=>"001110110",
  29371=>"011101000",
  29372=>"001101110",
  29373=>"001000011",
  29374=>"000001101",
  29375=>"110100100",
  29376=>"110000011",
  29377=>"011111101",
  29378=>"101111100",
  29379=>"110000011",
  29380=>"111110111",
  29381=>"001001111",
  29382=>"101001100",
  29383=>"111001111",
  29384=>"110101011",
  29385=>"000001001",
  29386=>"100011010",
  29387=>"100101101",
  29388=>"111011100",
  29389=>"111001001",
  29390=>"010101111",
  29391=>"110000101",
  29392=>"110111000",
  29393=>"011100011",
  29394=>"111100110",
  29395=>"000110011",
  29396=>"001111101",
  29397=>"001010111",
  29398=>"100101000",
  29399=>"000110111",
  29400=>"111111011",
  29401=>"110100111",
  29402=>"011000001",
  29403=>"010001011",
  29404=>"111010100",
  29405=>"010110100",
  29406=>"110110110",
  29407=>"100100011",
  29408=>"111111110",
  29409=>"101101011",
  29410=>"011111100",
  29411=>"100111100",
  29412=>"101111110",
  29413=>"000101010",
  29414=>"010011001",
  29415=>"000110010",
  29416=>"001001000",
  29417=>"010111000",
  29418=>"011101110",
  29419=>"000000011",
  29420=>"000011101",
  29421=>"010011010",
  29422=>"111010111",
  29423=>"010110101",
  29424=>"111110000",
  29425=>"110101001",
  29426=>"110010010",
  29427=>"110000010",
  29428=>"100111100",
  29429=>"111000100",
  29430=>"010100101",
  29431=>"011000101",
  29432=>"100011100",
  29433=>"001101101",
  29434=>"110100000",
  29435=>"001001001",
  29436=>"111110101",
  29437=>"011111001",
  29438=>"110011111",
  29439=>"101011111",
  29440=>"101001101",
  29441=>"001010111",
  29442=>"011110101",
  29443=>"010001001",
  29444=>"101100010",
  29445=>"101000000",
  29446=>"110101010",
  29447=>"110110101",
  29448=>"111101111",
  29449=>"001001011",
  29450=>"010011011",
  29451=>"101101001",
  29452=>"111100101",
  29453=>"110100101",
  29454=>"111101100",
  29455=>"000011111",
  29456=>"000110100",
  29457=>"001001011",
  29458=>"001011011",
  29459=>"010110001",
  29460=>"000010111",
  29461=>"000111111",
  29462=>"000001001",
  29463=>"000010000",
  29464=>"001001101",
  29465=>"101000101",
  29466=>"000011100",
  29467=>"110000010",
  29468=>"110111110",
  29469=>"110001011",
  29470=>"101001111",
  29471=>"110001010",
  29472=>"000101100",
  29473=>"110011001",
  29474=>"110010110",
  29475=>"111111001",
  29476=>"011000110",
  29477=>"010010110",
  29478=>"100011011",
  29479=>"101111000",
  29480=>"001101100",
  29481=>"100111011",
  29482=>"100001110",
  29483=>"101101110",
  29484=>"111101101",
  29485=>"111001001",
  29486=>"001111111",
  29487=>"000100011",
  29488=>"111111111",
  29489=>"111111010",
  29490=>"000110011",
  29491=>"000110111",
  29492=>"001000000",
  29493=>"111001011",
  29494=>"101100000",
  29495=>"010010101",
  29496=>"011011110",
  29497=>"100110001",
  29498=>"000010110",
  29499=>"011101101",
  29500=>"000100110",
  29501=>"001011101",
  29502=>"001111101",
  29503=>"101000010",
  29504=>"010000000",
  29505=>"101100001",
  29506=>"010111111",
  29507=>"100110101",
  29508=>"010000001",
  29509=>"111111110",
  29510=>"011100000",
  29511=>"101000011",
  29512=>"011011110",
  29513=>"000000001",
  29514=>"101111011",
  29515=>"010101101",
  29516=>"011010101",
  29517=>"101111000",
  29518=>"110001001",
  29519=>"010011001",
  29520=>"100110110",
  29521=>"010110110",
  29522=>"001000000",
  29523=>"000011001",
  29524=>"000101000",
  29525=>"110100011",
  29526=>"100110110",
  29527=>"010101110",
  29528=>"000111010",
  29529=>"011101010",
  29530=>"001101101",
  29531=>"111100100",
  29532=>"110111011",
  29533=>"000010001",
  29534=>"001111111",
  29535=>"111101001",
  29536=>"011000110",
  29537=>"000001101",
  29538=>"110111100",
  29539=>"010101100",
  29540=>"101100111",
  29541=>"001111000",
  29542=>"111100010",
  29543=>"000000001",
  29544=>"110110110",
  29545=>"110111011",
  29546=>"111110110",
  29547=>"011000100",
  29548=>"011001110",
  29549=>"011000010",
  29550=>"010101110",
  29551=>"100110111",
  29552=>"000010000",
  29553=>"110111110",
  29554=>"101110011",
  29555=>"001001011",
  29556=>"010100001",
  29557=>"000000001",
  29558=>"111001100",
  29559=>"011000000",
  29560=>"101001110",
  29561=>"010001001",
  29562=>"000010010",
  29563=>"101111010",
  29564=>"001011011",
  29565=>"001010011",
  29566=>"001111111",
  29567=>"010010111",
  29568=>"001110101",
  29569=>"011001011",
  29570=>"001000000",
  29571=>"100110100",
  29572=>"100000010",
  29573=>"000111011",
  29574=>"110111100",
  29575=>"001111010",
  29576=>"000101111",
  29577=>"000101000",
  29578=>"111101011",
  29579=>"010000011",
  29580=>"111110110",
  29581=>"110101111",
  29582=>"000000110",
  29583=>"010001010",
  29584=>"010101001",
  29585=>"011001110",
  29586=>"001111110",
  29587=>"101011001",
  29588=>"100110111",
  29589=>"000011000",
  29590=>"100101101",
  29591=>"000000110",
  29592=>"100111110",
  29593=>"001010011",
  29594=>"111100110",
  29595=>"001110101",
  29596=>"000011011",
  29597=>"001111111",
  29598=>"111000001",
  29599=>"010100001",
  29600=>"011111011",
  29601=>"100000000",
  29602=>"110110111",
  29603=>"111011000",
  29604=>"100001011",
  29605=>"010101111",
  29606=>"010100111",
  29607=>"101000001",
  29608=>"100101010",
  29609=>"111100111",
  29610=>"100001000",
  29611=>"100001010",
  29612=>"010011001",
  29613=>"101110001",
  29614=>"011110110",
  29615=>"100101111",
  29616=>"100110100",
  29617=>"110011101",
  29618=>"101011010",
  29619=>"010010010",
  29620=>"001101100",
  29621=>"110011101",
  29622=>"100010011",
  29623=>"010101011",
  29624=>"001001101",
  29625=>"000111001",
  29626=>"000010000",
  29627=>"111110000",
  29628=>"011101001",
  29629=>"101110011",
  29630=>"000100111",
  29631=>"000001010",
  29632=>"110111100",
  29633=>"100100100",
  29634=>"110110100",
  29635=>"100001000",
  29636=>"001101101",
  29637=>"011111100",
  29638=>"101000011",
  29639=>"111010101",
  29640=>"111111101",
  29641=>"010110100",
  29642=>"001100001",
  29643=>"100001011",
  29644=>"001101011",
  29645=>"000111100",
  29646=>"000100000",
  29647=>"111011011",
  29648=>"001111001",
  29649=>"010001001",
  29650=>"000000010",
  29651=>"000000111",
  29652=>"000000011",
  29653=>"111111010",
  29654=>"011001001",
  29655=>"111001010",
  29656=>"100100011",
  29657=>"110110100",
  29658=>"110101000",
  29659=>"111000000",
  29660=>"101000000",
  29661=>"010110000",
  29662=>"001001001",
  29663=>"010001100",
  29664=>"110100001",
  29665=>"001001010",
  29666=>"111100100",
  29667=>"001010111",
  29668=>"111110111",
  29669=>"000010010",
  29670=>"000001100",
  29671=>"000111110",
  29672=>"101001001",
  29673=>"100101010",
  29674=>"000111110",
  29675=>"000000111",
  29676=>"101011100",
  29677=>"011000101",
  29678=>"101110011",
  29679=>"011001011",
  29680=>"100000111",
  29681=>"010000000",
  29682=>"001110110",
  29683=>"111010110",
  29684=>"100001110",
  29685=>"000011111",
  29686=>"010100110",
  29687=>"111100001",
  29688=>"101001000",
  29689=>"001110001",
  29690=>"001100101",
  29691=>"100000101",
  29692=>"001010101",
  29693=>"010101111",
  29694=>"101111111",
  29695=>"101011001",
  29696=>"010011010",
  29697=>"101101111",
  29698=>"000100111",
  29699=>"111001010",
  29700=>"010010101",
  29701=>"101011001",
  29702=>"110000000",
  29703=>"111001000",
  29704=>"110100011",
  29705=>"010000101",
  29706=>"110000100",
  29707=>"110010011",
  29708=>"110000110",
  29709=>"100100100",
  29710=>"001111111",
  29711=>"000111011",
  29712=>"010100010",
  29713=>"001101100",
  29714=>"000011010",
  29715=>"110000001",
  29716=>"000000001",
  29717=>"101010101",
  29718=>"011100110",
  29719=>"100000001",
  29720=>"010100010",
  29721=>"000010000",
  29722=>"110010000",
  29723=>"111110100",
  29724=>"100000001",
  29725=>"100001000",
  29726=>"011000010",
  29727=>"010100110",
  29728=>"111111001",
  29729=>"110101010",
  29730=>"111000111",
  29731=>"100100000",
  29732=>"011010101",
  29733=>"100101100",
  29734=>"111100001",
  29735=>"000110000",
  29736=>"010101111",
  29737=>"101000101",
  29738=>"000101101",
  29739=>"001001111",
  29740=>"011010111",
  29741=>"111110111",
  29742=>"111000010",
  29743=>"100110111",
  29744=>"101101101",
  29745=>"010111110",
  29746=>"111110001",
  29747=>"010011101",
  29748=>"100101010",
  29749=>"100101101",
  29750=>"101111110",
  29751=>"111111111",
  29752=>"011110010",
  29753=>"001000011",
  29754=>"110000110",
  29755=>"111000101",
  29756=>"000100010",
  29757=>"000100000",
  29758=>"110000110",
  29759=>"100000111",
  29760=>"001111000",
  29761=>"100001111",
  29762=>"010010101",
  29763=>"011101000",
  29764=>"001010100",
  29765=>"111011010",
  29766=>"001110000",
  29767=>"010101111",
  29768=>"111000000",
  29769=>"001100000",
  29770=>"011101111",
  29771=>"111000010",
  29772=>"010011010",
  29773=>"011111111",
  29774=>"101100011",
  29775=>"011101011",
  29776=>"011100000",
  29777=>"010010101",
  29778=>"000011111",
  29779=>"001110001",
  29780=>"101001100",
  29781=>"000000010",
  29782=>"011011100",
  29783=>"100101000",
  29784=>"101100011",
  29785=>"101111010",
  29786=>"001000111",
  29787=>"010010011",
  29788=>"010000001",
  29789=>"100101010",
  29790=>"100001011",
  29791=>"100100100",
  29792=>"111000111",
  29793=>"100010000",
  29794=>"100000101",
  29795=>"111110110",
  29796=>"010100010",
  29797=>"110101010",
  29798=>"111111011",
  29799=>"001101111",
  29800=>"100111001",
  29801=>"111011111",
  29802=>"011001111",
  29803=>"000100001",
  29804=>"000000000",
  29805=>"001111110",
  29806=>"011011110",
  29807=>"010010101",
  29808=>"110110000",
  29809=>"001011001",
  29810=>"011001000",
  29811=>"110001101",
  29812=>"011000011",
  29813=>"000110010",
  29814=>"011010011",
  29815=>"110001110",
  29816=>"100101100",
  29817=>"111010011",
  29818=>"111110111",
  29819=>"011000000",
  29820=>"101100101",
  29821=>"000100000",
  29822=>"010001010",
  29823=>"000100001",
  29824=>"011010111",
  29825=>"100000010",
  29826=>"000101101",
  29827=>"010111011",
  29828=>"101110111",
  29829=>"110011010",
  29830=>"011011001",
  29831=>"011110001",
  29832=>"111011110",
  29833=>"001100111",
  29834=>"110011111",
  29835=>"111001010",
  29836=>"100000000",
  29837=>"011110100",
  29838=>"110110101",
  29839=>"011111110",
  29840=>"110101010",
  29841=>"110110000",
  29842=>"110111000",
  29843=>"110101111",
  29844=>"001010110",
  29845=>"110111001",
  29846=>"001000110",
  29847=>"010100111",
  29848=>"100100000",
  29849=>"100011111",
  29850=>"011101111",
  29851=>"100111010",
  29852=>"100111110",
  29853=>"110011011",
  29854=>"000010100",
  29855=>"010101010",
  29856=>"100000010",
  29857=>"100100000",
  29858=>"111010100",
  29859=>"101001101",
  29860=>"100001011",
  29861=>"000101000",
  29862=>"010010010",
  29863=>"100001001",
  29864=>"001110100",
  29865=>"100000111",
  29866=>"011110000",
  29867=>"011011010",
  29868=>"111111010",
  29869=>"101001000",
  29870=>"001100000",
  29871=>"011111010",
  29872=>"001010000",
  29873=>"011111100",
  29874=>"100000101",
  29875=>"000010010",
  29876=>"000100011",
  29877=>"101111000",
  29878=>"000000101",
  29879=>"111011111",
  29880=>"111001001",
  29881=>"111101011",
  29882=>"000110000",
  29883=>"001001110",
  29884=>"111110010",
  29885=>"011110010",
  29886=>"101101111",
  29887=>"110010010",
  29888=>"101111001",
  29889=>"010100000",
  29890=>"000100001",
  29891=>"011110001",
  29892=>"100011000",
  29893=>"100101010",
  29894=>"111001111",
  29895=>"111010101",
  29896=>"110110111",
  29897=>"110100000",
  29898=>"111111011",
  29899=>"001011010",
  29900=>"111000101",
  29901=>"100110100",
  29902=>"010110100",
  29903=>"000001010",
  29904=>"111001000",
  29905=>"000101101",
  29906=>"001010101",
  29907=>"101111000",
  29908=>"101010111",
  29909=>"001011011",
  29910=>"101011011",
  29911=>"001010010",
  29912=>"001110000",
  29913=>"001011001",
  29914=>"000111101",
  29915=>"101110101",
  29916=>"110100001",
  29917=>"011110000",
  29918=>"000111110",
  29919=>"101101111",
  29920=>"100001010",
  29921=>"000001010",
  29922=>"100011101",
  29923=>"000000011",
  29924=>"001111011",
  29925=>"000001001",
  29926=>"100100110",
  29927=>"011100010",
  29928=>"001110010",
  29929=>"101101010",
  29930=>"001101101",
  29931=>"101110111",
  29932=>"011001001",
  29933=>"100010110",
  29934=>"001001111",
  29935=>"010110000",
  29936=>"101101001",
  29937=>"100100010",
  29938=>"011110110",
  29939=>"011110011",
  29940=>"000110011",
  29941=>"011000100",
  29942=>"011101011",
  29943=>"100000001",
  29944=>"100000001",
  29945=>"100011101",
  29946=>"011001110",
  29947=>"101100010",
  29948=>"001100001",
  29949=>"100010000",
  29950=>"110011011",
  29951=>"000101111",
  29952=>"010011110",
  29953=>"000100010",
  29954=>"111101001",
  29955=>"011001000",
  29956=>"001110011",
  29957=>"110110000",
  29958=>"010010010",
  29959=>"000110011",
  29960=>"101111111",
  29961=>"011101000",
  29962=>"110011110",
  29963=>"111111001",
  29964=>"101011101",
  29965=>"000111011",
  29966=>"100100111",
  29967=>"000100110",
  29968=>"000110010",
  29969=>"111110111",
  29970=>"110111110",
  29971=>"101001101",
  29972=>"100101100",
  29973=>"011101001",
  29974=>"001011100",
  29975=>"100000000",
  29976=>"000110011",
  29977=>"110110011",
  29978=>"011111001",
  29979=>"010011000",
  29980=>"011011000",
  29981=>"010000001",
  29982=>"000010100",
  29983=>"001000111",
  29984=>"000010101",
  29985=>"101110100",
  29986=>"000011000",
  29987=>"010011101",
  29988=>"101110111",
  29989=>"111001000",
  29990=>"011101101",
  29991=>"101010011",
  29992=>"010010000",
  29993=>"001000000",
  29994=>"001111101",
  29995=>"101110010",
  29996=>"000100010",
  29997=>"111111111",
  29998=>"111010101",
  29999=>"101011000",
  30000=>"111100001",
  30001=>"101001001",
  30002=>"000001000",
  30003=>"000000100",
  30004=>"010010011",
  30005=>"010100000",
  30006=>"101001000",
  30007=>"100010011",
  30008=>"111101111",
  30009=>"001100110",
  30010=>"000101100",
  30011=>"000011000",
  30012=>"101110111",
  30013=>"111111011",
  30014=>"010101011",
  30015=>"110010001",
  30016=>"111001001",
  30017=>"101101101",
  30018=>"000101000",
  30019=>"011000011",
  30020=>"111110001",
  30021=>"001011001",
  30022=>"111000110",
  30023=>"001101010",
  30024=>"111010111",
  30025=>"100100100",
  30026=>"000100001",
  30027=>"000010100",
  30028=>"100010110",
  30029=>"111001010",
  30030=>"000101011",
  30031=>"101111101",
  30032=>"111010110",
  30033=>"110110011",
  30034=>"010001101",
  30035=>"100010101",
  30036=>"000011101",
  30037=>"010100001",
  30038=>"001011101",
  30039=>"100000101",
  30040=>"100001011",
  30041=>"000000000",
  30042=>"111101101",
  30043=>"100010010",
  30044=>"000001100",
  30045=>"000001111",
  30046=>"110100010",
  30047=>"110001001",
  30048=>"001010110",
  30049=>"010011110",
  30050=>"000000000",
  30051=>"010110001",
  30052=>"101111110",
  30053=>"011111111",
  30054=>"001101111",
  30055=>"101111100",
  30056=>"000111110",
  30057=>"000000101",
  30058=>"111011011",
  30059=>"010010110",
  30060=>"010101100",
  30061=>"000111101",
  30062=>"000101001",
  30063=>"001111101",
  30064=>"100000110",
  30065=>"100010100",
  30066=>"000010000",
  30067=>"101011001",
  30068=>"111110111",
  30069=>"010111110",
  30070=>"010000110",
  30071=>"110111001",
  30072=>"001000110",
  30073=>"100101000",
  30074=>"101001010",
  30075=>"011111011",
  30076=>"000111111",
  30077=>"110110010",
  30078=>"001111011",
  30079=>"111101111",
  30080=>"000111100",
  30081=>"010000000",
  30082=>"001000110",
  30083=>"100001101",
  30084=>"100000110",
  30085=>"111000100",
  30086=>"011111110",
  30087=>"110110101",
  30088=>"110010110",
  30089=>"101001000",
  30090=>"001011100",
  30091=>"001110101",
  30092=>"011011010",
  30093=>"100110111",
  30094=>"101001001",
  30095=>"001000010",
  30096=>"000110010",
  30097=>"110000101",
  30098=>"001011100",
  30099=>"100000010",
  30100=>"011101000",
  30101=>"100011110",
  30102=>"111001011",
  30103=>"111101011",
  30104=>"101010111",
  30105=>"001100111",
  30106=>"010011001",
  30107=>"000001001",
  30108=>"001010101",
  30109=>"101010011",
  30110=>"000110000",
  30111=>"000000100",
  30112=>"010110011",
  30113=>"111101110",
  30114=>"110110100",
  30115=>"111010011",
  30116=>"101001001",
  30117=>"111100010",
  30118=>"000101001",
  30119=>"001011000",
  30120=>"001100101",
  30121=>"111001011",
  30122=>"000010111",
  30123=>"101100111",
  30124=>"001011101",
  30125=>"011111001",
  30126=>"000011010",
  30127=>"111000101",
  30128=>"000001111",
  30129=>"111001101",
  30130=>"111111111",
  30131=>"110101101",
  30132=>"010000010",
  30133=>"111000000",
  30134=>"010000110",
  30135=>"010000101",
  30136=>"101000011",
  30137=>"000000111",
  30138=>"001000110",
  30139=>"111010001",
  30140=>"111100001",
  30141=>"111110110",
  30142=>"000010111",
  30143=>"011110100",
  30144=>"011100111",
  30145=>"000000000",
  30146=>"101001100",
  30147=>"001101100",
  30148=>"010100100",
  30149=>"011011101",
  30150=>"010100010",
  30151=>"010010100",
  30152=>"111111110",
  30153=>"010111011",
  30154=>"000001100",
  30155=>"000001000",
  30156=>"100000100",
  30157=>"001111000",
  30158=>"110111110",
  30159=>"001001110",
  30160=>"100111010",
  30161=>"010110101",
  30162=>"101110000",
  30163=>"011000100",
  30164=>"110010011",
  30165=>"110101011",
  30166=>"101110010",
  30167=>"110000000",
  30168=>"001011101",
  30169=>"001000011",
  30170=>"000010111",
  30171=>"101001101",
  30172=>"100011111",
  30173=>"101100011",
  30174=>"011101000",
  30175=>"101011000",
  30176=>"010011110",
  30177=>"011010111",
  30178=>"110101010",
  30179=>"010100100",
  30180=>"111100000",
  30181=>"111001011",
  30182=>"000100100",
  30183=>"000010111",
  30184=>"110001111",
  30185=>"011001110",
  30186=>"111011100",
  30187=>"111001010",
  30188=>"111110001",
  30189=>"011110000",
  30190=>"111101110",
  30191=>"101100110",
  30192=>"000100101",
  30193=>"011111010",
  30194=>"010100011",
  30195=>"110111110",
  30196=>"000111111",
  30197=>"000100100",
  30198=>"000101011",
  30199=>"100011111",
  30200=>"010000000",
  30201=>"101110100",
  30202=>"000001011",
  30203=>"000110000",
  30204=>"010010110",
  30205=>"000110001",
  30206=>"000110011",
  30207=>"110101000",
  30208=>"010000010",
  30209=>"000101101",
  30210=>"101110100",
  30211=>"000000000",
  30212=>"110010111",
  30213=>"000101011",
  30214=>"110100010",
  30215=>"101111001",
  30216=>"101010111",
  30217=>"100010111",
  30218=>"110100100",
  30219=>"100110010",
  30220=>"111101001",
  30221=>"010001000",
  30222=>"000110010",
  30223=>"000101011",
  30224=>"111111000",
  30225=>"011001001",
  30226=>"100010101",
  30227=>"111101110",
  30228=>"101000001",
  30229=>"111011110",
  30230=>"011100011",
  30231=>"110000100",
  30232=>"110010001",
  30233=>"101100101",
  30234=>"001100101",
  30235=>"110110010",
  30236=>"101011111",
  30237=>"001100010",
  30238=>"101111111",
  30239=>"111111000",
  30240=>"101101100",
  30241=>"111100000",
  30242=>"110010100",
  30243=>"010110001",
  30244=>"000011011",
  30245=>"011101100",
  30246=>"001010101",
  30247=>"000010000",
  30248=>"001111011",
  30249=>"000100111",
  30250=>"110110110",
  30251=>"100100000",
  30252=>"101110110",
  30253=>"000001010",
  30254=>"000111010",
  30255=>"110111101",
  30256=>"101011010",
  30257=>"001110010",
  30258=>"111111111",
  30259=>"101111001",
  30260=>"010010000",
  30261=>"001101111",
  30262=>"000110000",
  30263=>"111110010",
  30264=>"111101110",
  30265=>"001001011",
  30266=>"100011100",
  30267=>"111000101",
  30268=>"010001110",
  30269=>"010010111",
  30270=>"000010010",
  30271=>"000010111",
  30272=>"011000000",
  30273=>"100101010",
  30274=>"011001011",
  30275=>"000001110",
  30276=>"101001011",
  30277=>"100000110",
  30278=>"110001111",
  30279=>"000001001",
  30280=>"111010011",
  30281=>"010000111",
  30282=>"001010000",
  30283=>"001001110",
  30284=>"110101110",
  30285=>"001110111",
  30286=>"100011111",
  30287=>"100000010",
  30288=>"111111110",
  30289=>"101110111",
  30290=>"111000100",
  30291=>"010100111",
  30292=>"000010000",
  30293=>"111100100",
  30294=>"100000010",
  30295=>"001010011",
  30296=>"100110100",
  30297=>"111111101",
  30298=>"010011010",
  30299=>"000000111",
  30300=>"101000110",
  30301=>"010111001",
  30302=>"110101011",
  30303=>"011011111",
  30304=>"001101100",
  30305=>"101101000",
  30306=>"001000101",
  30307=>"101101000",
  30308=>"110111101",
  30309=>"000110011",
  30310=>"110101000",
  30311=>"010010101",
  30312=>"101110100",
  30313=>"100100001",
  30314=>"100100011",
  30315=>"111000101",
  30316=>"110011011",
  30317=>"011100000",
  30318=>"100011010",
  30319=>"100100111",
  30320=>"001100110",
  30321=>"101000011",
  30322=>"101110000",
  30323=>"010010110",
  30324=>"111111010",
  30325=>"100100001",
  30326=>"000001001",
  30327=>"101101010",
  30328=>"001011001",
  30329=>"110000101",
  30330=>"101110010",
  30331=>"101001100",
  30332=>"011000101",
  30333=>"111101111",
  30334=>"000101001",
  30335=>"010010011",
  30336=>"101000100",
  30337=>"110100101",
  30338=>"111001110",
  30339=>"101001010",
  30340=>"011011100",
  30341=>"100010000",
  30342=>"111001111",
  30343=>"100110011",
  30344=>"000000011",
  30345=>"001111101",
  30346=>"001000111",
  30347=>"101110111",
  30348=>"000101101",
  30349=>"011011011",
  30350=>"011010000",
  30351=>"001000101",
  30352=>"001001111",
  30353=>"101110110",
  30354=>"010001000",
  30355=>"001001010",
  30356=>"000110011",
  30357=>"101111001",
  30358=>"010100001",
  30359=>"101100110",
  30360=>"101110111",
  30361=>"110011101",
  30362=>"001100101",
  30363=>"110111100",
  30364=>"001000000",
  30365=>"101100101",
  30366=>"111001000",
  30367=>"101000001",
  30368=>"110000001",
  30369=>"111000000",
  30370=>"111111000",
  30371=>"100001110",
  30372=>"000110101",
  30373=>"010001111",
  30374=>"101111001",
  30375=>"100000100",
  30376=>"101100111",
  30377=>"010001111",
  30378=>"111010101",
  30379=>"010110110",
  30380=>"100000110",
  30381=>"010100110",
  30382=>"110010011",
  30383=>"110000111",
  30384=>"000111010",
  30385=>"001100010",
  30386=>"000100001",
  30387=>"001001111",
  30388=>"010011000",
  30389=>"110110010",
  30390=>"011001000",
  30391=>"011001110",
  30392=>"101010010",
  30393=>"111000111",
  30394=>"100100111",
  30395=>"010111110",
  30396=>"001010000",
  30397=>"011001000",
  30398=>"011100101",
  30399=>"000110000",
  30400=>"111010001",
  30401=>"010010111",
  30402=>"100010010",
  30403=>"000111011",
  30404=>"111010110",
  30405=>"011110000",
  30406=>"001011100",
  30407=>"010011101",
  30408=>"011010010",
  30409=>"011111100",
  30410=>"011100100",
  30411=>"100101010",
  30412=>"000111001",
  30413=>"011011011",
  30414=>"110100111",
  30415=>"101001010",
  30416=>"100000010",
  30417=>"111100101",
  30418=>"001111000",
  30419=>"111001110",
  30420=>"111111110",
  30421=>"110110110",
  30422=>"010110011",
  30423=>"000001111",
  30424=>"100101011",
  30425=>"000110101",
  30426=>"111010010",
  30427=>"011110000",
  30428=>"000011100",
  30429=>"101101010",
  30430=>"000000001",
  30431=>"000111100",
  30432=>"110010101",
  30433=>"010101011",
  30434=>"000011000",
  30435=>"100010010",
  30436=>"111001101",
  30437=>"000011110",
  30438=>"101011100",
  30439=>"000001010",
  30440=>"000011100",
  30441=>"010011110",
  30442=>"111101010",
  30443=>"001010110",
  30444=>"000000110",
  30445=>"001110010",
  30446=>"010010001",
  30447=>"000010100",
  30448=>"000011000",
  30449=>"001111000",
  30450=>"101011101",
  30451=>"001110011",
  30452=>"111000011",
  30453=>"110000111",
  30454=>"110110111",
  30455=>"101001101",
  30456=>"110100101",
  30457=>"001001011",
  30458=>"000000001",
  30459=>"100101011",
  30460=>"110101001",
  30461=>"111100000",
  30462=>"001011111",
  30463=>"101011001",
  30464=>"110110011",
  30465=>"000101111",
  30466=>"111001000",
  30467=>"010111011",
  30468=>"110001101",
  30469=>"011000110",
  30470=>"111011010",
  30471=>"011101011",
  30472=>"100111110",
  30473=>"011111111",
  30474=>"011000001",
  30475=>"001000111",
  30476=>"001110101",
  30477=>"010110001",
  30478=>"101101011",
  30479=>"001010011",
  30480=>"011000110",
  30481=>"000111000",
  30482=>"111100110",
  30483=>"111101011",
  30484=>"111111110",
  30485=>"011010011",
  30486=>"100010100",
  30487=>"110011001",
  30488=>"110010101",
  30489=>"010110010",
  30490=>"000001111",
  30491=>"111101111",
  30492=>"101111000",
  30493=>"101100010",
  30494=>"001000111",
  30495=>"001101110",
  30496=>"011011110",
  30497=>"000110111",
  30498=>"100110010",
  30499=>"011110011",
  30500=>"010010001",
  30501=>"111101111",
  30502=>"100001010",
  30503=>"011001101",
  30504=>"010010100",
  30505=>"100000101",
  30506=>"011000101",
  30507=>"011111100",
  30508=>"010110111",
  30509=>"110010100",
  30510=>"011101111",
  30511=>"011111001",
  30512=>"000010010",
  30513=>"101111001",
  30514=>"001101001",
  30515=>"010001100",
  30516=>"001100010",
  30517=>"010000101",
  30518=>"110111111",
  30519=>"010000010",
  30520=>"111111000",
  30521=>"110001101",
  30522=>"011001011",
  30523=>"000100110",
  30524=>"100110101",
  30525=>"101001001",
  30526=>"001111011",
  30527=>"111100010",
  30528=>"010110101",
  30529=>"110111110",
  30530=>"001000110",
  30531=>"011011110",
  30532=>"010100101",
  30533=>"000000000",
  30534=>"101100110",
  30535=>"100100001",
  30536=>"101010101",
  30537=>"010000101",
  30538=>"000101001",
  30539=>"011111100",
  30540=>"011001110",
  30541=>"111010110",
  30542=>"010101100",
  30543=>"101001101",
  30544=>"000010110",
  30545=>"101111010",
  30546=>"100000000",
  30547=>"101100010",
  30548=>"000001000",
  30549=>"111100100",
  30550=>"111001111",
  30551=>"000011110",
  30552=>"101100110",
  30553=>"111000100",
  30554=>"000001100",
  30555=>"111101000",
  30556=>"110010111",
  30557=>"011010100",
  30558=>"011101100",
  30559=>"010000000",
  30560=>"000110100",
  30561=>"110000010",
  30562=>"000011111",
  30563=>"110001111",
  30564=>"011100011",
  30565=>"011010001",
  30566=>"111100011",
  30567=>"100001010",
  30568=>"000111001",
  30569=>"000001110",
  30570=>"010111001",
  30571=>"111110101",
  30572=>"111111101",
  30573=>"000010010",
  30574=>"110100011",
  30575=>"110000010",
  30576=>"100001100",
  30577=>"111011100",
  30578=>"111100101",
  30579=>"011100000",
  30580=>"111000001",
  30581=>"001011111",
  30582=>"001001010",
  30583=>"011110111",
  30584=>"100100100",
  30585=>"000101010",
  30586=>"111001100",
  30587=>"000100100",
  30588=>"011001110",
  30589=>"101101110",
  30590=>"010111100",
  30591=>"101000000",
  30592=>"110101101",
  30593=>"110110101",
  30594=>"111110010",
  30595=>"101000101",
  30596=>"011010000",
  30597=>"101111010",
  30598=>"000011001",
  30599=>"111011110",
  30600=>"111000111",
  30601=>"010000100",
  30602=>"111000000",
  30603=>"000111010",
  30604=>"111111101",
  30605=>"000010011",
  30606=>"101111100",
  30607=>"110101011",
  30608=>"010101110",
  30609=>"110101011",
  30610=>"000110001",
  30611=>"011110010",
  30612=>"111111101",
  30613=>"000111010",
  30614=>"110001101",
  30615=>"000111101",
  30616=>"000010100",
  30617=>"100110110",
  30618=>"000000100",
  30619=>"111000010",
  30620=>"101001001",
  30621=>"011101110",
  30622=>"001111001",
  30623=>"111101001",
  30624=>"010110000",
  30625=>"001110101",
  30626=>"000010111",
  30627=>"111111011",
  30628=>"010100101",
  30629=>"011010010",
  30630=>"100100000",
  30631=>"011101011",
  30632=>"011101111",
  30633=>"000000001",
  30634=>"010110010",
  30635=>"111101011",
  30636=>"010001100",
  30637=>"000011111",
  30638=>"111111011",
  30639=>"001100101",
  30640=>"101100101",
  30641=>"110100110",
  30642=>"011111100",
  30643=>"101001000",
  30644=>"100100010",
  30645=>"000111101",
  30646=>"100100110",
  30647=>"000001101",
  30648=>"101011110",
  30649=>"000110010",
  30650=>"100001101",
  30651=>"111010001",
  30652=>"010101111",
  30653=>"010010010",
  30654=>"010000000",
  30655=>"010011000",
  30656=>"001001000",
  30657=>"100000000",
  30658=>"101111110",
  30659=>"101100101",
  30660=>"110010110",
  30661=>"101110001",
  30662=>"100110011",
  30663=>"101110100",
  30664=>"010101110",
  30665=>"001111011",
  30666=>"100111011",
  30667=>"111111011",
  30668=>"011001000",
  30669=>"110100000",
  30670=>"101110110",
  30671=>"000101000",
  30672=>"110001000",
  30673=>"100000110",
  30674=>"010010010",
  30675=>"101101100",
  30676=>"101011100",
  30677=>"110001010",
  30678=>"011111111",
  30679=>"010111111",
  30680=>"011010011",
  30681=>"100111001",
  30682=>"101010010",
  30683=>"110000100",
  30684=>"010010010",
  30685=>"000011001",
  30686=>"110101011",
  30687=>"100111010",
  30688=>"100110101",
  30689=>"100111111",
  30690=>"011010111",
  30691=>"010100111",
  30692=>"001100010",
  30693=>"100010000",
  30694=>"001100011",
  30695=>"000011000",
  30696=>"100100000",
  30697=>"010011011",
  30698=>"110001110",
  30699=>"001100111",
  30700=>"000101111",
  30701=>"011111001",
  30702=>"011000000",
  30703=>"000101110",
  30704=>"111101101",
  30705=>"011010001",
  30706=>"001101100",
  30707=>"000010001",
  30708=>"000100011",
  30709=>"110000011",
  30710=>"001101111",
  30711=>"001101000",
  30712=>"000001010",
  30713=>"100000010",
  30714=>"000100101",
  30715=>"011100101",
  30716=>"001101011",
  30717=>"110001000",
  30718=>"110000100",
  30719=>"100010010",
  30720=>"101001000",
  30721=>"010000111",
  30722=>"011011101",
  30723=>"001000000",
  30724=>"001001110",
  30725=>"101110000",
  30726=>"001001100",
  30727=>"010011000",
  30728=>"011110000",
  30729=>"000100010",
  30730=>"111010100",
  30731=>"000110001",
  30732=>"110011010",
  30733=>"011111111",
  30734=>"101010011",
  30735=>"001100000",
  30736=>"001100111",
  30737=>"111100100",
  30738=>"111101001",
  30739=>"110001111",
  30740=>"011000000",
  30741=>"011111001",
  30742=>"111100100",
  30743=>"000110000",
  30744=>"100000011",
  30745=>"100001010",
  30746=>"011111011",
  30747=>"001000101",
  30748=>"101101001",
  30749=>"111010110",
  30750=>"110001000",
  30751=>"100001010",
  30752=>"001010111",
  30753=>"011100100",
  30754=>"111100010",
  30755=>"001001101",
  30756=>"101100000",
  30757=>"100011010",
  30758=>"010000001",
  30759=>"001000010",
  30760=>"000001000",
  30761=>"010110100",
  30762=>"001110010",
  30763=>"110000001",
  30764=>"101011100",
  30765=>"110111100",
  30766=>"100100000",
  30767=>"001100111",
  30768=>"001101001",
  30769=>"010010010",
  30770=>"011100011",
  30771=>"011001100",
  30772=>"110001001",
  30773=>"100011100",
  30774=>"011101100",
  30775=>"100110100",
  30776=>"101010000",
  30777=>"011000001",
  30778=>"010000010",
  30779=>"100000101",
  30780=>"100110100",
  30781=>"101100011",
  30782=>"101000110",
  30783=>"000101101",
  30784=>"011110101",
  30785=>"000110011",
  30786=>"010010010",
  30787=>"101011000",
  30788=>"010110011",
  30789=>"111000100",
  30790=>"000110101",
  30791=>"000001001",
  30792=>"100000010",
  30793=>"111110100",
  30794=>"000000011",
  30795=>"000110001",
  30796=>"000101101",
  30797=>"100110011",
  30798=>"110001000",
  30799=>"101010011",
  30800=>"001100101",
  30801=>"000010000",
  30802=>"111101011",
  30803=>"010001011",
  30804=>"010011111",
  30805=>"111100011",
  30806=>"110001101",
  30807=>"011010110",
  30808=>"000001110",
  30809=>"011011000",
  30810=>"011000100",
  30811=>"000000100",
  30812=>"100110101",
  30813=>"000010101",
  30814=>"000000011",
  30815=>"000001011",
  30816=>"101110101",
  30817=>"110001001",
  30818=>"001000111",
  30819=>"000010011",
  30820=>"000000001",
  30821=>"010001101",
  30822=>"000011010",
  30823=>"010001001",
  30824=>"100000000",
  30825=>"001010111",
  30826=>"000000100",
  30827=>"011111100",
  30828=>"001010000",
  30829=>"001111001",
  30830=>"000110001",
  30831=>"000000110",
  30832=>"010000001",
  30833=>"110110001",
  30834=>"010000010",
  30835=>"001111110",
  30836=>"001010000",
  30837=>"001011011",
  30838=>"100111001",
  30839=>"001100010",
  30840=>"001100010",
  30841=>"001010101",
  30842=>"101010111",
  30843=>"010100010",
  30844=>"101110101",
  30845=>"110011100",
  30846=>"101000100",
  30847=>"011010000",
  30848=>"100000001",
  30849=>"101111000",
  30850=>"100000010",
  30851=>"001101111",
  30852=>"111000001",
  30853=>"001011000",
  30854=>"010101011",
  30855=>"000000111",
  30856=>"001100110",
  30857=>"110010000",
  30858=>"010001100",
  30859=>"100000000",
  30860=>"100110111",
  30861=>"100101000",
  30862=>"010011110",
  30863=>"011101001",
  30864=>"010101010",
  30865=>"000000110",
  30866=>"010100001",
  30867=>"001101001",
  30868=>"111111011",
  30869=>"110100110",
  30870=>"100000011",
  30871=>"100111010",
  30872=>"010011110",
  30873=>"101101011",
  30874=>"001001011",
  30875=>"010000000",
  30876=>"011011010",
  30877=>"110001011",
  30878=>"011110001",
  30879=>"011000011",
  30880=>"001000111",
  30881=>"100110000",
  30882=>"111010100",
  30883=>"100001000",
  30884=>"100111000",
  30885=>"101111010",
  30886=>"000100010",
  30887=>"101001011",
  30888=>"101101001",
  30889=>"100011100",
  30890=>"100000011",
  30891=>"111001100",
  30892=>"110001110",
  30893=>"101111000",
  30894=>"001010101",
  30895=>"000001110",
  30896=>"001101001",
  30897=>"000110010",
  30898=>"111010100",
  30899=>"010100111",
  30900=>"101010001",
  30901=>"101010100",
  30902=>"001111111",
  30903=>"001000011",
  30904=>"000000110",
  30905=>"011111001",
  30906=>"000001000",
  30907=>"011010001",
  30908=>"100001101",
  30909=>"111000000",
  30910=>"001011011",
  30911=>"000110000",
  30912=>"100010010",
  30913=>"010111000",
  30914=>"000110010",
  30915=>"010100010",
  30916=>"001011101",
  30917=>"011100111",
  30918=>"110001010",
  30919=>"110100101",
  30920=>"111001011",
  30921=>"000101100",
  30922=>"101101011",
  30923=>"010110110",
  30924=>"010011110",
  30925=>"011001001",
  30926=>"101001000",
  30927=>"110000000",
  30928=>"111000000",
  30929=>"000000010",
  30930=>"101000001",
  30931=>"101101001",
  30932=>"000001110",
  30933=>"101011001",
  30934=>"110011000",
  30935=>"111101111",
  30936=>"000000110",
  30937=>"111101000",
  30938=>"000000000",
  30939=>"011110011",
  30940=>"010100001",
  30941=>"110011100",
  30942=>"000001101",
  30943=>"001110111",
  30944=>"010111011",
  30945=>"011011010",
  30946=>"011110111",
  30947=>"101001100",
  30948=>"000100000",
  30949=>"000101000",
  30950=>"010000110",
  30951=>"001110111",
  30952=>"000000101",
  30953=>"011101111",
  30954=>"000111100",
  30955=>"111001110",
  30956=>"100001001",
  30957=>"100101000",
  30958=>"011011001",
  30959=>"011111110",
  30960=>"101001110",
  30961=>"001100110",
  30962=>"010001111",
  30963=>"000110110",
  30964=>"111111111",
  30965=>"111010000",
  30966=>"011010101",
  30967=>"110110000",
  30968=>"111110010",
  30969=>"101001010",
  30970=>"000000111",
  30971=>"110000001",
  30972=>"011101010",
  30973=>"101011111",
  30974=>"011110011",
  30975=>"000001110",
  30976=>"101101001",
  30977=>"110111010",
  30978=>"101100100",
  30979=>"000010001",
  30980=>"001001101",
  30981=>"101011010",
  30982=>"000110100",
  30983=>"001100011",
  30984=>"010100000",
  30985=>"001010011",
  30986=>"001001110",
  30987=>"100110110",
  30988=>"010001101",
  30989=>"110110001",
  30990=>"011010111",
  30991=>"110111010",
  30992=>"010100110",
  30993=>"000100110",
  30994=>"101010011",
  30995=>"000001110",
  30996=>"100110110",
  30997=>"000000100",
  30998=>"011100000",
  30999=>"001000000",
  31000=>"101000000",
  31001=>"101101001",
  31002=>"000101111",
  31003=>"000010010",
  31004=>"001000100",
  31005=>"011110001",
  31006=>"011001001",
  31007=>"000001001",
  31008=>"001110111",
  31009=>"110111011",
  31010=>"010101010",
  31011=>"011100001",
  31012=>"010110001",
  31013=>"111111010",
  31014=>"101101101",
  31015=>"110111110",
  31016=>"111110110",
  31017=>"111111011",
  31018=>"101101111",
  31019=>"101000100",
  31020=>"111101110",
  31021=>"100001010",
  31022=>"110110110",
  31023=>"001000001",
  31024=>"111111111",
  31025=>"101111000",
  31026=>"111111000",
  31027=>"100100001",
  31028=>"111101001",
  31029=>"011001011",
  31030=>"101010000",
  31031=>"000010011",
  31032=>"111101111",
  31033=>"111011110",
  31034=>"001010011",
  31035=>"110000000",
  31036=>"100111001",
  31037=>"101000101",
  31038=>"000110000",
  31039=>"000101110",
  31040=>"100100100",
  31041=>"100110111",
  31042=>"001010010",
  31043=>"010000100",
  31044=>"011010001",
  31045=>"011000110",
  31046=>"011000000",
  31047=>"000110000",
  31048=>"000100110",
  31049=>"111011101",
  31050=>"000111000",
  31051=>"000011110",
  31052=>"101001100",
  31053=>"000000000",
  31054=>"100001101",
  31055=>"011100110",
  31056=>"011000101",
  31057=>"001001100",
  31058=>"000000101",
  31059=>"100000010",
  31060=>"001100010",
  31061=>"001011110",
  31062=>"001111111",
  31063=>"111001000",
  31064=>"000100101",
  31065=>"111111111",
  31066=>"011101011",
  31067=>"001110111",
  31068=>"001101001",
  31069=>"000010011",
  31070=>"100111000",
  31071=>"101111111",
  31072=>"011100011",
  31073=>"010001110",
  31074=>"011101110",
  31075=>"000110111",
  31076=>"101110011",
  31077=>"111111100",
  31078=>"001110011",
  31079=>"111111000",
  31080=>"001100001",
  31081=>"011000010",
  31082=>"110011100",
  31083=>"011111011",
  31084=>"100011001",
  31085=>"011000010",
  31086=>"110000011",
  31087=>"111010001",
  31088=>"000111000",
  31089=>"100101001",
  31090=>"010000011",
  31091=>"001000111",
  31092=>"101100110",
  31093=>"000010101",
  31094=>"100110010",
  31095=>"110000010",
  31096=>"110101010",
  31097=>"010100100",
  31098=>"100001001",
  31099=>"111101011",
  31100=>"111010010",
  31101=>"100101001",
  31102=>"110101001",
  31103=>"100100110",
  31104=>"011011011",
  31105=>"000101110",
  31106=>"110111110",
  31107=>"101100000",
  31108=>"011110010",
  31109=>"001001101",
  31110=>"111001101",
  31111=>"011010110",
  31112=>"101010011",
  31113=>"001100001",
  31114=>"101001011",
  31115=>"111111101",
  31116=>"100111110",
  31117=>"010111110",
  31118=>"110011101",
  31119=>"001010011",
  31120=>"010011110",
  31121=>"011101110",
  31122=>"000000000",
  31123=>"010111101",
  31124=>"101100101",
  31125=>"010001011",
  31126=>"000001011",
  31127=>"011001111",
  31128=>"111000111",
  31129=>"111111100",
  31130=>"101011011",
  31131=>"000000110",
  31132=>"011001011",
  31133=>"010000000",
  31134=>"100000010",
  31135=>"111101111",
  31136=>"011001011",
  31137=>"110101110",
  31138=>"000111100",
  31139=>"001001010",
  31140=>"111100000",
  31141=>"100000011",
  31142=>"010010000",
  31143=>"001001100",
  31144=>"110011111",
  31145=>"111100000",
  31146=>"110101100",
  31147=>"111110000",
  31148=>"111011101",
  31149=>"110010000",
  31150=>"001110110",
  31151=>"010001100",
  31152=>"011011010",
  31153=>"100111000",
  31154=>"101100010",
  31155=>"111001011",
  31156=>"000011111",
  31157=>"100010011",
  31158=>"111011101",
  31159=>"000100010",
  31160=>"111101011",
  31161=>"011001000",
  31162=>"110101100",
  31163=>"011011110",
  31164=>"111010110",
  31165=>"001010101",
  31166=>"011110100",
  31167=>"010110111",
  31168=>"000001111",
  31169=>"001111001",
  31170=>"110100011",
  31171=>"010110001",
  31172=>"100110001",
  31173=>"111001100",
  31174=>"001111101",
  31175=>"000100001",
  31176=>"000101110",
  31177=>"101110101",
  31178=>"100011010",
  31179=>"110111110",
  31180=>"111001001",
  31181=>"000001110",
  31182=>"111111100",
  31183=>"101100110",
  31184=>"011000110",
  31185=>"010000001",
  31186=>"000111011",
  31187=>"101110111",
  31188=>"101100011",
  31189=>"101100101",
  31190=>"001011101",
  31191=>"000100011",
  31192=>"101011010",
  31193=>"000000010",
  31194=>"001010100",
  31195=>"010000100",
  31196=>"111111111",
  31197=>"000111000",
  31198=>"111111111",
  31199=>"110001101",
  31200=>"110011101",
  31201=>"001110000",
  31202=>"111110100",
  31203=>"101010101",
  31204=>"010100110",
  31205=>"111101111",
  31206=>"011101011",
  31207=>"000001000",
  31208=>"010111111",
  31209=>"111010101",
  31210=>"110010011",
  31211=>"111100100",
  31212=>"101100011",
  31213=>"110110011",
  31214=>"101011000",
  31215=>"000101000",
  31216=>"100011010",
  31217=>"010000010",
  31218=>"101110000",
  31219=>"000000101",
  31220=>"011000100",
  31221=>"010100001",
  31222=>"111011011",
  31223=>"011011101",
  31224=>"010001010",
  31225=>"001010100",
  31226=>"101000010",
  31227=>"101101011",
  31228=>"111000100",
  31229=>"100011101",
  31230=>"000101001",
  31231=>"100000001",
  31232=>"111011001",
  31233=>"111101110",
  31234=>"010000111",
  31235=>"101011010",
  31236=>"101010011",
  31237=>"000110111",
  31238=>"001101100",
  31239=>"000000110",
  31240=>"001100011",
  31241=>"100011110",
  31242=>"000110110",
  31243=>"100111110",
  31244=>"101110100",
  31245=>"101101001",
  31246=>"000100000",
  31247=>"011010100",
  31248=>"010011010",
  31249=>"010101100",
  31250=>"111111110",
  31251=>"100110001",
  31252=>"110010111",
  31253=>"100011101",
  31254=>"001010100",
  31255=>"111110011",
  31256=>"111001100",
  31257=>"111000011",
  31258=>"001100011",
  31259=>"101010000",
  31260=>"011111100",
  31261=>"101100100",
  31262=>"110000011",
  31263=>"010100101",
  31264=>"001000000",
  31265=>"011001111",
  31266=>"110100101",
  31267=>"111001011",
  31268=>"010111101",
  31269=>"001101011",
  31270=>"001100010",
  31271=>"011000000",
  31272=>"110111101",
  31273=>"011111000",
  31274=>"111011001",
  31275=>"101100000",
  31276=>"000011100",
  31277=>"111101001",
  31278=>"101000000",
  31279=>"000000001",
  31280=>"101011001",
  31281=>"110001010",
  31282=>"010101000",
  31283=>"000001000",
  31284=>"101110101",
  31285=>"111110011",
  31286=>"101110010",
  31287=>"010111001",
  31288=>"101100110",
  31289=>"100010010",
  31290=>"011011100",
  31291=>"111000010",
  31292=>"010110111",
  31293=>"010001010",
  31294=>"010100000",
  31295=>"111100111",
  31296=>"011111011",
  31297=>"100000111",
  31298=>"100011111",
  31299=>"101110011",
  31300=>"011000100",
  31301=>"001110100",
  31302=>"110110011",
  31303=>"000000000",
  31304=>"001101101",
  31305=>"101111011",
  31306=>"000010000",
  31307=>"000110000",
  31308=>"100010010",
  31309=>"011011001",
  31310=>"101100000",
  31311=>"111101011",
  31312=>"100100111",
  31313=>"100010101",
  31314=>"111000101",
  31315=>"100111110",
  31316=>"001001000",
  31317=>"111011110",
  31318=>"110101011",
  31319=>"111101100",
  31320=>"010100100",
  31321=>"001001110",
  31322=>"010011100",
  31323=>"100110101",
  31324=>"000000000",
  31325=>"101111011",
  31326=>"001000111",
  31327=>"110110101",
  31328=>"101110111",
  31329=>"100001100",
  31330=>"010111101",
  31331=>"001010011",
  31332=>"111011001",
  31333=>"110110100",
  31334=>"101001010",
  31335=>"010000000",
  31336=>"101100011",
  31337=>"001010100",
  31338=>"011101000",
  31339=>"001101100",
  31340=>"110011001",
  31341=>"111100001",
  31342=>"100001110",
  31343=>"000101111",
  31344=>"001110011",
  31345=>"111111111",
  31346=>"011001011",
  31347=>"001111101",
  31348=>"000101111",
  31349=>"001000010",
  31350=>"000111110",
  31351=>"000101100",
  31352=>"110001010",
  31353=>"110010011",
  31354=>"101010000",
  31355=>"101101111",
  31356=>"100111011",
  31357=>"000000101",
  31358=>"010101111",
  31359=>"001011010",
  31360=>"011100110",
  31361=>"000010110",
  31362=>"101110010",
  31363=>"101011010",
  31364=>"001010111",
  31365=>"101001110",
  31366=>"101011100",
  31367=>"100001010",
  31368=>"100100101",
  31369=>"001101000",
  31370=>"001111101",
  31371=>"001011100",
  31372=>"100010100",
  31373=>"001101111",
  31374=>"000001110",
  31375=>"001000110",
  31376=>"011000100",
  31377=>"101011110",
  31378=>"001101100",
  31379=>"001111111",
  31380=>"001100101",
  31381=>"000111010",
  31382=>"000001000",
  31383=>"111100100",
  31384=>"111101110",
  31385=>"101101111",
  31386=>"110011100",
  31387=>"011100011",
  31388=>"110001111",
  31389=>"101000000",
  31390=>"101100010",
  31391=>"101000100",
  31392=>"000000101",
  31393=>"111110000",
  31394=>"010100111",
  31395=>"010110000",
  31396=>"000011001",
  31397=>"111101110",
  31398=>"000010000",
  31399=>"100101001",
  31400=>"010001011",
  31401=>"111000111",
  31402=>"110100001",
  31403=>"010101100",
  31404=>"000010000",
  31405=>"000011010",
  31406=>"111101111",
  31407=>"110100111",
  31408=>"110010010",
  31409=>"001001011",
  31410=>"101110110",
  31411=>"011100011",
  31412=>"001001011",
  31413=>"100101011",
  31414=>"010111010",
  31415=>"111001000",
  31416=>"000101011",
  31417=>"001100110",
  31418=>"100011011",
  31419=>"000101000",
  31420=>"100100011",
  31421=>"110000010",
  31422=>"001101000",
  31423=>"100110101",
  31424=>"011111101",
  31425=>"100001001",
  31426=>"001000011",
  31427=>"110110111",
  31428=>"101110101",
  31429=>"001100110",
  31430=>"101111010",
  31431=>"001000110",
  31432=>"010110011",
  31433=>"110110100",
  31434=>"001111111",
  31435=>"010010011",
  31436=>"001011110",
  31437=>"100011101",
  31438=>"100000100",
  31439=>"111100000",
  31440=>"111111000",
  31441=>"001001001",
  31442=>"100101111",
  31443=>"010001100",
  31444=>"001100000",
  31445=>"110100011",
  31446=>"001100011",
  31447=>"100010000",
  31448=>"111000000",
  31449=>"101100001",
  31450=>"000101010",
  31451=>"100001011",
  31452=>"111110100",
  31453=>"100110101",
  31454=>"101010000",
  31455=>"001111110",
  31456=>"010001110",
  31457=>"010001111",
  31458=>"011000110",
  31459=>"011011111",
  31460=>"011011100",
  31461=>"111011001",
  31462=>"111100100",
  31463=>"010100110",
  31464=>"110101011",
  31465=>"001011001",
  31466=>"100101000",
  31467=>"011001010",
  31468=>"000000010",
  31469=>"100110111",
  31470=>"110100101",
  31471=>"111110101",
  31472=>"001001111",
  31473=>"010100000",
  31474=>"101010010",
  31475=>"010011011",
  31476=>"100111010",
  31477=>"000110000",
  31478=>"101100111",
  31479=>"010111100",
  31480=>"110110100",
  31481=>"110111100",
  31482=>"101101010",
  31483=>"111100110",
  31484=>"001011110",
  31485=>"000100010",
  31486=>"010110010",
  31487=>"111000100",
  31488=>"001001101",
  31489=>"111010110",
  31490=>"000011001",
  31491=>"110100100",
  31492=>"010010100",
  31493=>"001001111",
  31494=>"101111011",
  31495=>"000100000",
  31496=>"011001110",
  31497=>"100100011",
  31498=>"011101000",
  31499=>"100100000",
  31500=>"000111101",
  31501=>"111110111",
  31502=>"010000101",
  31503=>"010100010",
  31504=>"111110000",
  31505=>"011000011",
  31506=>"101010010",
  31507=>"100111111",
  31508=>"110000110",
  31509=>"001101100",
  31510=>"010110100",
  31511=>"101011110",
  31512=>"000011011",
  31513=>"110110001",
  31514=>"000010000",
  31515=>"111010010",
  31516=>"101110110",
  31517=>"000011000",
  31518=>"100110100",
  31519=>"100000111",
  31520=>"010011110",
  31521=>"000100010",
  31522=>"110111111",
  31523=>"100010010",
  31524=>"111000010",
  31525=>"010101010",
  31526=>"101000101",
  31527=>"011011011",
  31528=>"010100001",
  31529=>"011101010",
  31530=>"011011000",
  31531=>"100011110",
  31532=>"111010101",
  31533=>"100100010",
  31534=>"010010010",
  31535=>"001101000",
  31536=>"101010011",
  31537=>"111111011",
  31538=>"101111111",
  31539=>"000101100",
  31540=>"111010001",
  31541=>"101000111",
  31542=>"100001100",
  31543=>"010010000",
  31544=>"101010000",
  31545=>"001010111",
  31546=>"101101010",
  31547=>"111111011",
  31548=>"001001000",
  31549=>"100000001",
  31550=>"100000111",
  31551=>"001110000",
  31552=>"000101001",
  31553=>"101000100",
  31554=>"000001011",
  31555=>"001100110",
  31556=>"000011000",
  31557=>"101011111",
  31558=>"000101001",
  31559=>"001100011",
  31560=>"010000111",
  31561=>"011110000",
  31562=>"111001011",
  31563=>"000100001",
  31564=>"010000010",
  31565=>"011110001",
  31566=>"011011001",
  31567=>"110010100",
  31568=>"100001110",
  31569=>"101101111",
  31570=>"100011111",
  31571=>"101101100",
  31572=>"110111101",
  31573=>"100011010",
  31574=>"100000100",
  31575=>"100010011",
  31576=>"100011011",
  31577=>"111010010",
  31578=>"010110010",
  31579=>"001011001",
  31580=>"100000001",
  31581=>"011111110",
  31582=>"000010010",
  31583=>"100001101",
  31584=>"100100010",
  31585=>"111010000",
  31586=>"101000100",
  31587=>"001000011",
  31588=>"001000000",
  31589=>"101111111",
  31590=>"111111000",
  31591=>"110010100",
  31592=>"000000010",
  31593=>"100101111",
  31594=>"011101110",
  31595=>"101101100",
  31596=>"101111010",
  31597=>"101011001",
  31598=>"111011100",
  31599=>"001101001",
  31600=>"000011010",
  31601=>"101110011",
  31602=>"100010000",
  31603=>"011101010",
  31604=>"110010101",
  31605=>"101110100",
  31606=>"001101001",
  31607=>"100100011",
  31608=>"001011001",
  31609=>"000010000",
  31610=>"111100000",
  31611=>"101011111",
  31612=>"110100001",
  31613=>"110111010",
  31614=>"110100110",
  31615=>"111111111",
  31616=>"011000000",
  31617=>"011101001",
  31618=>"110100101",
  31619=>"110101000",
  31620=>"100111011",
  31621=>"110111011",
  31622=>"011111001",
  31623=>"011000000",
  31624=>"010010011",
  31625=>"011100111",
  31626=>"101101010",
  31627=>"100011110",
  31628=>"001001001",
  31629=>"011101010",
  31630=>"001101010",
  31631=>"110100000",
  31632=>"010010111",
  31633=>"101110100",
  31634=>"100011000",
  31635=>"011100000",
  31636=>"100101001",
  31637=>"011110111",
  31638=>"000001000",
  31639=>"110001111",
  31640=>"101001000",
  31641=>"010010010",
  31642=>"011011110",
  31643=>"011010001",
  31644=>"111111011",
  31645=>"001101111",
  31646=>"001111110",
  31647=>"110111110",
  31648=>"110110111",
  31649=>"000000110",
  31650=>"000010001",
  31651=>"101010111",
  31652=>"100110111",
  31653=>"111010000",
  31654=>"001000011",
  31655=>"000011100",
  31656=>"011011110",
  31657=>"000001100",
  31658=>"011001111",
  31659=>"000001011",
  31660=>"101001010",
  31661=>"011000101",
  31662=>"010001000",
  31663=>"011100111",
  31664=>"111100000",
  31665=>"111011111",
  31666=>"010111000",
  31667=>"001001001",
  31668=>"010100010",
  31669=>"101010110",
  31670=>"000111101",
  31671=>"000011000",
  31672=>"001111101",
  31673=>"000011100",
  31674=>"111101000",
  31675=>"110000110",
  31676=>"001001110",
  31677=>"001000011",
  31678=>"000100000",
  31679=>"011000011",
  31680=>"011001001",
  31681=>"111101110",
  31682=>"100010000",
  31683=>"000000010",
  31684=>"110010000",
  31685=>"001010101",
  31686=>"100010001",
  31687=>"011101000",
  31688=>"000000010",
  31689=>"001011011",
  31690=>"000001000",
  31691=>"110011111",
  31692=>"010101001",
  31693=>"011100011",
  31694=>"010110101",
  31695=>"101001011",
  31696=>"000001101",
  31697=>"100110101",
  31698=>"001101100",
  31699=>"011100100",
  31700=>"000010101",
  31701=>"000100000",
  31702=>"011010011",
  31703=>"011101001",
  31704=>"000000000",
  31705=>"111000100",
  31706=>"011101011",
  31707=>"000110101",
  31708=>"110011110",
  31709=>"010010000",
  31710=>"111100110",
  31711=>"010110111",
  31712=>"111110000",
  31713=>"001000010",
  31714=>"100101000",
  31715=>"001100000",
  31716=>"000111000",
  31717=>"111000001",
  31718=>"100111101",
  31719=>"001000010",
  31720=>"110011011",
  31721=>"110010100",
  31722=>"000011101",
  31723=>"011001000",
  31724=>"001001010",
  31725=>"101100011",
  31726=>"110111100",
  31727=>"011101111",
  31728=>"010110000",
  31729=>"001001101",
  31730=>"101001110",
  31731=>"111011100",
  31732=>"000011001",
  31733=>"110000111",
  31734=>"110101000",
  31735=>"110111101",
  31736=>"101111110",
  31737=>"000111101",
  31738=>"110000111",
  31739=>"010100110",
  31740=>"011010110",
  31741=>"101100110",
  31742=>"100111110",
  31743=>"100011001",
  31744=>"111000001",
  31745=>"010111110",
  31746=>"100110000",
  31747=>"110110001",
  31748=>"001011011",
  31749=>"010010000",
  31750=>"000100101",
  31751=>"100011011",
  31752=>"101000011",
  31753=>"100010101",
  31754=>"101100001",
  31755=>"110010110",
  31756=>"101100001",
  31757=>"010011110",
  31758=>"110111010",
  31759=>"000000100",
  31760=>"101111011",
  31761=>"111111100",
  31762=>"100011000",
  31763=>"110011011",
  31764=>"001110001",
  31765=>"001010111",
  31766=>"001111101",
  31767=>"000011111",
  31768=>"010010000",
  31769=>"010000010",
  31770=>"101100000",
  31771=>"101010111",
  31772=>"110001100",
  31773=>"101000011",
  31774=>"011110101",
  31775=>"000100000",
  31776=>"010011001",
  31777=>"101011001",
  31778=>"000101100",
  31779=>"100000001",
  31780=>"010100111",
  31781=>"010110110",
  31782=>"000101001",
  31783=>"010011010",
  31784=>"000011011",
  31785=>"100010101",
  31786=>"001010011",
  31787=>"001111101",
  31788=>"111101001",
  31789=>"001101100",
  31790=>"111101011",
  31791=>"011100001",
  31792=>"000010001",
  31793=>"100110011",
  31794=>"100111111",
  31795=>"101101111",
  31796=>"111001001",
  31797=>"000001110",
  31798=>"100110100",
  31799=>"110001100",
  31800=>"010001110",
  31801=>"110110110",
  31802=>"100111010",
  31803=>"011100011",
  31804=>"010010000",
  31805=>"111110001",
  31806=>"111011100",
  31807=>"011001000",
  31808=>"010110100",
  31809=>"100101101",
  31810=>"010010000",
  31811=>"011100001",
  31812=>"010111101",
  31813=>"110101001",
  31814=>"010000100",
  31815=>"001011000",
  31816=>"000100110",
  31817=>"111100000",
  31818=>"001000010",
  31819=>"001001100",
  31820=>"010110000",
  31821=>"111111100",
  31822=>"111110110",
  31823=>"000010001",
  31824=>"100110010",
  31825=>"111100111",
  31826=>"110100000",
  31827=>"010011100",
  31828=>"101011010",
  31829=>"101001001",
  31830=>"110100011",
  31831=>"101010100",
  31832=>"011101110",
  31833=>"011111111",
  31834=>"011111110",
  31835=>"101110011",
  31836=>"000000001",
  31837=>"000010011",
  31838=>"000000010",
  31839=>"011011100",
  31840=>"111001100",
  31841=>"111010000",
  31842=>"001001011",
  31843=>"010100011",
  31844=>"100100110",
  31845=>"000101111",
  31846=>"111010100",
  31847=>"000001100",
  31848=>"001011100",
  31849=>"011011110",
  31850=>"110001010",
  31851=>"001011100",
  31852=>"100100111",
  31853=>"101000111",
  31854=>"110111010",
  31855=>"111011110",
  31856=>"001000111",
  31857=>"001110001",
  31858=>"011111010",
  31859=>"110010100",
  31860=>"011110111",
  31861=>"110110111",
  31862=>"011111010",
  31863=>"011111110",
  31864=>"100101101",
  31865=>"011100101",
  31866=>"001010011",
  31867=>"011110101",
  31868=>"101101100",
  31869=>"000001110",
  31870=>"001001110",
  31871=>"100011000",
  31872=>"100110011",
  31873=>"010111110",
  31874=>"001010100",
  31875=>"101100001",
  31876=>"011011110",
  31877=>"000001000",
  31878=>"101010100",
  31879=>"111110001",
  31880=>"111101110",
  31881=>"001100001",
  31882=>"110011111",
  31883=>"011001101",
  31884=>"111101101",
  31885=>"011001100",
  31886=>"100110111",
  31887=>"001111001",
  31888=>"001001011",
  31889=>"110001110",
  31890=>"101010001",
  31891=>"110001110",
  31892=>"001000011",
  31893=>"001110001",
  31894=>"100001010",
  31895=>"000100100",
  31896=>"001100110",
  31897=>"100011011",
  31898=>"001011001",
  31899=>"110001011",
  31900=>"010000110",
  31901=>"100100010",
  31902=>"000100100",
  31903=>"100110000",
  31904=>"010110001",
  31905=>"111110000",
  31906=>"101001111",
  31907=>"111001000",
  31908=>"000011110",
  31909=>"111010101",
  31910=>"000000101",
  31911=>"001110100",
  31912=>"111011010",
  31913=>"100010101",
  31914=>"001000100",
  31915=>"101000111",
  31916=>"011010101",
  31917=>"110010010",
  31918=>"101001001",
  31919=>"100110011",
  31920=>"000001011",
  31921=>"111011111",
  31922=>"000010100",
  31923=>"001000000",
  31924=>"010100101",
  31925=>"010101000",
  31926=>"000001010",
  31927=>"111000000",
  31928=>"100010101",
  31929=>"100000110",
  31930=>"001111001",
  31931=>"001010101",
  31932=>"001111011",
  31933=>"100000100",
  31934=>"010111111",
  31935=>"011011001",
  31936=>"011010110",
  31937=>"001110100",
  31938=>"001010111",
  31939=>"100101100",
  31940=>"100010101",
  31941=>"111101111",
  31942=>"100110111",
  31943=>"110010010",
  31944=>"100100000",
  31945=>"110001001",
  31946=>"101011011",
  31947=>"001010110",
  31948=>"000110010",
  31949=>"101111111",
  31950=>"010010111",
  31951=>"100101000",
  31952=>"000101010",
  31953=>"001000110",
  31954=>"000100111",
  31955=>"100011010",
  31956=>"111000001",
  31957=>"000111001",
  31958=>"101101101",
  31959=>"010000010",
  31960=>"011001101",
  31961=>"000010100",
  31962=>"101011100",
  31963=>"110110101",
  31964=>"111000011",
  31965=>"110000010",
  31966=>"000000011",
  31967=>"111101111",
  31968=>"000000111",
  31969=>"001000110",
  31970=>"110001001",
  31971=>"000101110",
  31972=>"011011110",
  31973=>"100110001",
  31974=>"110010100",
  31975=>"001000001",
  31976=>"000000100",
  31977=>"000011001",
  31978=>"001111001",
  31979=>"100111001",
  31980=>"111101011",
  31981=>"010100011",
  31982=>"010000100",
  31983=>"100010100",
  31984=>"110010110",
  31985=>"101101110",
  31986=>"010101111",
  31987=>"101111100",
  31988=>"111000001",
  31989=>"110010100",
  31990=>"010111101",
  31991=>"011010010",
  31992=>"001001110",
  31993=>"101111000",
  31994=>"001101111",
  31995=>"010100000",
  31996=>"010111010",
  31997=>"111001110",
  31998=>"011101101",
  31999=>"000010001",
  32000=>"110010100",
  32001=>"010001010",
  32002=>"110111110",
  32003=>"001101011",
  32004=>"011001111",
  32005=>"111111001",
  32006=>"100001000",
  32007=>"100111011",
  32008=>"010010011",
  32009=>"110000111",
  32010=>"001000001",
  32011=>"011110011",
  32012=>"000000010",
  32013=>"101010011",
  32014=>"001000101",
  32015=>"111110011",
  32016=>"100001010",
  32017=>"010010111",
  32018=>"011101000",
  32019=>"111011110",
  32020=>"111001100",
  32021=>"011110011",
  32022=>"000111010",
  32023=>"001001111",
  32024=>"101101000",
  32025=>"100011110",
  32026=>"110110101",
  32027=>"011000010",
  32028=>"101100011",
  32029=>"100010110",
  32030=>"100001000",
  32031=>"000100110",
  32032=>"010111010",
  32033=>"000011001",
  32034=>"100110101",
  32035=>"000110110",
  32036=>"011110110",
  32037=>"110000000",
  32038=>"100110100",
  32039=>"100111000",
  32040=>"100111000",
  32041=>"111111010",
  32042=>"011000110",
  32043=>"001100100",
  32044=>"101100101",
  32045=>"011010001",
  32046=>"011100110",
  32047=>"010000111",
  32048=>"111001110",
  32049=>"000000001",
  32050=>"001100110",
  32051=>"010110000",
  32052=>"111001010",
  32053=>"110001000",
  32054=>"100111000",
  32055=>"010010111",
  32056=>"100000100",
  32057=>"111110110",
  32058=>"011010110",
  32059=>"010111010",
  32060=>"010101001",
  32061=>"010111101",
  32062=>"000000010",
  32063=>"010101111",
  32064=>"100010111",
  32065=>"100101011",
  32066=>"100100110",
  32067=>"110000110",
  32068=>"001000110",
  32069=>"010110010",
  32070=>"000111100",
  32071=>"010001010",
  32072=>"110011010",
  32073=>"110100000",
  32074=>"100000000",
  32075=>"010001011",
  32076=>"010100101",
  32077=>"001111011",
  32078=>"000000010",
  32079=>"001101100",
  32080=>"001110101",
  32081=>"100000111",
  32082=>"100000100",
  32083=>"111010111",
  32084=>"100001111",
  32085=>"001101000",
  32086=>"001111111",
  32087=>"001100011",
  32088=>"100001101",
  32089=>"100110110",
  32090=>"001001101",
  32091=>"010100001",
  32092=>"000100000",
  32093=>"011100101",
  32094=>"100100010",
  32095=>"101000000",
  32096=>"100100110",
  32097=>"101101100",
  32098=>"101001000",
  32099=>"010110010",
  32100=>"000100111",
  32101=>"111111101",
  32102=>"100100011",
  32103=>"111010010",
  32104=>"100111111",
  32105=>"101101001",
  32106=>"001001100",
  32107=>"110111010",
  32108=>"000101010",
  32109=>"110101101",
  32110=>"000001110",
  32111=>"010010000",
  32112=>"011000001",
  32113=>"010100001",
  32114=>"000011011",
  32115=>"101011110",
  32116=>"000100100",
  32117=>"010011010",
  32118=>"000101110",
  32119=>"100101010",
  32120=>"111100100",
  32121=>"011110111",
  32122=>"110011011",
  32123=>"101111101",
  32124=>"111101111",
  32125=>"111100011",
  32126=>"000111011",
  32127=>"110111110",
  32128=>"001101011",
  32129=>"011011100",
  32130=>"000001011",
  32131=>"000001010",
  32132=>"111101000",
  32133=>"010101101",
  32134=>"101111101",
  32135=>"100110000",
  32136=>"000000000",
  32137=>"101010111",
  32138=>"001001100",
  32139=>"110101010",
  32140=>"000110000",
  32141=>"001110111",
  32142=>"111001100",
  32143=>"010111110",
  32144=>"010110010",
  32145=>"010101101",
  32146=>"010111100",
  32147=>"000101111",
  32148=>"001000100",
  32149=>"011000000",
  32150=>"001001110",
  32151=>"110001111",
  32152=>"100011110",
  32153=>"001100011",
  32154=>"000010100",
  32155=>"111100110",
  32156=>"110100111",
  32157=>"100001011",
  32158=>"001101100",
  32159=>"010111001",
  32160=>"111011000",
  32161=>"001010001",
  32162=>"111010001",
  32163=>"000000000",
  32164=>"011000001",
  32165=>"010100001",
  32166=>"100111010",
  32167=>"111011111",
  32168=>"101100001",
  32169=>"010010110",
  32170=>"000111010",
  32171=>"000010001",
  32172=>"010000010",
  32173=>"101010111",
  32174=>"111101110",
  32175=>"010011011",
  32176=>"000001111",
  32177=>"100100010",
  32178=>"010100001",
  32179=>"101101011",
  32180=>"101000100",
  32181=>"100110110",
  32182=>"110111110",
  32183=>"001000011",
  32184=>"111100010",
  32185=>"001001010",
  32186=>"000111011",
  32187=>"101010010",
  32188=>"110100111",
  32189=>"100101000",
  32190=>"110100010",
  32191=>"010111010",
  32192=>"000000010",
  32193=>"100111001",
  32194=>"010100101",
  32195=>"101111001",
  32196=>"101101001",
  32197=>"000011011",
  32198=>"110000110",
  32199=>"110111111",
  32200=>"111110111",
  32201=>"000000011",
  32202=>"000000100",
  32203=>"110010011",
  32204=>"011010100",
  32205=>"101110101",
  32206=>"011001000",
  32207=>"001011101",
  32208=>"111100001",
  32209=>"000000000",
  32210=>"010101101",
  32211=>"011000000",
  32212=>"011111101",
  32213=>"100110100",
  32214=>"011001111",
  32215=>"011111000",
  32216=>"110001110",
  32217=>"101011111",
  32218=>"010001111",
  32219=>"011100011",
  32220=>"111010110",
  32221=>"111101101",
  32222=>"101010001",
  32223=>"101100101",
  32224=>"101100100",
  32225=>"000101010",
  32226=>"010011100",
  32227=>"110011010",
  32228=>"110001011",
  32229=>"110000101",
  32230=>"110110000",
  32231=>"111101001",
  32232=>"111010100",
  32233=>"100110000",
  32234=>"101110111",
  32235=>"000001111",
  32236=>"000000001",
  32237=>"001100010",
  32238=>"010000100",
  32239=>"111010000",
  32240=>"001110110",
  32241=>"010011100",
  32242=>"100010011",
  32243=>"010100000",
  32244=>"101000010",
  32245=>"111101101",
  32246=>"100110011",
  32247=>"101111100",
  32248=>"011000010",
  32249=>"000111010",
  32250=>"111010110",
  32251=>"100111101",
  32252=>"100101001",
  32253=>"100110011",
  32254=>"010101100",
  32255=>"010001100",
  32256=>"100000000",
  32257=>"111101111",
  32258=>"000011000",
  32259=>"010000000",
  32260=>"111100001",
  32261=>"010000010",
  32262=>"101000101",
  32263=>"000111110",
  32264=>"001010001",
  32265=>"100000110",
  32266=>"110101101",
  32267=>"000011010",
  32268=>"101001100",
  32269=>"111111001",
  32270=>"100000111",
  32271=>"001001000",
  32272=>"010100100",
  32273=>"000011111",
  32274=>"100110010",
  32275=>"001001000",
  32276=>"010100011",
  32277=>"111100100",
  32278=>"010101111",
  32279=>"010001110",
  32280=>"101110100",
  32281=>"000010100",
  32282=>"000010001",
  32283=>"000001000",
  32284=>"010111000",
  32285=>"111101101",
  32286=>"110011001",
  32287=>"001011011",
  32288=>"101010100",
  32289=>"100001100",
  32290=>"001111101",
  32291=>"001000000",
  32292=>"100101111",
  32293=>"001110010",
  32294=>"011101101",
  32295=>"000000110",
  32296=>"000111111",
  32297=>"000001101",
  32298=>"100100100",
  32299=>"001100100",
  32300=>"111001110",
  32301=>"111101111",
  32302=>"110011001",
  32303=>"101111001",
  32304=>"010001110",
  32305=>"001000111",
  32306=>"000110100",
  32307=>"110101010",
  32308=>"000010000",
  32309=>"101000001",
  32310=>"101110000",
  32311=>"111010111",
  32312=>"100000110",
  32313=>"111101000",
  32314=>"101001101",
  32315=>"111110010",
  32316=>"010111011",
  32317=>"011110110",
  32318=>"100001000",
  32319=>"101100001",
  32320=>"110000010",
  32321=>"001000001",
  32322=>"111001000",
  32323=>"001010111",
  32324=>"110001000",
  32325=>"110101001",
  32326=>"111101110",
  32327=>"100010010",
  32328=>"011000001",
  32329=>"100111000",
  32330=>"010110100",
  32331=>"001101100",
  32332=>"111001110",
  32333=>"000100100",
  32334=>"000000010",
  32335=>"000101110",
  32336=>"100111010",
  32337=>"000000111",
  32338=>"111011100",
  32339=>"011100001",
  32340=>"100111000",
  32341=>"111010100",
  32342=>"000100010",
  32343=>"100011010",
  32344=>"010010110",
  32345=>"010001101",
  32346=>"001101000",
  32347=>"010101101",
  32348=>"011010100",
  32349=>"001010110",
  32350=>"101001001",
  32351=>"010110000",
  32352=>"110111011",
  32353=>"000101100",
  32354=>"100100100",
  32355=>"110100000",
  32356=>"101010001",
  32357=>"101110101",
  32358=>"011111010",
  32359=>"010010011",
  32360=>"100000010",
  32361=>"010100110",
  32362=>"011001000",
  32363=>"101100101",
  32364=>"001111111",
  32365=>"000011111",
  32366=>"110001111",
  32367=>"011000111",
  32368=>"000010110",
  32369=>"010101101",
  32370=>"001111110",
  32371=>"101100111",
  32372=>"010001010",
  32373=>"111111111",
  32374=>"000110001",
  32375=>"101000100",
  32376=>"110111000",
  32377=>"001010100",
  32378=>"110100110",
  32379=>"101001110",
  32380=>"101100110",
  32381=>"111110011",
  32382=>"110011001",
  32383=>"011001011",
  32384=>"010010010",
  32385=>"011111010",
  32386=>"100000010",
  32387=>"100011101",
  32388=>"010000001",
  32389=>"101000110",
  32390=>"100100010",
  32391=>"010111100",
  32392=>"000111110",
  32393=>"000000000",
  32394=>"111000010",
  32395=>"010010100",
  32396=>"000101111",
  32397=>"111111110",
  32398=>"001000000",
  32399=>"111101010",
  32400=>"100011010",
  32401=>"111011100",
  32402=>"011100000",
  32403=>"000010101",
  32404=>"100000101",
  32405=>"101011111",
  32406=>"100111111",
  32407=>"011100011",
  32408=>"001010001",
  32409=>"111110100",
  32410=>"011101111",
  32411=>"000001001",
  32412=>"111000100",
  32413=>"111111111",
  32414=>"011101010",
  32415=>"001101111",
  32416=>"010101010",
  32417=>"001000001",
  32418=>"101110000",
  32419=>"000010100",
  32420=>"010101111",
  32421=>"100111100",
  32422=>"110001111",
  32423=>"001110111",
  32424=>"101101111",
  32425=>"001111000",
  32426=>"111010010",
  32427=>"101101011",
  32428=>"101011011",
  32429=>"111101011",
  32430=>"111110100",
  32431=>"001000010",
  32432=>"110011010",
  32433=>"100000111",
  32434=>"100011010",
  32435=>"011101100",
  32436=>"011000010",
  32437=>"000001011",
  32438=>"110000110",
  32439=>"001100101",
  32440=>"110011111",
  32441=>"000101000",
  32442=>"101011111",
  32443=>"000110100",
  32444=>"000000101",
  32445=>"100110110",
  32446=>"000010010",
  32447=>"110110000",
  32448=>"111101111",
  32449=>"110111111",
  32450=>"110111001",
  32451=>"001100011",
  32452=>"101000010",
  32453=>"011011000",
  32454=>"111010010",
  32455=>"011110110",
  32456=>"101110100",
  32457=>"110011101",
  32458=>"000010011",
  32459=>"001000001",
  32460=>"110110010",
  32461=>"011110001",
  32462=>"101110010",
  32463=>"010010000",
  32464=>"110011001",
  32465=>"101110001",
  32466=>"010100000",
  32467=>"011000110",
  32468=>"110111000",
  32469=>"000010100",
  32470=>"000010001",
  32471=>"110000000",
  32472=>"000111011",
  32473=>"101110110",
  32474=>"111100100",
  32475=>"010111111",
  32476=>"110001010",
  32477=>"111111101",
  32478=>"111110000",
  32479=>"001101100",
  32480=>"000000100",
  32481=>"100000110",
  32482=>"001100100",
  32483=>"111000110",
  32484=>"100000000",
  32485=>"000101101",
  32486=>"010010010",
  32487=>"101010011",
  32488=>"010011101",
  32489=>"011111110",
  32490=>"110001000",
  32491=>"000110011",
  32492=>"100110110",
  32493=>"001101010",
  32494=>"111000100",
  32495=>"111101011",
  32496=>"011011010",
  32497=>"000100000",
  32498=>"000001111",
  32499=>"101100100",
  32500=>"110000010",
  32501=>"011100010",
  32502=>"111111101",
  32503=>"000100101",
  32504=>"111001000",
  32505=>"000101101",
  32506=>"011100000",
  32507=>"000100101",
  32508=>"111111100",
  32509=>"101111101",
  32510=>"001010110",
  32511=>"011111111",
  32512=>"111110111",
  32513=>"001110100",
  32514=>"010110011",
  32515=>"010101110",
  32516=>"110101110",
  32517=>"000000110",
  32518=>"001101110",
  32519=>"001110011",
  32520=>"000101001",
  32521=>"111011001",
  32522=>"100111101",
  32523=>"000111110",
  32524=>"110111001",
  32525=>"001000111",
  32526=>"111010100",
  32527=>"001000010",
  32528=>"001011111",
  32529=>"001000010",
  32530=>"101101010",
  32531=>"001010111",
  32532=>"110010000",
  32533=>"010101010",
  32534=>"001000011",
  32535=>"111000100",
  32536=>"100010110",
  32537=>"110101111",
  32538=>"011101111",
  32539=>"000000110",
  32540=>"111111010",
  32541=>"011011111",
  32542=>"001001000",
  32543=>"101110110",
  32544=>"111110010",
  32545=>"111111000",
  32546=>"000011111",
  32547=>"011001110",
  32548=>"001001001",
  32549=>"001000111",
  32550=>"111110111",
  32551=>"000001010",
  32552=>"110010010",
  32553=>"111010100",
  32554=>"011011101",
  32555=>"000001110",
  32556=>"011000100",
  32557=>"000000010",
  32558=>"100101111",
  32559=>"000000000",
  32560=>"101001110",
  32561=>"111110000",
  32562=>"010000001",
  32563=>"111010110",
  32564=>"111101100",
  32565=>"101010001",
  32566=>"000000010",
  32567=>"010011111",
  32568=>"101101000",
  32569=>"101111001",
  32570=>"000100010",
  32571=>"111100000",
  32572=>"010111100",
  32573=>"111101100",
  32574=>"001110101",
  32575=>"111101000",
  32576=>"010100000",
  32577=>"101101010",
  32578=>"001111101",
  32579=>"101001111",
  32580=>"110010111",
  32581=>"101001001",
  32582=>"110101111",
  32583=>"000110100",
  32584=>"011000111",
  32585=>"110010111",
  32586=>"000101000",
  32587=>"100100111",
  32588=>"100000110",
  32589=>"001110010",
  32590=>"110011110",
  32591=>"001101001",
  32592=>"111111110",
  32593=>"000001100",
  32594=>"101001001",
  32595=>"100001101",
  32596=>"001011101",
  32597=>"011100010",
  32598=>"110111011",
  32599=>"010110011",
  32600=>"110000000",
  32601=>"011011100",
  32602=>"011010011",
  32603=>"110100100",
  32604=>"111111100",
  32605=>"111100100",
  32606=>"111101010",
  32607=>"101001001",
  32608=>"110000110",
  32609=>"111111101",
  32610=>"011010011",
  32611=>"000100001",
  32612=>"110101011",
  32613=>"001110101",
  32614=>"001101000",
  32615=>"100111111",
  32616=>"111000111",
  32617=>"011010001",
  32618=>"001010000",
  32619=>"101101001",
  32620=>"101010101",
  32621=>"100001110",
  32622=>"100010100",
  32623=>"011100000",
  32624=>"100110100",
  32625=>"001001001",
  32626=>"110000100",
  32627=>"000011100",
  32628=>"100110110",
  32629=>"010001010",
  32630=>"100111010",
  32631=>"000101100",
  32632=>"111100111",
  32633=>"100110011",
  32634=>"101000010",
  32635=>"101000101",
  32636=>"111010010",
  32637=>"011000011",
  32638=>"001010100",
  32639=>"011000100",
  32640=>"000010001",
  32641=>"000010111",
  32642=>"010010100",
  32643=>"000000100",
  32644=>"100010110",
  32645=>"011100100",
  32646=>"000100100",
  32647=>"110011001",
  32648=>"010101010",
  32649=>"011011001",
  32650=>"111111000",
  32651=>"000000100",
  32652=>"100101001",
  32653=>"110100100",
  32654=>"010101001",
  32655=>"110010100",
  32656=>"111111101",
  32657=>"110101001",
  32658=>"110110101",
  32659=>"101010111",
  32660=>"101110111",
  32661=>"010010101",
  32662=>"010000001",
  32663=>"101011101",
  32664=>"111001011",
  32665=>"001010101",
  32666=>"000010000",
  32667=>"011001100",
  32668=>"011011101",
  32669=>"011001111",
  32670=>"101001011",
  32671=>"110011101",
  32672=>"111101001",
  32673=>"011110111",
  32674=>"001001001",
  32675=>"100000010",
  32676=>"000001010",
  32677=>"010110101",
  32678=>"000100010",
  32679=>"111001001",
  32680=>"011010110",
  32681=>"000110100",
  32682=>"010111110",
  32683=>"000000111",
  32684=>"011110111",
  32685=>"011100101",
  32686=>"100101010",
  32687=>"010011001",
  32688=>"001000101",
  32689=>"100011111",
  32690=>"000001111",
  32691=>"100110111",
  32692=>"111111101",
  32693=>"010101000",
  32694=>"000010011",
  32695=>"111010001",
  32696=>"000010100",
  32697=>"011101101",
  32698=>"110101011",
  32699=>"110111110",
  32700=>"100000010",
  32701=>"101000010",
  32702=>"100010101",
  32703=>"001010000",
  32704=>"000100011",
  32705=>"101100011",
  32706=>"000010000",
  32707=>"000111010",
  32708=>"111111010",
  32709=>"100101110",
  32710=>"110000101",
  32711=>"101100110",
  32712=>"111001010",
  32713=>"101101010",
  32714=>"001010000",
  32715=>"011011010",
  32716=>"101011000",
  32717=>"011000011",
  32718=>"010111001",
  32719=>"100101010",
  32720=>"111111101",
  32721=>"000000010",
  32722=>"101001000",
  32723=>"011101001",
  32724=>"111101111",
  32725=>"111101011",
  32726=>"010011001",
  32727=>"010110101",
  32728=>"010100101",
  32729=>"101101111",
  32730=>"001000001",
  32731=>"100000101",
  32732=>"111000011",
  32733=>"111011010",
  32734=>"111001111",
  32735=>"000000001",
  32736=>"001000101",
  32737=>"111001110",
  32738=>"111000110",
  32739=>"010001100",
  32740=>"100100101",
  32741=>"111000110",
  32742=>"001001101",
  32743=>"100111011",
  32744=>"001100101",
  32745=>"011100000",
  32746=>"001101001",
  32747=>"110101001",
  32748=>"111001011",
  32749=>"000100000",
  32750=>"001101001",
  32751=>"111110010",
  32752=>"110000011",
  32753=>"101100100",
  32754=>"101011100",
  32755=>"001101110",
  32756=>"000110001",
  32757=>"111111111",
  32758=>"111101011",
  32759=>"000001000",
  32760=>"011000101",
  32761=>"101101011",
  32762=>"110101100",
  32763=>"111000000",
  32764=>"011011000",
  32765=>"101100110",
  32766=>"111100010",
  32767=>"010100010",
  32768=>"010010110",
  32769=>"000101000",
  32770=>"111011011",
  32771=>"100100110",
  32772=>"111011010",
  32773=>"000011001",
  32774=>"001101000",
  32775=>"111101010",
  32776=>"011000110",
  32777=>"000000001",
  32778=>"010101110",
  32779=>"011001000",
  32780=>"010001100",
  32781=>"001110001",
  32782=>"010110000",
  32783=>"011011011",
  32784=>"000001100",
  32785=>"000100010",
  32786=>"000101110",
  32787=>"000001111",
  32788=>"110011100",
  32789=>"100110011",
  32790=>"100110001",
  32791=>"110101110",
  32792=>"100101100",
  32793=>"000010100",
  32794=>"011000011",
  32795=>"011011110",
  32796=>"100000010",
  32797=>"111000101",
  32798=>"011110011",
  32799=>"010000101",
  32800=>"101100001",
  32801=>"111110111",
  32802=>"011000010",
  32803=>"111101010",
  32804=>"110001111",
  32805=>"010100100",
  32806=>"111000011",
  32807=>"110101010",
  32808=>"010101101",
  32809=>"010011111",
  32810=>"111010110",
  32811=>"101001010",
  32812=>"110111100",
  32813=>"100000110",
  32814=>"010000001",
  32815=>"011000000",
  32816=>"001010100",
  32817=>"001000111",
  32818=>"110001000",
  32819=>"011111101",
  32820=>"111011100",
  32821=>"011011001",
  32822=>"100111001",
  32823=>"001111011",
  32824=>"011001100",
  32825=>"110000101",
  32826=>"000000110",
  32827=>"000101010",
  32828=>"100100001",
  32829=>"100110111",
  32830=>"000001100",
  32831=>"111110011",
  32832=>"010000011",
  32833=>"000011010",
  32834=>"011101001",
  32835=>"110010011",
  32836=>"011000100",
  32837=>"001100111",
  32838=>"101011101",
  32839=>"001111010",
  32840=>"100110011",
  32841=>"101000000",
  32842=>"000100001",
  32843=>"000010011",
  32844=>"110111111",
  32845=>"100101101",
  32846=>"001110110",
  32847=>"101101110",
  32848=>"110100001",
  32849=>"101110001",
  32850=>"110101011",
  32851=>"111000001",
  32852=>"101110000",
  32853=>"011000011",
  32854=>"101100001",
  32855=>"111111101",
  32856=>"101011011",
  32857=>"100001011",
  32858=>"001100001",
  32859=>"000100110",
  32860=>"110000111",
  32861=>"111001010",
  32862=>"001000000",
  32863=>"110001010",
  32864=>"011011101",
  32865=>"001011001",
  32866=>"010010010",
  32867=>"011101101",
  32868=>"011101000",
  32869=>"011010010",
  32870=>"011110111",
  32871=>"001101000",
  32872=>"011100001",
  32873=>"111110101",
  32874=>"111000111",
  32875=>"011111110",
  32876=>"010000001",
  32877=>"010011101",
  32878=>"001110100",
  32879=>"101101000",
  32880=>"011001001",
  32881=>"001001110",
  32882=>"011001000",
  32883=>"111011111",
  32884=>"101000100",
  32885=>"000101010",
  32886=>"000101101",
  32887=>"001111100",
  32888=>"111001000",
  32889=>"001111001",
  32890=>"000101101",
  32891=>"000010011",
  32892=>"001010100",
  32893=>"000000101",
  32894=>"010000111",
  32895=>"011110010",
  32896=>"110100101",
  32897=>"011011001",
  32898=>"000000010",
  32899=>"000001100",
  32900=>"011111000",
  32901=>"001000010",
  32902=>"111100110",
  32903=>"010011111",
  32904=>"001011011",
  32905=>"011000001",
  32906=>"111101011",
  32907=>"000111110",
  32908=>"011010101",
  32909=>"011000001",
  32910=>"001011110",
  32911=>"000000110",
  32912=>"110110001",
  32913=>"111010001",
  32914=>"011111100",
  32915=>"111110000",
  32916=>"111000110",
  32917=>"110111101",
  32918=>"100110111",
  32919=>"100111110",
  32920=>"111110100",
  32921=>"000110000",
  32922=>"110000100",
  32923=>"110011000",
  32924=>"100110101",
  32925=>"011001010",
  32926=>"111111110",
  32927=>"101111100",
  32928=>"000101110",
  32929=>"101011010",
  32930=>"010100101",
  32931=>"100101011",
  32932=>"011011001",
  32933=>"001010110",
  32934=>"100110010",
  32935=>"100000011",
  32936=>"101001110",
  32937=>"101100100",
  32938=>"101011000",
  32939=>"010010000",
  32940=>"111101111",
  32941=>"111110111",
  32942=>"100110110",
  32943=>"100111110",
  32944=>"000011000",
  32945=>"000000000",
  32946=>"100110111",
  32947=>"100011010",
  32948=>"110010011",
  32949=>"101111111",
  32950=>"001011111",
  32951=>"001110100",
  32952=>"100101011",
  32953=>"010110010",
  32954=>"001111011",
  32955=>"001000110",
  32956=>"110001011",
  32957=>"000100111",
  32958=>"010001011",
  32959=>"111011011",
  32960=>"000111001",
  32961=>"000010101",
  32962=>"011000100",
  32963=>"001010001",
  32964=>"110010111",
  32965=>"000100011",
  32966=>"100101110",
  32967=>"100010100",
  32968=>"011000011",
  32969=>"100110111",
  32970=>"001110100",
  32971=>"100101100",
  32972=>"011100111",
  32973=>"111011111",
  32974=>"000000001",
  32975=>"001100010",
  32976=>"110001100",
  32977=>"100001001",
  32978=>"011001110",
  32979=>"111010010",
  32980=>"001101100",
  32981=>"011010011",
  32982=>"110010101",
  32983=>"000111001",
  32984=>"010000000",
  32985=>"000000011",
  32986=>"101010011",
  32987=>"000011100",
  32988=>"101010101",
  32989=>"010001000",
  32990=>"110100111",
  32991=>"100111110",
  32992=>"100001000",
  32993=>"101101111",
  32994=>"010010010",
  32995=>"111011001",
  32996=>"100101000",
  32997=>"101110110",
  32998=>"001011010",
  32999=>"000111010",
  33000=>"000010111",
  33001=>"011010000",
  33002=>"000111001",
  33003=>"110110010",
  33004=>"111111010",
  33005=>"100011000",
  33006=>"101100101",
  33007=>"001011001",
  33008=>"101001100",
  33009=>"111011100",
  33010=>"010001100",
  33011=>"111010110",
  33012=>"100101000",
  33013=>"000100101",
  33014=>"000111101",
  33015=>"000011110",
  33016=>"100010101",
  33017=>"010100100",
  33018=>"000001111",
  33019=>"010010100",
  33020=>"010010000",
  33021=>"101110110",
  33022=>"000101001",
  33023=>"011100110",
  33024=>"111001000",
  33025=>"011111111",
  33026=>"000000101",
  33027=>"000010000",
  33028=>"101010110",
  33029=>"101010010",
  33030=>"111011101",
  33031=>"100000101",
  33032=>"001000100",
  33033=>"100001100",
  33034=>"111111011",
  33035=>"100100000",
  33036=>"001001001",
  33037=>"001101001",
  33038=>"000010001",
  33039=>"111110000",
  33040=>"000010001",
  33041=>"111001110",
  33042=>"010001111",
  33043=>"100100011",
  33044=>"110011100",
  33045=>"001101000",
  33046=>"001111000",
  33047=>"111101000",
  33048=>"101111101",
  33049=>"010010111",
  33050=>"110101111",
  33051=>"000010110",
  33052=>"011110010",
  33053=>"110110100",
  33054=>"010000100",
  33055=>"000011110",
  33056=>"011001100",
  33057=>"011100101",
  33058=>"010001100",
  33059=>"000000001",
  33060=>"001000111",
  33061=>"011111001",
  33062=>"110000010",
  33063=>"111011100",
  33064=>"010100010",
  33065=>"101001011",
  33066=>"001111001",
  33067=>"001001001",
  33068=>"011000100",
  33069=>"001111111",
  33070=>"011001010",
  33071=>"100100110",
  33072=>"101110100",
  33073=>"111001001",
  33074=>"001101111",
  33075=>"000011110",
  33076=>"000010110",
  33077=>"010001111",
  33078=>"011011001",
  33079=>"010011101",
  33080=>"100110000",
  33081=>"001111010",
  33082=>"000000110",
  33083=>"111101000",
  33084=>"011111010",
  33085=>"000011110",
  33086=>"011000100",
  33087=>"001110001",
  33088=>"111011000",
  33089=>"001001110",
  33090=>"010101111",
  33091=>"111110010",
  33092=>"101101100",
  33093=>"000010100",
  33094=>"110110000",
  33095=>"101010110",
  33096=>"111010001",
  33097=>"100010011",
  33098=>"101000000",
  33099=>"011110110",
  33100=>"101101101",
  33101=>"010110101",
  33102=>"101101100",
  33103=>"010011001",
  33104=>"110000010",
  33105=>"010110011",
  33106=>"001101010",
  33107=>"100010100",
  33108=>"110011011",
  33109=>"100101000",
  33110=>"000000010",
  33111=>"111110110",
  33112=>"101011000",
  33113=>"010010010",
  33114=>"000111100",
  33115=>"100010101",
  33116=>"110101100",
  33117=>"010110101",
  33118=>"101001001",
  33119=>"000110000",
  33120=>"100001011",
  33121=>"010100000",
  33122=>"010010110",
  33123=>"110100001",
  33124=>"001110001",
  33125=>"010011000",
  33126=>"000001010",
  33127=>"100001100",
  33128=>"001010010",
  33129=>"011101101",
  33130=>"111111000",
  33131=>"000101000",
  33132=>"011101010",
  33133=>"011100110",
  33134=>"100100011",
  33135=>"110100000",
  33136=>"001100101",
  33137=>"011011101",
  33138=>"101100101",
  33139=>"111100101",
  33140=>"011111000",
  33141=>"011001100",
  33142=>"010010011",
  33143=>"000111111",
  33144=>"001011110",
  33145=>"100010110",
  33146=>"011100000",
  33147=>"011110101",
  33148=>"101100011",
  33149=>"001000100",
  33150=>"000010000",
  33151=>"101010100",
  33152=>"101110010",
  33153=>"010101110",
  33154=>"111001110",
  33155=>"111001001",
  33156=>"100010111",
  33157=>"001011111",
  33158=>"010111010",
  33159=>"000111000",
  33160=>"010100100",
  33161=>"000101010",
  33162=>"010011111",
  33163=>"111001011",
  33164=>"010111011",
  33165=>"011011111",
  33166=>"000101101",
  33167=>"101010100",
  33168=>"001011111",
  33169=>"011100000",
  33170=>"111111110",
  33171=>"010001100",
  33172=>"100010110",
  33173=>"000000100",
  33174=>"101001111",
  33175=>"010100101",
  33176=>"000001111",
  33177=>"110000001",
  33178=>"111001111",
  33179=>"010010111",
  33180=>"111001010",
  33181=>"100110001",
  33182=>"100001101",
  33183=>"101100101",
  33184=>"111111010",
  33185=>"000001110",
  33186=>"111001101",
  33187=>"010100011",
  33188=>"000011000",
  33189=>"000011100",
  33190=>"110100110",
  33191=>"100101111",
  33192=>"101101101",
  33193=>"101111101",
  33194=>"001101010",
  33195=>"100000011",
  33196=>"011010101",
  33197=>"000000111",
  33198=>"110010000",
  33199=>"110110101",
  33200=>"110100100",
  33201=>"001001100",
  33202=>"010110000",
  33203=>"110001010",
  33204=>"011001001",
  33205=>"110001101",
  33206=>"101110111",
  33207=>"101111011",
  33208=>"001001001",
  33209=>"000100011",
  33210=>"110111110",
  33211=>"100111111",
  33212=>"100000010",
  33213=>"100100111",
  33214=>"001101010",
  33215=>"111000000",
  33216=>"110010001",
  33217=>"011001011",
  33218=>"111010010",
  33219=>"001001100",
  33220=>"011100110",
  33221=>"010100000",
  33222=>"110111100",
  33223=>"010010010",
  33224=>"101001000",
  33225=>"011110000",
  33226=>"000001101",
  33227=>"001000001",
  33228=>"110011111",
  33229=>"001011100",
  33230=>"101101011",
  33231=>"110011011",
  33232=>"011110101",
  33233=>"110110110",
  33234=>"011001111",
  33235=>"010110011",
  33236=>"111100110",
  33237=>"111010110",
  33238=>"111110010",
  33239=>"001000011",
  33240=>"010101001",
  33241=>"000110111",
  33242=>"100101010",
  33243=>"111000111",
  33244=>"001010110",
  33245=>"000110111",
  33246=>"101100001",
  33247=>"101000001",
  33248=>"100100110",
  33249=>"011101110",
  33250=>"101110111",
  33251=>"001000111",
  33252=>"010011111",
  33253=>"101001111",
  33254=>"101010110",
  33255=>"110011110",
  33256=>"010010110",
  33257=>"111011000",
  33258=>"100011010",
  33259=>"000111101",
  33260=>"100000100",
  33261=>"100010001",
  33262=>"011110100",
  33263=>"001001001",
  33264=>"101101001",
  33265=>"001001101",
  33266=>"010111111",
  33267=>"100100010",
  33268=>"001101111",
  33269=>"010110000",
  33270=>"111111100",
  33271=>"010010001",
  33272=>"000001000",
  33273=>"101101010",
  33274=>"011010110",
  33275=>"101001010",
  33276=>"010101001",
  33277=>"100011110",
  33278=>"100010110",
  33279=>"001001101",
  33280=>"011110011",
  33281=>"001000001",
  33282=>"111100110",
  33283=>"000011011",
  33284=>"110011001",
  33285=>"110100000",
  33286=>"011110111",
  33287=>"100000010",
  33288=>"000010000",
  33289=>"110100101",
  33290=>"001110000",
  33291=>"100101110",
  33292=>"100011101",
  33293=>"100100101",
  33294=>"000010101",
  33295=>"000000011",
  33296=>"100110110",
  33297=>"100111101",
  33298=>"010001100",
  33299=>"000001011",
  33300=>"110011101",
  33301=>"001000010",
  33302=>"011011101",
  33303=>"111001100",
  33304=>"011100100",
  33305=>"010000000",
  33306=>"000001101",
  33307=>"100001101",
  33308=>"000100111",
  33309=>"010011111",
  33310=>"010010011",
  33311=>"010110000",
  33312=>"000001011",
  33313=>"101010000",
  33314=>"101011111",
  33315=>"011000101",
  33316=>"111010110",
  33317=>"000001010",
  33318=>"101001011",
  33319=>"000111000",
  33320=>"000101100",
  33321=>"101101110",
  33322=>"000010010",
  33323=>"000100000",
  33324=>"010000101",
  33325=>"101100011",
  33326=>"000111000",
  33327=>"110110111",
  33328=>"000001100",
  33329=>"100110001",
  33330=>"000001111",
  33331=>"110001111",
  33332=>"000100101",
  33333=>"000011011",
  33334=>"001110111",
  33335=>"000101111",
  33336=>"100111110",
  33337=>"000000101",
  33338=>"011010000",
  33339=>"010011000",
  33340=>"100011011",
  33341=>"111001100",
  33342=>"011010000",
  33343=>"000001110",
  33344=>"000011010",
  33345=>"110010100",
  33346=>"010011100",
  33347=>"101100101",
  33348=>"111110010",
  33349=>"011000000",
  33350=>"001010101",
  33351=>"000001101",
  33352=>"100000110",
  33353=>"001111100",
  33354=>"111011100",
  33355=>"110000011",
  33356=>"101111001",
  33357=>"001110000",
  33358=>"010010011",
  33359=>"111100001",
  33360=>"010110111",
  33361=>"010110001",
  33362=>"111110010",
  33363=>"000001001",
  33364=>"010000001",
  33365=>"110111001",
  33366=>"111110110",
  33367=>"101101011",
  33368=>"001011000",
  33369=>"110111100",
  33370=>"100010011",
  33371=>"110110000",
  33372=>"000001011",
  33373=>"011100100",
  33374=>"011111000",
  33375=>"010111011",
  33376=>"000100100",
  33377=>"110100011",
  33378=>"111001110",
  33379=>"101000111",
  33380=>"111001111",
  33381=>"001101110",
  33382=>"010100010",
  33383=>"111000010",
  33384=>"011000100",
  33385=>"100101110",
  33386=>"101110101",
  33387=>"000101010",
  33388=>"111111000",
  33389=>"110111111",
  33390=>"101110101",
  33391=>"110100000",
  33392=>"000010111",
  33393=>"011101000",
  33394=>"011111001",
  33395=>"111110001",
  33396=>"111100011",
  33397=>"011101100",
  33398=>"111011011",
  33399=>"001011011",
  33400=>"010010000",
  33401=>"001110110",
  33402=>"001100011",
  33403=>"110001111",
  33404=>"100010100",
  33405=>"010101111",
  33406=>"010010010",
  33407=>"001001001",
  33408=>"111111010",
  33409=>"001011010",
  33410=>"000010010",
  33411=>"000101101",
  33412=>"111100100",
  33413=>"010101100",
  33414=>"010101111",
  33415=>"011000100",
  33416=>"011000010",
  33417=>"100000000",
  33418=>"010011110",
  33419=>"010110000",
  33420=>"010000011",
  33421=>"101101000",
  33422=>"100001111",
  33423=>"100001010",
  33424=>"101111111",
  33425=>"010010100",
  33426=>"110110011",
  33427=>"101101101",
  33428=>"110100000",
  33429=>"110111100",
  33430=>"000000101",
  33431=>"111010100",
  33432=>"110001000",
  33433=>"101010010",
  33434=>"110000011",
  33435=>"100000001",
  33436=>"010001100",
  33437=>"110011100",
  33438=>"101110011",
  33439=>"101100001",
  33440=>"100000011",
  33441=>"100000110",
  33442=>"001100110",
  33443=>"001011100",
  33444=>"100101101",
  33445=>"101010110",
  33446=>"000011110",
  33447=>"101001111",
  33448=>"001011110",
  33449=>"011010101",
  33450=>"001110000",
  33451=>"110011000",
  33452=>"000101111",
  33453=>"111011101",
  33454=>"001010010",
  33455=>"010110000",
  33456=>"010100110",
  33457=>"010111010",
  33458=>"101100010",
  33459=>"000011010",
  33460=>"101100100",
  33461=>"011100000",
  33462=>"000111101",
  33463=>"100101010",
  33464=>"011000110",
  33465=>"101010001",
  33466=>"111111101",
  33467=>"010111010",
  33468=>"011010101",
  33469=>"100101110",
  33470=>"010000001",
  33471=>"011001000",
  33472=>"101111110",
  33473=>"110001110",
  33474=>"100111000",
  33475=>"011101001",
  33476=>"010111110",
  33477=>"011001110",
  33478=>"101110001",
  33479=>"001111010",
  33480=>"110110100",
  33481=>"110001100",
  33482=>"011111010",
  33483=>"110010010",
  33484=>"000110001",
  33485=>"000001011",
  33486=>"101001000",
  33487=>"101111011",
  33488=>"010000011",
  33489=>"011011011",
  33490=>"001010110",
  33491=>"110101110",
  33492=>"001111011",
  33493=>"100100100",
  33494=>"101001000",
  33495=>"010101110",
  33496=>"011111010",
  33497=>"111101010",
  33498=>"100010000",
  33499=>"111011111",
  33500=>"111001111",
  33501=>"101101000",
  33502=>"011010010",
  33503=>"010010110",
  33504=>"111001101",
  33505=>"101001100",
  33506=>"110011000",
  33507=>"000101001",
  33508=>"111110010",
  33509=>"111110111",
  33510=>"000000001",
  33511=>"010001010",
  33512=>"010011100",
  33513=>"011000001",
  33514=>"111110111",
  33515=>"110110001",
  33516=>"110110100",
  33517=>"111010000",
  33518=>"101001111",
  33519=>"110101111",
  33520=>"100001111",
  33521=>"011011110",
  33522=>"111000110",
  33523=>"010010110",
  33524=>"111010010",
  33525=>"111111110",
  33526=>"011101110",
  33527=>"000100101",
  33528=>"000000110",
  33529=>"010010000",
  33530=>"101000110",
  33531=>"100001101",
  33532=>"001101011",
  33533=>"001000110",
  33534=>"001001110",
  33535=>"111011000",
  33536=>"000100111",
  33537=>"100111111",
  33538=>"111111011",
  33539=>"111011000",
  33540=>"111000001",
  33541=>"010101001",
  33542=>"000101001",
  33543=>"000101100",
  33544=>"111110000",
  33545=>"010110011",
  33546=>"111100110",
  33547=>"110000101",
  33548=>"000000001",
  33549=>"101000011",
  33550=>"011100100",
  33551=>"001101011",
  33552=>"110110100",
  33553=>"000111100",
  33554=>"101001101",
  33555=>"100110100",
  33556=>"100011110",
  33557=>"000100111",
  33558=>"011000110",
  33559=>"010011000",
  33560=>"010001110",
  33561=>"100000011",
  33562=>"111000110",
  33563=>"000000011",
  33564=>"101100111",
  33565=>"101111010",
  33566=>"010100101",
  33567=>"010011011",
  33568=>"111001101",
  33569=>"101000000",
  33570=>"001011100",
  33571=>"100011100",
  33572=>"000111001",
  33573=>"100001000",
  33574=>"100111010",
  33575=>"101101001",
  33576=>"011010010",
  33577=>"001111100",
  33578=>"010010101",
  33579=>"101001000",
  33580=>"010110001",
  33581=>"001111010",
  33582=>"010000000",
  33583=>"110010000",
  33584=>"111111011",
  33585=>"111100001",
  33586=>"111100000",
  33587=>"011000111",
  33588=>"110110010",
  33589=>"100011010",
  33590=>"110101000",
  33591=>"110000111",
  33592=>"100001110",
  33593=>"110010000",
  33594=>"101000001",
  33595=>"101001000",
  33596=>"100000100",
  33597=>"011010010",
  33598=>"101010100",
  33599=>"111011111",
  33600=>"110001101",
  33601=>"010101001",
  33602=>"110001100",
  33603=>"110110110",
  33604=>"001110011",
  33605=>"101101100",
  33606=>"101000011",
  33607=>"110111000",
  33608=>"110100111",
  33609=>"111010101",
  33610=>"010100010",
  33611=>"101000011",
  33612=>"111011011",
  33613=>"101000001",
  33614=>"111100010",
  33615=>"000110111",
  33616=>"011111000",
  33617=>"010000101",
  33618=>"110010010",
  33619=>"001001101",
  33620=>"111001001",
  33621=>"110111110",
  33622=>"000010111",
  33623=>"001000110",
  33624=>"011011010",
  33625=>"000010011",
  33626=>"010110011",
  33627=>"100001011",
  33628=>"111000011",
  33629=>"100000111",
  33630=>"101000100",
  33631=>"001001011",
  33632=>"000001110",
  33633=>"010111001",
  33634=>"110101110",
  33635=>"110101001",
  33636=>"010011110",
  33637=>"000000100",
  33638=>"110111000",
  33639=>"100010000",
  33640=>"010100010",
  33641=>"011101111",
  33642=>"110000110",
  33643=>"010000011",
  33644=>"100101011",
  33645=>"111111100",
  33646=>"001001110",
  33647=>"110110011",
  33648=>"010000111",
  33649=>"100010001",
  33650=>"110010000",
  33651=>"001110011",
  33652=>"010010111",
  33653=>"000001101",
  33654=>"010101111",
  33655=>"100010001",
  33656=>"110100111",
  33657=>"110100100",
  33658=>"100010110",
  33659=>"010000000",
  33660=>"010001010",
  33661=>"010100110",
  33662=>"001010111",
  33663=>"101111011",
  33664=>"101010000",
  33665=>"110111111",
  33666=>"000010010",
  33667=>"111111010",
  33668=>"100000101",
  33669=>"011100000",
  33670=>"100001111",
  33671=>"001000110",
  33672=>"100010011",
  33673=>"011110110",
  33674=>"000001001",
  33675=>"110100011",
  33676=>"010101111",
  33677=>"111100111",
  33678=>"001010111",
  33679=>"010010111",
  33680=>"000000110",
  33681=>"100111101",
  33682=>"000100110",
  33683=>"011000110",
  33684=>"101000110",
  33685=>"001001000",
  33686=>"000101111",
  33687=>"101111101",
  33688=>"111111000",
  33689=>"000101010",
  33690=>"101111001",
  33691=>"001001110",
  33692=>"110001100",
  33693=>"101101001",
  33694=>"000010010",
  33695=>"101011111",
  33696=>"011100011",
  33697=>"001100001",
  33698=>"000100100",
  33699=>"010011000",
  33700=>"101010111",
  33701=>"111010110",
  33702=>"000010111",
  33703=>"011000011",
  33704=>"001100110",
  33705=>"101010001",
  33706=>"111101010",
  33707=>"001010000",
  33708=>"010001000",
  33709=>"101111000",
  33710=>"110000111",
  33711=>"100010101",
  33712=>"111001010",
  33713=>"111110110",
  33714=>"011010100",
  33715=>"110101010",
  33716=>"111001100",
  33717=>"000100101",
  33718=>"111111000",
  33719=>"001010101",
  33720=>"000100000",
  33721=>"001001111",
  33722=>"010011011",
  33723=>"111010010",
  33724=>"100011010",
  33725=>"111000011",
  33726=>"001110101",
  33727=>"010011110",
  33728=>"010000000",
  33729=>"000000001",
  33730=>"110101010",
  33731=>"111111000",
  33732=>"001101110",
  33733=>"011001001",
  33734=>"011000001",
  33735=>"101110000",
  33736=>"000001001",
  33737=>"101110010",
  33738=>"100010010",
  33739=>"110000011",
  33740=>"111111110",
  33741=>"101111011",
  33742=>"010010110",
  33743=>"001111100",
  33744=>"001010011",
  33745=>"010101010",
  33746=>"000011110",
  33747=>"000100000",
  33748=>"101111101",
  33749=>"111010001",
  33750=>"001101101",
  33751=>"100101111",
  33752=>"100101101",
  33753=>"011011011",
  33754=>"100010011",
  33755=>"111000100",
  33756=>"001000110",
  33757=>"111011101",
  33758=>"001101110",
  33759=>"100001111",
  33760=>"111110111",
  33761=>"011011011",
  33762=>"111011000",
  33763=>"001010000",
  33764=>"111001000",
  33765=>"110110011",
  33766=>"000010011",
  33767=>"101011011",
  33768=>"111010010",
  33769=>"000011010",
  33770=>"001011000",
  33771=>"100110000",
  33772=>"101110001",
  33773=>"110110000",
  33774=>"100011010",
  33775=>"000011011",
  33776=>"110011111",
  33777=>"000111011",
  33778=>"100000110",
  33779=>"010000011",
  33780=>"101011100",
  33781=>"000110010",
  33782=>"100011010",
  33783=>"000010000",
  33784=>"000000010",
  33785=>"100000000",
  33786=>"010101100",
  33787=>"000000000",
  33788=>"100000011",
  33789=>"111100011",
  33790=>"010110000",
  33791=>"111100110",
  33792=>"011111000",
  33793=>"100011001",
  33794=>"011101011",
  33795=>"100010111",
  33796=>"101111111",
  33797=>"100001001",
  33798=>"110101001",
  33799=>"001101001",
  33800=>"100111001",
  33801=>"110111100",
  33802=>"011100010",
  33803=>"000110010",
  33804=>"111110101",
  33805=>"101110010",
  33806=>"110111110",
  33807=>"000011111",
  33808=>"101100010",
  33809=>"001111110",
  33810=>"000100110",
  33811=>"111010010",
  33812=>"110101110",
  33813=>"110001010",
  33814=>"010101010",
  33815=>"001011111",
  33816=>"001001011",
  33817=>"111100011",
  33818=>"110000010",
  33819=>"111101110",
  33820=>"011000000",
  33821=>"101001011",
  33822=>"001111010",
  33823=>"011000001",
  33824=>"110100101",
  33825=>"000100100",
  33826=>"100111000",
  33827=>"100111000",
  33828=>"001111111",
  33829=>"001000111",
  33830=>"111110101",
  33831=>"111111010",
  33832=>"101110100",
  33833=>"011001001",
  33834=>"010011100",
  33835=>"111110101",
  33836=>"111001010",
  33837=>"110100101",
  33838=>"000110101",
  33839=>"010001000",
  33840=>"111111011",
  33841=>"101110111",
  33842=>"001111010",
  33843=>"011011000",
  33844=>"111101000",
  33845=>"000011100",
  33846=>"111011000",
  33847=>"111101111",
  33848=>"001100110",
  33849=>"000000101",
  33850=>"000110011",
  33851=>"010100111",
  33852=>"010001111",
  33853=>"110111100",
  33854=>"000010110",
  33855=>"100101100",
  33856=>"100001111",
  33857=>"010101000",
  33858=>"011011100",
  33859=>"001011111",
  33860=>"001011001",
  33861=>"110110000",
  33862=>"010001111",
  33863=>"111001100",
  33864=>"111110111",
  33865=>"000001100",
  33866=>"011011010",
  33867=>"111001101",
  33868=>"101101100",
  33869=>"110100001",
  33870=>"101001101",
  33871=>"001010100",
  33872=>"101110000",
  33873=>"101101000",
  33874=>"111101001",
  33875=>"000110011",
  33876=>"111010100",
  33877=>"000001110",
  33878=>"100011111",
  33879=>"110100111",
  33880=>"000101111",
  33881=>"111101010",
  33882=>"101001110",
  33883=>"001101100",
  33884=>"111111100",
  33885=>"100001111",
  33886=>"111110011",
  33887=>"011001000",
  33888=>"111100000",
  33889=>"101110000",
  33890=>"111011001",
  33891=>"010101001",
  33892=>"101110011",
  33893=>"100110001",
  33894=>"100010000",
  33895=>"101111111",
  33896=>"111001101",
  33897=>"110110110",
  33898=>"000101010",
  33899=>"111100010",
  33900=>"001101101",
  33901=>"011111100",
  33902=>"010111001",
  33903=>"001100100",
  33904=>"101010110",
  33905=>"111111110",
  33906=>"010001110",
  33907=>"011101000",
  33908=>"001111100",
  33909=>"001010010",
  33910=>"010110001",
  33911=>"000000011",
  33912=>"000100001",
  33913=>"111001010",
  33914=>"001100100",
  33915=>"010001011",
  33916=>"000000100",
  33917=>"010100001",
  33918=>"100101000",
  33919=>"110001001",
  33920=>"000110100",
  33921=>"011001010",
  33922=>"000010100",
  33923=>"010001101",
  33924=>"001101101",
  33925=>"000111001",
  33926=>"011101100",
  33927=>"100010111",
  33928=>"000101101",
  33929=>"110011010",
  33930=>"000001001",
  33931=>"111111111",
  33932=>"001100100",
  33933=>"110011010",
  33934=>"000101011",
  33935=>"100011011",
  33936=>"010011111",
  33937=>"101100000",
  33938=>"000101011",
  33939=>"110000011",
  33940=>"001101000",
  33941=>"110111010",
  33942=>"101011101",
  33943=>"001000101",
  33944=>"111101101",
  33945=>"101101111",
  33946=>"010000100",
  33947=>"111001000",
  33948=>"110001100",
  33949=>"000100100",
  33950=>"000000001",
  33951=>"111111000",
  33952=>"010111110",
  33953=>"001001101",
  33954=>"010001111",
  33955=>"111001110",
  33956=>"000001110",
  33957=>"110011110",
  33958=>"011011111",
  33959=>"101100010",
  33960=>"100000001",
  33961=>"001011010",
  33962=>"010100001",
  33963=>"100001011",
  33964=>"110000111",
  33965=>"000000111",
  33966=>"001100101",
  33967=>"111001111",
  33968=>"110100011",
  33969=>"010011101",
  33970=>"000011101",
  33971=>"011111001",
  33972=>"010001101",
  33973=>"010001000",
  33974=>"001100000",
  33975=>"000100010",
  33976=>"000110000",
  33977=>"111010110",
  33978=>"000000001",
  33979=>"000011100",
  33980=>"100010000",
  33981=>"010000101",
  33982=>"010011001",
  33983=>"111010010",
  33984=>"100001110",
  33985=>"111011110",
  33986=>"100000000",
  33987=>"110000111",
  33988=>"101110011",
  33989=>"111101110",
  33990=>"101100110",
  33991=>"010100100",
  33992=>"101100001",
  33993=>"001001100",
  33994=>"100001000",
  33995=>"110011001",
  33996=>"001000010",
  33997=>"000001111",
  33998=>"110111110",
  33999=>"011001110",
  34000=>"001100001",
  34001=>"100010101",
  34002=>"010100000",
  34003=>"001001010",
  34004=>"111001010",
  34005=>"001011111",
  34006=>"001101010",
  34007=>"000010100",
  34008=>"111001101",
  34009=>"000010101",
  34010=>"101111111",
  34011=>"110000110",
  34012=>"100111100",
  34013=>"111110001",
  34014=>"000001000",
  34015=>"111000010",
  34016=>"100000110",
  34017=>"000110111",
  34018=>"100001000",
  34019=>"011001101",
  34020=>"101001111",
  34021=>"110000111",
  34022=>"010001001",
  34023=>"111101011",
  34024=>"001111101",
  34025=>"010000011",
  34026=>"110101110",
  34027=>"001001001",
  34028=>"011101000",
  34029=>"100000111",
  34030=>"101111100",
  34031=>"100010000",
  34032=>"011010000",
  34033=>"111100101",
  34034=>"111010100",
  34035=>"111011100",
  34036=>"100100111",
  34037=>"111101010",
  34038=>"100111001",
  34039=>"011010110",
  34040=>"000001001",
  34041=>"110111000",
  34042=>"011111100",
  34043=>"011100000",
  34044=>"111100000",
  34045=>"100000111",
  34046=>"010010000",
  34047=>"011010101",
  34048=>"011110110",
  34049=>"000101010",
  34050=>"010000111",
  34051=>"000011001",
  34052=>"000000001",
  34053=>"010111011",
  34054=>"011100011",
  34055=>"010111101",
  34056=>"101000111",
  34057=>"111000100",
  34058=>"001010000",
  34059=>"110001100",
  34060=>"110110010",
  34061=>"110011010",
  34062=>"100000011",
  34063=>"001001110",
  34064=>"100111101",
  34065=>"000111011",
  34066=>"001101110",
  34067=>"000100100",
  34068=>"110011100",
  34069=>"111111111",
  34070=>"010101111",
  34071=>"101000010",
  34072=>"111100111",
  34073=>"001101111",
  34074=>"100000010",
  34075=>"111110100",
  34076=>"100000011",
  34077=>"110001100",
  34078=>"111000110",
  34079=>"000111000",
  34080=>"101011101",
  34081=>"110100001",
  34082=>"110110110",
  34083=>"110100110",
  34084=>"110010111",
  34085=>"110001111",
  34086=>"110011000",
  34087=>"101010110",
  34088=>"101101011",
  34089=>"101111110",
  34090=>"101010001",
  34091=>"011110101",
  34092=>"101100111",
  34093=>"011001001",
  34094=>"000011000",
  34095=>"010110100",
  34096=>"110001001",
  34097=>"010001001",
  34098=>"001010011",
  34099=>"000001011",
  34100=>"001000000",
  34101=>"000101101",
  34102=>"011100000",
  34103=>"101110000",
  34104=>"010100110",
  34105=>"110011110",
  34106=>"010011010",
  34107=>"001100000",
  34108=>"010011101",
  34109=>"110110001",
  34110=>"111011110",
  34111=>"010000110",
  34112=>"100010110",
  34113=>"110101011",
  34114=>"101011011",
  34115=>"010101111",
  34116=>"000001111",
  34117=>"110111010",
  34118=>"001101001",
  34119=>"111001011",
  34120=>"011010000",
  34121=>"010011011",
  34122=>"100100000",
  34123=>"010100111",
  34124=>"001011110",
  34125=>"010010010",
  34126=>"010110010",
  34127=>"001100111",
  34128=>"111011010",
  34129=>"011100000",
  34130=>"001100011",
  34131=>"100111111",
  34132=>"010000111",
  34133=>"110001011",
  34134=>"101010100",
  34135=>"110110010",
  34136=>"110011111",
  34137=>"110000110",
  34138=>"100011111",
  34139=>"111000001",
  34140=>"010100001",
  34141=>"100100111",
  34142=>"100000011",
  34143=>"011111110",
  34144=>"110000000",
  34145=>"110101011",
  34146=>"010100100",
  34147=>"101101011",
  34148=>"100000001",
  34149=>"100110110",
  34150=>"100101101",
  34151=>"101010010",
  34152=>"101011111",
  34153=>"111010010",
  34154=>"010001110",
  34155=>"010000011",
  34156=>"001101011",
  34157=>"000100000",
  34158=>"111001000",
  34159=>"001000111",
  34160=>"100001110",
  34161=>"111010001",
  34162=>"000000000",
  34163=>"100100000",
  34164=>"001001110",
  34165=>"011001000",
  34166=>"111101001",
  34167=>"000101011",
  34168=>"100010110",
  34169=>"001010011",
  34170=>"011001000",
  34171=>"111110011",
  34172=>"011001001",
  34173=>"110011011",
  34174=>"001001110",
  34175=>"010101010",
  34176=>"001110001",
  34177=>"000101111",
  34178=>"010110100",
  34179=>"110110010",
  34180=>"100001100",
  34181=>"111010001",
  34182=>"101110000",
  34183=>"010000010",
  34184=>"111101011",
  34185=>"101011011",
  34186=>"110010111",
  34187=>"011111101",
  34188=>"001011010",
  34189=>"111100110",
  34190=>"100001000",
  34191=>"111111000",
  34192=>"100000011",
  34193=>"111001101",
  34194=>"101010110",
  34195=>"010111000",
  34196=>"000011100",
  34197=>"000001001",
  34198=>"000110101",
  34199=>"100110100",
  34200=>"001101100",
  34201=>"001101011",
  34202=>"010001000",
  34203=>"110000111",
  34204=>"010101101",
  34205=>"101010011",
  34206=>"100000000",
  34207=>"010001010",
  34208=>"001111001",
  34209=>"101001101",
  34210=>"101010010",
  34211=>"001111101",
  34212=>"010101001",
  34213=>"001110111",
  34214=>"101001110",
  34215=>"001110111",
  34216=>"110110010",
  34217=>"000000110",
  34218=>"101000111",
  34219=>"011000010",
  34220=>"000011010",
  34221=>"011110110",
  34222=>"110111100",
  34223=>"111010000",
  34224=>"011010001",
  34225=>"000000111",
  34226=>"101111110",
  34227=>"011011111",
  34228=>"100100001",
  34229=>"000010010",
  34230=>"110010111",
  34231=>"001101110",
  34232=>"111101101",
  34233=>"001001000",
  34234=>"110110010",
  34235=>"010110001",
  34236=>"001100010",
  34237=>"000011111",
  34238=>"010110111",
  34239=>"000101100",
  34240=>"011011001",
  34241=>"000000111",
  34242=>"101101000",
  34243=>"101101110",
  34244=>"000000010",
  34245=>"010100001",
  34246=>"111110000",
  34247=>"111000000",
  34248=>"011110111",
  34249=>"000101100",
  34250=>"100000100",
  34251=>"001011010",
  34252=>"101100101",
  34253=>"000101100",
  34254=>"000001011",
  34255=>"000010001",
  34256=>"010100110",
  34257=>"011011100",
  34258=>"010010001",
  34259=>"001111001",
  34260=>"001111000",
  34261=>"010000010",
  34262=>"100001000",
  34263=>"001011100",
  34264=>"000100001",
  34265=>"111101010",
  34266=>"101000111",
  34267=>"110001111",
  34268=>"101000001",
  34269=>"101001110",
  34270=>"011100100",
  34271=>"010000111",
  34272=>"001110000",
  34273=>"000001111",
  34274=>"011001000",
  34275=>"110000100",
  34276=>"000111001",
  34277=>"101001011",
  34278=>"111111001",
  34279=>"010011110",
  34280=>"111101001",
  34281=>"111100000",
  34282=>"011010000",
  34283=>"101011001",
  34284=>"100111000",
  34285=>"011100000",
  34286=>"111101110",
  34287=>"011010101",
  34288=>"000111001",
  34289=>"110101010",
  34290=>"100000111",
  34291=>"001110100",
  34292=>"100110100",
  34293=>"011010010",
  34294=>"011010010",
  34295=>"111101011",
  34296=>"000010001",
  34297=>"011101010",
  34298=>"100110100",
  34299=>"001000011",
  34300=>"000010111",
  34301=>"010000001",
  34302=>"000101010",
  34303=>"011000000",
  34304=>"010101011",
  34305=>"010010111",
  34306=>"011010000",
  34307=>"010100100",
  34308=>"101011000",
  34309=>"001011011",
  34310=>"111111001",
  34311=>"000011010",
  34312=>"010101100",
  34313=>"000101101",
  34314=>"111111101",
  34315=>"000010100",
  34316=>"000100100",
  34317=>"111101111",
  34318=>"101001110",
  34319=>"101101001",
  34320=>"010100100",
  34321=>"110101101",
  34322=>"111101110",
  34323=>"000010010",
  34324=>"111100000",
  34325=>"101111010",
  34326=>"001010001",
  34327=>"000110010",
  34328=>"111110100",
  34329=>"111110111",
  34330=>"100111100",
  34331=>"110000111",
  34332=>"010011011",
  34333=>"000000010",
  34334=>"101001111",
  34335=>"000000110",
  34336=>"110000101",
  34337=>"110101110",
  34338=>"111100101",
  34339=>"111101110",
  34340=>"111000111",
  34341=>"000000001",
  34342=>"111111000",
  34343=>"110011000",
  34344=>"111101011",
  34345=>"001011011",
  34346=>"010010011",
  34347=>"001001011",
  34348=>"111111110",
  34349=>"001001011",
  34350=>"010000010",
  34351=>"100110011",
  34352=>"001111111",
  34353=>"000100000",
  34354=>"010000100",
  34355=>"101011111",
  34356=>"000101101",
  34357=>"011110111",
  34358=>"100110100",
  34359=>"111011110",
  34360=>"011010101",
  34361=>"010000000",
  34362=>"101010100",
  34363=>"101100011",
  34364=>"011001100",
  34365=>"011011011",
  34366=>"110100010",
  34367=>"110100100",
  34368=>"101101010",
  34369=>"010001011",
  34370=>"001101001",
  34371=>"000110000",
  34372=>"011111101",
  34373=>"100001100",
  34374=>"100100110",
  34375=>"110110100",
  34376=>"000110011",
  34377=>"011000011",
  34378=>"110101001",
  34379=>"010001000",
  34380=>"100001010",
  34381=>"101000000",
  34382=>"011011011",
  34383=>"111110011",
  34384=>"110101111",
  34385=>"010000100",
  34386=>"011001000",
  34387=>"111001100",
  34388=>"011101100",
  34389=>"000010001",
  34390=>"111000001",
  34391=>"000011010",
  34392=>"110110010",
  34393=>"000111101",
  34394=>"100001010",
  34395=>"111110001",
  34396=>"111101011",
  34397=>"101000010",
  34398=>"000101000",
  34399=>"001011111",
  34400=>"011110101",
  34401=>"101001011",
  34402=>"011100000",
  34403=>"110101001",
  34404=>"111011000",
  34405=>"010011011",
  34406=>"010110101",
  34407=>"111011100",
  34408=>"111010010",
  34409=>"011001110",
  34410=>"010101100",
  34411=>"001110001",
  34412=>"101101110",
  34413=>"100111111",
  34414=>"101001001",
  34415=>"001000000",
  34416=>"111000001",
  34417=>"100101111",
  34418=>"111000000",
  34419=>"000011010",
  34420=>"000001011",
  34421=>"100111101",
  34422=>"110111000",
  34423=>"010000100",
  34424=>"011110111",
  34425=>"100011110",
  34426=>"011110100",
  34427=>"110100110",
  34428=>"010001001",
  34429=>"000001111",
  34430=>"001000001",
  34431=>"001100000",
  34432=>"000001101",
  34433=>"000101010",
  34434=>"011101001",
  34435=>"111110111",
  34436=>"001010110",
  34437=>"110010111",
  34438=>"011010101",
  34439=>"010111100",
  34440=>"111010110",
  34441=>"101110010",
  34442=>"111001101",
  34443=>"111111000",
  34444=>"111111001",
  34445=>"000100000",
  34446=>"101011110",
  34447=>"110011000",
  34448=>"000111110",
  34449=>"111011111",
  34450=>"010000101",
  34451=>"011111011",
  34452=>"010001010",
  34453=>"010101110",
  34454=>"101010110",
  34455=>"101100101",
  34456=>"110111001",
  34457=>"100110001",
  34458=>"001111100",
  34459=>"100001110",
  34460=>"001011111",
  34461=>"001011001",
  34462=>"010000001",
  34463=>"111001010",
  34464=>"011001100",
  34465=>"111010110",
  34466=>"000100000",
  34467=>"110110110",
  34468=>"111011100",
  34469=>"000000101",
  34470=>"101001001",
  34471=>"011111111",
  34472=>"111100011",
  34473=>"001110111",
  34474=>"101001010",
  34475=>"100011110",
  34476=>"111111001",
  34477=>"101001100",
  34478=>"010100100",
  34479=>"111111000",
  34480=>"110001101",
  34481=>"000111101",
  34482=>"111111100",
  34483=>"001000101",
  34484=>"101010101",
  34485=>"010000101",
  34486=>"000101011",
  34487=>"010101100",
  34488=>"110100101",
  34489=>"010100010",
  34490=>"110100011",
  34491=>"001001101",
  34492=>"101001100",
  34493=>"111111001",
  34494=>"001000011",
  34495=>"111001011",
  34496=>"010001100",
  34497=>"010001011",
  34498=>"000101000",
  34499=>"011011010",
  34500=>"110000000",
  34501=>"001010011",
  34502=>"011101000",
  34503=>"100100001",
  34504=>"010110110",
  34505=>"110000001",
  34506=>"111000101",
  34507=>"000010001",
  34508=>"110111000",
  34509=>"111000111",
  34510=>"011100001",
  34511=>"010000000",
  34512=>"000001100",
  34513=>"000110110",
  34514=>"111000100",
  34515=>"110001110",
  34516=>"110111111",
  34517=>"110001000",
  34518=>"111110011",
  34519=>"100001011",
  34520=>"011110011",
  34521=>"111011110",
  34522=>"001001100",
  34523=>"110010010",
  34524=>"011011001",
  34525=>"111000000",
  34526=>"101110110",
  34527=>"110100110",
  34528=>"110000011",
  34529=>"010100001",
  34530=>"110110011",
  34531=>"010101111",
  34532=>"110111100",
  34533=>"111101000",
  34534=>"011100111",
  34535=>"000000111",
  34536=>"000101000",
  34537=>"101011001",
  34538=>"100110001",
  34539=>"010100011",
  34540=>"100000010",
  34541=>"110001011",
  34542=>"111010010",
  34543=>"010011000",
  34544=>"100101010",
  34545=>"000011001",
  34546=>"011010110",
  34547=>"000000000",
  34548=>"010010000",
  34549=>"011010100",
  34550=>"000110001",
  34551=>"101111011",
  34552=>"011100001",
  34553=>"110100111",
  34554=>"010100001",
  34555=>"100000000",
  34556=>"101100110",
  34557=>"010011010",
  34558=>"101101010",
  34559=>"100110000",
  34560=>"101010010",
  34561=>"011010100",
  34562=>"011001111",
  34563=>"000100001",
  34564=>"011111100",
  34565=>"101110111",
  34566=>"110111100",
  34567=>"001010101",
  34568=>"010100001",
  34569=>"101110001",
  34570=>"111100010",
  34571=>"000010100",
  34572=>"101010000",
  34573=>"110000001",
  34574=>"000011100",
  34575=>"110010100",
  34576=>"001110011",
  34577=>"011001000",
  34578=>"001000001",
  34579=>"110100101",
  34580=>"100010000",
  34581=>"111111101",
  34582=>"110100100",
  34583=>"001101011",
  34584=>"101111010",
  34585=>"001001011",
  34586=>"000111111",
  34587=>"100010100",
  34588=>"011110110",
  34589=>"001010010",
  34590=>"000110011",
  34591=>"110101001",
  34592=>"010011010",
  34593=>"100011000",
  34594=>"001011101",
  34595=>"000001001",
  34596=>"001100101",
  34597=>"001000000",
  34598=>"110110100",
  34599=>"010000110",
  34600=>"010111001",
  34601=>"100101010",
  34602=>"000011101",
  34603=>"101000110",
  34604=>"001000001",
  34605=>"000010000",
  34606=>"001001101",
  34607=>"000011000",
  34608=>"000100111",
  34609=>"010111100",
  34610=>"000011101",
  34611=>"101110111",
  34612=>"001010000",
  34613=>"110111100",
  34614=>"111000011",
  34615=>"010011100",
  34616=>"100010010",
  34617=>"010001111",
  34618=>"111100010",
  34619=>"100100000",
  34620=>"010011111",
  34621=>"000000101",
  34622=>"101000010",
  34623=>"111110101",
  34624=>"101110111",
  34625=>"101100100",
  34626=>"101011110",
  34627=>"010011000",
  34628=>"011101100",
  34629=>"111111101",
  34630=>"111101010",
  34631=>"010001011",
  34632=>"010001101",
  34633=>"101011101",
  34634=>"010011111",
  34635=>"011000001",
  34636=>"011000111",
  34637=>"111010000",
  34638=>"011001111",
  34639=>"010100100",
  34640=>"100011001",
  34641=>"100100110",
  34642=>"111101100",
  34643=>"101011111",
  34644=>"111110110",
  34645=>"111000111",
  34646=>"101101011",
  34647=>"010100111",
  34648=>"011011100",
  34649=>"101000010",
  34650=>"000101001",
  34651=>"011010101",
  34652=>"100111001",
  34653=>"111011110",
  34654=>"010001101",
  34655=>"001111011",
  34656=>"100101001",
  34657=>"010000001",
  34658=>"101100101",
  34659=>"101110100",
  34660=>"111011110",
  34661=>"001001011",
  34662=>"000000010",
  34663=>"000100110",
  34664=>"001000110",
  34665=>"000011111",
  34666=>"100101000",
  34667=>"011100110",
  34668=>"100111100",
  34669=>"100010110",
  34670=>"001100000",
  34671=>"110000000",
  34672=>"101011001",
  34673=>"000111010",
  34674=>"110000000",
  34675=>"101001000",
  34676=>"000100000",
  34677=>"100111011",
  34678=>"010100010",
  34679=>"101001100",
  34680=>"001101101",
  34681=>"000111101",
  34682=>"011101010",
  34683=>"100101011",
  34684=>"001010000",
  34685=>"111000110",
  34686=>"110010001",
  34687=>"011110111",
  34688=>"000011101",
  34689=>"110000010",
  34690=>"101111011",
  34691=>"011111111",
  34692=>"100000000",
  34693=>"110111000",
  34694=>"011111011",
  34695=>"010011001",
  34696=>"100110011",
  34697=>"100000100",
  34698=>"000100001",
  34699=>"001000001",
  34700=>"100001000",
  34701=>"110001000",
  34702=>"001010000",
  34703=>"001010100",
  34704=>"101101011",
  34705=>"110000101",
  34706=>"111000111",
  34707=>"000001000",
  34708=>"101101110",
  34709=>"101101001",
  34710=>"001011101",
  34711=>"001011000",
  34712=>"011111001",
  34713=>"110011001",
  34714=>"011111101",
  34715=>"001011100",
  34716=>"001001010",
  34717=>"001110110",
  34718=>"000101101",
  34719=>"101000111",
  34720=>"101110111",
  34721=>"110011101",
  34722=>"100001000",
  34723=>"101100101",
  34724=>"100101000",
  34725=>"101010100",
  34726=>"011011010",
  34727=>"000010111",
  34728=>"101011101",
  34729=>"000101011",
  34730=>"110110010",
  34731=>"101001001",
  34732=>"111110111",
  34733=>"110010011",
  34734=>"011001011",
  34735=>"110010001",
  34736=>"011100010",
  34737=>"001111111",
  34738=>"001000000",
  34739=>"100100011",
  34740=>"111111100",
  34741=>"010010100",
  34742=>"011001010",
  34743=>"101110011",
  34744=>"000001001",
  34745=>"101100111",
  34746=>"000111000",
  34747=>"110110101",
  34748=>"100100001",
  34749=>"010000100",
  34750=>"010110110",
  34751=>"001001001",
  34752=>"111000101",
  34753=>"010000011",
  34754=>"010100000",
  34755=>"010100100",
  34756=>"000111010",
  34757=>"111101011",
  34758=>"001000100",
  34759=>"000111101",
  34760=>"101100010",
  34761=>"010100000",
  34762=>"011011100",
  34763=>"001001100",
  34764=>"111001011",
  34765=>"100000111",
  34766=>"110001001",
  34767=>"001111111",
  34768=>"001010111",
  34769=>"111100011",
  34770=>"100011000",
  34771=>"010001111",
  34772=>"111100001",
  34773=>"101101100",
  34774=>"011111010",
  34775=>"101000100",
  34776=>"111111100",
  34777=>"111000111",
  34778=>"111110111",
  34779=>"100000001",
  34780=>"001001101",
  34781=>"100110011",
  34782=>"111011100",
  34783=>"001110000",
  34784=>"001111010",
  34785=>"011001101",
  34786=>"101000110",
  34787=>"000001111",
  34788=>"000011010",
  34789=>"111100111",
  34790=>"100000111",
  34791=>"011111110",
  34792=>"100110111",
  34793=>"110111111",
  34794=>"010011111",
  34795=>"001110011",
  34796=>"010011110",
  34797=>"000111110",
  34798=>"000110110",
  34799=>"101101001",
  34800=>"100100111",
  34801=>"111101101",
  34802=>"011011110",
  34803=>"011101101",
  34804=>"011001111",
  34805=>"000010000",
  34806=>"111110011",
  34807=>"011101100",
  34808=>"000011100",
  34809=>"101110000",
  34810=>"110000110",
  34811=>"111111110",
  34812=>"110000011",
  34813=>"100101011",
  34814=>"101011111",
  34815=>"011000111",
  34816=>"110101001",
  34817=>"000111000",
  34818=>"001010101",
  34819=>"010110011",
  34820=>"111010110",
  34821=>"000101100",
  34822=>"011001111",
  34823=>"100000010",
  34824=>"011101000",
  34825=>"110000101",
  34826=>"010100000",
  34827=>"110001011",
  34828=>"110011010",
  34829=>"110000001",
  34830=>"110111111",
  34831=>"010000001",
  34832=>"011000101",
  34833=>"011110101",
  34834=>"000001110",
  34835=>"100100010",
  34836=>"110010001",
  34837=>"010000001",
  34838=>"011011101",
  34839=>"101000011",
  34840=>"001001110",
  34841=>"010110011",
  34842=>"001000100",
  34843=>"011101100",
  34844=>"101101001",
  34845=>"011011011",
  34846=>"110111011",
  34847=>"110101100",
  34848=>"000000100",
  34849=>"111101111",
  34850=>"100111001",
  34851=>"101110010",
  34852=>"011000010",
  34853=>"011110111",
  34854=>"111110111",
  34855=>"101010101",
  34856=>"011111000",
  34857=>"110111000",
  34858=>"010000011",
  34859=>"111111101",
  34860=>"111101111",
  34861=>"111101110",
  34862=>"111110001",
  34863=>"001111010",
  34864=>"111000101",
  34865=>"110000001",
  34866=>"001011001",
  34867=>"111000001",
  34868=>"101000100",
  34869=>"000110111",
  34870=>"000111101",
  34871=>"100110000",
  34872=>"000010001",
  34873=>"111101101",
  34874=>"000000110",
  34875=>"011010110",
  34876=>"010010100",
  34877=>"000011001",
  34878=>"111000100",
  34879=>"100001110",
  34880=>"101100011",
  34881=>"100110000",
  34882=>"100101100",
  34883=>"011011110",
  34884=>"011111101",
  34885=>"011010010",
  34886=>"001011010",
  34887=>"111110111",
  34888=>"100100111",
  34889=>"100100010",
  34890=>"011010110",
  34891=>"011000011",
  34892=>"100000101",
  34893=>"011110000",
  34894=>"011000001",
  34895=>"010100010",
  34896=>"111101010",
  34897=>"000100110",
  34898=>"101010111",
  34899=>"101010001",
  34900=>"010111011",
  34901=>"010101000",
  34902=>"110100010",
  34903=>"101100110",
  34904=>"011101011",
  34905=>"110011010",
  34906=>"010110000",
  34907=>"010000100",
  34908=>"001011111",
  34909=>"110100111",
  34910=>"111001100",
  34911=>"100000000",
  34912=>"100100111",
  34913=>"010000010",
  34914=>"111010011",
  34915=>"110011011",
  34916=>"001100011",
  34917=>"011111111",
  34918=>"100101100",
  34919=>"000110111",
  34920=>"011010110",
  34921=>"010110000",
  34922=>"000001100",
  34923=>"100101001",
  34924=>"000100101",
  34925=>"000010100",
  34926=>"110000000",
  34927=>"001111010",
  34928=>"000001010",
  34929=>"011100110",
  34930=>"010100000",
  34931=>"010011110",
  34932=>"001111100",
  34933=>"000001010",
  34934=>"101001011",
  34935=>"000110111",
  34936=>"000110011",
  34937=>"110110011",
  34938=>"110000010",
  34939=>"100101110",
  34940=>"010110101",
  34941=>"000100100",
  34942=>"010111001",
  34943=>"101001111",
  34944=>"111010000",
  34945=>"111010010",
  34946=>"011011100",
  34947=>"110001011",
  34948=>"001000010",
  34949=>"111101101",
  34950=>"001011000",
  34951=>"000001100",
  34952=>"111100100",
  34953=>"010101110",
  34954=>"101010010",
  34955=>"001010110",
  34956=>"100110011",
  34957=>"100001000",
  34958=>"011110100",
  34959=>"011000101",
  34960=>"000110000",
  34961=>"000000001",
  34962=>"101101011",
  34963=>"111110011",
  34964=>"000000101",
  34965=>"110100101",
  34966=>"010010000",
  34967=>"000010101",
  34968=>"010010100",
  34969=>"001000001",
  34970=>"111010011",
  34971=>"000111101",
  34972=>"110110011",
  34973=>"000011001",
  34974=>"011011011",
  34975=>"001000010",
  34976=>"111100000",
  34977=>"100110000",
  34978=>"001011110",
  34979=>"001011011",
  34980=>"110111000",
  34981=>"000001110",
  34982=>"100110110",
  34983=>"011001011",
  34984=>"110101100",
  34985=>"000111110",
  34986=>"100011110",
  34987=>"011011001",
  34988=>"000011111",
  34989=>"110101000",
  34990=>"000000001",
  34991=>"101110011",
  34992=>"000011010",
  34993=>"101101101",
  34994=>"100001010",
  34995=>"010000110",
  34996=>"100110001",
  34997=>"101101110",
  34998=>"001111100",
  34999=>"010100101",
  35000=>"000111000",
  35001=>"001110011",
  35002=>"001000100",
  35003=>"100111101",
  35004=>"010001110",
  35005=>"110001010",
  35006=>"100100001",
  35007=>"101000001",
  35008=>"000100110",
  35009=>"000010110",
  35010=>"110001000",
  35011=>"100101101",
  35012=>"001011001",
  35013=>"001111010",
  35014=>"001011110",
  35015=>"111110011",
  35016=>"100110010",
  35017=>"011001101",
  35018=>"010001000",
  35019=>"011001001",
  35020=>"100110010",
  35021=>"010110010",
  35022=>"111100101",
  35023=>"011000111",
  35024=>"100001101",
  35025=>"000101010",
  35026=>"000000010",
  35027=>"001001110",
  35028=>"100000011",
  35029=>"001010101",
  35030=>"000111011",
  35031=>"100111000",
  35032=>"110100000",
  35033=>"100000101",
  35034=>"001101011",
  35035=>"000000010",
  35036=>"001000011",
  35037=>"101100000",
  35038=>"010010000",
  35039=>"100111111",
  35040=>"001001010",
  35041=>"001000010",
  35042=>"101010100",
  35043=>"010001111",
  35044=>"111001010",
  35045=>"101011100",
  35046=>"111101010",
  35047=>"001001000",
  35048=>"111001111",
  35049=>"111011011",
  35050=>"100011011",
  35051=>"010111011",
  35052=>"011100111",
  35053=>"110110101",
  35054=>"000100111",
  35055=>"011010100",
  35056=>"101101111",
  35057=>"011111110",
  35058=>"100101011",
  35059=>"011111101",
  35060=>"101000101",
  35061=>"110100100",
  35062=>"100111000",
  35063=>"100110011",
  35064=>"011101001",
  35065=>"001110110",
  35066=>"011111001",
  35067=>"001000000",
  35068=>"111101101",
  35069=>"100110001",
  35070=>"001100111",
  35071=>"111001011",
  35072=>"010110001",
  35073=>"110001001",
  35074=>"011101111",
  35075=>"011001111",
  35076=>"100010100",
  35077=>"011110100",
  35078=>"010000000",
  35079=>"110001111",
  35080=>"111110011",
  35081=>"111111110",
  35082=>"111001011",
  35083=>"101010110",
  35084=>"100100001",
  35085=>"011111110",
  35086=>"011011011",
  35087=>"000001010",
  35088=>"000000000",
  35089=>"111111100",
  35090=>"110101000",
  35091=>"000001100",
  35092=>"100101111",
  35093=>"000100010",
  35094=>"011011101",
  35095=>"111001001",
  35096=>"111001001",
  35097=>"100010101",
  35098=>"110001110",
  35099=>"000000000",
  35100=>"110000110",
  35101=>"101100101",
  35102=>"010000111",
  35103=>"000111000",
  35104=>"001010100",
  35105=>"011100111",
  35106=>"001111111",
  35107=>"100100111",
  35108=>"000100000",
  35109=>"101100011",
  35110=>"110100101",
  35111=>"101101100",
  35112=>"100000100",
  35113=>"110101000",
  35114=>"011011100",
  35115=>"000011101",
  35116=>"010111110",
  35117=>"110000001",
  35118=>"000000010",
  35119=>"000100100",
  35120=>"011110110",
  35121=>"001010000",
  35122=>"110011110",
  35123=>"100010011",
  35124=>"101001010",
  35125=>"001110000",
  35126=>"111010010",
  35127=>"010000111",
  35128=>"110000010",
  35129=>"010110011",
  35130=>"000010111",
  35131=>"110110001",
  35132=>"100000101",
  35133=>"101011100",
  35134=>"010111001",
  35135=>"111000110",
  35136=>"000011100",
  35137=>"101100100",
  35138=>"100000011",
  35139=>"110110010",
  35140=>"110000111",
  35141=>"010010100",
  35142=>"000000000",
  35143=>"000011000",
  35144=>"010011000",
  35145=>"011010000",
  35146=>"001000110",
  35147=>"100101011",
  35148=>"010110000",
  35149=>"010111110",
  35150=>"001011010",
  35151=>"011011011",
  35152=>"010001101",
  35153=>"110001100",
  35154=>"111111001",
  35155=>"010110100",
  35156=>"110110010",
  35157=>"111000000",
  35158=>"110101111",
  35159=>"110010010",
  35160=>"001101001",
  35161=>"100001111",
  35162=>"011001001",
  35163=>"010001000",
  35164=>"111110110",
  35165=>"100110111",
  35166=>"100001110",
  35167=>"001110011",
  35168=>"111010000",
  35169=>"101010011",
  35170=>"000000010",
  35171=>"000001001",
  35172=>"011001010",
  35173=>"010001111",
  35174=>"001010100",
  35175=>"001110001",
  35176=>"000110110",
  35177=>"011111000",
  35178=>"111011101",
  35179=>"001100101",
  35180=>"001010001",
  35181=>"100001101",
  35182=>"101001010",
  35183=>"010100001",
  35184=>"110110111",
  35185=>"000110101",
  35186=>"000000000",
  35187=>"110101111",
  35188=>"110011010",
  35189=>"010101000",
  35190=>"110010010",
  35191=>"000111111",
  35192=>"000000000",
  35193=>"100010011",
  35194=>"101101011",
  35195=>"001001100",
  35196=>"100101001",
  35197=>"011001101",
  35198=>"000011000",
  35199=>"101111010",
  35200=>"101001110",
  35201=>"000011111",
  35202=>"000110110",
  35203=>"011010010",
  35204=>"110100001",
  35205=>"001001001",
  35206=>"111101110",
  35207=>"110011000",
  35208=>"001001000",
  35209=>"011101001",
  35210=>"111011000",
  35211=>"010010101",
  35212=>"100000100",
  35213=>"010110010",
  35214=>"110111101",
  35215=>"001010111",
  35216=>"110001111",
  35217=>"110110010",
  35218=>"110110010",
  35219=>"111111111",
  35220=>"111000000",
  35221=>"001000101",
  35222=>"000010011",
  35223=>"101100011",
  35224=>"011001110",
  35225=>"001111010",
  35226=>"000010011",
  35227=>"111011000",
  35228=>"001001100",
  35229=>"000110100",
  35230=>"001100110",
  35231=>"111101100",
  35232=>"110010000",
  35233=>"110101110",
  35234=>"010101111",
  35235=>"100100100",
  35236=>"011010101",
  35237=>"000100100",
  35238=>"000101111",
  35239=>"011111001",
  35240=>"110000100",
  35241=>"111010100",
  35242=>"000101011",
  35243=>"110100000",
  35244=>"010111110",
  35245=>"110000011",
  35246=>"101110111",
  35247=>"101010110",
  35248=>"010101111",
  35249=>"000001010",
  35250=>"101000000",
  35251=>"101010010",
  35252=>"111111010",
  35253=>"110010011",
  35254=>"000100101",
  35255=>"100001111",
  35256=>"101110101",
  35257=>"001001000",
  35258=>"010010010",
  35259=>"010100101",
  35260=>"100111010",
  35261=>"001010010",
  35262=>"101000011",
  35263=>"100000111",
  35264=>"100010110",
  35265=>"000001011",
  35266=>"111000011",
  35267=>"101001000",
  35268=>"111101100",
  35269=>"001011011",
  35270=>"011001101",
  35271=>"110010110",
  35272=>"110101101",
  35273=>"001001001",
  35274=>"101111011",
  35275=>"000011110",
  35276=>"110011001",
  35277=>"100100011",
  35278=>"110001001",
  35279=>"000001101",
  35280=>"010001001",
  35281=>"001001001",
  35282=>"010000000",
  35283=>"001010001",
  35284=>"111001001",
  35285=>"101010110",
  35286=>"101010011",
  35287=>"011000011",
  35288=>"110010111",
  35289=>"111110101",
  35290=>"101111010",
  35291=>"101001010",
  35292=>"110100101",
  35293=>"101101011",
  35294=>"001001010",
  35295=>"100100111",
  35296=>"101100100",
  35297=>"011011000",
  35298=>"001001001",
  35299=>"101101111",
  35300=>"110101001",
  35301=>"011110000",
  35302=>"111110100",
  35303=>"010001011",
  35304=>"001001010",
  35305=>"010010011",
  35306=>"001111111",
  35307=>"010111000",
  35308=>"011000100",
  35309=>"101010001",
  35310=>"110010011",
  35311=>"101111111",
  35312=>"010001000",
  35313=>"111010010",
  35314=>"101111010",
  35315=>"000000011",
  35316=>"000001010",
  35317=>"101111000",
  35318=>"101110110",
  35319=>"100000111",
  35320=>"011001010",
  35321=>"101000010",
  35322=>"011110110",
  35323=>"000010010",
  35324=>"100000000",
  35325=>"010010001",
  35326=>"010111101",
  35327=>"001101110",
  35328=>"011001110",
  35329=>"101010100",
  35330=>"000101101",
  35331=>"010110000",
  35332=>"100011000",
  35333=>"001110111",
  35334=>"011101010",
  35335=>"001101101",
  35336=>"010100111",
  35337=>"010000101",
  35338=>"100010000",
  35339=>"001011011",
  35340=>"111111110",
  35341=>"010101010",
  35342=>"000001100",
  35343=>"100010001",
  35344=>"001000100",
  35345=>"001001100",
  35346=>"000010000",
  35347=>"111000011",
  35348=>"100101100",
  35349=>"010001110",
  35350=>"101111101",
  35351=>"001101110",
  35352=>"100110001",
  35353=>"110001101",
  35354=>"010000110",
  35355=>"110011000",
  35356=>"000000100",
  35357=>"101010000",
  35358=>"100001101",
  35359=>"001010110",
  35360=>"101111010",
  35361=>"010000010",
  35362=>"000101111",
  35363=>"000001001",
  35364=>"100100010",
  35365=>"101000100",
  35366=>"100001110",
  35367=>"110011000",
  35368=>"111011110",
  35369=>"011000111",
  35370=>"101101000",
  35371=>"001011110",
  35372=>"111010010",
  35373=>"001010111",
  35374=>"100101101",
  35375=>"000011001",
  35376=>"100010000",
  35377=>"101011011",
  35378=>"110110000",
  35379=>"110111111",
  35380=>"011001010",
  35381=>"000111001",
  35382=>"011011000",
  35383=>"101101010",
  35384=>"110010111",
  35385=>"010100101",
  35386=>"000010001",
  35387=>"100010000",
  35388=>"000011001",
  35389=>"000001010",
  35390=>"010011110",
  35391=>"101000001",
  35392=>"010000000",
  35393=>"010000010",
  35394=>"100000100",
  35395=>"111011011",
  35396=>"100001110",
  35397=>"011100101",
  35398=>"000000001",
  35399=>"001001010",
  35400=>"011110111",
  35401=>"000100001",
  35402=>"010011101",
  35403=>"000100010",
  35404=>"111010010",
  35405=>"011010010",
  35406=>"011010100",
  35407=>"000001011",
  35408=>"010111011",
  35409=>"101011110",
  35410=>"110110100",
  35411=>"001101100",
  35412=>"111000001",
  35413=>"101100101",
  35414=>"111100101",
  35415=>"000101011",
  35416=>"000010111",
  35417=>"100110110",
  35418=>"101101111",
  35419=>"110110110",
  35420=>"100100110",
  35421=>"100011100",
  35422=>"101001111",
  35423=>"000011101",
  35424=>"001100101",
  35425=>"000010111",
  35426=>"101000001",
  35427=>"111001011",
  35428=>"000010011",
  35429=>"111110000",
  35430=>"000111100",
  35431=>"000011110",
  35432=>"110100101",
  35433=>"001001101",
  35434=>"110101100",
  35435=>"000000101",
  35436=>"101110011",
  35437=>"001010000",
  35438=>"000100101",
  35439=>"001111100",
  35440=>"001110010",
  35441=>"100000010",
  35442=>"111011010",
  35443=>"111010011",
  35444=>"011111110",
  35445=>"111101011",
  35446=>"110010110",
  35447=>"001101010",
  35448=>"010000011",
  35449=>"100010101",
  35450=>"001101010",
  35451=>"010111101",
  35452=>"100000110",
  35453=>"100110100",
  35454=>"000110101",
  35455=>"000010000",
  35456=>"110011110",
  35457=>"000110011",
  35458=>"010000000",
  35459=>"111000101",
  35460=>"010101011",
  35461=>"001010101",
  35462=>"110010011",
  35463=>"101111101",
  35464=>"101000111",
  35465=>"010010010",
  35466=>"101011000",
  35467=>"100110101",
  35468=>"100000101",
  35469=>"101001111",
  35470=>"000110010",
  35471=>"101011000",
  35472=>"101100010",
  35473=>"010100000",
  35474=>"000110010",
  35475=>"101000010",
  35476=>"010101001",
  35477=>"101111100",
  35478=>"010101011",
  35479=>"011111101",
  35480=>"001110111",
  35481=>"110011101",
  35482=>"110111000",
  35483=>"111110011",
  35484=>"110100000",
  35485=>"100110001",
  35486=>"110101111",
  35487=>"101000000",
  35488=>"010011100",
  35489=>"111100110",
  35490=>"110001101",
  35491=>"010011101",
  35492=>"010110110",
  35493=>"100000111",
  35494=>"100101111",
  35495=>"001001001",
  35496=>"111111111",
  35497=>"010101010",
  35498=>"101110110",
  35499=>"111000101",
  35500=>"011000011",
  35501=>"111111001",
  35502=>"100110100",
  35503=>"010000101",
  35504=>"000000110",
  35505=>"100001010",
  35506=>"010010010",
  35507=>"010101001",
  35508=>"001100000",
  35509=>"110000110",
  35510=>"001001101",
  35511=>"000011001",
  35512=>"010111010",
  35513=>"010000001",
  35514=>"111100110",
  35515=>"111000011",
  35516=>"001000010",
  35517=>"110010000",
  35518=>"000010100",
  35519=>"000010111",
  35520=>"100110101",
  35521=>"001101111",
  35522=>"001110001",
  35523=>"111001111",
  35524=>"111010110",
  35525=>"100011011",
  35526=>"011001100",
  35527=>"010010111",
  35528=>"100001100",
  35529=>"101010011",
  35530=>"100010001",
  35531=>"010011000",
  35532=>"001111000",
  35533=>"000100100",
  35534=>"010110010",
  35535=>"001101010",
  35536=>"100000000",
  35537=>"100001000",
  35538=>"110010101",
  35539=>"001100010",
  35540=>"101100101",
  35541=>"001100100",
  35542=>"000110001",
  35543=>"010011010",
  35544=>"000111111",
  35545=>"001001100",
  35546=>"011101001",
  35547=>"010011111",
  35548=>"100101101",
  35549=>"110001110",
  35550=>"100001010",
  35551=>"000010110",
  35552=>"010100100",
  35553=>"100110001",
  35554=>"010110111",
  35555=>"101101001",
  35556=>"101010000",
  35557=>"110110000",
  35558=>"000011000",
  35559=>"010000011",
  35560=>"010001000",
  35561=>"101011110",
  35562=>"111111111",
  35563=>"110010101",
  35564=>"000101101",
  35565=>"011000001",
  35566=>"111110000",
  35567=>"011001011",
  35568=>"111100000",
  35569=>"010100011",
  35570=>"001100101",
  35571=>"110001010",
  35572=>"100000000",
  35573=>"010101111",
  35574=>"010111010",
  35575=>"010001110",
  35576=>"110000001",
  35577=>"011010111",
  35578=>"010010000",
  35579=>"000001111",
  35580=>"111101000",
  35581=>"111001111",
  35582=>"001000100",
  35583=>"001000001",
  35584=>"010110000",
  35585=>"111101000",
  35586=>"000111101",
  35587=>"010001011",
  35588=>"111111101",
  35589=>"010101001",
  35590=>"001111111",
  35591=>"000000000",
  35592=>"011000101",
  35593=>"111110110",
  35594=>"001000100",
  35595=>"010010111",
  35596=>"000011111",
  35597=>"110101011",
  35598=>"100011111",
  35599=>"011100001",
  35600=>"001100010",
  35601=>"011110011",
  35602=>"011011101",
  35603=>"111110011",
  35604=>"000100101",
  35605=>"100110011",
  35606=>"100001011",
  35607=>"101111001",
  35608=>"011110001",
  35609=>"101011000",
  35610=>"001100001",
  35611=>"100111111",
  35612=>"111111111",
  35613=>"011101001",
  35614=>"111010000",
  35615=>"011011010",
  35616=>"111001011",
  35617=>"101010010",
  35618=>"010100111",
  35619=>"110110011",
  35620=>"000111101",
  35621=>"101111101",
  35622=>"010101000",
  35623=>"000000101",
  35624=>"100001010",
  35625=>"111011000",
  35626=>"010101101",
  35627=>"000010001",
  35628=>"010001100",
  35629=>"000000100",
  35630=>"111011011",
  35631=>"100001111",
  35632=>"000000000",
  35633=>"100001100",
  35634=>"111010101",
  35635=>"011010000",
  35636=>"110101001",
  35637=>"000111100",
  35638=>"110010010",
  35639=>"000000000",
  35640=>"110010000",
  35641=>"010111101",
  35642=>"101100011",
  35643=>"011101111",
  35644=>"110010001",
  35645=>"010011101",
  35646=>"010101010",
  35647=>"101110010",
  35648=>"010010010",
  35649=>"011001101",
  35650=>"011000100",
  35651=>"101011010",
  35652=>"110110010",
  35653=>"001000110",
  35654=>"111010011",
  35655=>"100010010",
  35656=>"110011100",
  35657=>"010001010",
  35658=>"110010110",
  35659=>"001011111",
  35660=>"000110001",
  35661=>"000010111",
  35662=>"011111000",
  35663=>"110011111",
  35664=>"101111011",
  35665=>"011000100",
  35666=>"110100001",
  35667=>"001010111",
  35668=>"111001111",
  35669=>"010000001",
  35670=>"101000001",
  35671=>"101011000",
  35672=>"111001001",
  35673=>"010111011",
  35674=>"100010001",
  35675=>"111001101",
  35676=>"110100111",
  35677=>"000010000",
  35678=>"001000100",
  35679=>"101111101",
  35680=>"010100110",
  35681=>"010111001",
  35682=>"100011110",
  35683=>"010110000",
  35684=>"101100110",
  35685=>"101001100",
  35686=>"010010110",
  35687=>"000110001",
  35688=>"101101001",
  35689=>"000001111",
  35690=>"001001110",
  35691=>"001111110",
  35692=>"001101110",
  35693=>"001010000",
  35694=>"101001101",
  35695=>"011001000",
  35696=>"010001010",
  35697=>"011011110",
  35698=>"111101011",
  35699=>"100011010",
  35700=>"010101100",
  35701=>"100100010",
  35702=>"111110101",
  35703=>"110010010",
  35704=>"001111110",
  35705=>"111001001",
  35706=>"001100100",
  35707=>"101000100",
  35708=>"110111001",
  35709=>"000000011",
  35710=>"011110111",
  35711=>"001111110",
  35712=>"001011110",
  35713=>"011111000",
  35714=>"111001011",
  35715=>"000111001",
  35716=>"001011000",
  35717=>"100001100",
  35718=>"110111011",
  35719=>"010100111",
  35720=>"010111111",
  35721=>"110111001",
  35722=>"100010111",
  35723=>"000000010",
  35724=>"011101100",
  35725=>"000001000",
  35726=>"101001010",
  35727=>"100111100",
  35728=>"010010111",
  35729=>"001100001",
  35730=>"010010001",
  35731=>"011011000",
  35732=>"110101111",
  35733=>"101001110",
  35734=>"100101001",
  35735=>"011111100",
  35736=>"010110111",
  35737=>"000100111",
  35738=>"000000001",
  35739=>"110010011",
  35740=>"011101010",
  35741=>"101010011",
  35742=>"011010000",
  35743=>"101000101",
  35744=>"110111100",
  35745=>"000110000",
  35746=>"110101001",
  35747=>"100001111",
  35748=>"011010100",
  35749=>"011001110",
  35750=>"110101011",
  35751=>"111110100",
  35752=>"000100111",
  35753=>"110111000",
  35754=>"010110011",
  35755=>"100101010",
  35756=>"011011010",
  35757=>"100001101",
  35758=>"110100011",
  35759=>"101101001",
  35760=>"001100111",
  35761=>"111010000",
  35762=>"100000001",
  35763=>"011110001",
  35764=>"101010111",
  35765=>"101010111",
  35766=>"110000001",
  35767=>"011001000",
  35768=>"000010110",
  35769=>"000010110",
  35770=>"010001110",
  35771=>"011001101",
  35772=>"001101100",
  35773=>"110100000",
  35774=>"000100010",
  35775=>"101010100",
  35776=>"010111010",
  35777=>"011101010",
  35778=>"111011000",
  35779=>"010100101",
  35780=>"000110110",
  35781=>"011011110",
  35782=>"110010010",
  35783=>"000011100",
  35784=>"110000000",
  35785=>"110010110",
  35786=>"011110010",
  35787=>"110010011",
  35788=>"100000101",
  35789=>"100000011",
  35790=>"011010111",
  35791=>"001111001",
  35792=>"010110001",
  35793=>"000000111",
  35794=>"001100000",
  35795=>"000110110",
  35796=>"111000111",
  35797=>"100100101",
  35798=>"110000010",
  35799=>"110101000",
  35800=>"011110011",
  35801=>"001001001",
  35802=>"100000001",
  35803=>"001111110",
  35804=>"011100100",
  35805=>"010111010",
  35806=>"101101111",
  35807=>"000001000",
  35808=>"101111100",
  35809=>"110010111",
  35810=>"000101110",
  35811=>"101110101",
  35812=>"000110100",
  35813=>"011111010",
  35814=>"001000101",
  35815=>"110100110",
  35816=>"000011001",
  35817=>"110100111",
  35818=>"101111100",
  35819=>"100101010",
  35820=>"010111110",
  35821=>"111001011",
  35822=>"000000001",
  35823=>"000100101",
  35824=>"111001000",
  35825=>"011100100",
  35826=>"101101110",
  35827=>"100111010",
  35828=>"011011011",
  35829=>"100101001",
  35830=>"001000100",
  35831=>"000100110",
  35832=>"011001101",
  35833=>"111111000",
  35834=>"000010111",
  35835=>"001011001",
  35836=>"100111001",
  35837=>"000000011",
  35838=>"100101111",
  35839=>"010010010",
  35840=>"010100101",
  35841=>"011000000",
  35842=>"111000000",
  35843=>"101000001",
  35844=>"101111110",
  35845=>"111010110",
  35846=>"101001101",
  35847=>"000000100",
  35848=>"001011111",
  35849=>"001000100",
  35850=>"101001111",
  35851=>"001011100",
  35852=>"110010001",
  35853=>"001001010",
  35854=>"011010011",
  35855=>"001101111",
  35856=>"010000111",
  35857=>"101000011",
  35858=>"000001100",
  35859=>"100110110",
  35860=>"101000010",
  35861=>"010100001",
  35862=>"101011000",
  35863=>"000000000",
  35864=>"000110110",
  35865=>"111011111",
  35866=>"011011000",
  35867=>"000011100",
  35868=>"111001010",
  35869=>"111011000",
  35870=>"011010101",
  35871=>"011010001",
  35872=>"100110111",
  35873=>"000101111",
  35874=>"110000000",
  35875=>"110110010",
  35876=>"001011100",
  35877=>"111011101",
  35878=>"110101000",
  35879=>"101100111",
  35880=>"111101000",
  35881=>"000110110",
  35882=>"100001101",
  35883=>"000110101",
  35884=>"100100010",
  35885=>"111010111",
  35886=>"011011101",
  35887=>"100010111",
  35888=>"000010010",
  35889=>"001110110",
  35890=>"100101110",
  35891=>"101000011",
  35892=>"011100111",
  35893=>"001000110",
  35894=>"001110101",
  35895=>"100010010",
  35896=>"010001111",
  35897=>"010100010",
  35898=>"000001011",
  35899=>"101110111",
  35900=>"100001011",
  35901=>"101010010",
  35902=>"010100011",
  35903=>"010101011",
  35904=>"101101001",
  35905=>"010111100",
  35906=>"010101000",
  35907=>"000100011",
  35908=>"101111101",
  35909=>"100001001",
  35910=>"011010000",
  35911=>"110010000",
  35912=>"100001000",
  35913=>"001100011",
  35914=>"100010101",
  35915=>"110000111",
  35916=>"001100011",
  35917=>"010000100",
  35918=>"110111110",
  35919=>"110110100",
  35920=>"100011110",
  35921=>"000011100",
  35922=>"110001000",
  35923=>"011010101",
  35924=>"101000111",
  35925=>"001001100",
  35926=>"100010000",
  35927=>"001001011",
  35928=>"111010010",
  35929=>"111100001",
  35930=>"011001101",
  35931=>"011100111",
  35932=>"111010111",
  35933=>"110001011",
  35934=>"000101101",
  35935=>"110110100",
  35936=>"010110100",
  35937=>"010111110",
  35938=>"001111011",
  35939=>"101000001",
  35940=>"010100010",
  35941=>"111001100",
  35942=>"000101000",
  35943=>"100011111",
  35944=>"111100100",
  35945=>"000010111",
  35946=>"111010011",
  35947=>"001110111",
  35948=>"010000000",
  35949=>"000010011",
  35950=>"001011101",
  35951=>"000100010",
  35952=>"101111010",
  35953=>"010001001",
  35954=>"110010011",
  35955=>"101110111",
  35956=>"010100110",
  35957=>"011010100",
  35958=>"010111111",
  35959=>"110000011",
  35960=>"100010110",
  35961=>"000001101",
  35962=>"100110000",
  35963=>"011100001",
  35964=>"001000110",
  35965=>"010100010",
  35966=>"000001011",
  35967=>"110000011",
  35968=>"001111011",
  35969=>"011111101",
  35970=>"101110111",
  35971=>"010001101",
  35972=>"001011111",
  35973=>"001111000",
  35974=>"100010110",
  35975=>"010000100",
  35976=>"011101100",
  35977=>"100001000",
  35978=>"010000000",
  35979=>"011110001",
  35980=>"101000100",
  35981=>"001000100",
  35982=>"101011111",
  35983=>"000100101",
  35984=>"000111010",
  35985=>"110001111",
  35986=>"100110100",
  35987=>"011001110",
  35988=>"110111100",
  35989=>"001001110",
  35990=>"101000011",
  35991=>"011001000",
  35992=>"011010000",
  35993=>"010010001",
  35994=>"100100111",
  35995=>"101111011",
  35996=>"111110110",
  35997=>"000100100",
  35998=>"110001010",
  35999=>"001011101",
  36000=>"000101100",
  36001=>"011100111",
  36002=>"001000011",
  36003=>"010110100",
  36004=>"111110000",
  36005=>"000110100",
  36006=>"101000010",
  36007=>"000101101",
  36008=>"010111110",
  36009=>"100110100",
  36010=>"011010110",
  36011=>"010000111",
  36012=>"001001101",
  36013=>"010010000",
  36014=>"010100110",
  36015=>"000100011",
  36016=>"011110100",
  36017=>"000100110",
  36018=>"111011011",
  36019=>"000011111",
  36020=>"001110101",
  36021=>"000100100",
  36022=>"101000001",
  36023=>"000101100",
  36024=>"000101010",
  36025=>"011110000",
  36026=>"010011111",
  36027=>"001110100",
  36028=>"110001110",
  36029=>"111100010",
  36030=>"101101110",
  36031=>"111011011",
  36032=>"000100011",
  36033=>"101010000",
  36034=>"110101110",
  36035=>"001111010",
  36036=>"110110010",
  36037=>"011100000",
  36038=>"000100010",
  36039=>"010001010",
  36040=>"100110011",
  36041=>"111110101",
  36042=>"010011100",
  36043=>"000010101",
  36044=>"100011011",
  36045=>"000111111",
  36046=>"101101000",
  36047=>"011010011",
  36048=>"011000011",
  36049=>"011101001",
  36050=>"001100000",
  36051=>"111101001",
  36052=>"011000101",
  36053=>"000011110",
  36054=>"001011000",
  36055=>"010110101",
  36056=>"111000100",
  36057=>"110101110",
  36058=>"001000100",
  36059=>"110010010",
  36060=>"110010011",
  36061=>"100000110",
  36062=>"100100011",
  36063=>"011001100",
  36064=>"101001100",
  36065=>"010001100",
  36066=>"010011101",
  36067=>"010101001",
  36068=>"101101011",
  36069=>"010100001",
  36070=>"110111110",
  36071=>"100010101",
  36072=>"000100000",
  36073=>"010010001",
  36074=>"101011011",
  36075=>"110011110",
  36076=>"101010111",
  36077=>"110111000",
  36078=>"010101101",
  36079=>"001001100",
  36080=>"011110100",
  36081=>"010101110",
  36082=>"110100010",
  36083=>"111111000",
  36084=>"101110100",
  36085=>"000100010",
  36086=>"110001000",
  36087=>"111000101",
  36088=>"100011101",
  36089=>"100000011",
  36090=>"010110000",
  36091=>"101001101",
  36092=>"001110111",
  36093=>"000001011",
  36094=>"001111111",
  36095=>"000100101",
  36096=>"111001011",
  36097=>"010001111",
  36098=>"100100110",
  36099=>"111010010",
  36100=>"100100000",
  36101=>"100000011",
  36102=>"101001101",
  36103=>"111011100",
  36104=>"100001100",
  36105=>"111100000",
  36106=>"111100010",
  36107=>"000000111",
  36108=>"101100011",
  36109=>"111011100",
  36110=>"010101010",
  36111=>"111001100",
  36112=>"001101101",
  36113=>"100111001",
  36114=>"100110110",
  36115=>"011101111",
  36116=>"111000001",
  36117=>"001000100",
  36118=>"101011101",
  36119=>"100100100",
  36120=>"011011110",
  36121=>"000000000",
  36122=>"111110000",
  36123=>"101110001",
  36124=>"011001101",
  36125=>"100100011",
  36126=>"101110110",
  36127=>"000000100",
  36128=>"010111110",
  36129=>"110011110",
  36130=>"011011010",
  36131=>"011100111",
  36132=>"101110101",
  36133=>"000000101",
  36134=>"101110011",
  36135=>"110101111",
  36136=>"011111011",
  36137=>"001100111",
  36138=>"111011111",
  36139=>"111010111",
  36140=>"000011000",
  36141=>"111111111",
  36142=>"110111000",
  36143=>"000011001",
  36144=>"010010011",
  36145=>"000001111",
  36146=>"011001101",
  36147=>"111001011",
  36148=>"011010111",
  36149=>"000011111",
  36150=>"100000000",
  36151=>"001011001",
  36152=>"110000001",
  36153=>"001000010",
  36154=>"100111111",
  36155=>"011011111",
  36156=>"011000101",
  36157=>"010011111",
  36158=>"111000000",
  36159=>"001101001",
  36160=>"101001111",
  36161=>"000010111",
  36162=>"101101110",
  36163=>"011001001",
  36164=>"101111010",
  36165=>"010100110",
  36166=>"011110000",
  36167=>"101110011",
  36168=>"110011000",
  36169=>"010101010",
  36170=>"111111110",
  36171=>"101010100",
  36172=>"100100101",
  36173=>"000110110",
  36174=>"011111101",
  36175=>"011011111",
  36176=>"000110011",
  36177=>"001110011",
  36178=>"011011101",
  36179=>"100001101",
  36180=>"101011001",
  36181=>"001010011",
  36182=>"100000100",
  36183=>"011101011",
  36184=>"001101010",
  36185=>"111110100",
  36186=>"111111110",
  36187=>"110010011",
  36188=>"100011101",
  36189=>"000000001",
  36190=>"010000110",
  36191=>"111010110",
  36192=>"110011100",
  36193=>"100110010",
  36194=>"100100011",
  36195=>"001111110",
  36196=>"110101010",
  36197=>"010101100",
  36198=>"011101111",
  36199=>"111111101",
  36200=>"010111011",
  36201=>"100111111",
  36202=>"000000010",
  36203=>"000011001",
  36204=>"100101010",
  36205=>"111000000",
  36206=>"100001011",
  36207=>"011101000",
  36208=>"000101001",
  36209=>"110011110",
  36210=>"010011010",
  36211=>"000001011",
  36212=>"110000101",
  36213=>"010000110",
  36214=>"110110101",
  36215=>"101001110",
  36216=>"100110000",
  36217=>"001110110",
  36218=>"110010101",
  36219=>"111110001",
  36220=>"010010100",
  36221=>"000011101",
  36222=>"010111011",
  36223=>"010001111",
  36224=>"000011010",
  36225=>"000101100",
  36226=>"010011001",
  36227=>"110111110",
  36228=>"011100011",
  36229=>"111011011",
  36230=>"000011110",
  36231=>"111101110",
  36232=>"001001110",
  36233=>"000000111",
  36234=>"111010011",
  36235=>"011000000",
  36236=>"100100111",
  36237=>"001001111",
  36238=>"110011111",
  36239=>"100010111",
  36240=>"101010000",
  36241=>"100111100",
  36242=>"111111010",
  36243=>"111000001",
  36244=>"101101111",
  36245=>"010011100",
  36246=>"000011001",
  36247=>"011010001",
  36248=>"111110101",
  36249=>"111011001",
  36250=>"001100111",
  36251=>"110010000",
  36252=>"010001101",
  36253=>"111010111",
  36254=>"000101111",
  36255=>"011100101",
  36256=>"101011011",
  36257=>"010110011",
  36258=>"110110110",
  36259=>"101000001",
  36260=>"010110010",
  36261=>"110111111",
  36262=>"100001001",
  36263=>"000111001",
  36264=>"110010000",
  36265=>"111110110",
  36266=>"011001011",
  36267=>"101111101",
  36268=>"111111001",
  36269=>"001001111",
  36270=>"110011001",
  36271=>"101101111",
  36272=>"010000110",
  36273=>"010110101",
  36274=>"100010010",
  36275=>"000111010",
  36276=>"110110011",
  36277=>"101110100",
  36278=>"101000000",
  36279=>"001000010",
  36280=>"111110011",
  36281=>"100110111",
  36282=>"011000000",
  36283=>"110111101",
  36284=>"100100100",
  36285=>"010000100",
  36286=>"111001010",
  36287=>"010101100",
  36288=>"000110110",
  36289=>"011001110",
  36290=>"110111000",
  36291=>"100110100",
  36292=>"100000000",
  36293=>"000011000",
  36294=>"000001101",
  36295=>"001001001",
  36296=>"000011000",
  36297=>"011100010",
  36298=>"000010010",
  36299=>"001010110",
  36300=>"001001101",
  36301=>"000001100",
  36302=>"000010100",
  36303=>"011011110",
  36304=>"010111001",
  36305=>"001110100",
  36306=>"010000001",
  36307=>"010000010",
  36308=>"001100110",
  36309=>"000000100",
  36310=>"011101111",
  36311=>"001101111",
  36312=>"011010110",
  36313=>"111111001",
  36314=>"100000000",
  36315=>"001000100",
  36316=>"000011000",
  36317=>"101101010",
  36318=>"001111011",
  36319=>"010010100",
  36320=>"111110101",
  36321=>"000111010",
  36322=>"111000110",
  36323=>"100011110",
  36324=>"100011100",
  36325=>"100101100",
  36326=>"001010001",
  36327=>"111010001",
  36328=>"010000110",
  36329=>"111111001",
  36330=>"111111010",
  36331=>"101000010",
  36332=>"100001000",
  36333=>"010001001",
  36334=>"011101110",
  36335=>"010011110",
  36336=>"110000011",
  36337=>"111110000",
  36338=>"101001011",
  36339=>"010000000",
  36340=>"001000110",
  36341=>"110010001",
  36342=>"001100001",
  36343=>"011110010",
  36344=>"100100010",
  36345=>"110010111",
  36346=>"010100011",
  36347=>"110100100",
  36348=>"001011001",
  36349=>"100100100",
  36350=>"011001010",
  36351=>"110101101",
  36352=>"001101110",
  36353=>"111110000",
  36354=>"000010100",
  36355=>"100101011",
  36356=>"001000110",
  36357=>"000010110",
  36358=>"100000001",
  36359=>"010011101",
  36360=>"101000011",
  36361=>"101100010",
  36362=>"100101001",
  36363=>"000110101",
  36364=>"001100100",
  36365=>"101001010",
  36366=>"100001101",
  36367=>"111010010",
  36368=>"000101100",
  36369=>"000100010",
  36370=>"001000110",
  36371=>"000011101",
  36372=>"000010111",
  36373=>"100101011",
  36374=>"111011011",
  36375=>"111101111",
  36376=>"000110011",
  36377=>"101010011",
  36378=>"011000000",
  36379=>"101011101",
  36380=>"010000110",
  36381=>"011001110",
  36382=>"011000011",
  36383=>"100101101",
  36384=>"110110110",
  36385=>"110111101",
  36386=>"000100101",
  36387=>"010011111",
  36388=>"100110110",
  36389=>"000001101",
  36390=>"000101011",
  36391=>"110010111",
  36392=>"111100001",
  36393=>"101001000",
  36394=>"101001000",
  36395=>"100111011",
  36396=>"010100100",
  36397=>"101111100",
  36398=>"100000010",
  36399=>"000010001",
  36400=>"001110110",
  36401=>"000111011",
  36402=>"111000011",
  36403=>"111110011",
  36404=>"100011000",
  36405=>"010010101",
  36406=>"111001001",
  36407=>"000101001",
  36408=>"110011111",
  36409=>"100100111",
  36410=>"001000101",
  36411=>"011000010",
  36412=>"001101001",
  36413=>"011001000",
  36414=>"001110111",
  36415=>"011110110",
  36416=>"111110100",
  36417=>"101100101",
  36418=>"000110000",
  36419=>"000100101",
  36420=>"010010111",
  36421=>"100100101",
  36422=>"001010111",
  36423=>"100010111",
  36424=>"111001001",
  36425=>"101101100",
  36426=>"011011001",
  36427=>"010011100",
  36428=>"011111101",
  36429=>"000000001",
  36430=>"011001011",
  36431=>"001000101",
  36432=>"001101110",
  36433=>"101101001",
  36434=>"010111001",
  36435=>"010110110",
  36436=>"111011100",
  36437=>"011001010",
  36438=>"100100100",
  36439=>"100011011",
  36440=>"010100100",
  36441=>"010110101",
  36442=>"001100101",
  36443=>"111011101",
  36444=>"001110001",
  36445=>"000000010",
  36446=>"000011000",
  36447=>"000111010",
  36448=>"101111110",
  36449=>"100101010",
  36450=>"100001011",
  36451=>"000101000",
  36452=>"010110100",
  36453=>"010110011",
  36454=>"010111000",
  36455=>"110101110",
  36456=>"010100010",
  36457=>"101000110",
  36458=>"111111101",
  36459=>"101100001",
  36460=>"011101001",
  36461=>"011001010",
  36462=>"101111001",
  36463=>"100011100",
  36464=>"000100001",
  36465=>"010001000",
  36466=>"011010101",
  36467=>"100010101",
  36468=>"010111101",
  36469=>"000101011",
  36470=>"111010111",
  36471=>"100000001",
  36472=>"010111111",
  36473=>"101010010",
  36474=>"001001110",
  36475=>"100101010",
  36476=>"111111001",
  36477=>"100111000",
  36478=>"000110110",
  36479=>"010100001",
  36480=>"001100010",
  36481=>"001111101",
  36482=>"111100111",
  36483=>"001100110",
  36484=>"010000010",
  36485=>"100100010",
  36486=>"111011010",
  36487=>"010000110",
  36488=>"111110000",
  36489=>"010101000",
  36490=>"010011110",
  36491=>"011111000",
  36492=>"110111111",
  36493=>"110011000",
  36494=>"011011001",
  36495=>"110101101",
  36496=>"001000000",
  36497=>"110010010",
  36498=>"010110011",
  36499=>"011010100",
  36500=>"101100010",
  36501=>"101111011",
  36502=>"010111111",
  36503=>"001110011",
  36504=>"101111111",
  36505=>"010101101",
  36506=>"100011101",
  36507=>"011111111",
  36508=>"010110110",
  36509=>"111001000",
  36510=>"011111101",
  36511=>"010111101",
  36512=>"100011010",
  36513=>"101000111",
  36514=>"110011011",
  36515=>"000100010",
  36516=>"111010100",
  36517=>"011111011",
  36518=>"000101100",
  36519=>"001000000",
  36520=>"010010011",
  36521=>"001110111",
  36522=>"100111011",
  36523=>"001101101",
  36524=>"011011110",
  36525=>"111011100",
  36526=>"110000110",
  36527=>"101000000",
  36528=>"100001010",
  36529=>"110100100",
  36530=>"101010101",
  36531=>"000100111",
  36532=>"101010010",
  36533=>"110111110",
  36534=>"100000000",
  36535=>"101101001",
  36536=>"011100101",
  36537=>"010001110",
  36538=>"001111011",
  36539=>"000011100",
  36540=>"100100111",
  36541=>"011001111",
  36542=>"100100111",
  36543=>"110110000",
  36544=>"010000111",
  36545=>"001001101",
  36546=>"110111100",
  36547=>"111000010",
  36548=>"110001100",
  36549=>"110010111",
  36550=>"100001100",
  36551=>"001110110",
  36552=>"011011010",
  36553=>"111001001",
  36554=>"010110101",
  36555=>"101001010",
  36556=>"110000110",
  36557=>"100110100",
  36558=>"001001010",
  36559=>"110001111",
  36560=>"100000000",
  36561=>"101101001",
  36562=>"110001010",
  36563=>"000111111",
  36564=>"110000101",
  36565=>"000001011",
  36566=>"011110011",
  36567=>"100100101",
  36568=>"011110010",
  36569=>"101111111",
  36570=>"111101010",
  36571=>"000010011",
  36572=>"000101101",
  36573=>"010001101",
  36574=>"101110111",
  36575=>"000100001",
  36576=>"001010100",
  36577=>"010000100",
  36578=>"100100001",
  36579=>"100000000",
  36580=>"010011101",
  36581=>"101011011",
  36582=>"011000110",
  36583=>"101000000",
  36584=>"010101011",
  36585=>"110110101",
  36586=>"111001010",
  36587=>"111100000",
  36588=>"010001101",
  36589=>"011110011",
  36590=>"010000101",
  36591=>"100101100",
  36592=>"001101000",
  36593=>"000010101",
  36594=>"111011001",
  36595=>"011111111",
  36596=>"010101100",
  36597=>"111011110",
  36598=>"101000100",
  36599=>"111001001",
  36600=>"010011000",
  36601=>"100100011",
  36602=>"111111110",
  36603=>"110110100",
  36604=>"101101011",
  36605=>"111001011",
  36606=>"010011101",
  36607=>"010001000",
  36608=>"001010110",
  36609=>"001001111",
  36610=>"110011011",
  36611=>"001010001",
  36612=>"010001010",
  36613=>"100011100",
  36614=>"110110001",
  36615=>"110001110",
  36616=>"101011010",
  36617=>"100001110",
  36618=>"100111100",
  36619=>"101111111",
  36620=>"010011001",
  36621=>"001101101",
  36622=>"101111010",
  36623=>"100111110",
  36624=>"110101011",
  36625=>"000000111",
  36626=>"001000111",
  36627=>"010110000",
  36628=>"111100101",
  36629=>"100111110",
  36630=>"111110100",
  36631=>"000000000",
  36632=>"111011110",
  36633=>"011010001",
  36634=>"101101110",
  36635=>"100010100",
  36636=>"000010100",
  36637=>"100000110",
  36638=>"111110110",
  36639=>"110101101",
  36640=>"110101001",
  36641=>"111110101",
  36642=>"111110011",
  36643=>"011101000",
  36644=>"100000101",
  36645=>"111111011",
  36646=>"110100101",
  36647=>"101111110",
  36648=>"100001011",
  36649=>"100000100",
  36650=>"110001110",
  36651=>"100101111",
  36652=>"111010101",
  36653=>"000000001",
  36654=>"000111110",
  36655=>"011011001",
  36656=>"001100000",
  36657=>"100000100",
  36658=>"100101110",
  36659=>"101100111",
  36660=>"001111000",
  36661=>"011001001",
  36662=>"000100111",
  36663=>"000110000",
  36664=>"100011111",
  36665=>"101000101",
  36666=>"000100011",
  36667=>"100100000",
  36668=>"000101010",
  36669=>"101111101",
  36670=>"001010010",
  36671=>"111001110",
  36672=>"110000001",
  36673=>"001010010",
  36674=>"111111011",
  36675=>"110010011",
  36676=>"100111011",
  36677=>"010000011",
  36678=>"000000100",
  36679=>"110101010",
  36680=>"001111000",
  36681=>"010100000",
  36682=>"011010001",
  36683=>"010011000",
  36684=>"100010000",
  36685=>"100010100",
  36686=>"011101000",
  36687=>"101001000",
  36688=>"111111000",
  36689=>"001011001",
  36690=>"000100000",
  36691=>"011100111",
  36692=>"110100101",
  36693=>"001011010",
  36694=>"110110101",
  36695=>"010100110",
  36696=>"101010101",
  36697=>"111011111",
  36698=>"111011101",
  36699=>"101000100",
  36700=>"100101100",
  36701=>"010111100",
  36702=>"111011010",
  36703=>"010011010",
  36704=>"101011011",
  36705=>"100010000",
  36706=>"000000010",
  36707=>"101110111",
  36708=>"000100000",
  36709=>"111000001",
  36710=>"000000000",
  36711=>"010000111",
  36712=>"001010111",
  36713=>"000000111",
  36714=>"000011101",
  36715=>"111011101",
  36716=>"000111010",
  36717=>"100000011",
  36718=>"001000100",
  36719=>"001000100",
  36720=>"000001100",
  36721=>"110110110",
  36722=>"010101100",
  36723=>"010001011",
  36724=>"100001001",
  36725=>"001100111",
  36726=>"001001001",
  36727=>"001000001",
  36728=>"101111010",
  36729=>"101101001",
  36730=>"011010111",
  36731=>"010011100",
  36732=>"010000111",
  36733=>"001000001",
  36734=>"100010010",
  36735=>"111011101",
  36736=>"101010111",
  36737=>"100111000",
  36738=>"000001011",
  36739=>"100110111",
  36740=>"001101010",
  36741=>"100011010",
  36742=>"011111001",
  36743=>"000001100",
  36744=>"101111111",
  36745=>"000011110",
  36746=>"101001100",
  36747=>"000010000",
  36748=>"000100001",
  36749=>"101100111",
  36750=>"100110000",
  36751=>"110110010",
  36752=>"010111000",
  36753=>"101111110",
  36754=>"110001000",
  36755=>"100110101",
  36756=>"000011110",
  36757=>"101101111",
  36758=>"110000101",
  36759=>"010000110",
  36760=>"111101111",
  36761=>"000000111",
  36762=>"100101000",
  36763=>"111101111",
  36764=>"100001110",
  36765=>"101111110",
  36766=>"111100110",
  36767=>"010000011",
  36768=>"101101001",
  36769=>"011001101",
  36770=>"011100101",
  36771=>"010001110",
  36772=>"100101010",
  36773=>"111010110",
  36774=>"001011111",
  36775=>"011100110",
  36776=>"010101001",
  36777=>"001101011",
  36778=>"110111100",
  36779=>"111001001",
  36780=>"000001111",
  36781=>"001110001",
  36782=>"100010010",
  36783=>"111100001",
  36784=>"111111111",
  36785=>"110110111",
  36786=>"110100101",
  36787=>"100111010",
  36788=>"111001011",
  36789=>"010011100",
  36790=>"010110100",
  36791=>"101001101",
  36792=>"010110110",
  36793=>"101100101",
  36794=>"000101101",
  36795=>"001100011",
  36796=>"000001010",
  36797=>"110110100",
  36798=>"011101001",
  36799=>"001000110",
  36800=>"111000011",
  36801=>"110111000",
  36802=>"010101000",
  36803=>"111001010",
  36804=>"010001110",
  36805=>"001000100",
  36806=>"011101110",
  36807=>"011001111",
  36808=>"000011011",
  36809=>"000010111",
  36810=>"111100111",
  36811=>"000101010",
  36812=>"011100000",
  36813=>"101100001",
  36814=>"111010111",
  36815=>"001010001",
  36816=>"110101000",
  36817=>"000101111",
  36818=>"111010111",
  36819=>"000011110",
  36820=>"000001001",
  36821=>"000000101",
  36822=>"101101111",
  36823=>"101010001",
  36824=>"001100011",
  36825=>"010000000",
  36826=>"101010011",
  36827=>"101000001",
  36828=>"111100011",
  36829=>"101101010",
  36830=>"110101010",
  36831=>"100100111",
  36832=>"101001001",
  36833=>"101010101",
  36834=>"100111001",
  36835=>"001001110",
  36836=>"011011001",
  36837=>"000110000",
  36838=>"101111011",
  36839=>"111010011",
  36840=>"010100101",
  36841=>"100100110",
  36842=>"100110001",
  36843=>"000010111",
  36844=>"000011110",
  36845=>"111001011",
  36846=>"110001100",
  36847=>"111100001",
  36848=>"011010011",
  36849=>"100110110",
  36850=>"111101110",
  36851=>"100000010",
  36852=>"010111011",
  36853=>"000001110",
  36854=>"101100011",
  36855=>"010100001",
  36856=>"100101111",
  36857=>"101110000",
  36858=>"101011101",
  36859=>"101111110",
  36860=>"111001011",
  36861=>"000011000",
  36862=>"101110111",
  36863=>"101100000",
  36864=>"000111011",
  36865=>"111111011",
  36866=>"100110010",
  36867=>"100001101",
  36868=>"001100111",
  36869=>"000011100",
  36870=>"001101101",
  36871=>"000101100",
  36872=>"010000011",
  36873=>"101100010",
  36874=>"011111011",
  36875=>"100011010",
  36876=>"001000001",
  36877=>"111110111",
  36878=>"011011011",
  36879=>"011011101",
  36880=>"011100101",
  36881=>"110111011",
  36882=>"100011010",
  36883=>"010010110",
  36884=>"111101110",
  36885=>"110010011",
  36886=>"000010010",
  36887=>"011101101",
  36888=>"010011110",
  36889=>"001001011",
  36890=>"011111111",
  36891=>"000101000",
  36892=>"111011110",
  36893=>"111011000",
  36894=>"100010000",
  36895=>"000110101",
  36896=>"110011111",
  36897=>"000111100",
  36898=>"111010000",
  36899=>"000100000",
  36900=>"000101100",
  36901=>"011010101",
  36902=>"000011101",
  36903=>"100010101",
  36904=>"111101001",
  36905=>"111110101",
  36906=>"110000000",
  36907=>"100100000",
  36908=>"011111101",
  36909=>"101110101",
  36910=>"111000111",
  36911=>"101000000",
  36912=>"110000110",
  36913=>"000101000",
  36914=>"110010001",
  36915=>"100110111",
  36916=>"111001110",
  36917=>"000111100",
  36918=>"000111100",
  36919=>"000010110",
  36920=>"100111000",
  36921=>"111111110",
  36922=>"001100011",
  36923=>"101110011",
  36924=>"001011110",
  36925=>"011001101",
  36926=>"100110010",
  36927=>"111100111",
  36928=>"011000111",
  36929=>"010000010",
  36930=>"111101110",
  36931=>"110111100",
  36932=>"001011011",
  36933=>"101010110",
  36934=>"010111100",
  36935=>"101011001",
  36936=>"010011111",
  36937=>"110011101",
  36938=>"011101111",
  36939=>"111100001",
  36940=>"111011111",
  36941=>"011001010",
  36942=>"100001001",
  36943=>"101010101",
  36944=>"100110011",
  36945=>"011111111",
  36946=>"101001011",
  36947=>"101100001",
  36948=>"110000010",
  36949=>"100000111",
  36950=>"101110010",
  36951=>"111111111",
  36952=>"001100101",
  36953=>"111101011",
  36954=>"011100000",
  36955=>"000111011",
  36956=>"101101110",
  36957=>"101011111",
  36958=>"111110111",
  36959=>"101100111",
  36960=>"111111111",
  36961=>"010001000",
  36962=>"111110010",
  36963=>"011100111",
  36964=>"101010101",
  36965=>"111010100",
  36966=>"100001111",
  36967=>"111110010",
  36968=>"000001001",
  36969=>"000100000",
  36970=>"111111010",
  36971=>"110110111",
  36972=>"111001001",
  36973=>"101111100",
  36974=>"010110101",
  36975=>"111010010",
  36976=>"100110010",
  36977=>"000110101",
  36978=>"011111011",
  36979=>"010010100",
  36980=>"111100111",
  36981=>"011010111",
  36982=>"111010000",
  36983=>"101001111",
  36984=>"001111011",
  36985=>"110000001",
  36986=>"111010011",
  36987=>"101001000",
  36988=>"011100101",
  36989=>"100101100",
  36990=>"101000111",
  36991=>"000010001",
  36992=>"101100110",
  36993=>"101101100",
  36994=>"110001101",
  36995=>"011010100",
  36996=>"101010110",
  36997=>"100110000",
  36998=>"000101100",
  36999=>"101001001",
  37000=>"001010110",
  37001=>"000111110",
  37002=>"101100111",
  37003=>"111111111",
  37004=>"001010101",
  37005=>"010101000",
  37006=>"101001001",
  37007=>"001100100",
  37008=>"101111101",
  37009=>"011110001",
  37010=>"010100100",
  37011=>"111011001",
  37012=>"111011011",
  37013=>"011100111",
  37014=>"001111111",
  37015=>"100000111",
  37016=>"010110110",
  37017=>"111010110",
  37018=>"100111010",
  37019=>"011110000",
  37020=>"010001001",
  37021=>"000100010",
  37022=>"000001001",
  37023=>"000000011",
  37024=>"010001101",
  37025=>"011011001",
  37026=>"000000101",
  37027=>"011000101",
  37028=>"111010100",
  37029=>"110000010",
  37030=>"111010001",
  37031=>"011111010",
  37032=>"111101101",
  37033=>"010111101",
  37034=>"001011100",
  37035=>"010111100",
  37036=>"001110011",
  37037=>"001000111",
  37038=>"110101100",
  37039=>"111101000",
  37040=>"111011010",
  37041=>"111001011",
  37042=>"111111000",
  37043=>"110111111",
  37044=>"001011011",
  37045=>"111111001",
  37046=>"111111110",
  37047=>"101010100",
  37048=>"011111100",
  37049=>"100101111",
  37050=>"111110101",
  37051=>"111111000",
  37052=>"011001101",
  37053=>"011101111",
  37054=>"101010011",
  37055=>"000001101",
  37056=>"110001100",
  37057=>"011001001",
  37058=>"101101110",
  37059=>"111101111",
  37060=>"000010000",
  37061=>"001001111",
  37062=>"110101111",
  37063=>"101011000",
  37064=>"000111111",
  37065=>"011110101",
  37066=>"000110000",
  37067=>"110011110",
  37068=>"000011101",
  37069=>"000111000",
  37070=>"111100010",
  37071=>"110000011",
  37072=>"110000100",
  37073=>"001001001",
  37074=>"101010001",
  37075=>"011000001",
  37076=>"101110101",
  37077=>"001011101",
  37078=>"011011111",
  37079=>"110010000",
  37080=>"110000000",
  37081=>"100101100",
  37082=>"110010101",
  37083=>"011011011",
  37084=>"101011010",
  37085=>"000110001",
  37086=>"100101100",
  37087=>"110000010",
  37088=>"010010110",
  37089=>"011001101",
  37090=>"101011000",
  37091=>"101011001",
  37092=>"111010101",
  37093=>"001101111",
  37094=>"011011111",
  37095=>"101111001",
  37096=>"100110010",
  37097=>"101101000",
  37098=>"100111111",
  37099=>"111011110",
  37100=>"001101010",
  37101=>"010010100",
  37102=>"111101110",
  37103=>"010110000",
  37104=>"111110000",
  37105=>"011011001",
  37106=>"111100111",
  37107=>"111001010",
  37108=>"110111001",
  37109=>"011010110",
  37110=>"100111100",
  37111=>"001011011",
  37112=>"011001101",
  37113=>"110000000",
  37114=>"111011001",
  37115=>"001111101",
  37116=>"010000001",
  37117=>"110101011",
  37118=>"011110011",
  37119=>"001101000",
  37120=>"011000001",
  37121=>"010100110",
  37122=>"110100100",
  37123=>"111111100",
  37124=>"001111011",
  37125=>"101001011",
  37126=>"110111111",
  37127=>"000101101",
  37128=>"110000001",
  37129=>"100111111",
  37130=>"000011100",
  37131=>"111100110",
  37132=>"011011111",
  37133=>"000100011",
  37134=>"101001111",
  37135=>"111001101",
  37136=>"011011011",
  37137=>"011011110",
  37138=>"000011110",
  37139=>"100010100",
  37140=>"101111010",
  37141=>"010111111",
  37142=>"000101001",
  37143=>"100101101",
  37144=>"111100101",
  37145=>"010101101",
  37146=>"111111001",
  37147=>"101000111",
  37148=>"111111110",
  37149=>"010000111",
  37150=>"110010101",
  37151=>"001011111",
  37152=>"101111110",
  37153=>"111101001",
  37154=>"101100001",
  37155=>"000010011",
  37156=>"001000000",
  37157=>"100010111",
  37158=>"001000011",
  37159=>"111111110",
  37160=>"111011000",
  37161=>"100000010",
  37162=>"110100010",
  37163=>"111111111",
  37164=>"001101010",
  37165=>"100111100",
  37166=>"100110111",
  37167=>"001100010",
  37168=>"001111110",
  37169=>"100010001",
  37170=>"011011100",
  37171=>"110110110",
  37172=>"000100001",
  37173=>"111011010",
  37174=>"011001101",
  37175=>"100100100",
  37176=>"101110111",
  37177=>"101001010",
  37178=>"111011111",
  37179=>"011010101",
  37180=>"111011111",
  37181=>"100000111",
  37182=>"010001001",
  37183=>"000110001",
  37184=>"101101100",
  37185=>"101110010",
  37186=>"011101011",
  37187=>"000001011",
  37188=>"011011101",
  37189=>"110011011",
  37190=>"110100001",
  37191=>"011001111",
  37192=>"000000101",
  37193=>"001101111",
  37194=>"000000011",
  37195=>"111100000",
  37196=>"010000110",
  37197=>"111101100",
  37198=>"001010100",
  37199=>"110101011",
  37200=>"100010110",
  37201=>"110101101",
  37202=>"011001001",
  37203=>"101000101",
  37204=>"001011111",
  37205=>"100010000",
  37206=>"101110000",
  37207=>"001101011",
  37208=>"111100011",
  37209=>"011101011",
  37210=>"001000010",
  37211=>"011100111",
  37212=>"000001100",
  37213=>"100000011",
  37214=>"000101010",
  37215=>"100110111",
  37216=>"110100001",
  37217=>"011011111",
  37218=>"011011101",
  37219=>"110101101",
  37220=>"000111111",
  37221=>"001000111",
  37222=>"110111001",
  37223=>"011010010",
  37224=>"011011001",
  37225=>"000100101",
  37226=>"110100000",
  37227=>"110101100",
  37228=>"001110010",
  37229=>"000101111",
  37230=>"110101101",
  37231=>"010011110",
  37232=>"010011111",
  37233=>"001110110",
  37234=>"111000000",
  37235=>"100000010",
  37236=>"101100001",
  37237=>"011100101",
  37238=>"011110111",
  37239=>"100010011",
  37240=>"111000101",
  37241=>"011111110",
  37242=>"100010010",
  37243=>"011000000",
  37244=>"111110010",
  37245=>"101111000",
  37246=>"011111001",
  37247=>"011111101",
  37248=>"100001101",
  37249=>"111111100",
  37250=>"011000000",
  37251=>"011011110",
  37252=>"000101111",
  37253=>"110111010",
  37254=>"110101000",
  37255=>"010111011",
  37256=>"001111101",
  37257=>"110000010",
  37258=>"010111001",
  37259=>"111101001",
  37260=>"001001001",
  37261=>"011110111",
  37262=>"100110001",
  37263=>"000000000",
  37264=>"111000101",
  37265=>"011111100",
  37266=>"111110110",
  37267=>"100110010",
  37268=>"111010000",
  37269=>"101010001",
  37270=>"001001111",
  37271=>"011000001",
  37272=>"100101001",
  37273=>"111110111",
  37274=>"110001010",
  37275=>"011010100",
  37276=>"110001101",
  37277=>"011101001",
  37278=>"111010101",
  37279=>"101110010",
  37280=>"100100100",
  37281=>"010011111",
  37282=>"000001110",
  37283=>"110111100",
  37284=>"111000001",
  37285=>"100000001",
  37286=>"010010011",
  37287=>"111010100",
  37288=>"011000110",
  37289=>"101001000",
  37290=>"011100111",
  37291=>"001100111",
  37292=>"101011101",
  37293=>"010110111",
  37294=>"101010111",
  37295=>"101101001",
  37296=>"001011001",
  37297=>"010011011",
  37298=>"001100000",
  37299=>"111111000",
  37300=>"110111111",
  37301=>"111100000",
  37302=>"110111011",
  37303=>"010010101",
  37304=>"100100110",
  37305=>"000001100",
  37306=>"111100111",
  37307=>"110011100",
  37308=>"000000100",
  37309=>"111011011",
  37310=>"000000111",
  37311=>"010011011",
  37312=>"000011010",
  37313=>"001000010",
  37314=>"011000110",
  37315=>"110001110",
  37316=>"000011111",
  37317=>"010000010",
  37318=>"111101111",
  37319=>"100001011",
  37320=>"100101110",
  37321=>"010101110",
  37322=>"000000100",
  37323=>"111100011",
  37324=>"011110101",
  37325=>"000001010",
  37326=>"111010101",
  37327=>"000100000",
  37328=>"110000000",
  37329=>"011011011",
  37330=>"111101010",
  37331=>"001110010",
  37332=>"001100100",
  37333=>"110001001",
  37334=>"001111011",
  37335=>"011001111",
  37336=>"010110100",
  37337=>"000001010",
  37338=>"111001000",
  37339=>"101000101",
  37340=>"111100110",
  37341=>"000101100",
  37342=>"100101000",
  37343=>"100110111",
  37344=>"100001000",
  37345=>"001110111",
  37346=>"001000011",
  37347=>"110110110",
  37348=>"101011101",
  37349=>"011111111",
  37350=>"000000111",
  37351=>"011000111",
  37352=>"111111100",
  37353=>"010111001",
  37354=>"110010101",
  37355=>"010111100",
  37356=>"111010010",
  37357=>"110001101",
  37358=>"000101100",
  37359=>"101111011",
  37360=>"000010000",
  37361=>"011001010",
  37362=>"111111110",
  37363=>"010010100",
  37364=>"110010100",
  37365=>"111011100",
  37366=>"011110110",
  37367=>"101110000",
  37368=>"011110111",
  37369=>"010100010",
  37370=>"100000100",
  37371=>"010110111",
  37372=>"001111000",
  37373=>"110101111",
  37374=>"000110101",
  37375=>"000101111",
  37376=>"101100010",
  37377=>"000011000",
  37378=>"000011011",
  37379=>"101011011",
  37380=>"101001000",
  37381=>"001011111",
  37382=>"010110010",
  37383=>"111111010",
  37384=>"100001111",
  37385=>"110000010",
  37386=>"101101110",
  37387=>"110111110",
  37388=>"010101010",
  37389=>"101101010",
  37390=>"000000011",
  37391=>"101011000",
  37392=>"101111001",
  37393=>"110101111",
  37394=>"100111010",
  37395=>"110101100",
  37396=>"011110101",
  37397=>"001011001",
  37398=>"001001110",
  37399=>"011110010",
  37400=>"001001111",
  37401=>"001111111",
  37402=>"101111111",
  37403=>"110100001",
  37404=>"000111011",
  37405=>"011011101",
  37406=>"001000001",
  37407=>"010010110",
  37408=>"011101001",
  37409=>"000011010",
  37410=>"101110110",
  37411=>"011111010",
  37412=>"001001011",
  37413=>"000100010",
  37414=>"010001011",
  37415=>"001011010",
  37416=>"101100000",
  37417=>"101111101",
  37418=>"100011100",
  37419=>"101101110",
  37420=>"110110101",
  37421=>"011010110",
  37422=>"010000000",
  37423=>"101111011",
  37424=>"001011011",
  37425=>"011010101",
  37426=>"000100101",
  37427=>"101101110",
  37428=>"110101111",
  37429=>"001100000",
  37430=>"010010101",
  37431=>"110000111",
  37432=>"010100101",
  37433=>"101011010",
  37434=>"110100001",
  37435=>"100110110",
  37436=>"111110110",
  37437=>"001010110",
  37438=>"110101001",
  37439=>"000100000",
  37440=>"010000100",
  37441=>"011000011",
  37442=>"010001110",
  37443=>"110011111",
  37444=>"110101110",
  37445=>"101111100",
  37446=>"001010001",
  37447=>"011000101",
  37448=>"010111011",
  37449=>"011111000",
  37450=>"010011000",
  37451=>"011001011",
  37452=>"100101010",
  37453=>"101011110",
  37454=>"000010010",
  37455=>"100011111",
  37456=>"111000001",
  37457=>"110010100",
  37458=>"000101000",
  37459=>"110111111",
  37460=>"001111000",
  37461=>"100101000",
  37462=>"001000100",
  37463=>"100000100",
  37464=>"100110011",
  37465=>"111001101",
  37466=>"100100100",
  37467=>"100111100",
  37468=>"001001111",
  37469=>"000100001",
  37470=>"111101111",
  37471=>"011000001",
  37472=>"000110010",
  37473=>"010011110",
  37474=>"100001010",
  37475=>"000001000",
  37476=>"110111111",
  37477=>"111111100",
  37478=>"111100001",
  37479=>"010100111",
  37480=>"111101111",
  37481=>"001011011",
  37482=>"101000010",
  37483=>"100011111",
  37484=>"110011100",
  37485=>"000010010",
  37486=>"100001000",
  37487=>"101000100",
  37488=>"010101010",
  37489=>"110010011",
  37490=>"111010100",
  37491=>"010100000",
  37492=>"001111101",
  37493=>"000100110",
  37494=>"000010000",
  37495=>"000011001",
  37496=>"000110110",
  37497=>"000011110",
  37498=>"010101100",
  37499=>"010001111",
  37500=>"110111110",
  37501=>"000011101",
  37502=>"000000100",
  37503=>"000001010",
  37504=>"000111111",
  37505=>"110110001",
  37506=>"001111001",
  37507=>"101010011",
  37508=>"111111111",
  37509=>"111000110",
  37510=>"110111110",
  37511=>"000011111",
  37512=>"111011010",
  37513=>"011101101",
  37514=>"010100100",
  37515=>"101110011",
  37516=>"100000111",
  37517=>"101101001",
  37518=>"000010001",
  37519=>"001001000",
  37520=>"011110111",
  37521=>"011001011",
  37522=>"100011011",
  37523=>"010011011",
  37524=>"110101101",
  37525=>"110110101",
  37526=>"011010010",
  37527=>"010110100",
  37528=>"101111011",
  37529=>"001111000",
  37530=>"011111110",
  37531=>"101100010",
  37532=>"011101111",
  37533=>"110011001",
  37534=>"110000011",
  37535=>"001011001",
  37536=>"111011011",
  37537=>"001110001",
  37538=>"111111100",
  37539=>"100000111",
  37540=>"001001111",
  37541=>"001101001",
  37542=>"010100010",
  37543=>"011011001",
  37544=>"101111111",
  37545=>"100111000",
  37546=>"101100010",
  37547=>"011000101",
  37548=>"111100100",
  37549=>"111001100",
  37550=>"011111110",
  37551=>"111110000",
  37552=>"111011101",
  37553=>"001110110",
  37554=>"000111111",
  37555=>"011011001",
  37556=>"111100011",
  37557=>"111111101",
  37558=>"101101011",
  37559=>"101000100",
  37560=>"000011111",
  37561=>"010100101",
  37562=>"101000000",
  37563=>"100011110",
  37564=>"101100000",
  37565=>"001011101",
  37566=>"100001110",
  37567=>"001100111",
  37568=>"010010101",
  37569=>"110100110",
  37570=>"010011001",
  37571=>"101101111",
  37572=>"111110101",
  37573=>"001000100",
  37574=>"100100110",
  37575=>"000111111",
  37576=>"000000011",
  37577=>"111111001",
  37578=>"110101101",
  37579=>"110110100",
  37580=>"101111110",
  37581=>"110010000",
  37582=>"110101110",
  37583=>"111001101",
  37584=>"010110111",
  37585=>"100100001",
  37586=>"011110101",
  37587=>"001011101",
  37588=>"110110111",
  37589=>"111111001",
  37590=>"100010000",
  37591=>"111011001",
  37592=>"101011000",
  37593=>"111101111",
  37594=>"000010111",
  37595=>"001101101",
  37596=>"111111000",
  37597=>"100000100",
  37598=>"100110011",
  37599=>"001110100",
  37600=>"010110101",
  37601=>"000001110",
  37602=>"001100101",
  37603=>"110101010",
  37604=>"111111101",
  37605=>"000000100",
  37606=>"011101001",
  37607=>"001010101",
  37608=>"010011001",
  37609=>"101001001",
  37610=>"111000010",
  37611=>"000010010",
  37612=>"000110110",
  37613=>"011011010",
  37614=>"111100100",
  37615=>"011011000",
  37616=>"000100011",
  37617=>"011001001",
  37618=>"101100101",
  37619=>"000010110",
  37620=>"110110000",
  37621=>"110110110",
  37622=>"110101001",
  37623=>"011010101",
  37624=>"010010100",
  37625=>"111001111",
  37626=>"111101000",
  37627=>"110111100",
  37628=>"100101101",
  37629=>"001101110",
  37630=>"111110010",
  37631=>"111011111",
  37632=>"110111111",
  37633=>"111100111",
  37634=>"110110111",
  37635=>"111010010",
  37636=>"110101011",
  37637=>"001010010",
  37638=>"101111000",
  37639=>"100001001",
  37640=>"111101101",
  37641=>"101110110",
  37642=>"000100000",
  37643=>"000101111",
  37644=>"000100100",
  37645=>"111111111",
  37646=>"010010010",
  37647=>"001011001",
  37648=>"111111101",
  37649=>"011001011",
  37650=>"101000101",
  37651=>"110110000",
  37652=>"001110101",
  37653=>"100000011",
  37654=>"000010001",
  37655=>"010111100",
  37656=>"101101101",
  37657=>"000111011",
  37658=>"111111010",
  37659=>"100001101",
  37660=>"100111010",
  37661=>"110010111",
  37662=>"010010111",
  37663=>"101101110",
  37664=>"101000000",
  37665=>"101001110",
  37666=>"110000110",
  37667=>"100001011",
  37668=>"011100001",
  37669=>"101000011",
  37670=>"110101110",
  37671=>"001101011",
  37672=>"101000111",
  37673=>"110110001",
  37674=>"100011000",
  37675=>"001000111",
  37676=>"111000011",
  37677=>"111111101",
  37678=>"101101111",
  37679=>"000001111",
  37680=>"111111111",
  37681=>"001001110",
  37682=>"010100000",
  37683=>"100100000",
  37684=>"001010000",
  37685=>"000111110",
  37686=>"110001100",
  37687=>"100110100",
  37688=>"111110001",
  37689=>"001011001",
  37690=>"010110000",
  37691=>"011000110",
  37692=>"000111110",
  37693=>"101011100",
  37694=>"100110011",
  37695=>"110011011",
  37696=>"000000010",
  37697=>"110001110",
  37698=>"001000001",
  37699=>"000110100",
  37700=>"001001101",
  37701=>"010011110",
  37702=>"100011101",
  37703=>"001011011",
  37704=>"110110101",
  37705=>"011100111",
  37706=>"111010001",
  37707=>"010111101",
  37708=>"110100110",
  37709=>"110001010",
  37710=>"111001010",
  37711=>"111000010",
  37712=>"100011000",
  37713=>"111111111",
  37714=>"011111011",
  37715=>"000101101",
  37716=>"100100111",
  37717=>"110010101",
  37718=>"111110111",
  37719=>"000000011",
  37720=>"110001111",
  37721=>"011100101",
  37722=>"110001111",
  37723=>"001111111",
  37724=>"111111011",
  37725=>"101101100",
  37726=>"001011101",
  37727=>"011011101",
  37728=>"100010100",
  37729=>"011001111",
  37730=>"111111011",
  37731=>"101011100",
  37732=>"010100110",
  37733=>"011100101",
  37734=>"101101001",
  37735=>"100100000",
  37736=>"001101101",
  37737=>"110000100",
  37738=>"111100111",
  37739=>"011001001",
  37740=>"111101111",
  37741=>"010001001",
  37742=>"000100000",
  37743=>"001101111",
  37744=>"111111101",
  37745=>"100111111",
  37746=>"001000010",
  37747=>"001111111",
  37748=>"101011001",
  37749=>"100000001",
  37750=>"100101001",
  37751=>"110001001",
  37752=>"111001010",
  37753=>"101011110",
  37754=>"011111101",
  37755=>"000101111",
  37756=>"011011011",
  37757=>"111101101",
  37758=>"111000110",
  37759=>"000000000",
  37760=>"111011110",
  37761=>"111111110",
  37762=>"000100000",
  37763=>"010111011",
  37764=>"011111010",
  37765=>"111111111",
  37766=>"110011001",
  37767=>"011001110",
  37768=>"011000001",
  37769=>"111111110",
  37770=>"100100110",
  37771=>"011001110",
  37772=>"010010111",
  37773=>"001001100",
  37774=>"100000000",
  37775=>"100010011",
  37776=>"000000000",
  37777=>"110011010",
  37778=>"000010111",
  37779=>"000111000",
  37780=>"100000001",
  37781=>"010010111",
  37782=>"001011001",
  37783=>"000111110",
  37784=>"001100110",
  37785=>"001000011",
  37786=>"100001110",
  37787=>"101001101",
  37788=>"010001000",
  37789=>"111011110",
  37790=>"111110111",
  37791=>"001010101",
  37792=>"001111101",
  37793=>"011000010",
  37794=>"111011101",
  37795=>"011101111",
  37796=>"001001111",
  37797=>"110101001",
  37798=>"001010010",
  37799=>"100000100",
  37800=>"001101011",
  37801=>"101100000",
  37802=>"101010000",
  37803=>"101111101",
  37804=>"101011001",
  37805=>"001001011",
  37806=>"000101000",
  37807=>"000000000",
  37808=>"111010111",
  37809=>"110000101",
  37810=>"110100001",
  37811=>"110000100",
  37812=>"110010001",
  37813=>"100111110",
  37814=>"000010000",
  37815=>"000100111",
  37816=>"000011000",
  37817=>"000000100",
  37818=>"100100011",
  37819=>"011011111",
  37820=>"100100110",
  37821=>"100001101",
  37822=>"001010011",
  37823=>"101011001",
  37824=>"100100010",
  37825=>"010111100",
  37826=>"110110111",
  37827=>"000101100",
  37828=>"000000001",
  37829=>"000100001",
  37830=>"011000011",
  37831=>"011111100",
  37832=>"111111110",
  37833=>"011111001",
  37834=>"101000010",
  37835=>"100100100",
  37836=>"010111000",
  37837=>"011001110",
  37838=>"110001100",
  37839=>"100101011",
  37840=>"001100110",
  37841=>"101000001",
  37842=>"111001000",
  37843=>"011110111",
  37844=>"101000001",
  37845=>"111100111",
  37846=>"011010000",
  37847=>"011100111",
  37848=>"111111100",
  37849=>"011100110",
  37850=>"011000111",
  37851=>"101000111",
  37852=>"100011110",
  37853=>"001000110",
  37854=>"010111111",
  37855=>"111111110",
  37856=>"111110100",
  37857=>"101001110",
  37858=>"000001010",
  37859=>"011001111",
  37860=>"001011011",
  37861=>"001000111",
  37862=>"000000000",
  37863=>"000101011",
  37864=>"100100110",
  37865=>"101111001",
  37866=>"000010101",
  37867=>"001101101",
  37868=>"010011000",
  37869=>"100110101",
  37870=>"100011100",
  37871=>"000100110",
  37872=>"111000100",
  37873=>"011001000",
  37874=>"010100110",
  37875=>"110101100",
  37876=>"110000110",
  37877=>"111100111",
  37878=>"000001001",
  37879=>"010110111",
  37880=>"110001010",
  37881=>"100100010",
  37882=>"100110001",
  37883=>"111110010",
  37884=>"001001011",
  37885=>"100011110",
  37886=>"011101101",
  37887=>"101011010",
  37888=>"100010111",
  37889=>"111111100",
  37890=>"100011101",
  37891=>"101110101",
  37892=>"110101010",
  37893=>"010010110",
  37894=>"010001111",
  37895=>"111100100",
  37896=>"110000011",
  37897=>"001101001",
  37898=>"101100001",
  37899=>"001111011",
  37900=>"000010001",
  37901=>"110100000",
  37902=>"111101011",
  37903=>"111101111",
  37904=>"010001000",
  37905=>"111111101",
  37906=>"110000110",
  37907=>"110100100",
  37908=>"111010101",
  37909=>"111100011",
  37910=>"101001101",
  37911=>"000010000",
  37912=>"111101001",
  37913=>"100001010",
  37914=>"110011110",
  37915=>"101001111",
  37916=>"100001001",
  37917=>"010101010",
  37918=>"001000111",
  37919=>"000001001",
  37920=>"110111010",
  37921=>"011000011",
  37922=>"100110000",
  37923=>"100000010",
  37924=>"100101100",
  37925=>"011000100",
  37926=>"100101011",
  37927=>"001111111",
  37928=>"000100110",
  37929=>"000010000",
  37930=>"010110000",
  37931=>"011001110",
  37932=>"111110001",
  37933=>"010001001",
  37934=>"011100000",
  37935=>"100010011",
  37936=>"010000000",
  37937=>"010010110",
  37938=>"010111010",
  37939=>"010010000",
  37940=>"101000100",
  37941=>"001101000",
  37942=>"101000000",
  37943=>"111010010",
  37944=>"100111101",
  37945=>"001001000",
  37946=>"110010011",
  37947=>"100110011",
  37948=>"001010100",
  37949=>"101111010",
  37950=>"011101000",
  37951=>"010111100",
  37952=>"010110001",
  37953=>"001000001",
  37954=>"010111111",
  37955=>"001011100",
  37956=>"111110111",
  37957=>"101100000",
  37958=>"101111010",
  37959=>"101001101",
  37960=>"111101001",
  37961=>"100000011",
  37962=>"111100110",
  37963=>"111000101",
  37964=>"110011110",
  37965=>"111001100",
  37966=>"110001010",
  37967=>"111001010",
  37968=>"001011000",
  37969=>"100100011",
  37970=>"111001101",
  37971=>"011101100",
  37972=>"011111000",
  37973=>"001000000",
  37974=>"011001001",
  37975=>"100000000",
  37976=>"001011111",
  37977=>"010110010",
  37978=>"101011101",
  37979=>"111011010",
  37980=>"010110000",
  37981=>"000110000",
  37982=>"111110101",
  37983=>"001100101",
  37984=>"000000110",
  37985=>"001110010",
  37986=>"100000100",
  37987=>"110110001",
  37988=>"100001101",
  37989=>"010000000",
  37990=>"101011111",
  37991=>"010101000",
  37992=>"111000001",
  37993=>"110010110",
  37994=>"101001101",
  37995=>"000100010",
  37996=>"101000001",
  37997=>"010000101",
  37998=>"111000010",
  37999=>"011110101",
  38000=>"011110010",
  38001=>"010000101",
  38002=>"111001010",
  38003=>"010110011",
  38004=>"011111010",
  38005=>"111100011",
  38006=>"011000110",
  38007=>"100110001",
  38008=>"100101100",
  38009=>"001011111",
  38010=>"111101010",
  38011=>"110010011",
  38012=>"011110011",
  38013=>"101010100",
  38014=>"010010110",
  38015=>"001110101",
  38016=>"101111010",
  38017=>"111111100",
  38018=>"000101000",
  38019=>"001000100",
  38020=>"010011000",
  38021=>"001011100",
  38022=>"110001000",
  38023=>"011001000",
  38024=>"011110101",
  38025=>"010100101",
  38026=>"001011000",
  38027=>"101000000",
  38028=>"101101111",
  38029=>"010100110",
  38030=>"110111000",
  38031=>"111000100",
  38032=>"010100100",
  38033=>"110100001",
  38034=>"001000101",
  38035=>"101001111",
  38036=>"111101100",
  38037=>"100011010",
  38038=>"010110101",
  38039=>"010010101",
  38040=>"110111010",
  38041=>"000000101",
  38042=>"010000001",
  38043=>"100010011",
  38044=>"011011100",
  38045=>"110100110",
  38046=>"101110110",
  38047=>"101111001",
  38048=>"111100000",
  38049=>"001111101",
  38050=>"000101110",
  38051=>"010110110",
  38052=>"111001110",
  38053=>"111110000",
  38054=>"011001100",
  38055=>"001010100",
  38056=>"110001000",
  38057=>"011111001",
  38058=>"010110001",
  38059=>"010110110",
  38060=>"101000101",
  38061=>"101111111",
  38062=>"101010111",
  38063=>"001101010",
  38064=>"111001000",
  38065=>"000110100",
  38066=>"110111010",
  38067=>"011100010",
  38068=>"001011111",
  38069=>"001001111",
  38070=>"000001000",
  38071=>"110111111",
  38072=>"101000000",
  38073=>"011000011",
  38074=>"000111011",
  38075=>"100000110",
  38076=>"001001011",
  38077=>"001111011",
  38078=>"111111110",
  38079=>"110011111",
  38080=>"010011111",
  38081=>"110010101",
  38082=>"110011000",
  38083=>"011001111",
  38084=>"000001110",
  38085=>"101001000",
  38086=>"010000011",
  38087=>"110001101",
  38088=>"000111000",
  38089=>"101011100",
  38090=>"001001111",
  38091=>"010000010",
  38092=>"100100001",
  38093=>"001010010",
  38094=>"001010101",
  38095=>"010001100",
  38096=>"011110000",
  38097=>"100111101",
  38098=>"010010000",
  38099=>"100100100",
  38100=>"011001001",
  38101=>"111111001",
  38102=>"111100001",
  38103=>"101101001",
  38104=>"101011001",
  38105=>"000110001",
  38106=>"110100010",
  38107=>"111011000",
  38108=>"000101100",
  38109=>"011000010",
  38110=>"111001110",
  38111=>"001111110",
  38112=>"110101010",
  38113=>"010000011",
  38114=>"111001111",
  38115=>"111100000",
  38116=>"001001110",
  38117=>"110011101",
  38118=>"110001011",
  38119=>"101100011",
  38120=>"001100100",
  38121=>"000110010",
  38122=>"100000011",
  38123=>"000000000",
  38124=>"101011110",
  38125=>"111111101",
  38126=>"000000010",
  38127=>"100000000",
  38128=>"111000101",
  38129=>"011010000",
  38130=>"110110111",
  38131=>"000011100",
  38132=>"110101101",
  38133=>"110011001",
  38134=>"001101111",
  38135=>"101100001",
  38136=>"110110100",
  38137=>"100001101",
  38138=>"101001100",
  38139=>"000001111",
  38140=>"010010111",
  38141=>"011000110",
  38142=>"001110001",
  38143=>"010100001",
  38144=>"011111000",
  38145=>"111000100",
  38146=>"000110000",
  38147=>"001111101",
  38148=>"011001001",
  38149=>"110011111",
  38150=>"110110111",
  38151=>"011010101",
  38152=>"100011101",
  38153=>"011010000",
  38154=>"110001110",
  38155=>"110001110",
  38156=>"011000101",
  38157=>"100001010",
  38158=>"101110011",
  38159=>"001101001",
  38160=>"110010111",
  38161=>"111010101",
  38162=>"010101110",
  38163=>"000000010",
  38164=>"110001100",
  38165=>"101111101",
  38166=>"111100010",
  38167=>"011110010",
  38168=>"011111111",
  38169=>"101011011",
  38170=>"000000011",
  38171=>"011101000",
  38172=>"011000111",
  38173=>"011001000",
  38174=>"111111100",
  38175=>"000111100",
  38176=>"111001001",
  38177=>"000001011",
  38178=>"001000100",
  38179=>"101101101",
  38180=>"111010101",
  38181=>"000111100",
  38182=>"111000100",
  38183=>"011100010",
  38184=>"001111011",
  38185=>"011111010",
  38186=>"000010101",
  38187=>"000001111",
  38188=>"100111000",
  38189=>"110011110",
  38190=>"110111100",
  38191=>"011100111",
  38192=>"111010011",
  38193=>"101011110",
  38194=>"110100111",
  38195=>"110010010",
  38196=>"100100000",
  38197=>"111100011",
  38198=>"000000011",
  38199=>"000101111",
  38200=>"000010011",
  38201=>"111000100",
  38202=>"010101111",
  38203=>"000111111",
  38204=>"010011000",
  38205=>"000000001",
  38206=>"010100011",
  38207=>"010010001",
  38208=>"100101111",
  38209=>"110110111",
  38210=>"111110000",
  38211=>"010000011",
  38212=>"001110010",
  38213=>"111011111",
  38214=>"101101100",
  38215=>"001001101",
  38216=>"110100110",
  38217=>"000110011",
  38218=>"110111010",
  38219=>"101010011",
  38220=>"110111111",
  38221=>"010101011",
  38222=>"011110001",
  38223=>"100010110",
  38224=>"011111011",
  38225=>"011111100",
  38226=>"001011001",
  38227=>"000110011",
  38228=>"110111111",
  38229=>"001010000",
  38230=>"010101001",
  38231=>"010011011",
  38232=>"100011010",
  38233=>"001001100",
  38234=>"101011010",
  38235=>"101010101",
  38236=>"111111001",
  38237=>"001100000",
  38238=>"111101101",
  38239=>"000111001",
  38240=>"101000010",
  38241=>"101111111",
  38242=>"110110010",
  38243=>"100111000",
  38244=>"100010110",
  38245=>"011010000",
  38246=>"001001010",
  38247=>"001011000",
  38248=>"111100001",
  38249=>"101010110",
  38250=>"000000100",
  38251=>"100110000",
  38252=>"100001001",
  38253=>"110111000",
  38254=>"101110000",
  38255=>"001010000",
  38256=>"000011001",
  38257=>"101011101",
  38258=>"001001110",
  38259=>"110001111",
  38260=>"111111111",
  38261=>"011010111",
  38262=>"010010010",
  38263=>"000111001",
  38264=>"010001011",
  38265=>"100000101",
  38266=>"000101111",
  38267=>"001000110",
  38268=>"101010101",
  38269=>"111011111",
  38270=>"101010010",
  38271=>"110000100",
  38272=>"110010100",
  38273=>"010000000",
  38274=>"010111111",
  38275=>"010110111",
  38276=>"110010001",
  38277=>"000011111",
  38278=>"010000111",
  38279=>"011000001",
  38280=>"011100110",
  38281=>"100011101",
  38282=>"011011100",
  38283=>"001101101",
  38284=>"000111100",
  38285=>"110010000",
  38286=>"000100001",
  38287=>"101001101",
  38288=>"010000111",
  38289=>"000110110",
  38290=>"011011000",
  38291=>"110110100",
  38292=>"100011111",
  38293=>"110000001",
  38294=>"111001000",
  38295=>"000101010",
  38296=>"100101111",
  38297=>"100001001",
  38298=>"110100101",
  38299=>"001001111",
  38300=>"011000111",
  38301=>"000011010",
  38302=>"000011000",
  38303=>"001011100",
  38304=>"111100101",
  38305=>"101100010",
  38306=>"011010010",
  38307=>"110100000",
  38308=>"111100001",
  38309=>"011000111",
  38310=>"111000101",
  38311=>"110011000",
  38312=>"111100001",
  38313=>"001001101",
  38314=>"000011000",
  38315=>"000010001",
  38316=>"111110100",
  38317=>"010000010",
  38318=>"111000110",
  38319=>"001100110",
  38320=>"100010110",
  38321=>"011001011",
  38322=>"011111011",
  38323=>"011010011",
  38324=>"100000111",
  38325=>"110001111",
  38326=>"011011101",
  38327=>"000100001",
  38328=>"000110000",
  38329=>"001101110",
  38330=>"000101000",
  38331=>"100101001",
  38332=>"111111100",
  38333=>"111100001",
  38334=>"000100111",
  38335=>"111000111",
  38336=>"110110000",
  38337=>"001011001",
  38338=>"110100000",
  38339=>"000001000",
  38340=>"000111000",
  38341=>"001001111",
  38342=>"100111111",
  38343=>"111110100",
  38344=>"101100010",
  38345=>"100101011",
  38346=>"100011001",
  38347=>"011001111",
  38348=>"000011100",
  38349=>"011001110",
  38350=>"000000110",
  38351=>"000011101",
  38352=>"111101111",
  38353=>"011101000",
  38354=>"001000111",
  38355=>"000100101",
  38356=>"010000101",
  38357=>"100000111",
  38358=>"110010011",
  38359=>"101111010",
  38360=>"010111111",
  38361=>"101000110",
  38362=>"011010001",
  38363=>"001100101",
  38364=>"010011101",
  38365=>"111001100",
  38366=>"101110011",
  38367=>"111100101",
  38368=>"011110011",
  38369=>"101001001",
  38370=>"001010100",
  38371=>"100010001",
  38372=>"110001110",
  38373=>"010000100",
  38374=>"100111010",
  38375=>"011100010",
  38376=>"111101101",
  38377=>"101111111",
  38378=>"011101101",
  38379=>"111010100",
  38380=>"100001010",
  38381=>"010000100",
  38382=>"010001101",
  38383=>"101011101",
  38384=>"001111110",
  38385=>"101011000",
  38386=>"001100011",
  38387=>"100111000",
  38388=>"001100001",
  38389=>"110011000",
  38390=>"001000011",
  38391=>"110111011",
  38392=>"010010001",
  38393=>"101010000",
  38394=>"010011011",
  38395=>"110000101",
  38396=>"100000001",
  38397=>"100111111",
  38398=>"001111010",
  38399=>"010011011",
  38400=>"001010001",
  38401=>"101001001",
  38402=>"000100100",
  38403=>"010111000",
  38404=>"101101010",
  38405=>"100010101",
  38406=>"100001001",
  38407=>"011100111",
  38408=>"010010111",
  38409=>"011010010",
  38410=>"001100101",
  38411=>"011011101",
  38412=>"101111111",
  38413=>"011001100",
  38414=>"000100000",
  38415=>"111111000",
  38416=>"111101111",
  38417=>"011011111",
  38418=>"000000001",
  38419=>"010010001",
  38420=>"100111111",
  38421=>"011001010",
  38422=>"100110111",
  38423=>"100000111",
  38424=>"011010001",
  38425=>"010001010",
  38426=>"110000000",
  38427=>"110101001",
  38428=>"000001000",
  38429=>"000001111",
  38430=>"000110100",
  38431=>"100110110",
  38432=>"101101001",
  38433=>"001011110",
  38434=>"110000011",
  38435=>"101000100",
  38436=>"001100110",
  38437=>"001000011",
  38438=>"001010101",
  38439=>"110011110",
  38440=>"000000010",
  38441=>"001000100",
  38442=>"000001001",
  38443=>"000011010",
  38444=>"110000011",
  38445=>"001000010",
  38446=>"000100000",
  38447=>"111011010",
  38448=>"011111100",
  38449=>"000100101",
  38450=>"000000001",
  38451=>"110110011",
  38452=>"110110001",
  38453=>"010000000",
  38454=>"111000001",
  38455=>"000001000",
  38456=>"101101111",
  38457=>"100111111",
  38458=>"011101011",
  38459=>"011111000",
  38460=>"110110101",
  38461=>"010111110",
  38462=>"001010000",
  38463=>"000000010",
  38464=>"110101000",
  38465=>"101010110",
  38466=>"010011101",
  38467=>"111100001",
  38468=>"100001101",
  38469=>"010000100",
  38470=>"000010010",
  38471=>"110010110",
  38472=>"010100000",
  38473=>"001011101",
  38474=>"000101110",
  38475=>"000110110",
  38476=>"011101101",
  38477=>"001010101",
  38478=>"000001001",
  38479=>"000100001",
  38480=>"110100011",
  38481=>"100011100",
  38482=>"010011111",
  38483=>"110001011",
  38484=>"100001110",
  38485=>"011111111",
  38486=>"001111000",
  38487=>"110100010",
  38488=>"100000000",
  38489=>"111011011",
  38490=>"111111101",
  38491=>"000111110",
  38492=>"100011010",
  38493=>"010111100",
  38494=>"001101010",
  38495=>"111110010",
  38496=>"111001110",
  38497=>"001111001",
  38498=>"101000101",
  38499=>"000000010",
  38500=>"100011101",
  38501=>"010010011",
  38502=>"000010110",
  38503=>"011010111",
  38504=>"001011001",
  38505=>"111110111",
  38506=>"110000001",
  38507=>"011110100",
  38508=>"000011101",
  38509=>"011100000",
  38510=>"000011101",
  38511=>"001010101",
  38512=>"001100010",
  38513=>"011100011",
  38514=>"000010010",
  38515=>"000110101",
  38516=>"010000011",
  38517=>"000101100",
  38518=>"010010101",
  38519=>"000000110",
  38520=>"010110001",
  38521=>"101000101",
  38522=>"110010001",
  38523=>"100111001",
  38524=>"100100100",
  38525=>"010010000",
  38526=>"100001110",
  38527=>"000101100",
  38528=>"001000101",
  38529=>"111100000",
  38530=>"000000101",
  38531=>"100100111",
  38532=>"011100101",
  38533=>"101001111",
  38534=>"111001010",
  38535=>"111011000",
  38536=>"100000001",
  38537=>"110101000",
  38538=>"010111111",
  38539=>"111100100",
  38540=>"011100010",
  38541=>"001001000",
  38542=>"101010011",
  38543=>"001100000",
  38544=>"011111110",
  38545=>"011011100",
  38546=>"010101110",
  38547=>"001001000",
  38548=>"010011101",
  38549=>"101000001",
  38550=>"101101000",
  38551=>"010010000",
  38552=>"100010110",
  38553=>"111011101",
  38554=>"000011111",
  38555=>"111110111",
  38556=>"111001100",
  38557=>"000001011",
  38558=>"011111101",
  38559=>"111110101",
  38560=>"000000111",
  38561=>"110000111",
  38562=>"000000100",
  38563=>"010000001",
  38564=>"100000110",
  38565=>"000011100",
  38566=>"000011001",
  38567=>"000101000",
  38568=>"011110010",
  38569=>"101001111",
  38570=>"010100001",
  38571=>"010001011",
  38572=>"110111010",
  38573=>"010110001",
  38574=>"111111101",
  38575=>"101000110",
  38576=>"100000000",
  38577=>"111011101",
  38578=>"100011101",
  38579=>"011000001",
  38580=>"110101101",
  38581=>"001101111",
  38582=>"111001000",
  38583=>"011100001",
  38584=>"010100011",
  38585=>"000101101",
  38586=>"111111011",
  38587=>"011011000",
  38588=>"111001101",
  38589=>"010001001",
  38590=>"101100110",
  38591=>"101111001",
  38592=>"011011100",
  38593=>"101010101",
  38594=>"000001001",
  38595=>"101011000",
  38596=>"010001110",
  38597=>"011100110",
  38598=>"110011000",
  38599=>"101000111",
  38600=>"111111010",
  38601=>"000101010",
  38602=>"110001010",
  38603=>"100011001",
  38604=>"010000001",
  38605=>"100000011",
  38606=>"000010000",
  38607=>"011101111",
  38608=>"010011111",
  38609=>"101000011",
  38610=>"110011101",
  38611=>"000101010",
  38612=>"100010110",
  38613=>"100101100",
  38614=>"011010111",
  38615=>"010110101",
  38616=>"001101011",
  38617=>"001011011",
  38618=>"010110000",
  38619=>"011011111",
  38620=>"100111010",
  38621=>"100000001",
  38622=>"101111000",
  38623=>"100111000",
  38624=>"000100011",
  38625=>"000011000",
  38626=>"011110000",
  38627=>"110011000",
  38628=>"001001011",
  38629=>"010001000",
  38630=>"001000101",
  38631=>"000110001",
  38632=>"001110001",
  38633=>"111110000",
  38634=>"111111000",
  38635=>"011011110",
  38636=>"011111101",
  38637=>"100100000",
  38638=>"111110010",
  38639=>"110010110",
  38640=>"111001010",
  38641=>"100110110",
  38642=>"010010110",
  38643=>"001010010",
  38644=>"110010110",
  38645=>"111101110",
  38646=>"100011110",
  38647=>"010010111",
  38648=>"000100110",
  38649=>"001100101",
  38650=>"000100000",
  38651=>"001000101",
  38652=>"110000101",
  38653=>"010100011",
  38654=>"000010101",
  38655=>"110010000",
  38656=>"111000010",
  38657=>"110101110",
  38658=>"000110100",
  38659=>"100110100",
  38660=>"100001000",
  38661=>"101000011",
  38662=>"110000010",
  38663=>"100101100",
  38664=>"100000100",
  38665=>"100111010",
  38666=>"101111101",
  38667=>"101100001",
  38668=>"101001000",
  38669=>"100001110",
  38670=>"011000000",
  38671=>"110100000",
  38672=>"101101000",
  38673=>"110001110",
  38674=>"100111001",
  38675=>"101000101",
  38676=>"000100100",
  38677=>"100110010",
  38678=>"101110010",
  38679=>"100001111",
  38680=>"001001011",
  38681=>"001001000",
  38682=>"111101111",
  38683=>"011010110",
  38684=>"110100000",
  38685=>"110010001",
  38686=>"000111110",
  38687=>"111111100",
  38688=>"010101101",
  38689=>"101010111",
  38690=>"000000101",
  38691=>"000001011",
  38692=>"010111010",
  38693=>"111010000",
  38694=>"111111110",
  38695=>"100001110",
  38696=>"000101110",
  38697=>"101000101",
  38698=>"000110101",
  38699=>"100110001",
  38700=>"101001000",
  38701=>"010000000",
  38702=>"010010011",
  38703=>"110111011",
  38704=>"011001110",
  38705=>"110000001",
  38706=>"000101000",
  38707=>"111111101",
  38708=>"111100110",
  38709=>"010110001",
  38710=>"110011110",
  38711=>"100100010",
  38712=>"110111111",
  38713=>"100101100",
  38714=>"000101000",
  38715=>"001100101",
  38716=>"111100110",
  38717=>"001011000",
  38718=>"010011001",
  38719=>"001110101",
  38720=>"110011110",
  38721=>"101110001",
  38722=>"100111110",
  38723=>"001110010",
  38724=>"010000010",
  38725=>"111100101",
  38726=>"000111001",
  38727=>"111111100",
  38728=>"010000011",
  38729=>"000110001",
  38730=>"010000011",
  38731=>"001000010",
  38732=>"011010110",
  38733=>"100000100",
  38734=>"101100001",
  38735=>"110100100",
  38736=>"011100001",
  38737=>"001000010",
  38738=>"001011001",
  38739=>"000111111",
  38740=>"101101101",
  38741=>"101011011",
  38742=>"100110110",
  38743=>"101001010",
  38744=>"001100011",
  38745=>"010110100",
  38746=>"001011001",
  38747=>"000100010",
  38748=>"000001010",
  38749=>"110110100",
  38750=>"101011110",
  38751=>"001001100",
  38752=>"011011100",
  38753=>"011011000",
  38754=>"001000101",
  38755=>"111101110",
  38756=>"010110010",
  38757=>"110110111",
  38758=>"111110010",
  38759=>"111111000",
  38760=>"000101110",
  38761=>"010010010",
  38762=>"101100100",
  38763=>"101011001",
  38764=>"001111011",
  38765=>"110110111",
  38766=>"111101110",
  38767=>"101101101",
  38768=>"000000000",
  38769=>"100111010",
  38770=>"010100001",
  38771=>"111010101",
  38772=>"001010001",
  38773=>"001011110",
  38774=>"000000010",
  38775=>"111011010",
  38776=>"001001000",
  38777=>"110011110",
  38778=>"110001110",
  38779=>"011001001",
  38780=>"000001000",
  38781=>"010110111",
  38782=>"110000110",
  38783=>"011111110",
  38784=>"000010001",
  38785=>"001100011",
  38786=>"000010100",
  38787=>"111101001",
  38788=>"001010100",
  38789=>"000010100",
  38790=>"001010100",
  38791=>"110011011",
  38792=>"110101110",
  38793=>"000110010",
  38794=>"001111000",
  38795=>"100110111",
  38796=>"010000110",
  38797=>"111101110",
  38798=>"110011000",
  38799=>"110011100",
  38800=>"000001110",
  38801=>"111101100",
  38802=>"000000100",
  38803=>"001100000",
  38804=>"000010001",
  38805=>"110000110",
  38806=>"001111101",
  38807=>"011110001",
  38808=>"000011000",
  38809=>"000101001",
  38810=>"101111100",
  38811=>"110111100",
  38812=>"100100111",
  38813=>"001001100",
  38814=>"011000100",
  38815=>"000011011",
  38816=>"001010110",
  38817=>"110010101",
  38818=>"000010001",
  38819=>"000000100",
  38820=>"100011011",
  38821=>"010011000",
  38822=>"010000001",
  38823=>"001011111",
  38824=>"000011111",
  38825=>"000000000",
  38826=>"101101010",
  38827=>"000110000",
  38828=>"011000011",
  38829=>"000000010",
  38830=>"101100001",
  38831=>"110110100",
  38832=>"000000011",
  38833=>"111101100",
  38834=>"101110100",
  38835=>"110000001",
  38836=>"010000111",
  38837=>"000001111",
  38838=>"010101100",
  38839=>"011100011",
  38840=>"100000100",
  38841=>"010111101",
  38842=>"110101100",
  38843=>"101101001",
  38844=>"111101111",
  38845=>"011101001",
  38846=>"011000100",
  38847=>"101111010",
  38848=>"110111010",
  38849=>"011111101",
  38850=>"010100110",
  38851=>"010110100",
  38852=>"110010110",
  38853=>"110010101",
  38854=>"110100010",
  38855=>"111000000",
  38856=>"011011111",
  38857=>"100011110",
  38858=>"100110011",
  38859=>"000100010",
  38860=>"100110101",
  38861=>"100010001",
  38862=>"101011000",
  38863=>"111010001",
  38864=>"001100010",
  38865=>"001110000",
  38866=>"000000001",
  38867=>"101001000",
  38868=>"001000100",
  38869=>"010001110",
  38870=>"110100001",
  38871=>"011000001",
  38872=>"000100000",
  38873=>"001001001",
  38874=>"100000011",
  38875=>"100000101",
  38876=>"110010011",
  38877=>"111110111",
  38878=>"000010011",
  38879=>"110101000",
  38880=>"001001110",
  38881=>"100011000",
  38882=>"110011001",
  38883=>"101010000",
  38884=>"100001100",
  38885=>"110100111",
  38886=>"011010001",
  38887=>"000100110",
  38888=>"100110100",
  38889=>"001001111",
  38890=>"110111011",
  38891=>"010100101",
  38892=>"010000101",
  38893=>"000111011",
  38894=>"110100110",
  38895=>"101100100",
  38896=>"100011111",
  38897=>"011010101",
  38898=>"100101010",
  38899=>"100100000",
  38900=>"111000100",
  38901=>"101110010",
  38902=>"101110000",
  38903=>"111100011",
  38904=>"100110110",
  38905=>"111111100",
  38906=>"111000111",
  38907=>"011010011",
  38908=>"001001010",
  38909=>"001100001",
  38910=>"100110011",
  38911=>"100110000",
  38912=>"100011001",
  38913=>"000100000",
  38914=>"011011001",
  38915=>"111100011",
  38916=>"111110111",
  38917=>"101011111",
  38918=>"111101001",
  38919=>"011100111",
  38920=>"110101100",
  38921=>"000000110",
  38922=>"011100101",
  38923=>"011110001",
  38924=>"111100001",
  38925=>"100000000",
  38926=>"010100011",
  38927=>"001111111",
  38928=>"000100001",
  38929=>"111011111",
  38930=>"001111101",
  38931=>"110111111",
  38932=>"000100101",
  38933=>"101101000",
  38934=>"000111000",
  38935=>"010011011",
  38936=>"100011011",
  38937=>"000000001",
  38938=>"011110010",
  38939=>"101110000",
  38940=>"111111101",
  38941=>"110111111",
  38942=>"100101101",
  38943=>"100111100",
  38944=>"010001100",
  38945=>"011000101",
  38946=>"111011011",
  38947=>"101110001",
  38948=>"110010101",
  38949=>"011101100",
  38950=>"110010110",
  38951=>"010001001",
  38952=>"101001101",
  38953=>"000111110",
  38954=>"010001110",
  38955=>"000111100",
  38956=>"011101100",
  38957=>"100010010",
  38958=>"001001101",
  38959=>"001001100",
  38960=>"110001010",
  38961=>"001100100",
  38962=>"111101000",
  38963=>"010000101",
  38964=>"000011011",
  38965=>"010100110",
  38966=>"101001010",
  38967=>"010011111",
  38968=>"010000100",
  38969=>"100101000",
  38970=>"001010011",
  38971=>"000110011",
  38972=>"001110000",
  38973=>"110100000",
  38974=>"101000101",
  38975=>"010110110",
  38976=>"111011001",
  38977=>"100110101",
  38978=>"100101100",
  38979=>"001001000",
  38980=>"011001001",
  38981=>"101101111",
  38982=>"010001011",
  38983=>"001000001",
  38984=>"011111101",
  38985=>"111000111",
  38986=>"000001000",
  38987=>"000010011",
  38988=>"101101000",
  38989=>"001101010",
  38990=>"011000111",
  38991=>"111000000",
  38992=>"011011010",
  38993=>"011111001",
  38994=>"011111100",
  38995=>"111010100",
  38996=>"100011000",
  38997=>"101100101",
  38998=>"111000000",
  38999=>"101000011",
  39000=>"011101010",
  39001=>"000100101",
  39002=>"111011010",
  39003=>"010010000",
  39004=>"010000110",
  39005=>"010010001",
  39006=>"001000101",
  39007=>"000001000",
  39008=>"111101000",
  39009=>"001010001",
  39010=>"101000101",
  39011=>"101111011",
  39012=>"010100110",
  39013=>"110000001",
  39014=>"000000110",
  39015=>"000010101",
  39016=>"010010100",
  39017=>"010101001",
  39018=>"001110001",
  39019=>"100101011",
  39020=>"110011110",
  39021=>"000011100",
  39022=>"011111110",
  39023=>"100101101",
  39024=>"001011110",
  39025=>"111111010",
  39026=>"010000010",
  39027=>"000011100",
  39028=>"000111111",
  39029=>"100011100",
  39030=>"110010010",
  39031=>"111000110",
  39032=>"110011110",
  39033=>"110111111",
  39034=>"000000000",
  39035=>"010101111",
  39036=>"000000101",
  39037=>"001011000",
  39038=>"000110100",
  39039=>"100001001",
  39040=>"001101010",
  39041=>"000110100",
  39042=>"001111011",
  39043=>"110001000",
  39044=>"111101111",
  39045=>"010110111",
  39046=>"011011101",
  39047=>"001011011",
  39048=>"100110111",
  39049=>"001101100",
  39050=>"010101101",
  39051=>"001000100",
  39052=>"111101100",
  39053=>"010111011",
  39054=>"011100001",
  39055=>"101111111",
  39056=>"111101010",
  39057=>"110001000",
  39058=>"110000000",
  39059=>"000110100",
  39060=>"010110110",
  39061=>"100101010",
  39062=>"110010110",
  39063=>"000010101",
  39064=>"001110110",
  39065=>"101101100",
  39066=>"010001110",
  39067=>"000000010",
  39068=>"010001001",
  39069=>"000001100",
  39070=>"011100000",
  39071=>"010111010",
  39072=>"101100101",
  39073=>"111101001",
  39074=>"000110111",
  39075=>"011101000",
  39076=>"100010010",
  39077=>"101101010",
  39078=>"000010111",
  39079=>"100101111",
  39080=>"000000011",
  39081=>"011110110",
  39082=>"101100011",
  39083=>"110011001",
  39084=>"001011101",
  39085=>"110110110",
  39086=>"001101100",
  39087=>"011000001",
  39088=>"111010110",
  39089=>"111011001",
  39090=>"100001111",
  39091=>"111001010",
  39092=>"100000111",
  39093=>"010101011",
  39094=>"101000011",
  39095=>"101010101",
  39096=>"110101001",
  39097=>"100110001",
  39098=>"000000110",
  39099=>"110110111",
  39100=>"111011001",
  39101=>"010001111",
  39102=>"101000010",
  39103=>"001001100",
  39104=>"101010011",
  39105=>"100101000",
  39106=>"100110110",
  39107=>"011100011",
  39108=>"011011001",
  39109=>"111110100",
  39110=>"000011100",
  39111=>"111111000",
  39112=>"111101110",
  39113=>"111000101",
  39114=>"010010000",
  39115=>"101100100",
  39116=>"010010010",
  39117=>"001011000",
  39118=>"001011110",
  39119=>"110001111",
  39120=>"110001101",
  39121=>"101110010",
  39122=>"010011111",
  39123=>"110000110",
  39124=>"011000010",
  39125=>"000111110",
  39126=>"010001100",
  39127=>"001111101",
  39128=>"101110001",
  39129=>"111000010",
  39130=>"101101101",
  39131=>"111111111",
  39132=>"111001001",
  39133=>"010001000",
  39134=>"100001110",
  39135=>"101010101",
  39136=>"100011110",
  39137=>"001011101",
  39138=>"010111011",
  39139=>"110101100",
  39140=>"110110011",
  39141=>"100111001",
  39142=>"111010001",
  39143=>"011001010",
  39144=>"010010001",
  39145=>"011101011",
  39146=>"110011111",
  39147=>"010011000",
  39148=>"101100100",
  39149=>"000111100",
  39150=>"001010001",
  39151=>"001101110",
  39152=>"100100101",
  39153=>"101111110",
  39154=>"001101001",
  39155=>"001001000",
  39156=>"101000001",
  39157=>"111000011",
  39158=>"001011111",
  39159=>"001001110",
  39160=>"010010100",
  39161=>"100001000",
  39162=>"110101011",
  39163=>"000000111",
  39164=>"001100100",
  39165=>"011101100",
  39166=>"011110001",
  39167=>"001000010",
  39168=>"011100011",
  39169=>"001000101",
  39170=>"001111001",
  39171=>"000111001",
  39172=>"110001100",
  39173=>"001001011",
  39174=>"101011000",
  39175=>"011001111",
  39176=>"000111011",
  39177=>"010111010",
  39178=>"001011110",
  39179=>"101111101",
  39180=>"111010010",
  39181=>"001110110",
  39182=>"010011100",
  39183=>"101010000",
  39184=>"000000100",
  39185=>"100011100",
  39186=>"101110000",
  39187=>"110011110",
  39188=>"111010000",
  39189=>"001111100",
  39190=>"110110010",
  39191=>"000110101",
  39192=>"000000011",
  39193=>"010001000",
  39194=>"111110100",
  39195=>"100100001",
  39196=>"010010000",
  39197=>"101010000",
  39198=>"000001000",
  39199=>"101000110",
  39200=>"101010101",
  39201=>"000001111",
  39202=>"110010011",
  39203=>"100000100",
  39204=>"000001111",
  39205=>"000000011",
  39206=>"011100010",
  39207=>"001111010",
  39208=>"101101010",
  39209=>"010000011",
  39210=>"000011100",
  39211=>"001100000",
  39212=>"110111101",
  39213=>"011111110",
  39214=>"111100011",
  39215=>"100011001",
  39216=>"011100111",
  39217=>"111100100",
  39218=>"010011011",
  39219=>"000000010",
  39220=>"110100001",
  39221=>"010101000",
  39222=>"010010100",
  39223=>"010110000",
  39224=>"000000100",
  39225=>"100001011",
  39226=>"110010111",
  39227=>"110011001",
  39228=>"110000011",
  39229=>"001001011",
  39230=>"000000001",
  39231=>"010010001",
  39232=>"111101000",
  39233=>"101010010",
  39234=>"010010101",
  39235=>"100011001",
  39236=>"100110101",
  39237=>"000110000",
  39238=>"010000000",
  39239=>"011000011",
  39240=>"001010110",
  39241=>"110000010",
  39242=>"000000001",
  39243=>"000010001",
  39244=>"010010111",
  39245=>"101001110",
  39246=>"001100000",
  39247=>"010000111",
  39248=>"101001000",
  39249=>"010010111",
  39250=>"000011001",
  39251=>"000001111",
  39252=>"101000001",
  39253=>"100010110",
  39254=>"000010001",
  39255=>"001101101",
  39256=>"010111000",
  39257=>"011101101",
  39258=>"110110100",
  39259=>"011001101",
  39260=>"101011101",
  39261=>"111110111",
  39262=>"100000010",
  39263=>"011101110",
  39264=>"010110100",
  39265=>"011011000",
  39266=>"010011100",
  39267=>"100001100",
  39268=>"001001000",
  39269=>"100001000",
  39270=>"001011010",
  39271=>"011111000",
  39272=>"100101001",
  39273=>"110010111",
  39274=>"101000100",
  39275=>"110101001",
  39276=>"000001010",
  39277=>"010100110",
  39278=>"011010111",
  39279=>"011110111",
  39280=>"000101101",
  39281=>"110111110",
  39282=>"001101101",
  39283=>"110101111",
  39284=>"111001000",
  39285=>"000101010",
  39286=>"000000001",
  39287=>"101110001",
  39288=>"010010100",
  39289=>"010111000",
  39290=>"110000110",
  39291=>"001000010",
  39292=>"100010100",
  39293=>"111100111",
  39294=>"011011110",
  39295=>"001010100",
  39296=>"111111101",
  39297=>"100001111",
  39298=>"110101100",
  39299=>"101111101",
  39300=>"110100111",
  39301=>"101000110",
  39302=>"011100001",
  39303=>"111110101",
  39304=>"000110000",
  39305=>"111000011",
  39306=>"000101111",
  39307=>"010100110",
  39308=>"000011101",
  39309=>"101101101",
  39310=>"011001010",
  39311=>"010100100",
  39312=>"011011100",
  39313=>"010000100",
  39314=>"010000010",
  39315=>"110110000",
  39316=>"010000100",
  39317=>"000110011",
  39318=>"001000010",
  39319=>"000001101",
  39320=>"000101101",
  39321=>"000101000",
  39322=>"000010000",
  39323=>"001001011",
  39324=>"011110000",
  39325=>"111111111",
  39326=>"100100000",
  39327=>"010011000",
  39328=>"111110000",
  39329=>"111110100",
  39330=>"101000000",
  39331=>"011100110",
  39332=>"011010011",
  39333=>"000100000",
  39334=>"111011111",
  39335=>"001001001",
  39336=>"110101111",
  39337=>"100001001",
  39338=>"000100101",
  39339=>"000000010",
  39340=>"001000100",
  39341=>"111011100",
  39342=>"011111011",
  39343=>"000001010",
  39344=>"010110010",
  39345=>"000100001",
  39346=>"110100011",
  39347=>"001010011",
  39348=>"111110111",
  39349=>"011100001",
  39350=>"110011101",
  39351=>"100111001",
  39352=>"000100101",
  39353=>"010001111",
  39354=>"000100010",
  39355=>"101000101",
  39356=>"100010011",
  39357=>"001111100",
  39358=>"000000011",
  39359=>"110000110",
  39360=>"100100000",
  39361=>"000111100",
  39362=>"101100011",
  39363=>"100100111",
  39364=>"011010100",
  39365=>"111110110",
  39366=>"011100000",
  39367=>"000011011",
  39368=>"000101011",
  39369=>"000011000",
  39370=>"000011000",
  39371=>"100001010",
  39372=>"001101010",
  39373=>"111111001",
  39374=>"111011000",
  39375=>"010010010",
  39376=>"111110000",
  39377=>"010011110",
  39378=>"101100100",
  39379=>"001111110",
  39380=>"000000001",
  39381=>"001111011",
  39382=>"011011001",
  39383=>"100100000",
  39384=>"010010100",
  39385=>"110101001",
  39386=>"110010010",
  39387=>"101010100",
  39388=>"011110111",
  39389=>"110010100",
  39390=>"111001111",
  39391=>"011101000",
  39392=>"110010011",
  39393=>"100100100",
  39394=>"100010100",
  39395=>"000100101",
  39396=>"101110110",
  39397=>"101011111",
  39398=>"001110001",
  39399=>"110000011",
  39400=>"000001000",
  39401=>"011100011",
  39402=>"101011011",
  39403=>"010001100",
  39404=>"011010001",
  39405=>"001011100",
  39406=>"000010110",
  39407=>"001100011",
  39408=>"111000100",
  39409=>"000111011",
  39410=>"001011010",
  39411=>"010011000",
  39412=>"010101000",
  39413=>"101110011",
  39414=>"101000110",
  39415=>"010000111",
  39416=>"011101111",
  39417=>"110010001",
  39418=>"100110100",
  39419=>"101011001",
  39420=>"011000000",
  39421=>"000011111",
  39422=>"100101110",
  39423=>"011111000",
  39424=>"100111011",
  39425=>"100011110",
  39426=>"111111011",
  39427=>"010011111",
  39428=>"010110110",
  39429=>"011100010",
  39430=>"001101000",
  39431=>"101001000",
  39432=>"111101001",
  39433=>"011011111",
  39434=>"010000011",
  39435=>"101111110",
  39436=>"100001100",
  39437=>"010001100",
  39438=>"110100100",
  39439=>"001010110",
  39440=>"000110111",
  39441=>"101100111",
  39442=>"000010010",
  39443=>"111110011",
  39444=>"110001001",
  39445=>"101110111",
  39446=>"001011000",
  39447=>"010001000",
  39448=>"011001010",
  39449=>"000111010",
  39450=>"110001000",
  39451=>"111000100",
  39452=>"000011101",
  39453=>"011011111",
  39454=>"111111111",
  39455=>"000110100",
  39456=>"101100010",
  39457=>"000010010",
  39458=>"111110100",
  39459=>"000100011",
  39460=>"010001111",
  39461=>"011110011",
  39462=>"100110001",
  39463=>"000000000",
  39464=>"000110010",
  39465=>"001000010",
  39466=>"101011101",
  39467=>"110011010",
  39468=>"010100000",
  39469=>"100100000",
  39470=>"010100000",
  39471=>"111101111",
  39472=>"010101001",
  39473=>"010110111",
  39474=>"000110100",
  39475=>"100010001",
  39476=>"100101011",
  39477=>"001011101",
  39478=>"110100000",
  39479=>"010000000",
  39480=>"111001111",
  39481=>"101011010",
  39482=>"110100011",
  39483=>"000010001",
  39484=>"100011000",
  39485=>"101100000",
  39486=>"110111000",
  39487=>"001001011",
  39488=>"111000101",
  39489=>"011100110",
  39490=>"111010100",
  39491=>"000001100",
  39492=>"000100110",
  39493=>"111000000",
  39494=>"100001010",
  39495=>"010011110",
  39496=>"110001110",
  39497=>"101011110",
  39498=>"010111001",
  39499=>"101101000",
  39500=>"011011010",
  39501=>"000110100",
  39502=>"000100001",
  39503=>"001000110",
  39504=>"011100110",
  39505=>"000011111",
  39506=>"111010100",
  39507=>"011001001",
  39508=>"101100001",
  39509=>"010100111",
  39510=>"101011000",
  39511=>"000010110",
  39512=>"100001100",
  39513=>"101100110",
  39514=>"000001111",
  39515=>"111001010",
  39516=>"000001111",
  39517=>"000110000",
  39518=>"111010011",
  39519=>"100001101",
  39520=>"001010000",
  39521=>"010000011",
  39522=>"110010001",
  39523=>"011000100",
  39524=>"000010011",
  39525=>"010000110",
  39526=>"000101101",
  39527=>"100100100",
  39528=>"111001111",
  39529=>"100000010",
  39530=>"001001000",
  39531=>"110000000",
  39532=>"010010110",
  39533=>"100001001",
  39534=>"110111010",
  39535=>"011011001",
  39536=>"000110101",
  39537=>"100100101",
  39538=>"100110100",
  39539=>"001111000",
  39540=>"101111001",
  39541=>"000111010",
  39542=>"000111010",
  39543=>"100011111",
  39544=>"110110111",
  39545=>"000011101",
  39546=>"000100000",
  39547=>"111001000",
  39548=>"111010100",
  39549=>"110001111",
  39550=>"011011000",
  39551=>"110001101",
  39552=>"001000111",
  39553=>"001000111",
  39554=>"111111011",
  39555=>"110101001",
  39556=>"110010111",
  39557=>"110101101",
  39558=>"011000000",
  39559=>"101100000",
  39560=>"100001011",
  39561=>"011100001",
  39562=>"101000010",
  39563=>"111101111",
  39564=>"111100111",
  39565=>"101110110",
  39566=>"000000001",
  39567=>"000000000",
  39568=>"001100011",
  39569=>"111011000",
  39570=>"100000010",
  39571=>"001001001",
  39572=>"111001100",
  39573=>"111001011",
  39574=>"001111100",
  39575=>"010001010",
  39576=>"111011010",
  39577=>"111101001",
  39578=>"000000111",
  39579=>"010111100",
  39580=>"000001100",
  39581=>"100111111",
  39582=>"111110110",
  39583=>"100011011",
  39584=>"011010111",
  39585=>"101101111",
  39586=>"101101000",
  39587=>"100110011",
  39588=>"100011101",
  39589=>"101100010",
  39590=>"001100010",
  39591=>"010001111",
  39592=>"011001111",
  39593=>"011110010",
  39594=>"011001000",
  39595=>"010101101",
  39596=>"100000000",
  39597=>"111100100",
  39598=>"101011001",
  39599=>"111000111",
  39600=>"110001101",
  39601=>"111010011",
  39602=>"010000010",
  39603=>"000000010",
  39604=>"100100111",
  39605=>"010001101",
  39606=>"101010111",
  39607=>"110111111",
  39608=>"000100110",
  39609=>"010001101",
  39610=>"000010000",
  39611=>"001001010",
  39612=>"111111001",
  39613=>"111000101",
  39614=>"010000101",
  39615=>"101000011",
  39616=>"011111110",
  39617=>"100000000",
  39618=>"111000000",
  39619=>"010010000",
  39620=>"110011111",
  39621=>"101001101",
  39622=>"010011001",
  39623=>"001001100",
  39624=>"010010000",
  39625=>"110111001",
  39626=>"011111101",
  39627=>"000111001",
  39628=>"001001001",
  39629=>"001101001",
  39630=>"011000010",
  39631=>"001111010",
  39632=>"000100111",
  39633=>"001111111",
  39634=>"101011100",
  39635=>"010110011",
  39636=>"101111110",
  39637=>"001100101",
  39638=>"010101011",
  39639=>"000111000",
  39640=>"010000000",
  39641=>"010001000",
  39642=>"000010001",
  39643=>"010110000",
  39644=>"010110110",
  39645=>"100100111",
  39646=>"100101101",
  39647=>"110111000",
  39648=>"011100011",
  39649=>"010000001",
  39650=>"010011111",
  39651=>"010000011",
  39652=>"011100011",
  39653=>"010100000",
  39654=>"111001101",
  39655=>"001111011",
  39656=>"011011111",
  39657=>"010110010",
  39658=>"011111101",
  39659=>"010001101",
  39660=>"100010101",
  39661=>"001010110",
  39662=>"100110100",
  39663=>"001111011",
  39664=>"111000111",
  39665=>"011010101",
  39666=>"011001100",
  39667=>"110010100",
  39668=>"101101011",
  39669=>"011011001",
  39670=>"000011111",
  39671=>"011001000",
  39672=>"111001111",
  39673=>"011011101",
  39674=>"011100001",
  39675=>"001101001",
  39676=>"001111111",
  39677=>"000110010",
  39678=>"100001011",
  39679=>"101101000",
  39680=>"011110111",
  39681=>"101111000",
  39682=>"101100011",
  39683=>"000100010",
  39684=>"010000100",
  39685=>"000001011",
  39686=>"100001000",
  39687=>"010101100",
  39688=>"010001101",
  39689=>"011001110",
  39690=>"000110100",
  39691=>"010010011",
  39692=>"010000101",
  39693=>"010101011",
  39694=>"000100011",
  39695=>"001000001",
  39696=>"011100001",
  39697=>"000000101",
  39698=>"100110111",
  39699=>"001111010",
  39700=>"010111100",
  39701=>"001001111",
  39702=>"011111111",
  39703=>"100100011",
  39704=>"110000110",
  39705=>"000001111",
  39706=>"100001110",
  39707=>"101101100",
  39708=>"011000100",
  39709=>"100100010",
  39710=>"101111101",
  39711=>"101001000",
  39712=>"001010010",
  39713=>"111000101",
  39714=>"110001110",
  39715=>"110110110",
  39716=>"101011100",
  39717=>"101111010",
  39718=>"111100001",
  39719=>"011111111",
  39720=>"010110101",
  39721=>"101100001",
  39722=>"001101100",
  39723=>"011010111",
  39724=>"110101101",
  39725=>"101001000",
  39726=>"111100100",
  39727=>"101010110",
  39728=>"000000110",
  39729=>"100001100",
  39730=>"111111101",
  39731=>"000001010",
  39732=>"010111110",
  39733=>"100000100",
  39734=>"101001110",
  39735=>"110011111",
  39736=>"010011110",
  39737=>"100100111",
  39738=>"011100110",
  39739=>"001101011",
  39740=>"101111010",
  39741=>"101110001",
  39742=>"110001001",
  39743=>"100111011",
  39744=>"001011101",
  39745=>"011111010",
  39746=>"110100010",
  39747=>"000101000",
  39748=>"101101000",
  39749=>"010010001",
  39750=>"101001111",
  39751=>"010111111",
  39752=>"110100111",
  39753=>"100100001",
  39754=>"110101100",
  39755=>"011011011",
  39756=>"100000010",
  39757=>"101001011",
  39758=>"010100100",
  39759=>"011000000",
  39760=>"110110000",
  39761=>"100011111",
  39762=>"101111111",
  39763=>"100101101",
  39764=>"011010001",
  39765=>"110111111",
  39766=>"000011010",
  39767=>"011110010",
  39768=>"100100011",
  39769=>"010111010",
  39770=>"010001111",
  39771=>"000101101",
  39772=>"111110100",
  39773=>"011111111",
  39774=>"111000011",
  39775=>"001100111",
  39776=>"110100110",
  39777=>"100000000",
  39778=>"010111000",
  39779=>"000000100",
  39780=>"011000010",
  39781=>"010111011",
  39782=>"010100111",
  39783=>"010010101",
  39784=>"000100100",
  39785=>"101101101",
  39786=>"011100000",
  39787=>"000001110",
  39788=>"010010001",
  39789=>"101101011",
  39790=>"100110011",
  39791=>"011011110",
  39792=>"011011100",
  39793=>"110100101",
  39794=>"111010101",
  39795=>"011101000",
  39796=>"001110111",
  39797=>"010001101",
  39798=>"100110100",
  39799=>"110000110",
  39800=>"011010010",
  39801=>"011011101",
  39802=>"110111011",
  39803=>"001011011",
  39804=>"100000111",
  39805=>"011000011",
  39806=>"000001010",
  39807=>"100010011",
  39808=>"001010110",
  39809=>"000110010",
  39810=>"010101100",
  39811=>"110101000",
  39812=>"010100101",
  39813=>"100010000",
  39814=>"011110100",
  39815=>"000110101",
  39816=>"001010111",
  39817=>"111111011",
  39818=>"111010100",
  39819=>"000011100",
  39820=>"010110100",
  39821=>"101111011",
  39822=>"000011110",
  39823=>"111010010",
  39824=>"010000001",
  39825=>"111111101",
  39826=>"101000110",
  39827=>"010010001",
  39828=>"101101011",
  39829=>"111000101",
  39830=>"110010000",
  39831=>"100001000",
  39832=>"111001001",
  39833=>"111111111",
  39834=>"010101000",
  39835=>"110001001",
  39836=>"100001011",
  39837=>"110001110",
  39838=>"000000100",
  39839=>"100111101",
  39840=>"111011011",
  39841=>"001010001",
  39842=>"001100110",
  39843=>"010011110",
  39844=>"001010101",
  39845=>"101010000",
  39846=>"001000111",
  39847=>"110000100",
  39848=>"001110101",
  39849=>"010000111",
  39850=>"111100100",
  39851=>"000100000",
  39852=>"011010000",
  39853=>"110111001",
  39854=>"010000111",
  39855=>"011101010",
  39856=>"011011000",
  39857=>"001011011",
  39858=>"101111100",
  39859=>"001101000",
  39860=>"011100001",
  39861=>"111110001",
  39862=>"011000110",
  39863=>"001101011",
  39864=>"101011010",
  39865=>"000000010",
  39866=>"100010101",
  39867=>"011111101",
  39868=>"000011111",
  39869=>"100011011",
  39870=>"110110111",
  39871=>"001010001",
  39872=>"011010001",
  39873=>"001000000",
  39874=>"110001011",
  39875=>"000101111",
  39876=>"101010011",
  39877=>"111101000",
  39878=>"111110001",
  39879=>"100011010",
  39880=>"110010011",
  39881=>"100001010",
  39882=>"001010000",
  39883=>"001110110",
  39884=>"110110101",
  39885=>"000001011",
  39886=>"001000100",
  39887=>"010110101",
  39888=>"010000101",
  39889=>"000010011",
  39890=>"111001011",
  39891=>"000000000",
  39892=>"101011101",
  39893=>"011100111",
  39894=>"110001000",
  39895=>"000100110",
  39896=>"100100000",
  39897=>"000010000",
  39898=>"111000011",
  39899=>"110011100",
  39900=>"100011110",
  39901=>"101011010",
  39902=>"001101011",
  39903=>"001010100",
  39904=>"010110111",
  39905=>"011000011",
  39906=>"110110100",
  39907=>"110000010",
  39908=>"001001011",
  39909=>"111111011",
  39910=>"001101101",
  39911=>"000010001",
  39912=>"111111011",
  39913=>"111001111",
  39914=>"001010110",
  39915=>"101110011",
  39916=>"111111111",
  39917=>"010101101",
  39918=>"001101010",
  39919=>"100001110",
  39920=>"010010010",
  39921=>"101001111",
  39922=>"001101100",
  39923=>"101100010",
  39924=>"001010011",
  39925=>"101111110",
  39926=>"110101010",
  39927=>"101101111",
  39928=>"110000001",
  39929=>"101110010",
  39930=>"100010110",
  39931=>"100001110",
  39932=>"110110010",
  39933=>"100100001",
  39934=>"111111000",
  39935=>"101000000",
  39936=>"111000000",
  39937=>"000010110",
  39938=>"100011100",
  39939=>"000100100",
  39940=>"101010010",
  39941=>"110110110",
  39942=>"010010110",
  39943=>"101000101",
  39944=>"011001000",
  39945=>"111100010",
  39946=>"001010001",
  39947=>"011111101",
  39948=>"001011111",
  39949=>"010100110",
  39950=>"110010011",
  39951=>"111110110",
  39952=>"011101001",
  39953=>"010100110",
  39954=>"110101110",
  39955=>"110110110",
  39956=>"111101010",
  39957=>"111101100",
  39958=>"110001000",
  39959=>"000101110",
  39960=>"000011000",
  39961=>"000101100",
  39962=>"110101111",
  39963=>"111011011",
  39964=>"100100111",
  39965=>"101110000",
  39966=>"010101101",
  39967=>"100000010",
  39968=>"110011010",
  39969=>"011110111",
  39970=>"010100100",
  39971=>"100000010",
  39972=>"111001001",
  39973=>"101000011",
  39974=>"111111111",
  39975=>"010110010",
  39976=>"001111011",
  39977=>"111111000",
  39978=>"101011100",
  39979=>"110110110",
  39980=>"000010000",
  39981=>"101111101",
  39982=>"011111010",
  39983=>"101101111",
  39984=>"010011100",
  39985=>"001011000",
  39986=>"011101010",
  39987=>"111111110",
  39988=>"110011100",
  39989=>"100110110",
  39990=>"100110111",
  39991=>"001010100",
  39992=>"111110100",
  39993=>"011000110",
  39994=>"001111111",
  39995=>"100011011",
  39996=>"110100110",
  39997=>"010011011",
  39998=>"101001100",
  39999=>"010111001",
  40000=>"110110111",
  40001=>"010011111",
  40002=>"101001100",
  40003=>"000110111",
  40004=>"100110010",
  40005=>"111000001",
  40006=>"110111111",
  40007=>"111001110",
  40008=>"010111111",
  40009=>"101100100",
  40010=>"011110110",
  40011=>"000010001",
  40012=>"001101110",
  40013=>"010000011",
  40014=>"111110010",
  40015=>"010110010",
  40016=>"000001111",
  40017=>"101110111",
  40018=>"011111101",
  40019=>"010011001",
  40020=>"111011010",
  40021=>"111001010",
  40022=>"110011100",
  40023=>"111001101",
  40024=>"100011101",
  40025=>"001101110",
  40026=>"101010100",
  40027=>"001110110",
  40028=>"110101111",
  40029=>"011100000",
  40030=>"010110100",
  40031=>"000001110",
  40032=>"101010001",
  40033=>"110101001",
  40034=>"110111101",
  40035=>"110111101",
  40036=>"000001000",
  40037=>"010101001",
  40038=>"101011110",
  40039=>"010011111",
  40040=>"010011011",
  40041=>"010100100",
  40042=>"010001010",
  40043=>"010100001",
  40044=>"101110110",
  40045=>"001011001",
  40046=>"011010100",
  40047=>"100111111",
  40048=>"101100001",
  40049=>"111110001",
  40050=>"110011111",
  40051=>"011100111",
  40052=>"001100111",
  40053=>"000011011",
  40054=>"110101100",
  40055=>"101000100",
  40056=>"011001001",
  40057=>"011100110",
  40058=>"100100111",
  40059=>"001111011",
  40060=>"000001111",
  40061=>"001000110",
  40062=>"001010000",
  40063=>"000010010",
  40064=>"100100011",
  40065=>"011101101",
  40066=>"000110111",
  40067=>"010011010",
  40068=>"010100001",
  40069=>"101010101",
  40070=>"100100000",
  40071=>"001101100",
  40072=>"011111110",
  40073=>"100000110",
  40074=>"001000010",
  40075=>"011011100",
  40076=>"011011111",
  40077=>"111011100",
  40078=>"001100011",
  40079=>"100101010",
  40080=>"000001111",
  40081=>"111100101",
  40082=>"000101100",
  40083=>"110000101",
  40084=>"000000100",
  40085=>"011110011",
  40086=>"110100100",
  40087=>"000010110",
  40088=>"111110010",
  40089=>"111100101",
  40090=>"101110010",
  40091=>"110000101",
  40092=>"111100101",
  40093=>"011110111",
  40094=>"101010101",
  40095=>"101100111",
  40096=>"011111101",
  40097=>"110010000",
  40098=>"110000111",
  40099=>"011110101",
  40100=>"010100101",
  40101=>"000111100",
  40102=>"100001101",
  40103=>"010011111",
  40104=>"011011001",
  40105=>"000010110",
  40106=>"011110010",
  40107=>"111000110",
  40108=>"111100101",
  40109=>"111110011",
  40110=>"011111101",
  40111=>"000100010",
  40112=>"001000010",
  40113=>"110100000",
  40114=>"010001111",
  40115=>"001110101",
  40116=>"111000011",
  40117=>"011000111",
  40118=>"110010010",
  40119=>"110001100",
  40120=>"011100110",
  40121=>"000101011",
  40122=>"110101010",
  40123=>"001000100",
  40124=>"100001001",
  40125=>"010100100",
  40126=>"101000011",
  40127=>"000001000",
  40128=>"001100000",
  40129=>"000001000",
  40130=>"001010100",
  40131=>"001110000",
  40132=>"111011001",
  40133=>"110111101",
  40134=>"100011111",
  40135=>"000011000",
  40136=>"111101111",
  40137=>"111101001",
  40138=>"000101110",
  40139=>"011110000",
  40140=>"000110000",
  40141=>"011111001",
  40142=>"100011110",
  40143=>"001000000",
  40144=>"101011000",
  40145=>"011100010",
  40146=>"011010010",
  40147=>"000111001",
  40148=>"010010011",
  40149=>"000000011",
  40150=>"101111011",
  40151=>"010011001",
  40152=>"111111001",
  40153=>"010001101",
  40154=>"111110111",
  40155=>"101010100",
  40156=>"100000101",
  40157=>"101101010",
  40158=>"000010000",
  40159=>"010111011",
  40160=>"110110100",
  40161=>"100100110",
  40162=>"000000101",
  40163=>"101101111",
  40164=>"010101110",
  40165=>"110100111",
  40166=>"010111100",
  40167=>"011010101",
  40168=>"001111101",
  40169=>"100001110",
  40170=>"100100111",
  40171=>"010111000",
  40172=>"111011011",
  40173=>"011110110",
  40174=>"000000110",
  40175=>"100010000",
  40176=>"010011100",
  40177=>"101000010",
  40178=>"110011010",
  40179=>"100001010",
  40180=>"100100000",
  40181=>"010110011",
  40182=>"101101000",
  40183=>"101001110",
  40184=>"100110001",
  40185=>"110100010",
  40186=>"111010110",
  40187=>"100110011",
  40188=>"110011111",
  40189=>"100011110",
  40190=>"110011011",
  40191=>"101010010",
  40192=>"100110101",
  40193=>"001100000",
  40194=>"011001100",
  40195=>"011011101",
  40196=>"110100000",
  40197=>"011011001",
  40198=>"100001100",
  40199=>"111101111",
  40200=>"000111011",
  40201=>"001111001",
  40202=>"011011010",
  40203=>"110110101",
  40204=>"001111111",
  40205=>"000001110",
  40206=>"100110100",
  40207=>"100110111",
  40208=>"100011111",
  40209=>"001111111",
  40210=>"000000110",
  40211=>"111101100",
  40212=>"010101010",
  40213=>"010110111",
  40214=>"010011010",
  40215=>"011101011",
  40216=>"111100110",
  40217=>"110000100",
  40218=>"110011001",
  40219=>"010110010",
  40220=>"000100010",
  40221=>"111100100",
  40222=>"100001100",
  40223=>"000001000",
  40224=>"101110110",
  40225=>"001011100",
  40226=>"000101011",
  40227=>"100110111",
  40228=>"000011011",
  40229=>"110110001",
  40230=>"010000100",
  40231=>"100100010",
  40232=>"111100101",
  40233=>"010101010",
  40234=>"000101111",
  40235=>"011110001",
  40236=>"100101100",
  40237=>"100011111",
  40238=>"001100000",
  40239=>"111001110",
  40240=>"110110011",
  40241=>"100100000",
  40242=>"110001100",
  40243=>"110111100",
  40244=>"010100101",
  40245=>"011001100",
  40246=>"100010001",
  40247=>"001100101",
  40248=>"101111101",
  40249=>"000010101",
  40250=>"100010111",
  40251=>"011101110",
  40252=>"000010010",
  40253=>"000011011",
  40254=>"111110011",
  40255=>"011000000",
  40256=>"111011100",
  40257=>"000001101",
  40258=>"010110110",
  40259=>"111000010",
  40260=>"000111110",
  40261=>"111010010",
  40262=>"000101100",
  40263=>"011110011",
  40264=>"011000110",
  40265=>"001100000",
  40266=>"101010000",
  40267=>"001011111",
  40268=>"011001110",
  40269=>"011110001",
  40270=>"101000010",
  40271=>"111111010",
  40272=>"011111001",
  40273=>"111011010",
  40274=>"111100111",
  40275=>"101111000",
  40276=>"101001000",
  40277=>"111101110",
  40278=>"111100011",
  40279=>"111110100",
  40280=>"101111100",
  40281=>"101011001",
  40282=>"110000011",
  40283=>"000000100",
  40284=>"111101011",
  40285=>"000111001",
  40286=>"000001111",
  40287=>"101101110",
  40288=>"101101101",
  40289=>"001110001",
  40290=>"110111111",
  40291=>"111101111",
  40292=>"011110110",
  40293=>"111010100",
  40294=>"011100010",
  40295=>"101111100",
  40296=>"100011000",
  40297=>"111001101",
  40298=>"001001010",
  40299=>"111001001",
  40300=>"110110110",
  40301=>"101110101",
  40302=>"000100101",
  40303=>"010001001",
  40304=>"010111101",
  40305=>"110101000",
  40306=>"101010101",
  40307=>"110000111",
  40308=>"010100000",
  40309=>"000010000",
  40310=>"110101011",
  40311=>"001010010",
  40312=>"010100100",
  40313=>"111111100",
  40314=>"100111010",
  40315=>"001111011",
  40316=>"101100001",
  40317=>"000010100",
  40318=>"111011011",
  40319=>"110100001",
  40320=>"001010011",
  40321=>"011100010",
  40322=>"001101001",
  40323=>"111111111",
  40324=>"011000010",
  40325=>"101111111",
  40326=>"111010010",
  40327=>"101001010",
  40328=>"010000101",
  40329=>"010000101",
  40330=>"000010000",
  40331=>"101001001",
  40332=>"000001100",
  40333=>"111110110",
  40334=>"101110000",
  40335=>"001101011",
  40336=>"001001110",
  40337=>"010010110",
  40338=>"010110011",
  40339=>"111101101",
  40340=>"100001011",
  40341=>"111111000",
  40342=>"100010111",
  40343=>"001001100",
  40344=>"101100010",
  40345=>"110011000",
  40346=>"001110010",
  40347=>"001000110",
  40348=>"000000000",
  40349=>"011110001",
  40350=>"101100000",
  40351=>"111111111",
  40352=>"111110101",
  40353=>"110101000",
  40354=>"111011010",
  40355=>"111110011",
  40356=>"100111101",
  40357=>"111100000",
  40358=>"011010001",
  40359=>"101101110",
  40360=>"001010100",
  40361=>"001101111",
  40362=>"100101111",
  40363=>"010001011",
  40364=>"100111110",
  40365=>"001001011",
  40366=>"111111011",
  40367=>"111100001",
  40368=>"011011111",
  40369=>"000011110",
  40370=>"010110101",
  40371=>"111011110",
  40372=>"000010100",
  40373=>"100001000",
  40374=>"111010011",
  40375=>"010001011",
  40376=>"110000001",
  40377=>"010111001",
  40378=>"000000001",
  40379=>"110001000",
  40380=>"110100110",
  40381=>"100011111",
  40382=>"111101111",
  40383=>"100111011",
  40384=>"000110110",
  40385=>"001001111",
  40386=>"010000100",
  40387=>"001111001",
  40388=>"010100110",
  40389=>"100111010",
  40390=>"010110010",
  40391=>"001110111",
  40392=>"000111110",
  40393=>"111001111",
  40394=>"010000010",
  40395=>"101100101",
  40396=>"000100000",
  40397=>"101001101",
  40398=>"111001000",
  40399=>"111001111",
  40400=>"111011001",
  40401=>"110111110",
  40402=>"000100000",
  40403=>"001001001",
  40404=>"111101110",
  40405=>"110010111",
  40406=>"110000100",
  40407=>"111001111",
  40408=>"111001001",
  40409=>"110000000",
  40410=>"101000111",
  40411=>"100110000",
  40412=>"111001000",
  40413=>"011011010",
  40414=>"010010100",
  40415=>"110001001",
  40416=>"100100001",
  40417=>"001011010",
  40418=>"101110110",
  40419=>"111110001",
  40420=>"011011000",
  40421=>"110100011",
  40422=>"001101010",
  40423=>"011000100",
  40424=>"110100110",
  40425=>"011100101",
  40426=>"000010000",
  40427=>"110100001",
  40428=>"000000000",
  40429=>"100011101",
  40430=>"011101100",
  40431=>"101111011",
  40432=>"000111001",
  40433=>"010001011",
  40434=>"010010011",
  40435=>"001001011",
  40436=>"101000010",
  40437=>"001001001",
  40438=>"010011001",
  40439=>"101110001",
  40440=>"100001100",
  40441=>"110010010",
  40442=>"010010100",
  40443=>"011101010",
  40444=>"001001100",
  40445=>"110011011",
  40446=>"110011110",
  40447=>"101100111",
  40448=>"011110100",
  40449=>"100011111",
  40450=>"111101000",
  40451=>"100011000",
  40452=>"101110001",
  40453=>"001111000",
  40454=>"010011000",
  40455=>"011001001",
  40456=>"001000101",
  40457=>"000011101",
  40458=>"001110010",
  40459=>"001101000",
  40460=>"100011001",
  40461=>"011100101",
  40462=>"001100001",
  40463=>"010000111",
  40464=>"101001100",
  40465=>"000111010",
  40466=>"101000101",
  40467=>"101111100",
  40468=>"101101000",
  40469=>"100001001",
  40470=>"100000110",
  40471=>"100110010",
  40472=>"111111001",
  40473=>"100011111",
  40474=>"110011001",
  40475=>"000000110",
  40476=>"100110101",
  40477=>"111010111",
  40478=>"111101011",
  40479=>"001111101",
  40480=>"101010001",
  40481=>"110100111",
  40482=>"000001101",
  40483=>"100110110",
  40484=>"101110001",
  40485=>"001101000",
  40486=>"101001011",
  40487=>"100010100",
  40488=>"001111011",
  40489=>"000010001",
  40490=>"110110100",
  40491=>"011010010",
  40492=>"101101111",
  40493=>"010010000",
  40494=>"110100100",
  40495=>"101101100",
  40496=>"111000000",
  40497=>"110100100",
  40498=>"101100100",
  40499=>"110100011",
  40500=>"100111010",
  40501=>"001101001",
  40502=>"001011100",
  40503=>"011100110",
  40504=>"111100011",
  40505=>"010010101",
  40506=>"100100111",
  40507=>"010000000",
  40508=>"111111010",
  40509=>"110100101",
  40510=>"010100001",
  40511=>"011001010",
  40512=>"100110101",
  40513=>"001101001",
  40514=>"000001111",
  40515=>"111100010",
  40516=>"011101110",
  40517=>"000110101",
  40518=>"111000100",
  40519=>"000110100",
  40520=>"111110111",
  40521=>"010000100",
  40522=>"110100110",
  40523=>"110101111",
  40524=>"011101001",
  40525=>"011011100",
  40526=>"010011110",
  40527=>"010110110",
  40528=>"000010011",
  40529=>"010110111",
  40530=>"101110011",
  40531=>"010011110",
  40532=>"100111111",
  40533=>"000011110",
  40534=>"110100001",
  40535=>"111011011",
  40536=>"000110010",
  40537=>"111000000",
  40538=>"101101001",
  40539=>"101101100",
  40540=>"001100000",
  40541=>"111111100",
  40542=>"100100111",
  40543=>"010000101",
  40544=>"000110001",
  40545=>"010001011",
  40546=>"111010101",
  40547=>"001100111",
  40548=>"010111110",
  40549=>"000011111",
  40550=>"001101101",
  40551=>"100101001",
  40552=>"111111111",
  40553=>"100001100",
  40554=>"001001010",
  40555=>"001111011",
  40556=>"000111011",
  40557=>"111101001",
  40558=>"001001101",
  40559=>"100010100",
  40560=>"000001111",
  40561=>"001000111",
  40562=>"101000011",
  40563=>"000111111",
  40564=>"001011001",
  40565=>"100010101",
  40566=>"001100111",
  40567=>"101010100",
  40568=>"110011000",
  40569=>"111001010",
  40570=>"011100010",
  40571=>"111100010",
  40572=>"110000000",
  40573=>"101001000",
  40574=>"010100100",
  40575=>"001101110",
  40576=>"111111110",
  40577=>"101000011",
  40578=>"000111100",
  40579=>"101010110",
  40580=>"111011110",
  40581=>"001001000",
  40582=>"011001001",
  40583=>"001011010",
  40584=>"010010010",
  40585=>"001110111",
  40586=>"101000001",
  40587=>"111000001",
  40588=>"111110001",
  40589=>"111011011",
  40590=>"000100100",
  40591=>"111111110",
  40592=>"101010111",
  40593=>"011001101",
  40594=>"100001100",
  40595=>"010010111",
  40596=>"011101111",
  40597=>"011010011",
  40598=>"100010001",
  40599=>"001000101",
  40600=>"111000101",
  40601=>"001000001",
  40602=>"011010110",
  40603=>"011101111",
  40604=>"110111111",
  40605=>"000011010",
  40606=>"000100000",
  40607=>"111100110",
  40608=>"000110110",
  40609=>"101000010",
  40610=>"111010000",
  40611=>"100100100",
  40612=>"000010010",
  40613=>"000100011",
  40614=>"010000111",
  40615=>"111111101",
  40616=>"100111101",
  40617=>"100000000",
  40618=>"110100000",
  40619=>"000111000",
  40620=>"111011101",
  40621=>"110010111",
  40622=>"101101001",
  40623=>"100011010",
  40624=>"011100101",
  40625=>"001111110",
  40626=>"100100100",
  40627=>"010111111",
  40628=>"111110011",
  40629=>"001011000",
  40630=>"000100100",
  40631=>"111001010",
  40632=>"011011100",
  40633=>"100110011",
  40634=>"111101100",
  40635=>"011111011",
  40636=>"111010110",
  40637=>"011001001",
  40638=>"100111101",
  40639=>"100010101",
  40640=>"010001011",
  40641=>"111010101",
  40642=>"000101010",
  40643=>"101000001",
  40644=>"110001110",
  40645=>"101001000",
  40646=>"101010101",
  40647=>"001010011",
  40648=>"010111000",
  40649=>"101111111",
  40650=>"011011101",
  40651=>"000100011",
  40652=>"111111001",
  40653=>"000100101",
  40654=>"100000111",
  40655=>"100000000",
  40656=>"011111010",
  40657=>"000000001",
  40658=>"101010100",
  40659=>"011110000",
  40660=>"000011110",
  40661=>"101111101",
  40662=>"100011101",
  40663=>"101100011",
  40664=>"001001110",
  40665=>"100010001",
  40666=>"010100100",
  40667=>"100100011",
  40668=>"111001000",
  40669=>"100111011",
  40670=>"000111110",
  40671=>"011010111",
  40672=>"001111100",
  40673=>"101101001",
  40674=>"100110111",
  40675=>"111011110",
  40676=>"010111010",
  40677=>"111001100",
  40678=>"100111011",
  40679=>"110010111",
  40680=>"010000010",
  40681=>"101101011",
  40682=>"101110000",
  40683=>"011010100",
  40684=>"110111101",
  40685=>"100001111",
  40686=>"111100000",
  40687=>"101001001",
  40688=>"001011110",
  40689=>"111001100",
  40690=>"011101110",
  40691=>"111101100",
  40692=>"100110110",
  40693=>"111011010",
  40694=>"001000100",
  40695=>"011100001",
  40696=>"101110100",
  40697=>"001001110",
  40698=>"000010001",
  40699=>"100010101",
  40700=>"001001100",
  40701=>"101001011",
  40702=>"100011000",
  40703=>"000101001",
  40704=>"000001000",
  40705=>"100010110",
  40706=>"010011010",
  40707=>"100001111",
  40708=>"011010001",
  40709=>"101011111",
  40710=>"100100000",
  40711=>"110101111",
  40712=>"101100100",
  40713=>"000111101",
  40714=>"010000110",
  40715=>"110000000",
  40716=>"110101111",
  40717=>"110111100",
  40718=>"010001010",
  40719=>"110000010",
  40720=>"111111110",
  40721=>"100100111",
  40722=>"101101101",
  40723=>"111000010",
  40724=>"010101000",
  40725=>"000010100",
  40726=>"011010000",
  40727=>"000010101",
  40728=>"011001001",
  40729=>"111001100",
  40730=>"010111000",
  40731=>"111001111",
  40732=>"101111101",
  40733=>"100000100",
  40734=>"110111111",
  40735=>"000010110",
  40736=>"100010101",
  40737=>"110101000",
  40738=>"101111011",
  40739=>"111001101",
  40740=>"001011111",
  40741=>"110110110",
  40742=>"010011110",
  40743=>"010000000",
  40744=>"110100101",
  40745=>"011111011",
  40746=>"110001001",
  40747=>"100000110",
  40748=>"110001011",
  40749=>"111010010",
  40750=>"000001110",
  40751=>"100111001",
  40752=>"011101110",
  40753=>"110001111",
  40754=>"101111110",
  40755=>"101100101",
  40756=>"010000110",
  40757=>"000110010",
  40758=>"110010101",
  40759=>"011100111",
  40760=>"100000000",
  40761=>"111001010",
  40762=>"111110101",
  40763=>"100110000",
  40764=>"100010111",
  40765=>"111100010",
  40766=>"011101101",
  40767=>"101011101",
  40768=>"011010100",
  40769=>"010011100",
  40770=>"100101110",
  40771=>"111111110",
  40772=>"001101111",
  40773=>"110111111",
  40774=>"100101101",
  40775=>"111101011",
  40776=>"010100001",
  40777=>"101110101",
  40778=>"101111101",
  40779=>"111010001",
  40780=>"110100011",
  40781=>"111101110",
  40782=>"011000111",
  40783=>"000001010",
  40784=>"000100100",
  40785=>"101000111",
  40786=>"100001001",
  40787=>"011111110",
  40788=>"001101000",
  40789=>"110100011",
  40790=>"001110000",
  40791=>"111100100",
  40792=>"010111100",
  40793=>"011011110",
  40794=>"011000100",
  40795=>"011000101",
  40796=>"111100011",
  40797=>"011110011",
  40798=>"110010110",
  40799=>"000010100",
  40800=>"110001110",
  40801=>"101101100",
  40802=>"100011011",
  40803=>"101001001",
  40804=>"001000010",
  40805=>"111010111",
  40806=>"001110100",
  40807=>"010010001",
  40808=>"011110011",
  40809=>"001110110",
  40810=>"111010001",
  40811=>"000111010",
  40812=>"100101100",
  40813=>"110110101",
  40814=>"111110010",
  40815=>"101011000",
  40816=>"110000010",
  40817=>"111010110",
  40818=>"111001100",
  40819=>"101101000",
  40820=>"111110011",
  40821=>"000111111",
  40822=>"000111111",
  40823=>"111010011",
  40824=>"010010101",
  40825=>"111100001",
  40826=>"100101100",
  40827=>"000000000",
  40828=>"011011011",
  40829=>"010100001",
  40830=>"101110111",
  40831=>"101011111",
  40832=>"011010010",
  40833=>"011111011",
  40834=>"111111101",
  40835=>"011011111",
  40836=>"010110001",
  40837=>"011110100",
  40838=>"010010111",
  40839=>"010101011",
  40840=>"011011111",
  40841=>"101011011",
  40842=>"010110010",
  40843=>"100000010",
  40844=>"011111110",
  40845=>"010111110",
  40846=>"111010101",
  40847=>"110110011",
  40848=>"100010000",
  40849=>"101100101",
  40850=>"110011110",
  40851=>"000111000",
  40852=>"000011111",
  40853=>"000011000",
  40854=>"101001001",
  40855=>"001001110",
  40856=>"111010111",
  40857=>"110001110",
  40858=>"000000111",
  40859=>"011100111",
  40860=>"110000001",
  40861=>"001001110",
  40862=>"001110001",
  40863=>"100011100",
  40864=>"111111000",
  40865=>"111110111",
  40866=>"000111010",
  40867=>"010011111",
  40868=>"100001001",
  40869=>"001001110",
  40870=>"110111000",
  40871=>"001000000",
  40872=>"001010110",
  40873=>"100101001",
  40874=>"100010110",
  40875=>"001101101",
  40876=>"111100000",
  40877=>"110101010",
  40878=>"010110010",
  40879=>"001000101",
  40880=>"101000011",
  40881=>"110001101",
  40882=>"110011111",
  40883=>"011100110",
  40884=>"000100100",
  40885=>"100011101",
  40886=>"011001000",
  40887=>"010010010",
  40888=>"000100010",
  40889=>"000110100",
  40890=>"001100000",
  40891=>"101100000",
  40892=>"000001111",
  40893=>"010100010",
  40894=>"000000110",
  40895=>"001101110",
  40896=>"110101111",
  40897=>"101101101",
  40898=>"111000000",
  40899=>"000011010",
  40900=>"100100010",
  40901=>"101110000",
  40902=>"001000000",
  40903=>"001000010",
  40904=>"100010110",
  40905=>"000011010",
  40906=>"101011010",
  40907=>"000100100",
  40908=>"100100000",
  40909=>"010110111",
  40910=>"111010010",
  40911=>"111001001",
  40912=>"110110101",
  40913=>"001101101",
  40914=>"110011100",
  40915=>"000101001",
  40916=>"000011101",
  40917=>"001111111",
  40918=>"011110110",
  40919=>"111101100",
  40920=>"011001011",
  40921=>"100010100",
  40922=>"001101011",
  40923=>"100001100",
  40924=>"101000010",
  40925=>"011011001",
  40926=>"101000000",
  40927=>"101011001",
  40928=>"001110101",
  40929=>"111100010",
  40930=>"010101000",
  40931=>"110110000",
  40932=>"110000010",
  40933=>"010101011",
  40934=>"110110000",
  40935=>"100111101",
  40936=>"101010101",
  40937=>"000000111",
  40938=>"100110100",
  40939=>"101001100",
  40940=>"001111010",
  40941=>"001000001",
  40942=>"110000010",
  40943=>"111011000",
  40944=>"110111101",
  40945=>"000000000",
  40946=>"101001100",
  40947=>"011100110",
  40948=>"000011101",
  40949=>"110000001",
  40950=>"000110000",
  40951=>"100101011",
  40952=>"101111100",
  40953=>"011000011",
  40954=>"110000101",
  40955=>"000100100",
  40956=>"001000011",
  40957=>"000011010",
  40958=>"010001010",
  40959=>"010101010",
  40960=>"111101110",
  40961=>"111001000",
  40962=>"010101111",
  40963=>"111101111",
  40964=>"110111110",
  40965=>"100010010",
  40966=>"111111111",
  40967=>"110001101",
  40968=>"010111010",
  40969=>"000110110",
  40970=>"110111001",
  40971=>"011101011",
  40972=>"111001100",
  40973=>"110110001",
  40974=>"111110100",
  40975=>"111010011",
  40976=>"101000100",
  40977=>"101000011",
  40978=>"111001000",
  40979=>"100001111",
  40980=>"011010100",
  40981=>"101110010",
  40982=>"001110111",
  40983=>"001111110",
  40984=>"110000000",
  40985=>"011110100",
  40986=>"001000100",
  40987=>"101101101",
  40988=>"000011010",
  40989=>"011110010",
  40990=>"111001101",
  40991=>"000000110",
  40992=>"100001111",
  40993=>"101000001",
  40994=>"100110101",
  40995=>"010111111",
  40996=>"101000110",
  40997=>"011010101",
  40998=>"100000101",
  40999=>"000010001",
  41000=>"010100111",
  41001=>"100110111",
  41002=>"011110110",
  41003=>"010000111",
  41004=>"100100111",
  41005=>"111010000",
  41006=>"100111010",
  41007=>"101100110",
  41008=>"010101111",
  41009=>"000010010",
  41010=>"000010011",
  41011=>"100010000",
  41012=>"101111110",
  41013=>"011001001",
  41014=>"100011101",
  41015=>"110011111",
  41016=>"000000001",
  41017=>"010000010",
  41018=>"000000011",
  41019=>"101100011",
  41020=>"001001100",
  41021=>"111000000",
  41022=>"000000101",
  41023=>"101111101",
  41024=>"010000101",
  41025=>"000101010",
  41026=>"010001101",
  41027=>"000010111",
  41028=>"100010111",
  41029=>"111100000",
  41030=>"000001010",
  41031=>"111000000",
  41032=>"110101100",
  41033=>"110110001",
  41034=>"100111100",
  41035=>"000000101",
  41036=>"011111110",
  41037=>"011110001",
  41038=>"001111100",
  41039=>"110000011",
  41040=>"101010101",
  41041=>"110101111",
  41042=>"001000111",
  41043=>"100111000",
  41044=>"101101011",
  41045=>"111001111",
  41046=>"000100001",
  41047=>"110000011",
  41048=>"110111011",
  41049=>"010101111",
  41050=>"101100101",
  41051=>"111000000",
  41052=>"010111001",
  41053=>"101001101",
  41054=>"110011101",
  41055=>"001100100",
  41056=>"011001100",
  41057=>"011011000",
  41058=>"001101110",
  41059=>"001110011",
  41060=>"101000100",
  41061=>"110010111",
  41062=>"111010101",
  41063=>"001101100",
  41064=>"001010000",
  41065=>"111100000",
  41066=>"100001001",
  41067=>"010111001",
  41068=>"011011000",
  41069=>"111100000",
  41070=>"101001101",
  41071=>"001011000",
  41072=>"111010010",
  41073=>"010111100",
  41074=>"000110110",
  41075=>"011010100",
  41076=>"001001100",
  41077=>"010001010",
  41078=>"110010001",
  41079=>"010101001",
  41080=>"111000101",
  41081=>"000100111",
  41082=>"001111101",
  41083=>"010010110",
  41084=>"001000111",
  41085=>"110111110",
  41086=>"000010100",
  41087=>"001110010",
  41088=>"101100010",
  41089=>"111100011",
  41090=>"111001100",
  41091=>"100100101",
  41092=>"011000010",
  41093=>"001000011",
  41094=>"011100101",
  41095=>"010011101",
  41096=>"010001010",
  41097=>"101000001",
  41098=>"001110010",
  41099=>"111111011",
  41100=>"101011001",
  41101=>"101000100",
  41102=>"000001000",
  41103=>"100000001",
  41104=>"111100111",
  41105=>"011010001",
  41106=>"101010010",
  41107=>"011000110",
  41108=>"101010010",
  41109=>"101010000",
  41110=>"001110010",
  41111=>"100000111",
  41112=>"011101010",
  41113=>"101000101",
  41114=>"100001000",
  41115=>"100000001",
  41116=>"111011010",
  41117=>"011010011",
  41118=>"000110001",
  41119=>"010101011",
  41120=>"001010011",
  41121=>"101011000",
  41122=>"100111100",
  41123=>"100001010",
  41124=>"011100111",
  41125=>"000111110",
  41126=>"100110000",
  41127=>"100110110",
  41128=>"101000111",
  41129=>"001111011",
  41130=>"000000101",
  41131=>"110111100",
  41132=>"101111111",
  41133=>"111001001",
  41134=>"110100101",
  41135=>"000000111",
  41136=>"000001000",
  41137=>"110111100",
  41138=>"110110110",
  41139=>"010101111",
  41140=>"110111000",
  41141=>"011010010",
  41142=>"011010111",
  41143=>"000101110",
  41144=>"100100000",
  41145=>"101110101",
  41146=>"110111101",
  41147=>"001110010",
  41148=>"011101111",
  41149=>"000100011",
  41150=>"000011011",
  41151=>"011011101",
  41152=>"101001100",
  41153=>"100011111",
  41154=>"011010100",
  41155=>"000010111",
  41156=>"111001010",
  41157=>"000100000",
  41158=>"010101110",
  41159=>"000001001",
  41160=>"110010010",
  41161=>"011100001",
  41162=>"110001001",
  41163=>"001100000",
  41164=>"011101010",
  41165=>"110000110",
  41166=>"001111111",
  41167=>"101000100",
  41168=>"110110001",
  41169=>"001101101",
  41170=>"010000111",
  41171=>"000100001",
  41172=>"001101000",
  41173=>"100010101",
  41174=>"000010010",
  41175=>"011011010",
  41176=>"011111100",
  41177=>"101000010",
  41178=>"101101111",
  41179=>"010000011",
  41180=>"010111100",
  41181=>"101010010",
  41182=>"101011000",
  41183=>"111100111",
  41184=>"000101000",
  41185=>"100101111",
  41186=>"101111101",
  41187=>"101101011",
  41188=>"101110010",
  41189=>"101011010",
  41190=>"111110011",
  41191=>"100100110",
  41192=>"100001111",
  41193=>"111011000",
  41194=>"001100111",
  41195=>"100110101",
  41196=>"111000110",
  41197=>"110010100",
  41198=>"000110110",
  41199=>"010000000",
  41200=>"111110010",
  41201=>"111011001",
  41202=>"011110101",
  41203=>"001110011",
  41204=>"110101001",
  41205=>"000101010",
  41206=>"110011010",
  41207=>"111010000",
  41208=>"011101110",
  41209=>"000111011",
  41210=>"100100101",
  41211=>"110010101",
  41212=>"001001100",
  41213=>"011101001",
  41214=>"011010000",
  41215=>"111100001",
  41216=>"100001001",
  41217=>"001111000",
  41218=>"100001110",
  41219=>"100001110",
  41220=>"010111010",
  41221=>"111111111",
  41222=>"111100001",
  41223=>"011010110",
  41224=>"011011100",
  41225=>"100001010",
  41226=>"000000101",
  41227=>"011010111",
  41228=>"110101111",
  41229=>"111101001",
  41230=>"001000000",
  41231=>"100111001",
  41232=>"000110000",
  41233=>"110010010",
  41234=>"001000111",
  41235=>"100000100",
  41236=>"101001110",
  41237=>"000100111",
  41238=>"100111100",
  41239=>"000101100",
  41240=>"010101110",
  41241=>"011111000",
  41242=>"111001001",
  41243=>"011001011",
  41244=>"001011011",
  41245=>"110101000",
  41246=>"010001000",
  41247=>"011100100",
  41248=>"000011010",
  41249=>"001001011",
  41250=>"001001000",
  41251=>"010011110",
  41252=>"111111101",
  41253=>"011011111",
  41254=>"000111110",
  41255=>"110100100",
  41256=>"000011000",
  41257=>"111100111",
  41258=>"111001011",
  41259=>"111010101",
  41260=>"000011110",
  41261=>"011001101",
  41262=>"001000101",
  41263=>"000000010",
  41264=>"111100100",
  41265=>"000011011",
  41266=>"110010000",
  41267=>"000010010",
  41268=>"110001110",
  41269=>"110001111",
  41270=>"101011001",
  41271=>"011000100",
  41272=>"100110101",
  41273=>"110001001",
  41274=>"010101010",
  41275=>"111001011",
  41276=>"110001100",
  41277=>"101100101",
  41278=>"111110110",
  41279=>"100011001",
  41280=>"000101010",
  41281=>"000100001",
  41282=>"101111110",
  41283=>"110101101",
  41284=>"001111011",
  41285=>"000001001",
  41286=>"101011001",
  41287=>"001011100",
  41288=>"011010100",
  41289=>"011001000",
  41290=>"111111110",
  41291=>"001010010",
  41292=>"111110101",
  41293=>"001010000",
  41294=>"111000110",
  41295=>"010001100",
  41296=>"010010100",
  41297=>"011001101",
  41298=>"000100010",
  41299=>"010010100",
  41300=>"111101100",
  41301=>"101111011",
  41302=>"110110001",
  41303=>"111101101",
  41304=>"100110011",
  41305=>"110001100",
  41306=>"110110101",
  41307=>"110000000",
  41308=>"111001000",
  41309=>"001101110",
  41310=>"011100010",
  41311=>"000010000",
  41312=>"101111001",
  41313=>"101101001",
  41314=>"100111010",
  41315=>"011001001",
  41316=>"101101101",
  41317=>"010100011",
  41318=>"010000111",
  41319=>"111011101",
  41320=>"000001000",
  41321=>"111011001",
  41322=>"100011111",
  41323=>"100100001",
  41324=>"011000101",
  41325=>"110010011",
  41326=>"111110001",
  41327=>"100110111",
  41328=>"111100011",
  41329=>"001000000",
  41330=>"111100110",
  41331=>"110110011",
  41332=>"110011110",
  41333=>"010001000",
  41334=>"010111101",
  41335=>"111000100",
  41336=>"100100011",
  41337=>"011001000",
  41338=>"111110100",
  41339=>"000011111",
  41340=>"111000001",
  41341=>"111001111",
  41342=>"111111101",
  41343=>"110101011",
  41344=>"010010011",
  41345=>"101010010",
  41346=>"100000001",
  41347=>"100010111",
  41348=>"010101101",
  41349=>"100101010",
  41350=>"000110101",
  41351=>"100100001",
  41352=>"011010110",
  41353=>"111010001",
  41354=>"100110001",
  41355=>"101010001",
  41356=>"000100101",
  41357=>"111110111",
  41358=>"001010000",
  41359=>"100111001",
  41360=>"000110001",
  41361=>"100001111",
  41362=>"111110100",
  41363=>"001001101",
  41364=>"101011100",
  41365=>"001100100",
  41366=>"010101000",
  41367=>"011101001",
  41368=>"000010010",
  41369=>"100100010",
  41370=>"110000010",
  41371=>"100110000",
  41372=>"011100010",
  41373=>"010011100",
  41374=>"101111010",
  41375=>"001010000",
  41376=>"000110111",
  41377=>"101100101",
  41378=>"101000100",
  41379=>"101010000",
  41380=>"000110101",
  41381=>"101101000",
  41382=>"011011011",
  41383=>"011111111",
  41384=>"010111111",
  41385=>"000100011",
  41386=>"010100110",
  41387=>"100111001",
  41388=>"101111111",
  41389=>"101101010",
  41390=>"000001110",
  41391=>"110010101",
  41392=>"010010101",
  41393=>"100001011",
  41394=>"001101100",
  41395=>"101100101",
  41396=>"100100001",
  41397=>"101100010",
  41398=>"001001100",
  41399=>"001011011",
  41400=>"000000001",
  41401=>"000101110",
  41402=>"110110000",
  41403=>"110111100",
  41404=>"011111000",
  41405=>"010000110",
  41406=>"000100110",
  41407=>"110111010",
  41408=>"000000100",
  41409=>"111111111",
  41410=>"000010110",
  41411=>"011111100",
  41412=>"001100000",
  41413=>"000101010",
  41414=>"110100110",
  41415=>"000001000",
  41416=>"010000111",
  41417=>"001001101",
  41418=>"010000101",
  41419=>"110110000",
  41420=>"110101110",
  41421=>"100000011",
  41422=>"111100010",
  41423=>"010100100",
  41424=>"111111000",
  41425=>"011011110",
  41426=>"011001100",
  41427=>"001111110",
  41428=>"110000101",
  41429=>"101110111",
  41430=>"011111100",
  41431=>"110010111",
  41432=>"011001110",
  41433=>"010101110",
  41434=>"010111011",
  41435=>"010111011",
  41436=>"011010010",
  41437=>"100010010",
  41438=>"111011000",
  41439=>"000101011",
  41440=>"101100001",
  41441=>"110101001",
  41442=>"110011000",
  41443=>"110100100",
  41444=>"110000100",
  41445=>"101000000",
  41446=>"001101100",
  41447=>"111001110",
  41448=>"011101010",
  41449=>"000111110",
  41450=>"001101000",
  41451=>"001000010",
  41452=>"011010011",
  41453=>"000100010",
  41454=>"000011111",
  41455=>"001100100",
  41456=>"111001110",
  41457=>"101001000",
  41458=>"100000101",
  41459=>"111101011",
  41460=>"101100111",
  41461=>"001010100",
  41462=>"101000011",
  41463=>"110110001",
  41464=>"000110100",
  41465=>"111101110",
  41466=>"000100111",
  41467=>"100011011",
  41468=>"101001110",
  41469=>"100000000",
  41470=>"000010010",
  41471=>"001101000",
  41472=>"000101110",
  41473=>"010111010",
  41474=>"101100000",
  41475=>"011011001",
  41476=>"000010011",
  41477=>"100001010",
  41478=>"000000111",
  41479=>"000001101",
  41480=>"010011101",
  41481=>"101111010",
  41482=>"001000110",
  41483=>"111110010",
  41484=>"110100001",
  41485=>"001010000",
  41486=>"011100001",
  41487=>"101001110",
  41488=>"010000111",
  41489=>"101001101",
  41490=>"101101111",
  41491=>"001010111",
  41492=>"100100101",
  41493=>"111010011",
  41494=>"100101010",
  41495=>"101010000",
  41496=>"110010000",
  41497=>"001010001",
  41498=>"011101101",
  41499=>"110110011",
  41500=>"011110100",
  41501=>"111010111",
  41502=>"100111000",
  41503=>"000010000",
  41504=>"010000110",
  41505=>"011111101",
  41506=>"000111001",
  41507=>"001110111",
  41508=>"111010010",
  41509=>"001110111",
  41510=>"001100001",
  41511=>"011110110",
  41512=>"001000100",
  41513=>"101101000",
  41514=>"101000000",
  41515=>"101101101",
  41516=>"001011001",
  41517=>"110011111",
  41518=>"001001000",
  41519=>"011010110",
  41520=>"010110001",
  41521=>"101001010",
  41522=>"010001000",
  41523=>"011001110",
  41524=>"000100101",
  41525=>"100100110",
  41526=>"100000110",
  41527=>"000100100",
  41528=>"001000010",
  41529=>"101100000",
  41530=>"011100101",
  41531=>"000101001",
  41532=>"010100100",
  41533=>"000010101",
  41534=>"001011000",
  41535=>"101110001",
  41536=>"100111111",
  41537=>"110101101",
  41538=>"001100000",
  41539=>"101110111",
  41540=>"001001011",
  41541=>"001110101",
  41542=>"111111101",
  41543=>"100101101",
  41544=>"010001101",
  41545=>"011101000",
  41546=>"000001101",
  41547=>"011001101",
  41548=>"000111010",
  41549=>"100111111",
  41550=>"010100000",
  41551=>"011101000",
  41552=>"001011110",
  41553=>"000000010",
  41554=>"001101001",
  41555=>"101011111",
  41556=>"001011110",
  41557=>"001100101",
  41558=>"010011010",
  41559=>"110011011",
  41560=>"000000001",
  41561=>"011001100",
  41562=>"100011011",
  41563=>"000100011",
  41564=>"000001101",
  41565=>"110000110",
  41566=>"010010001",
  41567=>"111101000",
  41568=>"100110111",
  41569=>"111111101",
  41570=>"000101101",
  41571=>"000100001",
  41572=>"001010100",
  41573=>"000101000",
  41574=>"011000000",
  41575=>"000101110",
  41576=>"111000011",
  41577=>"000000000",
  41578=>"001101100",
  41579=>"111011111",
  41580=>"000100110",
  41581=>"111011101",
  41582=>"001111000",
  41583=>"111001111",
  41584=>"110010100",
  41585=>"111010000",
  41586=>"110111110",
  41587=>"110111111",
  41588=>"011111000",
  41589=>"000000000",
  41590=>"011111011",
  41591=>"001000110",
  41592=>"110011100",
  41593=>"101111111",
  41594=>"001001110",
  41595=>"000001001",
  41596=>"010000001",
  41597=>"100111000",
  41598=>"001100101",
  41599=>"011001010",
  41600=>"101001100",
  41601=>"000011001",
  41602=>"010100010",
  41603=>"100010000",
  41604=>"001111101",
  41605=>"011011000",
  41606=>"010110110",
  41607=>"000111111",
  41608=>"000001011",
  41609=>"011001010",
  41610=>"110111001",
  41611=>"010001010",
  41612=>"001000011",
  41613=>"000010101",
  41614=>"111011110",
  41615=>"000000001",
  41616=>"110010000",
  41617=>"110000000",
  41618=>"110100110",
  41619=>"011100010",
  41620=>"101100001",
  41621=>"001001011",
  41622=>"110101010",
  41623=>"001010000",
  41624=>"111100010",
  41625=>"000010010",
  41626=>"000000010",
  41627=>"001101010",
  41628=>"010101110",
  41629=>"110010001",
  41630=>"111101111",
  41631=>"111110111",
  41632=>"000001011",
  41633=>"010101001",
  41634=>"000011111",
  41635=>"010110111",
  41636=>"101101101",
  41637=>"110001000",
  41638=>"001001001",
  41639=>"110110101",
  41640=>"111100000",
  41641=>"110100111",
  41642=>"001011000",
  41643=>"111011011",
  41644=>"111011000",
  41645=>"110111110",
  41646=>"001111111",
  41647=>"000100111",
  41648=>"001101110",
  41649=>"001010000",
  41650=>"111011111",
  41651=>"110001011",
  41652=>"010010001",
  41653=>"000000110",
  41654=>"100011101",
  41655=>"111010010",
  41656=>"100101010",
  41657=>"001111101",
  41658=>"010111110",
  41659=>"001111010",
  41660=>"111100110",
  41661=>"111100101",
  41662=>"010001011",
  41663=>"010111110",
  41664=>"100111011",
  41665=>"001000001",
  41666=>"010110101",
  41667=>"010001001",
  41668=>"000010010",
  41669=>"100001010",
  41670=>"111100111",
  41671=>"000011101",
  41672=>"000001000",
  41673=>"110000111",
  41674=>"111001011",
  41675=>"111000101",
  41676=>"010111010",
  41677=>"011110011",
  41678=>"111110000",
  41679=>"101011010",
  41680=>"001000000",
  41681=>"000100010",
  41682=>"100000101",
  41683=>"011000111",
  41684=>"010111110",
  41685=>"111000000",
  41686=>"101111001",
  41687=>"110011111",
  41688=>"000010011",
  41689=>"100110000",
  41690=>"000010100",
  41691=>"011001101",
  41692=>"110000010",
  41693=>"100100000",
  41694=>"101110000",
  41695=>"111000111",
  41696=>"101111110",
  41697=>"101011101",
  41698=>"011110101",
  41699=>"110000110",
  41700=>"010001100",
  41701=>"101101011",
  41702=>"111011111",
  41703=>"000100010",
  41704=>"101011011",
  41705=>"100010001",
  41706=>"111111010",
  41707=>"110111010",
  41708=>"110111000",
  41709=>"101111011",
  41710=>"010100101",
  41711=>"000010010",
  41712=>"010110100",
  41713=>"101001100",
  41714=>"111000010",
  41715=>"011111100",
  41716=>"010001000",
  41717=>"100010101",
  41718=>"000010000",
  41719=>"100000001",
  41720=>"111111100",
  41721=>"101100001",
  41722=>"111101010",
  41723=>"101000111",
  41724=>"010110011",
  41725=>"111110001",
  41726=>"100101111",
  41727=>"101011010",
  41728=>"111011001",
  41729=>"100010011",
  41730=>"100101111",
  41731=>"000100101",
  41732=>"011001111",
  41733=>"001100010",
  41734=>"011100000",
  41735=>"001000011",
  41736=>"100100000",
  41737=>"010010010",
  41738=>"101001110",
  41739=>"011100000",
  41740=>"011010100",
  41741=>"110000000",
  41742=>"100010111",
  41743=>"110000010",
  41744=>"110111110",
  41745=>"001110001",
  41746=>"101000001",
  41747=>"100110111",
  41748=>"111111111",
  41749=>"111001011",
  41750=>"000001010",
  41751=>"111000100",
  41752=>"001001101",
  41753=>"101011111",
  41754=>"100010000",
  41755=>"100010111",
  41756=>"110000101",
  41757=>"011110000",
  41758=>"010011010",
  41759=>"001001011",
  41760=>"000001001",
  41761=>"000101111",
  41762=>"000111111",
  41763=>"011101101",
  41764=>"111110101",
  41765=>"000001000",
  41766=>"000110000",
  41767=>"101101111",
  41768=>"111001000",
  41769=>"011010110",
  41770=>"010111101",
  41771=>"001111101",
  41772=>"000110000",
  41773=>"001001111",
  41774=>"001001001",
  41775=>"110000001",
  41776=>"110100011",
  41777=>"100000000",
  41778=>"100000001",
  41779=>"100110101",
  41780=>"110110110",
  41781=>"011010100",
  41782=>"111101111",
  41783=>"101001111",
  41784=>"000110010",
  41785=>"000001110",
  41786=>"110001110",
  41787=>"101010001",
  41788=>"011010101",
  41789=>"101110111",
  41790=>"001000000",
  41791=>"000011000",
  41792=>"001001000",
  41793=>"010001011",
  41794=>"001110001",
  41795=>"110101111",
  41796=>"000110000",
  41797=>"000001011",
  41798=>"011010000",
  41799=>"001111011",
  41800=>"010000111",
  41801=>"011110000",
  41802=>"111001010",
  41803=>"010111100",
  41804=>"001011011",
  41805=>"110000111",
  41806=>"100000010",
  41807=>"011000011",
  41808=>"100110001",
  41809=>"101011101",
  41810=>"001001110",
  41811=>"000100010",
  41812=>"100111111",
  41813=>"101100011",
  41814=>"011110110",
  41815=>"001001100",
  41816=>"100110111",
  41817=>"111100110",
  41818=>"001100111",
  41819=>"111011001",
  41820=>"110011000",
  41821=>"111110111",
  41822=>"111100011",
  41823=>"010100001",
  41824=>"000011101",
  41825=>"001111011",
  41826=>"011011110",
  41827=>"100101000",
  41828=>"101000100",
  41829=>"100110000",
  41830=>"011001100",
  41831=>"000101100",
  41832=>"111101000",
  41833=>"100110101",
  41834=>"001101001",
  41835=>"111011110",
  41836=>"000111000",
  41837=>"110001110",
  41838=>"110110000",
  41839=>"011011101",
  41840=>"011001110",
  41841=>"010000000",
  41842=>"100100011",
  41843=>"000010010",
  41844=>"000111100",
  41845=>"110101001",
  41846=>"010001011",
  41847=>"010111100",
  41848=>"011100100",
  41849=>"001110011",
  41850=>"000100100",
  41851=>"001110001",
  41852=>"111110101",
  41853=>"100000001",
  41854=>"011011110",
  41855=>"011101101",
  41856=>"111110101",
  41857=>"001000010",
  41858=>"000011010",
  41859=>"101101011",
  41860=>"001011010",
  41861=>"110011001",
  41862=>"010010101",
  41863=>"000000100",
  41864=>"110001001",
  41865=>"110011010",
  41866=>"001100100",
  41867=>"001000001",
  41868=>"001000011",
  41869=>"111011101",
  41870=>"000101111",
  41871=>"100010001",
  41872=>"111101100",
  41873=>"001001000",
  41874=>"000101010",
  41875=>"101100010",
  41876=>"001011010",
  41877=>"000101100",
  41878=>"000111000",
  41879=>"000001000",
  41880=>"100100010",
  41881=>"000011111",
  41882=>"001111010",
  41883=>"100011101",
  41884=>"111010101",
  41885=>"101000011",
  41886=>"101111000",
  41887=>"000100000",
  41888=>"001111101",
  41889=>"101111111",
  41890=>"010111000",
  41891=>"110101111",
  41892=>"111100100",
  41893=>"001001011",
  41894=>"101111011",
  41895=>"000001011",
  41896=>"001000010",
  41897=>"010010010",
  41898=>"101010110",
  41899=>"101000001",
  41900=>"000000001",
  41901=>"001111100",
  41902=>"110100011",
  41903=>"111010100",
  41904=>"101101010",
  41905=>"101010011",
  41906=>"011100010",
  41907=>"101011110",
  41908=>"010111000",
  41909=>"001001000",
  41910=>"011100000",
  41911=>"001111100",
  41912=>"111111100",
  41913=>"111100111",
  41914=>"101100010",
  41915=>"011000110",
  41916=>"000101100",
  41917=>"111011010",
  41918=>"000001101",
  41919=>"001111011",
  41920=>"100100110",
  41921=>"011001001",
  41922=>"000011101",
  41923=>"001100000",
  41924=>"111101011",
  41925=>"110110101",
  41926=>"010001001",
  41927=>"011100100",
  41928=>"110011001",
  41929=>"101111110",
  41930=>"010100101",
  41931=>"010001001",
  41932=>"010011011",
  41933=>"000010111",
  41934=>"101010000",
  41935=>"001101101",
  41936=>"111111001",
  41937=>"111110011",
  41938=>"101000010",
  41939=>"011110001",
  41940=>"010101100",
  41941=>"110001110",
  41942=>"011010111",
  41943=>"011010010",
  41944=>"100011100",
  41945=>"011111001",
  41946=>"000000101",
  41947=>"101000011",
  41948=>"100001111",
  41949=>"000000111",
  41950=>"101100000",
  41951=>"001001000",
  41952=>"000011001",
  41953=>"010000100",
  41954=>"101010101",
  41955=>"100010000",
  41956=>"100110011",
  41957=>"011110110",
  41958=>"100001111",
  41959=>"101010111",
  41960=>"101000000",
  41961=>"101000011",
  41962=>"000101001",
  41963=>"110010001",
  41964=>"111111111",
  41965=>"010001110",
  41966=>"000110100",
  41967=>"010000101",
  41968=>"011101101",
  41969=>"000011100",
  41970=>"101001010",
  41971=>"100000100",
  41972=>"010101000",
  41973=>"110010010",
  41974=>"101111000",
  41975=>"000010111",
  41976=>"010110000",
  41977=>"110111110",
  41978=>"111110001",
  41979=>"101000010",
  41980=>"100011011",
  41981=>"100011001",
  41982=>"010000011",
  41983=>"111011111",
  41984=>"110011000",
  41985=>"001101010",
  41986=>"010000111",
  41987=>"000110011",
  41988=>"101001001",
  41989=>"101011001",
  41990=>"011000001",
  41991=>"001001100",
  41992=>"110010011",
  41993=>"100111110",
  41994=>"110010001",
  41995=>"010010101",
  41996=>"100100100",
  41997=>"110100010",
  41998=>"000000111",
  41999=>"101000000",
  42000=>"101101000",
  42001=>"000110110",
  42002=>"110101111",
  42003=>"110000101",
  42004=>"001011100",
  42005=>"100001011",
  42006=>"100100001",
  42007=>"101001001",
  42008=>"010111111",
  42009=>"101000010",
  42010=>"110010100",
  42011=>"100110101",
  42012=>"101111010",
  42013=>"110101001",
  42014=>"100101110",
  42015=>"110100010",
  42016=>"001010000",
  42017=>"011100001",
  42018=>"101101011",
  42019=>"011100011",
  42020=>"101000001",
  42021=>"111001111",
  42022=>"010100001",
  42023=>"100100101",
  42024=>"000110100",
  42025=>"111001000",
  42026=>"000011011",
  42027=>"101110100",
  42028=>"100011001",
  42029=>"100101001",
  42030=>"010111000",
  42031=>"111101001",
  42032=>"101100000",
  42033=>"101111110",
  42034=>"101100111",
  42035=>"011110110",
  42036=>"011001001",
  42037=>"000100110",
  42038=>"100000000",
  42039=>"001101110",
  42040=>"010001101",
  42041=>"111011100",
  42042=>"001011001",
  42043=>"100110111",
  42044=>"101101010",
  42045=>"001100011",
  42046=>"110100000",
  42047=>"000010111",
  42048=>"100000110",
  42049=>"001101010",
  42050=>"101111111",
  42051=>"010100011",
  42052=>"111011111",
  42053=>"111001111",
  42054=>"111110110",
  42055=>"011011110",
  42056=>"011100110",
  42057=>"000000111",
  42058=>"000010011",
  42059=>"101110111",
  42060=>"100011111",
  42061=>"111101011",
  42062=>"011001000",
  42063=>"011010111",
  42064=>"001000110",
  42065=>"110101010",
  42066=>"010101111",
  42067=>"100010000",
  42068=>"000100011",
  42069=>"100100011",
  42070=>"000110000",
  42071=>"000100100",
  42072=>"110000001",
  42073=>"110010011",
  42074=>"101100101",
  42075=>"010111010",
  42076=>"100000000",
  42077=>"111100101",
  42078=>"100000101",
  42079=>"011010100",
  42080=>"100010010",
  42081=>"011111000",
  42082=>"111011001",
  42083=>"010010110",
  42084=>"111000110",
  42085=>"110001010",
  42086=>"111110110",
  42087=>"110100110",
  42088=>"011011011",
  42089=>"011110001",
  42090=>"011111100",
  42091=>"101001110",
  42092=>"101111000",
  42093=>"001001010",
  42094=>"111110111",
  42095=>"010101001",
  42096=>"001000000",
  42097=>"100000011",
  42098=>"011110001",
  42099=>"000110100",
  42100=>"111001110",
  42101=>"111111010",
  42102=>"000010110",
  42103=>"111100010",
  42104=>"001001010",
  42105=>"110001101",
  42106=>"000000011",
  42107=>"000101111",
  42108=>"010000100",
  42109=>"001101000",
  42110=>"111101010",
  42111=>"101100011",
  42112=>"000110010",
  42113=>"000011111",
  42114=>"111111000",
  42115=>"000110110",
  42116=>"110000000",
  42117=>"001111110",
  42118=>"011100110",
  42119=>"001111101",
  42120=>"000101001",
  42121=>"110000011",
  42122=>"111111111",
  42123=>"101111100",
  42124=>"110010001",
  42125=>"000010110",
  42126=>"001000010",
  42127=>"011000100",
  42128=>"010100110",
  42129=>"101000000",
  42130=>"110110111",
  42131=>"110001010",
  42132=>"000100010",
  42133=>"111000110",
  42134=>"000110110",
  42135=>"010111000",
  42136=>"011001111",
  42137=>"011110101",
  42138=>"110000011",
  42139=>"100101110",
  42140=>"010001000",
  42141=>"100000100",
  42142=>"000010011",
  42143=>"010101100",
  42144=>"001101001",
  42145=>"001101011",
  42146=>"101110100",
  42147=>"101010100",
  42148=>"101011110",
  42149=>"101101111",
  42150=>"111101000",
  42151=>"010101000",
  42152=>"000001000",
  42153=>"000100010",
  42154=>"101111010",
  42155=>"111110101",
  42156=>"001100010",
  42157=>"111000100",
  42158=>"101100010",
  42159=>"110001101",
  42160=>"101110111",
  42161=>"010001101",
  42162=>"111001001",
  42163=>"111111010",
  42164=>"010010011",
  42165=>"101111110",
  42166=>"000100010",
  42167=>"111110010",
  42168=>"011111101",
  42169=>"011101011",
  42170=>"001010011",
  42171=>"111100111",
  42172=>"011001111",
  42173=>"101110010",
  42174=>"000111011",
  42175=>"011101100",
  42176=>"110100010",
  42177=>"110000001",
  42178=>"100110000",
  42179=>"000010001",
  42180=>"010100011",
  42181=>"111001101",
  42182=>"000010100",
  42183=>"011101101",
  42184=>"101010001",
  42185=>"000100111",
  42186=>"001101001",
  42187=>"010010000",
  42188=>"001000110",
  42189=>"110101110",
  42190=>"000000010",
  42191=>"110011011",
  42192=>"001101001",
  42193=>"110101001",
  42194=>"001011110",
  42195=>"000000101",
  42196=>"001010000",
  42197=>"111111101",
  42198=>"011001000",
  42199=>"100001010",
  42200=>"101010110",
  42201=>"100010010",
  42202=>"000000111",
  42203=>"010000011",
  42204=>"100100001",
  42205=>"011000000",
  42206=>"001001000",
  42207=>"011010000",
  42208=>"111101011",
  42209=>"110101111",
  42210=>"001100110",
  42211=>"001010011",
  42212=>"000110100",
  42213=>"101110001",
  42214=>"101100011",
  42215=>"111011011",
  42216=>"111111100",
  42217=>"111001001",
  42218=>"010000100",
  42219=>"100011110",
  42220=>"111010011",
  42221=>"101100110",
  42222=>"110000000",
  42223=>"011101100",
  42224=>"100100001",
  42225=>"011100011",
  42226=>"000100111",
  42227=>"100000011",
  42228=>"100111010",
  42229=>"110110111",
  42230=>"100101100",
  42231=>"000000011",
  42232=>"010110101",
  42233=>"111011001",
  42234=>"111110110",
  42235=>"001101010",
  42236=>"000001100",
  42237=>"011100110",
  42238=>"110010101",
  42239=>"011101001",
  42240=>"010110010",
  42241=>"110101001",
  42242=>"100011111",
  42243=>"110111101",
  42244=>"010111010",
  42245=>"011100110",
  42246=>"111000000",
  42247=>"000011111",
  42248=>"110010011",
  42249=>"010001010",
  42250=>"110001000",
  42251=>"000111011",
  42252=>"010101111",
  42253=>"111000010",
  42254=>"011100111",
  42255=>"011001011",
  42256=>"110110001",
  42257=>"100010000",
  42258=>"010000100",
  42259=>"010010001",
  42260=>"011000100",
  42261=>"100100001",
  42262=>"011010001",
  42263=>"110001010",
  42264=>"101111010",
  42265=>"011011000",
  42266=>"011000111",
  42267=>"010100000",
  42268=>"110000100",
  42269=>"111100111",
  42270=>"000100011",
  42271=>"000001100",
  42272=>"001010111",
  42273=>"100000101",
  42274=>"000101001",
  42275=>"110110001",
  42276=>"010010000",
  42277=>"101000101",
  42278=>"101001101",
  42279=>"011101001",
  42280=>"110000111",
  42281=>"110101011",
  42282=>"100111000",
  42283=>"011111010",
  42284=>"111111101",
  42285=>"001000101",
  42286=>"000010111",
  42287=>"111000000",
  42288=>"110001110",
  42289=>"001110000",
  42290=>"001101100",
  42291=>"110100010",
  42292=>"000111001",
  42293=>"111110011",
  42294=>"010111101",
  42295=>"111010001",
  42296=>"000101111",
  42297=>"001110101",
  42298=>"010011111",
  42299=>"101000001",
  42300=>"111010000",
  42301=>"000010001",
  42302=>"110101010",
  42303=>"010100100",
  42304=>"001010111",
  42305=>"101101000",
  42306=>"110111011",
  42307=>"010111000",
  42308=>"010010010",
  42309=>"010010111",
  42310=>"011100010",
  42311=>"101010000",
  42312=>"001111100",
  42313=>"101101101",
  42314=>"001001001",
  42315=>"011000010",
  42316=>"110001000",
  42317=>"101101011",
  42318=>"000110110",
  42319=>"011000011",
  42320=>"010000101",
  42321=>"001011000",
  42322=>"000001000",
  42323=>"110111010",
  42324=>"000111000",
  42325=>"101011001",
  42326=>"011111101",
  42327=>"000111011",
  42328=>"101010000",
  42329=>"000100011",
  42330=>"010100010",
  42331=>"011111101",
  42332=>"101000001",
  42333=>"111011011",
  42334=>"111111111",
  42335=>"101100001",
  42336=>"011100000",
  42337=>"011011100",
  42338=>"011000000",
  42339=>"110000010",
  42340=>"101101111",
  42341=>"111000000",
  42342=>"010110010",
  42343=>"101111100",
  42344=>"111100111",
  42345=>"110101010",
  42346=>"100110001",
  42347=>"000011001",
  42348=>"110000100",
  42349=>"000110010",
  42350=>"101001010",
  42351=>"010100001",
  42352=>"101110100",
  42353=>"010000111",
  42354=>"111110001",
  42355=>"110100110",
  42356=>"111010001",
  42357=>"111101010",
  42358=>"000010000",
  42359=>"100101101",
  42360=>"100000011",
  42361=>"101011011",
  42362=>"000110010",
  42363=>"111010100",
  42364=>"100011110",
  42365=>"001101001",
  42366=>"100011101",
  42367=>"101001111",
  42368=>"001010011",
  42369=>"010101100",
  42370=>"101001110",
  42371=>"000010111",
  42372=>"010011101",
  42373=>"000111010",
  42374=>"011101110",
  42375=>"001111100",
  42376=>"000001100",
  42377=>"111100001",
  42378=>"000101111",
  42379=>"011101110",
  42380=>"011101101",
  42381=>"110000010",
  42382=>"111010110",
  42383=>"000111010",
  42384=>"100111101",
  42385=>"110000100",
  42386=>"101011000",
  42387=>"100000011",
  42388=>"010111110",
  42389=>"100100101",
  42390=>"010110010",
  42391=>"010011010",
  42392=>"110001000",
  42393=>"101110111",
  42394=>"010100100",
  42395=>"100001000",
  42396=>"110111011",
  42397=>"000110001",
  42398=>"100011110",
  42399=>"000110000",
  42400=>"111100001",
  42401=>"100100100",
  42402=>"010001100",
  42403=>"001000111",
  42404=>"001010000",
  42405=>"100000001",
  42406=>"000001101",
  42407=>"111011011",
  42408=>"110010111",
  42409=>"000011010",
  42410=>"111100011",
  42411=>"001001000",
  42412=>"110001001",
  42413=>"011011000",
  42414=>"111100000",
  42415=>"100000010",
  42416=>"001101100",
  42417=>"011000010",
  42418=>"011001110",
  42419=>"000100100",
  42420=>"010001001",
  42421=>"101110100",
  42422=>"001101110",
  42423=>"000110100",
  42424=>"001010111",
  42425=>"000011001",
  42426=>"001000101",
  42427=>"101000010",
  42428=>"111100011",
  42429=>"100111011",
  42430=>"010000001",
  42431=>"011011000",
  42432=>"010000011",
  42433=>"011100010",
  42434=>"011001001",
  42435=>"111010001",
  42436=>"010010111",
  42437=>"110001001",
  42438=>"000101001",
  42439=>"001011110",
  42440=>"110011101",
  42441=>"000001101",
  42442=>"110111110",
  42443=>"000001001",
  42444=>"011001100",
  42445=>"001010000",
  42446=>"110011011",
  42447=>"000001110",
  42448=>"100001110",
  42449=>"010001010",
  42450=>"000110110",
  42451=>"101111000",
  42452=>"111110101",
  42453=>"111111100",
  42454=>"101100010",
  42455=>"010000000",
  42456=>"000011110",
  42457=>"001010000",
  42458=>"100001111",
  42459=>"111100101",
  42460=>"111001011",
  42461=>"001110110",
  42462=>"101001011",
  42463=>"011011110",
  42464=>"110011011",
  42465=>"001000100",
  42466=>"000101111",
  42467=>"101111101",
  42468=>"000011011",
  42469=>"001000101",
  42470=>"000110000",
  42471=>"111001001",
  42472=>"001111101",
  42473=>"111111101",
  42474=>"010010100",
  42475=>"111000111",
  42476=>"111110000",
  42477=>"010100010",
  42478=>"011001011",
  42479=>"011110001",
  42480=>"100110000",
  42481=>"101111110",
  42482=>"001001111",
  42483=>"001000001",
  42484=>"000001000",
  42485=>"111011001",
  42486=>"110101100",
  42487=>"100110101",
  42488=>"110010010",
  42489=>"100001111",
  42490=>"100101110",
  42491=>"110001110",
  42492=>"101110001",
  42493=>"101110000",
  42494=>"110011000",
  42495=>"011111011",
  42496=>"110010011",
  42497=>"001011011",
  42498=>"001001000",
  42499=>"110100110",
  42500=>"011111101",
  42501=>"101011110",
  42502=>"111111000",
  42503=>"101101100",
  42504=>"011000101",
  42505=>"100110011",
  42506=>"000110111",
  42507=>"001111000",
  42508=>"001110010",
  42509=>"010100010",
  42510=>"101001011",
  42511=>"001001001",
  42512=>"100100010",
  42513=>"010000011",
  42514=>"100001001",
  42515=>"001111110",
  42516=>"110001000",
  42517=>"110110000",
  42518=>"010110101",
  42519=>"101110100",
  42520=>"101000111",
  42521=>"110011011",
  42522=>"010100100",
  42523=>"100010101",
  42524=>"000000000",
  42525=>"000101100",
  42526=>"110010111",
  42527=>"100010110",
  42528=>"100000001",
  42529=>"110111011",
  42530=>"100011000",
  42531=>"000000101",
  42532=>"001001010",
  42533=>"000101110",
  42534=>"011110100",
  42535=>"000011010",
  42536=>"001101100",
  42537=>"101011100",
  42538=>"011001101",
  42539=>"010110101",
  42540=>"010100010",
  42541=>"011110010",
  42542=>"001110111",
  42543=>"011001010",
  42544=>"111110001",
  42545=>"001110001",
  42546=>"000110110",
  42547=>"011001000",
  42548=>"000011000",
  42549=>"011001001",
  42550=>"010110001",
  42551=>"011110001",
  42552=>"000111010",
  42553=>"000111111",
  42554=>"001111100",
  42555=>"100111100",
  42556=>"100100101",
  42557=>"001001000",
  42558=>"000101011",
  42559=>"111010000",
  42560=>"111111000",
  42561=>"100111001",
  42562=>"011100111",
  42563=>"011111101",
  42564=>"001000110",
  42565=>"101010010",
  42566=>"000010101",
  42567=>"101100110",
  42568=>"010000111",
  42569=>"010101011",
  42570=>"011101110",
  42571=>"001011001",
  42572=>"100100000",
  42573=>"100001000",
  42574=>"000000000",
  42575=>"110111010",
  42576=>"010110101",
  42577=>"000100111",
  42578=>"010110001",
  42579=>"101001000",
  42580=>"111100101",
  42581=>"010110011",
  42582=>"011010110",
  42583=>"001000111",
  42584=>"100011001",
  42585=>"110010110",
  42586=>"010010110",
  42587=>"010011010",
  42588=>"000000011",
  42589=>"101010010",
  42590=>"110001011",
  42591=>"110001100",
  42592=>"111110111",
  42593=>"101011001",
  42594=>"100000000",
  42595=>"001110111",
  42596=>"101101101",
  42597=>"001010100",
  42598=>"111001111",
  42599=>"010001101",
  42600=>"111101111",
  42601=>"100001100",
  42602=>"101100001",
  42603=>"101010111",
  42604=>"000000001",
  42605=>"001010000",
  42606=>"001001101",
  42607=>"000011111",
  42608=>"100100011",
  42609=>"110001100",
  42610=>"000010001",
  42611=>"011010001",
  42612=>"010010111",
  42613=>"100111110",
  42614=>"001000101",
  42615=>"010110001",
  42616=>"110001001",
  42617=>"100000001",
  42618=>"100111110",
  42619=>"111101010",
  42620=>"110110101",
  42621=>"000011000",
  42622=>"100000111",
  42623=>"000010111",
  42624=>"000011111",
  42625=>"110101011",
  42626=>"000101111",
  42627=>"000001010",
  42628=>"011111110",
  42629=>"010000111",
  42630=>"111010001",
  42631=>"000010000",
  42632=>"000011100",
  42633=>"001011110",
  42634=>"101100011",
  42635=>"100100100",
  42636=>"010000001",
  42637=>"001100010",
  42638=>"000100100",
  42639=>"010100110",
  42640=>"101101110",
  42641=>"101001000",
  42642=>"100110000",
  42643=>"010010111",
  42644=>"101101110",
  42645=>"001110011",
  42646=>"010101101",
  42647=>"000100101",
  42648=>"011101000",
  42649=>"111010111",
  42650=>"000110101",
  42651=>"001100001",
  42652=>"101011101",
  42653=>"000111010",
  42654=>"011111000",
  42655=>"110111001",
  42656=>"110001000",
  42657=>"000011000",
  42658=>"111011111",
  42659=>"011011000",
  42660=>"010100111",
  42661=>"011011001",
  42662=>"010101110",
  42663=>"110100101",
  42664=>"101001010",
  42665=>"001000001",
  42666=>"100000100",
  42667=>"011010100",
  42668=>"010101001",
  42669=>"100010001",
  42670=>"101011111",
  42671=>"101011101",
  42672=>"011001011",
  42673=>"001111111",
  42674=>"110011000",
  42675=>"111000100",
  42676=>"100010000",
  42677=>"100010011",
  42678=>"110000100",
  42679=>"100010001",
  42680=>"100100101",
  42681=>"110110100",
  42682=>"111010100",
  42683=>"110001001",
  42684=>"000110010",
  42685=>"000100110",
  42686=>"001000111",
  42687=>"011001101",
  42688=>"100111010",
  42689=>"001101111",
  42690=>"000110100",
  42691=>"100001001",
  42692=>"100011100",
  42693=>"001100000",
  42694=>"000101111",
  42695=>"110010110",
  42696=>"010100000",
  42697=>"101101011",
  42698=>"111110110",
  42699=>"001011111",
  42700=>"111111010",
  42701=>"010000101",
  42702=>"000000011",
  42703=>"111011000",
  42704=>"001100100",
  42705=>"100100111",
  42706=>"111100011",
  42707=>"111000111",
  42708=>"110100110",
  42709=>"011111010",
  42710=>"111011111",
  42711=>"010101110",
  42712=>"110011011",
  42713=>"111101101",
  42714=>"000011100",
  42715=>"001111011",
  42716=>"101111111",
  42717=>"000101000",
  42718=>"100001000",
  42719=>"100000010",
  42720=>"000001000",
  42721=>"000000001",
  42722=>"111001101",
  42723=>"110110011",
  42724=>"111100100",
  42725=>"000110010",
  42726=>"001101001",
  42727=>"111000011",
  42728=>"000111000",
  42729=>"111110100",
  42730=>"111000010",
  42731=>"010100110",
  42732=>"101110100",
  42733=>"100010101",
  42734=>"000100101",
  42735=>"001111011",
  42736=>"101110001",
  42737=>"001000011",
  42738=>"010111100",
  42739=>"100010000",
  42740=>"000111111",
  42741=>"001100000",
  42742=>"111000010",
  42743=>"010111010",
  42744=>"110100111",
  42745=>"010110111",
  42746=>"010010100",
  42747=>"000101111",
  42748=>"011011010",
  42749=>"011111000",
  42750=>"010001011",
  42751=>"011000000",
  42752=>"110001010",
  42753=>"000000110",
  42754=>"010100000",
  42755=>"111101111",
  42756=>"010111011",
  42757=>"010000110",
  42758=>"101010111",
  42759=>"001111000",
  42760=>"100110000",
  42761=>"111111010",
  42762=>"011110111",
  42763=>"010111000",
  42764=>"011110100",
  42765=>"011000100",
  42766=>"111101101",
  42767=>"110011101",
  42768=>"011001101",
  42769=>"001101100",
  42770=>"001010001",
  42771=>"111001001",
  42772=>"000010001",
  42773=>"111001101",
  42774=>"110011000",
  42775=>"010100000",
  42776=>"000100101",
  42777=>"100111101",
  42778=>"000001110",
  42779=>"000010110",
  42780=>"101011001",
  42781=>"011101010",
  42782=>"001001010",
  42783=>"100010100",
  42784=>"001100101",
  42785=>"001001011",
  42786=>"010110100",
  42787=>"000101000",
  42788=>"111110001",
  42789=>"010110101",
  42790=>"000000111",
  42791=>"000100000",
  42792=>"111010001",
  42793=>"110110101",
  42794=>"110001000",
  42795=>"010101000",
  42796=>"101110010",
  42797=>"000000110",
  42798=>"110101000",
  42799=>"100001110",
  42800=>"010100000",
  42801=>"011001100",
  42802=>"100110001",
  42803=>"011101100",
  42804=>"110110101",
  42805=>"011111101",
  42806=>"000010100",
  42807=>"100110000",
  42808=>"000010001",
  42809=>"010001011",
  42810=>"010100000",
  42811=>"001111000",
  42812=>"000000101",
  42813=>"000010001",
  42814=>"001110000",
  42815=>"010101000",
  42816=>"000010011",
  42817=>"100111111",
  42818=>"100001001",
  42819=>"000010101",
  42820=>"101000110",
  42821=>"111010011",
  42822=>"001100000",
  42823=>"010000001",
  42824=>"001010010",
  42825=>"000110101",
  42826=>"000011100",
  42827=>"001101110",
  42828=>"010011010",
  42829=>"101010010",
  42830=>"000110101",
  42831=>"000101001",
  42832=>"110110001",
  42833=>"001110111",
  42834=>"010110111",
  42835=>"010000101",
  42836=>"111100000",
  42837=>"110110100",
  42838=>"001010001",
  42839=>"011110101",
  42840=>"011001011",
  42841=>"010100000",
  42842=>"110010011",
  42843=>"000000010",
  42844=>"100110110",
  42845=>"111111101",
  42846=>"001110001",
  42847=>"101100011",
  42848=>"010111000",
  42849=>"110000101",
  42850=>"000010100",
  42851=>"000110001",
  42852=>"111011001",
  42853=>"111000101",
  42854=>"110001111",
  42855=>"001101100",
  42856=>"011000010",
  42857=>"001001101",
  42858=>"100001010",
  42859=>"110000100",
  42860=>"010100010",
  42861=>"101001011",
  42862=>"111011101",
  42863=>"110000011",
  42864=>"100101110",
  42865=>"011011111",
  42866=>"111001001",
  42867=>"001010010",
  42868=>"001011010",
  42869=>"011100100",
  42870=>"010001111",
  42871=>"110011100",
  42872=>"111100010",
  42873=>"111011101",
  42874=>"100010101",
  42875=>"000010100",
  42876=>"010111011",
  42877=>"111100011",
  42878=>"010000101",
  42879=>"100010101",
  42880=>"001000001",
  42881=>"011011011",
  42882=>"000000111",
  42883=>"101100111",
  42884=>"010101101",
  42885=>"110101100",
  42886=>"101101010",
  42887=>"111011111",
  42888=>"110001111",
  42889=>"110101101",
  42890=>"111100111",
  42891=>"011000001",
  42892=>"001010111",
  42893=>"001110001",
  42894=>"100011010",
  42895=>"001000110",
  42896=>"001101000",
  42897=>"111011001",
  42898=>"010001100",
  42899=>"101100011",
  42900=>"101001101",
  42901=>"111001111",
  42902=>"101010100",
  42903=>"000101101",
  42904=>"001111101",
  42905=>"010101111",
  42906=>"010111001",
  42907=>"100000000",
  42908=>"011111110",
  42909=>"111000011",
  42910=>"110111010",
  42911=>"001000101",
  42912=>"001111011",
  42913=>"000011110",
  42914=>"110101001",
  42915=>"011001011",
  42916=>"111001011",
  42917=>"000110000",
  42918=>"110010100",
  42919=>"101101000",
  42920=>"110101000",
  42921=>"000010010",
  42922=>"110011011",
  42923=>"110010101",
  42924=>"001100010",
  42925=>"100101011",
  42926=>"110111110",
  42927=>"111011000",
  42928=>"011000001",
  42929=>"000001101",
  42930=>"011111110",
  42931=>"111100111",
  42932=>"111000001",
  42933=>"111001100",
  42934=>"111111110",
  42935=>"001101111",
  42936=>"100111110",
  42937=>"001010010",
  42938=>"100011010",
  42939=>"000100101",
  42940=>"111001001",
  42941=>"011010011",
  42942=>"000111100",
  42943=>"010111010",
  42944=>"000000001",
  42945=>"011000111",
  42946=>"110010111",
  42947=>"000101010",
  42948=>"010000111",
  42949=>"001010000",
  42950=>"001111010",
  42951=>"110110000",
  42952=>"111001101",
  42953=>"001010000",
  42954=>"010010010",
  42955=>"110110100",
  42956=>"111110101",
  42957=>"000001001",
  42958=>"100110001",
  42959=>"001111001",
  42960=>"010110011",
  42961=>"000110000",
  42962=>"011010001",
  42963=>"101110100",
  42964=>"011111011",
  42965=>"110011101",
  42966=>"101100000",
  42967=>"010111010",
  42968=>"000111101",
  42969=>"101010011",
  42970=>"001110100",
  42971=>"110000010",
  42972=>"010100100",
  42973=>"110110111",
  42974=>"000000101",
  42975=>"110011010",
  42976=>"010111111",
  42977=>"000000111",
  42978=>"001101100",
  42979=>"100101011",
  42980=>"010001100",
  42981=>"111110111",
  42982=>"001110110",
  42983=>"011111010",
  42984=>"101011011",
  42985=>"010110000",
  42986=>"111101111",
  42987=>"111011011",
  42988=>"110000110",
  42989=>"011110110",
  42990=>"010110111",
  42991=>"011011001",
  42992=>"011000100",
  42993=>"111010111",
  42994=>"011011000",
  42995=>"111111110",
  42996=>"011011011",
  42997=>"101010011",
  42998=>"110001100",
  42999=>"010101101",
  43000=>"111011110",
  43001=>"111111110",
  43002=>"110110010",
  43003=>"001111001",
  43004=>"011011010",
  43005=>"110001000",
  43006=>"110110000",
  43007=>"110110000",
  43008=>"010001110",
  43009=>"011100101",
  43010=>"000111001",
  43011=>"010110101",
  43012=>"110000110",
  43013=>"111101110",
  43014=>"111100100",
  43015=>"010000000",
  43016=>"111011101",
  43017=>"101110101",
  43018=>"101000010",
  43019=>"101100100",
  43020=>"000110010",
  43021=>"000000000",
  43022=>"010111111",
  43023=>"100000101",
  43024=>"100011111",
  43025=>"111000000",
  43026=>"011101100",
  43027=>"110111011",
  43028=>"000000011",
  43029=>"101000101",
  43030=>"110010111",
  43031=>"000101010",
  43032=>"000101100",
  43033=>"000001101",
  43034=>"110000101",
  43035=>"011111111",
  43036=>"010000100",
  43037=>"110000111",
  43038=>"100011101",
  43039=>"101110100",
  43040=>"011101010",
  43041=>"101101101",
  43042=>"001011000",
  43043=>"011111001",
  43044=>"111110100",
  43045=>"111011100",
  43046=>"101100001",
  43047=>"100101100",
  43048=>"000100001",
  43049=>"110010111",
  43050=>"100110110",
  43051=>"001110001",
  43052=>"110101110",
  43053=>"110100010",
  43054=>"011011111",
  43055=>"001111010",
  43056=>"001001000",
  43057=>"110110101",
  43058=>"000110010",
  43059=>"111101001",
  43060=>"111110110",
  43061=>"001100101",
  43062=>"010000100",
  43063=>"011101011",
  43064=>"000111000",
  43065=>"000010001",
  43066=>"101011011",
  43067=>"111000110",
  43068=>"000001011",
  43069=>"101101101",
  43070=>"111000010",
  43071=>"000011100",
  43072=>"111000000",
  43073=>"010000010",
  43074=>"010001100",
  43075=>"101110101",
  43076=>"011011010",
  43077=>"011111101",
  43078=>"000110010",
  43079=>"011111100",
  43080=>"101100011",
  43081=>"010100000",
  43082=>"001100100",
  43083=>"010000011",
  43084=>"001000101",
  43085=>"101110010",
  43086=>"101011001",
  43087=>"101110101",
  43088=>"111100100",
  43089=>"010011010",
  43090=>"101100101",
  43091=>"111010000",
  43092=>"111100001",
  43093=>"011110110",
  43094=>"100000000",
  43095=>"010100000",
  43096=>"110111001",
  43097=>"011111010",
  43098=>"111100110",
  43099=>"001100011",
  43100=>"100111000",
  43101=>"010001100",
  43102=>"011000011",
  43103=>"010110111",
  43104=>"100001011",
  43105=>"010010001",
  43106=>"001110000",
  43107=>"000000101",
  43108=>"000100110",
  43109=>"111000101",
  43110=>"000111101",
  43111=>"011100111",
  43112=>"100100010",
  43113=>"001010000",
  43114=>"100100000",
  43115=>"100000111",
  43116=>"000101000",
  43117=>"010111111",
  43118=>"101100110",
  43119=>"010010011",
  43120=>"101011101",
  43121=>"011010010",
  43122=>"010000101",
  43123=>"101000010",
  43124=>"000010011",
  43125=>"111000111",
  43126=>"100101110",
  43127=>"011000111",
  43128=>"111110010",
  43129=>"100011101",
  43130=>"011011001",
  43131=>"010100001",
  43132=>"110001111",
  43133=>"100111100",
  43134=>"001000001",
  43135=>"010010111",
  43136=>"001011001",
  43137=>"101010110",
  43138=>"101110110",
  43139=>"100000110",
  43140=>"100000111",
  43141=>"011111000",
  43142=>"100111000",
  43143=>"001000100",
  43144=>"111001111",
  43145=>"101001010",
  43146=>"011001011",
  43147=>"010110001",
  43148=>"001111001",
  43149=>"111010011",
  43150=>"100100011",
  43151=>"100000010",
  43152=>"100110100",
  43153=>"000110001",
  43154=>"011001010",
  43155=>"111111111",
  43156=>"011001100",
  43157=>"010111000",
  43158=>"001001000",
  43159=>"011110000",
  43160=>"110110001",
  43161=>"010011010",
  43162=>"100000000",
  43163=>"110100001",
  43164=>"000000111",
  43165=>"011011100",
  43166=>"000011111",
  43167=>"010001110",
  43168=>"101011011",
  43169=>"001011010",
  43170=>"100111110",
  43171=>"110101111",
  43172=>"010010010",
  43173=>"101100011",
  43174=>"011100000",
  43175=>"101001001",
  43176=>"001001011",
  43177=>"011101000",
  43178=>"000100000",
  43179=>"110000101",
  43180=>"100101110",
  43181=>"000011001",
  43182=>"101111011",
  43183=>"110010000",
  43184=>"000001010",
  43185=>"101001010",
  43186=>"000110111",
  43187=>"000110001",
  43188=>"110000110",
  43189=>"000100000",
  43190=>"101000111",
  43191=>"111111110",
  43192=>"010100001",
  43193=>"100110101",
  43194=>"111101100",
  43195=>"000000101",
  43196=>"001110011",
  43197=>"000111000",
  43198=>"000001011",
  43199=>"001101001",
  43200=>"110111110",
  43201=>"001101010",
  43202=>"000001010",
  43203=>"011100001",
  43204=>"011111101",
  43205=>"001001011",
  43206=>"011010100",
  43207=>"100100011",
  43208=>"111100010",
  43209=>"110111101",
  43210=>"101010110",
  43211=>"011000011",
  43212=>"100100000",
  43213=>"011111001",
  43214=>"010001000",
  43215=>"000000110",
  43216=>"011010001",
  43217=>"111001000",
  43218=>"110111001",
  43219=>"010100000",
  43220=>"111001011",
  43221=>"100101100",
  43222=>"000110000",
  43223=>"011101011",
  43224=>"110100101",
  43225=>"110111000",
  43226=>"000010001",
  43227=>"110100100",
  43228=>"001010010",
  43229=>"011010100",
  43230=>"011100111",
  43231=>"110010111",
  43232=>"000011100",
  43233=>"000011100",
  43234=>"000101110",
  43235=>"000010111",
  43236=>"010111100",
  43237=>"101001000",
  43238=>"001000010",
  43239=>"110101011",
  43240=>"010110011",
  43241=>"011001000",
  43242=>"010011100",
  43243=>"001010000",
  43244=>"111000001",
  43245=>"001001011",
  43246=>"000001110",
  43247=>"001111000",
  43248=>"001001001",
  43249=>"010011100",
  43250=>"010000000",
  43251=>"100011111",
  43252=>"110001111",
  43253=>"111101000",
  43254=>"000000100",
  43255=>"001101011",
  43256=>"011100100",
  43257=>"001110000",
  43258=>"111111100",
  43259=>"010010011",
  43260=>"110001111",
  43261=>"101010000",
  43262=>"101010010",
  43263=>"100111111",
  43264=>"111101111",
  43265=>"100100011",
  43266=>"101010001",
  43267=>"100111010",
  43268=>"011110110",
  43269=>"001011011",
  43270=>"000110011",
  43271=>"100111011",
  43272=>"010110100",
  43273=>"100000011",
  43274=>"111010010",
  43275=>"011101011",
  43276=>"000001101",
  43277=>"111111111",
  43278=>"010011010",
  43279=>"110001111",
  43280=>"110100001",
  43281=>"000101111",
  43282=>"110101111",
  43283=>"010011001",
  43284=>"111110000",
  43285=>"111100101",
  43286=>"111101011",
  43287=>"110101000",
  43288=>"101100101",
  43289=>"000100010",
  43290=>"100101110",
  43291=>"111001100",
  43292=>"110010010",
  43293=>"000100111",
  43294=>"111000110",
  43295=>"010000100",
  43296=>"011100100",
  43297=>"100011000",
  43298=>"001000110",
  43299=>"111101111",
  43300=>"111100111",
  43301=>"111111101",
  43302=>"111001001",
  43303=>"110001000",
  43304=>"000010010",
  43305=>"010111000",
  43306=>"000111000",
  43307=>"010000100",
  43308=>"011011111",
  43309=>"000000100",
  43310=>"000101011",
  43311=>"010010010",
  43312=>"111100011",
  43313=>"101110001",
  43314=>"111110010",
  43315=>"000000001",
  43316=>"000101101",
  43317=>"100000011",
  43318=>"000111111",
  43319=>"111100100",
  43320=>"110011001",
  43321=>"000101000",
  43322=>"111101110",
  43323=>"000000100",
  43324=>"000001100",
  43325=>"111101110",
  43326=>"001100100",
  43327=>"001011010",
  43328=>"111101110",
  43329=>"111110111",
  43330=>"111011011",
  43331=>"110011100",
  43332=>"101100101",
  43333=>"010011010",
  43334=>"000101000",
  43335=>"011010000",
  43336=>"100000001",
  43337=>"111101001",
  43338=>"110010011",
  43339=>"000010101",
  43340=>"000000101",
  43341=>"101100001",
  43342=>"001010011",
  43343=>"110110011",
  43344=>"111011000",
  43345=>"100011011",
  43346=>"100100111",
  43347=>"100010001",
  43348=>"001011101",
  43349=>"011101010",
  43350=>"001001011",
  43351=>"010011101",
  43352=>"110101001",
  43353=>"000001001",
  43354=>"000101101",
  43355=>"101001011",
  43356=>"100111001",
  43357=>"100011111",
  43358=>"000001011",
  43359=>"111110101",
  43360=>"011010011",
  43361=>"101111111",
  43362=>"110010010",
  43363=>"000110111",
  43364=>"001111000",
  43365=>"101101011",
  43366=>"110101001",
  43367=>"111111111",
  43368=>"000011000",
  43369=>"011101001",
  43370=>"111111001",
  43371=>"000011100",
  43372=>"101100001",
  43373=>"000101010",
  43374=>"001001011",
  43375=>"001101100",
  43376=>"000011011",
  43377=>"101001010",
  43378=>"001110001",
  43379=>"001100000",
  43380=>"001000101",
  43381=>"111101011",
  43382=>"110100010",
  43383=>"111100100",
  43384=>"100110000",
  43385=>"101101100",
  43386=>"110000010",
  43387=>"011101010",
  43388=>"110110100",
  43389=>"000001101",
  43390=>"001111001",
  43391=>"001111111",
  43392=>"000100110",
  43393=>"010010101",
  43394=>"010110100",
  43395=>"011101111",
  43396=>"011101010",
  43397=>"011010111",
  43398=>"101111110",
  43399=>"001101100",
  43400=>"000110100",
  43401=>"011001111",
  43402=>"101100101",
  43403=>"000100100",
  43404=>"011100000",
  43405=>"001010010",
  43406=>"011001010",
  43407=>"010000110",
  43408=>"100001001",
  43409=>"000011001",
  43410=>"101111011",
  43411=>"011001101",
  43412=>"000111111",
  43413=>"100111010",
  43414=>"001101111",
  43415=>"111010101",
  43416=>"001111110",
  43417=>"100100101",
  43418=>"011101011",
  43419=>"000100000",
  43420=>"011101101",
  43421=>"111111111",
  43422=>"010100111",
  43423=>"010110100",
  43424=>"001100000",
  43425=>"001011111",
  43426=>"011110001",
  43427=>"000010101",
  43428=>"001110110",
  43429=>"101000000",
  43430=>"000001100",
  43431=>"110101111",
  43432=>"110110001",
  43433=>"111110110",
  43434=>"000000111",
  43435=>"100101001",
  43436=>"001100101",
  43437=>"100011110",
  43438=>"111000001",
  43439=>"001111111",
  43440=>"100101011",
  43441=>"101100100",
  43442=>"010100100",
  43443=>"011011000",
  43444=>"101101010",
  43445=>"110010010",
  43446=>"000010111",
  43447=>"100100110",
  43448=>"101110110",
  43449=>"001110110",
  43450=>"000000010",
  43451=>"110000010",
  43452=>"010011000",
  43453=>"101000000",
  43454=>"111100010",
  43455=>"010101110",
  43456=>"000001001",
  43457=>"000011010",
  43458=>"100100110",
  43459=>"110111001",
  43460=>"100100010",
  43461=>"100000010",
  43462=>"111000000",
  43463=>"000101100",
  43464=>"001101111",
  43465=>"010110011",
  43466=>"001000000",
  43467=>"100111101",
  43468=>"100000110",
  43469=>"110000110",
  43470=>"000111010",
  43471=>"000000000",
  43472=>"000110000",
  43473=>"001100000",
  43474=>"101110110",
  43475=>"001011000",
  43476=>"001111111",
  43477=>"000011010",
  43478=>"111111100",
  43479=>"011111110",
  43480=>"101001111",
  43481=>"101010100",
  43482=>"010100101",
  43483=>"011110110",
  43484=>"100111010",
  43485=>"111111001",
  43486=>"011100100",
  43487=>"101000100",
  43488=>"010101000",
  43489=>"001111011",
  43490=>"101101110",
  43491=>"100010010",
  43492=>"101001111",
  43493=>"100010111",
  43494=>"100100000",
  43495=>"000100011",
  43496=>"000100010",
  43497=>"110001001",
  43498=>"100011011",
  43499=>"110001001",
  43500=>"001010101",
  43501=>"111111001",
  43502=>"010010000",
  43503=>"011010100",
  43504=>"010111001",
  43505=>"111100100",
  43506=>"010101001",
  43507=>"101101010",
  43508=>"110010000",
  43509=>"101110101",
  43510=>"111110011",
  43511=>"110110000",
  43512=>"101010001",
  43513=>"100001011",
  43514=>"011000001",
  43515=>"111111111",
  43516=>"000001111",
  43517=>"110010101",
  43518=>"011111110",
  43519=>"101011000",
  43520=>"001110111",
  43521=>"010001111",
  43522=>"110100010",
  43523=>"101001101",
  43524=>"100100011",
  43525=>"000000111",
  43526=>"011110011",
  43527=>"011110010",
  43528=>"111010100",
  43529=>"100000110",
  43530=>"000101110",
  43531=>"101010000",
  43532=>"100000001",
  43533=>"001001001",
  43534=>"111000011",
  43535=>"001111111",
  43536=>"010000101",
  43537=>"111111110",
  43538=>"110100111",
  43539=>"011110101",
  43540=>"011110100",
  43541=>"110111100",
  43542=>"011110010",
  43543=>"110000001",
  43544=>"010100111",
  43545=>"101110111",
  43546=>"000000100",
  43547=>"000000010",
  43548=>"110001101",
  43549=>"100001111",
  43550=>"011110000",
  43551=>"001110111",
  43552=>"110000111",
  43553=>"010110100",
  43554=>"000000010",
  43555=>"010010011",
  43556=>"000011110",
  43557=>"111110100",
  43558=>"000001100",
  43559=>"111001100",
  43560=>"011110000",
  43561=>"000111110",
  43562=>"000001000",
  43563=>"110000011",
  43564=>"100101010",
  43565=>"101010000",
  43566=>"000000111",
  43567=>"111111100",
  43568=>"010100110",
  43569=>"100000111",
  43570=>"000000110",
  43571=>"000111100",
  43572=>"000100001",
  43573=>"010100000",
  43574=>"101110100",
  43575=>"100111101",
  43576=>"001111101",
  43577=>"001111000",
  43578=>"101100001",
  43579=>"110101010",
  43580=>"110110000",
  43581=>"011110110",
  43582=>"110110000",
  43583=>"110111101",
  43584=>"001011001",
  43585=>"000000100",
  43586=>"100000011",
  43587=>"110001010",
  43588=>"001100011",
  43589=>"111111011",
  43590=>"100100101",
  43591=>"010110111",
  43592=>"011100001",
  43593=>"011011100",
  43594=>"001111000",
  43595=>"110100111",
  43596=>"011101000",
  43597=>"010000001",
  43598=>"110010000",
  43599=>"111000101",
  43600=>"101110100",
  43601=>"000000000",
  43602=>"011001001",
  43603=>"101010100",
  43604=>"000111111",
  43605=>"000111110",
  43606=>"010001011",
  43607=>"110000010",
  43608=>"101111111",
  43609=>"111001110",
  43610=>"000001001",
  43611=>"001000111",
  43612=>"011010110",
  43613=>"101011010",
  43614=>"000011101",
  43615=>"111111010",
  43616=>"011001011",
  43617=>"111100001",
  43618=>"111010010",
  43619=>"000011001",
  43620=>"000100000",
  43621=>"000010101",
  43622=>"000110101",
  43623=>"000100101",
  43624=>"111000000",
  43625=>"000011101",
  43626=>"111100101",
  43627=>"001100101",
  43628=>"100111000",
  43629=>"111010100",
  43630=>"000011101",
  43631=>"100111111",
  43632=>"011010110",
  43633=>"100001000",
  43634=>"111011100",
  43635=>"100001111",
  43636=>"010000100",
  43637=>"010110010",
  43638=>"100001000",
  43639=>"010111000",
  43640=>"011000000",
  43641=>"101100111",
  43642=>"111100010",
  43643=>"101000001",
  43644=>"001010110",
  43645=>"111101011",
  43646=>"111011110",
  43647=>"100111010",
  43648=>"111101111",
  43649=>"001011011",
  43650=>"000001111",
  43651=>"000001001",
  43652=>"100100000",
  43653=>"010010100",
  43654=>"110000010",
  43655=>"110111001",
  43656=>"010010000",
  43657=>"001110001",
  43658=>"110101010",
  43659=>"101011010",
  43660=>"001100001",
  43661=>"010100111",
  43662=>"111001001",
  43663=>"001111010",
  43664=>"011000000",
  43665=>"100010001",
  43666=>"010110000",
  43667=>"010101000",
  43668=>"010110100",
  43669=>"101110110",
  43670=>"000100101",
  43671=>"100011001",
  43672=>"101100101",
  43673=>"111101000",
  43674=>"110010010",
  43675=>"001111110",
  43676=>"000100001",
  43677=>"111000000",
  43678=>"111110011",
  43679=>"101001010",
  43680=>"111110011",
  43681=>"110101101",
  43682=>"100101000",
  43683=>"111101110",
  43684=>"100110101",
  43685=>"111101110",
  43686=>"010000100",
  43687=>"010000101",
  43688=>"000101111",
  43689=>"101100001",
  43690=>"110101011",
  43691=>"110000010",
  43692=>"010101111",
  43693=>"101111100",
  43694=>"110110100",
  43695=>"010111111",
  43696=>"001000111",
  43697=>"110011001",
  43698=>"001100101",
  43699=>"010001001",
  43700=>"000110010",
  43701=>"100011100",
  43702=>"010001110",
  43703=>"000100110",
  43704=>"110100001",
  43705=>"101101101",
  43706=>"110100000",
  43707=>"001000101",
  43708=>"001100110",
  43709=>"011110110",
  43710=>"010001110",
  43711=>"010111101",
  43712=>"101011101",
  43713=>"100001110",
  43714=>"110111010",
  43715=>"110100011",
  43716=>"100010001",
  43717=>"011000100",
  43718=>"100001000",
  43719=>"100000111",
  43720=>"000101100",
  43721=>"101010001",
  43722=>"010101110",
  43723=>"101101100",
  43724=>"010110000",
  43725=>"101010100",
  43726=>"110010001",
  43727=>"101011010",
  43728=>"111000111",
  43729=>"011011010",
  43730=>"110010010",
  43731=>"101100001",
  43732=>"001100111",
  43733=>"100000001",
  43734=>"101101110",
  43735=>"010111011",
  43736=>"001101000",
  43737=>"010011100",
  43738=>"111101011",
  43739=>"000001101",
  43740=>"100110001",
  43741=>"111011000",
  43742=>"110011110",
  43743=>"000001101",
  43744=>"100000100",
  43745=>"000000100",
  43746=>"000011100",
  43747=>"010001111",
  43748=>"101000100",
  43749=>"011001011",
  43750=>"011011111",
  43751=>"001000010",
  43752=>"000100011",
  43753=>"100011111",
  43754=>"111101001",
  43755=>"010010111",
  43756=>"010100000",
  43757=>"101011100",
  43758=>"100001011",
  43759=>"000001000",
  43760=>"110100100",
  43761=>"100111010",
  43762=>"101001010",
  43763=>"101101100",
  43764=>"000111011",
  43765=>"111111101",
  43766=>"100111111",
  43767=>"111010100",
  43768=>"101001101",
  43769=>"111000101",
  43770=>"010101110",
  43771=>"101100111",
  43772=>"111001000",
  43773=>"011011111",
  43774=>"010001001",
  43775=>"000011011",
  43776=>"010000101",
  43777=>"000111100",
  43778=>"001011010",
  43779=>"010110000",
  43780=>"000001111",
  43781=>"111111001",
  43782=>"000110100",
  43783=>"110011101",
  43784=>"010100110",
  43785=>"110001010",
  43786=>"111111010",
  43787=>"101010111",
  43788=>"100110000",
  43789=>"110000101",
  43790=>"011100011",
  43791=>"000101011",
  43792=>"001110111",
  43793=>"101110010",
  43794=>"010000101",
  43795=>"001101110",
  43796=>"110001001",
  43797=>"000000000",
  43798=>"110000101",
  43799=>"000000010",
  43800=>"110101000",
  43801=>"001101100",
  43802=>"000100001",
  43803=>"100100110",
  43804=>"001000000",
  43805=>"100001000",
  43806=>"111101111",
  43807=>"011100011",
  43808=>"011110010",
  43809=>"111001000",
  43810=>"011011010",
  43811=>"011001100",
  43812=>"001001000",
  43813=>"110100111",
  43814=>"100010011",
  43815=>"110111101",
  43816=>"100000101",
  43817=>"101111010",
  43818=>"010110011",
  43819=>"110100011",
  43820=>"000010111",
  43821=>"001111000",
  43822=>"010011000",
  43823=>"010100100",
  43824=>"001011111",
  43825=>"110110101",
  43826=>"000000000",
  43827=>"000101000",
  43828=>"000101010",
  43829=>"011010011",
  43830=>"011110011",
  43831=>"101000010",
  43832=>"100111010",
  43833=>"011101110",
  43834=>"110010010",
  43835=>"010110101",
  43836=>"100100101",
  43837=>"000010101",
  43838=>"101101111",
  43839=>"011001000",
  43840=>"101010001",
  43841=>"101111011",
  43842=>"011111010",
  43843=>"000111010",
  43844=>"001111111",
  43845=>"100001111",
  43846=>"001000001",
  43847=>"101001101",
  43848=>"101011011",
  43849=>"010001010",
  43850=>"010010111",
  43851=>"101001100",
  43852=>"010001111",
  43853=>"011000101",
  43854=>"000100100",
  43855=>"111001010",
  43856=>"001001110",
  43857=>"000110111",
  43858=>"000101100",
  43859=>"011001100",
  43860=>"000001100",
  43861=>"001010010",
  43862=>"000110111",
  43863=>"001111100",
  43864=>"010101101",
  43865=>"110011101",
  43866=>"010000011",
  43867=>"111101000",
  43868=>"101000000",
  43869=>"000000010",
  43870=>"110011100",
  43871=>"100100001",
  43872=>"011001101",
  43873=>"101011010",
  43874=>"100001001",
  43875=>"110011100",
  43876=>"110110100",
  43877=>"101001111",
  43878=>"111110111",
  43879=>"110110100",
  43880=>"000011010",
  43881=>"110100011",
  43882=>"110100101",
  43883=>"101111011",
  43884=>"111100011",
  43885=>"111111110",
  43886=>"000101101",
  43887=>"100101100",
  43888=>"000101101",
  43889=>"001000101",
  43890=>"110011000",
  43891=>"011010000",
  43892=>"101001110",
  43893=>"100010000",
  43894=>"110010100",
  43895=>"100010101",
  43896=>"110111111",
  43897=>"111011011",
  43898=>"011011110",
  43899=>"101010100",
  43900=>"000011001",
  43901=>"100000110",
  43902=>"110011111",
  43903=>"010100000",
  43904=>"110000111",
  43905=>"001001000",
  43906=>"100011010",
  43907=>"111011000",
  43908=>"111000000",
  43909=>"011010100",
  43910=>"110110011",
  43911=>"100010000",
  43912=>"011110001",
  43913=>"011111001",
  43914=>"111111111",
  43915=>"000001110",
  43916=>"001101010",
  43917=>"001011100",
  43918=>"011001010",
  43919=>"010110011",
  43920=>"100001101",
  43921=>"101111101",
  43922=>"001110100",
  43923=>"011101001",
  43924=>"100010010",
  43925=>"000111110",
  43926=>"111001100",
  43927=>"001011111",
  43928=>"110100100",
  43929=>"101100001",
  43930=>"000000000",
  43931=>"011111001",
  43932=>"111110011",
  43933=>"110000011",
  43934=>"101101000",
  43935=>"000010110",
  43936=>"010100010",
  43937=>"001110110",
  43938=>"100011011",
  43939=>"000000000",
  43940=>"100110110",
  43941=>"101101001",
  43942=>"001000000",
  43943=>"111000010",
  43944=>"101100100",
  43945=>"000011100",
  43946=>"111010011",
  43947=>"100111111",
  43948=>"000001111",
  43949=>"101111000",
  43950=>"111000111",
  43951=>"000011110",
  43952=>"000100100",
  43953=>"010101111",
  43954=>"100110000",
  43955=>"111010010",
  43956=>"111101111",
  43957=>"111001011",
  43958=>"011011100",
  43959=>"000011001",
  43960=>"111100011",
  43961=>"011110111",
  43962=>"011110011",
  43963=>"011111100",
  43964=>"111010011",
  43965=>"001010010",
  43966=>"011011111",
  43967=>"100101000",
  43968=>"011100111",
  43969=>"111010000",
  43970=>"010111101",
  43971=>"111111111",
  43972=>"100100000",
  43973=>"010111110",
  43974=>"010101100",
  43975=>"010010101",
  43976=>"000011011",
  43977=>"101011100",
  43978=>"010100101",
  43979=>"001100100",
  43980=>"101100101",
  43981=>"010000000",
  43982=>"011001010",
  43983=>"010011000",
  43984=>"100100111",
  43985=>"101011101",
  43986=>"100101000",
  43987=>"001001110",
  43988=>"010110010",
  43989=>"100000101",
  43990=>"101000110",
  43991=>"000101110",
  43992=>"000000110",
  43993=>"000001001",
  43994=>"010100101",
  43995=>"101110000",
  43996=>"110100001",
  43997=>"111110001",
  43998=>"100101011",
  43999=>"001110111",
  44000=>"011100111",
  44001=>"110110000",
  44002=>"100111011",
  44003=>"110111110",
  44004=>"101000010",
  44005=>"100010100",
  44006=>"010111101",
  44007=>"110101110",
  44008=>"101111101",
  44009=>"011110101",
  44010=>"110001100",
  44011=>"000010000",
  44012=>"000011111",
  44013=>"110101100",
  44014=>"000001000",
  44015=>"111110100",
  44016=>"111111011",
  44017=>"010000000",
  44018=>"110001010",
  44019=>"011011011",
  44020=>"110100110",
  44021=>"011011001",
  44022=>"011101111",
  44023=>"011111001",
  44024=>"010100110",
  44025=>"011110100",
  44026=>"111010110",
  44027=>"010000110",
  44028=>"011101010",
  44029=>"110110110",
  44030=>"011000111",
  44031=>"000100010",
  44032=>"010001000",
  44033=>"100110111",
  44034=>"000110000",
  44035=>"010011100",
  44036=>"101000111",
  44037=>"101000101",
  44038=>"001010000",
  44039=>"010110010",
  44040=>"110001000",
  44041=>"000011111",
  44042=>"011010100",
  44043=>"110010011",
  44044=>"100100100",
  44045=>"011111100",
  44046=>"011001011",
  44047=>"110110111",
  44048=>"001001000",
  44049=>"110010101",
  44050=>"010110101",
  44051=>"001101110",
  44052=>"010111011",
  44053=>"001001010",
  44054=>"110100001",
  44055=>"010000111",
  44056=>"111001000",
  44057=>"110100011",
  44058=>"111000101",
  44059=>"100011101",
  44060=>"100111010",
  44061=>"011011111",
  44062=>"000110101",
  44063=>"001010011",
  44064=>"011011000",
  44065=>"101100000",
  44066=>"110100000",
  44067=>"011011001",
  44068=>"100010011",
  44069=>"001011100",
  44070=>"010001001",
  44071=>"111101111",
  44072=>"110000000",
  44073=>"000000111",
  44074=>"011101111",
  44075=>"000000100",
  44076=>"111110000",
  44077=>"111100111",
  44078=>"111011101",
  44079=>"010011000",
  44080=>"011101001",
  44081=>"111000100",
  44082=>"010011000",
  44083=>"111101011",
  44084=>"100000000",
  44085=>"010000100",
  44086=>"001100110",
  44087=>"000011111",
  44088=>"011111000",
  44089=>"000011011",
  44090=>"100011001",
  44091=>"111101010",
  44092=>"111100011",
  44093=>"101100101",
  44094=>"010111101",
  44095=>"001111010",
  44096=>"110001001",
  44097=>"011000110",
  44098=>"010011011",
  44099=>"101100111",
  44100=>"010101100",
  44101=>"011001101",
  44102=>"000101101",
  44103=>"101000101",
  44104=>"100101001",
  44105=>"010110100",
  44106=>"010101110",
  44107=>"000011101",
  44108=>"110000111",
  44109=>"110010011",
  44110=>"100101001",
  44111=>"010100010",
  44112=>"001001100",
  44113=>"000000001",
  44114=>"111010011",
  44115=>"001101011",
  44116=>"100000001",
  44117=>"100111101",
  44118=>"011101010",
  44119=>"001101111",
  44120=>"000010010",
  44121=>"001010111",
  44122=>"110110000",
  44123=>"100100111",
  44124=>"100111010",
  44125=>"111110000",
  44126=>"100010001",
  44127=>"001001010",
  44128=>"101010000",
  44129=>"111100110",
  44130=>"111001111",
  44131=>"111010111",
  44132=>"000111000",
  44133=>"111011010",
  44134=>"011110111",
  44135=>"001010111",
  44136=>"000010001",
  44137=>"111010111",
  44138=>"000010001",
  44139=>"010110100",
  44140=>"100001100",
  44141=>"000001101",
  44142=>"101100000",
  44143=>"110101110",
  44144=>"111101100",
  44145=>"100101100",
  44146=>"110001110",
  44147=>"110101011",
  44148=>"000010111",
  44149=>"111110111",
  44150=>"100011000",
  44151=>"011111001",
  44152=>"101010111",
  44153=>"010101100",
  44154=>"111010110",
  44155=>"010110110",
  44156=>"111010100",
  44157=>"001101100",
  44158=>"001001100",
  44159=>"010110000",
  44160=>"011000000",
  44161=>"111110100",
  44162=>"111011000",
  44163=>"100100001",
  44164=>"101110110",
  44165=>"110000110",
  44166=>"100010100",
  44167=>"011101110",
  44168=>"000001110",
  44169=>"111100001",
  44170=>"100101011",
  44171=>"101110001",
  44172=>"110010001",
  44173=>"010000010",
  44174=>"010001110",
  44175=>"000100000",
  44176=>"100001111",
  44177=>"110110011",
  44178=>"110111100",
  44179=>"100011100",
  44180=>"011000110",
  44181=>"001110110",
  44182=>"101101101",
  44183=>"111100001",
  44184=>"001010010",
  44185=>"101100010",
  44186=>"111100001",
  44187=>"110011001",
  44188=>"010110111",
  44189=>"000011101",
  44190=>"011110101",
  44191=>"100000001",
  44192=>"110011110",
  44193=>"100001001",
  44194=>"000010111",
  44195=>"111011110",
  44196=>"011110000",
  44197=>"001001000",
  44198=>"000010100",
  44199=>"000111111",
  44200=>"101011010",
  44201=>"101011100",
  44202=>"011000000",
  44203=>"011010101",
  44204=>"000000010",
  44205=>"111010111",
  44206=>"001001010",
  44207=>"100011101",
  44208=>"000011000",
  44209=>"010100011",
  44210=>"000010100",
  44211=>"110000010",
  44212=>"100110110",
  44213=>"000110010",
  44214=>"010100100",
  44215=>"011000100",
  44216=>"110000100",
  44217=>"001011111",
  44218=>"101000110",
  44219=>"000010001",
  44220=>"010011000",
  44221=>"110011110",
  44222=>"011111101",
  44223=>"011111011",
  44224=>"000110001",
  44225=>"000001101",
  44226=>"101011111",
  44227=>"000001011",
  44228=>"001101011",
  44229=>"000101001",
  44230=>"010010111",
  44231=>"001101101",
  44232=>"110011001",
  44233=>"001011011",
  44234=>"101011100",
  44235=>"100001110",
  44236=>"100110010",
  44237=>"101110000",
  44238=>"110100111",
  44239=>"011101001",
  44240=>"101101111",
  44241=>"101001110",
  44242=>"000011000",
  44243=>"111001001",
  44244=>"111011111",
  44245=>"101110011",
  44246=>"110001110",
  44247=>"011000101",
  44248=>"111111011",
  44249=>"010010000",
  44250=>"000001011",
  44251=>"011001111",
  44252=>"000110011",
  44253=>"001001011",
  44254=>"010101111",
  44255=>"100011000",
  44256=>"101110010",
  44257=>"000100000",
  44258=>"011110100",
  44259=>"011110101",
  44260=>"111111110",
  44261=>"110000111",
  44262=>"001100100",
  44263=>"100111000",
  44264=>"101100111",
  44265=>"110001011",
  44266=>"111111100",
  44267=>"010100011",
  44268=>"100011001",
  44269=>"001010110",
  44270=>"000000111",
  44271=>"000010000",
  44272=>"010101101",
  44273=>"000010010",
  44274=>"110000101",
  44275=>"001000100",
  44276=>"011001010",
  44277=>"010110010",
  44278=>"000101010",
  44279=>"111110101",
  44280=>"110101000",
  44281=>"000111111",
  44282=>"010001101",
  44283=>"100001100",
  44284=>"000100110",
  44285=>"001101000",
  44286=>"100000011",
  44287=>"010000111",
  44288=>"111110111",
  44289=>"101011000",
  44290=>"000110111",
  44291=>"110000100",
  44292=>"010110000",
  44293=>"000010111",
  44294=>"001110000",
  44295=>"101101110",
  44296=>"100110111",
  44297=>"011010110",
  44298=>"010000101",
  44299=>"001111011",
  44300=>"000010110",
  44301=>"001000111",
  44302=>"010100010",
  44303=>"010001000",
  44304=>"100101100",
  44305=>"111111111",
  44306=>"011001001",
  44307=>"111100000",
  44308=>"001001001",
  44309=>"101000111",
  44310=>"011010001",
  44311=>"011000011",
  44312=>"001001111",
  44313=>"101010010",
  44314=>"000011100",
  44315=>"011100001",
  44316=>"110101010",
  44317=>"110110111",
  44318=>"100111111",
  44319=>"100100001",
  44320=>"001101101",
  44321=>"110111000",
  44322=>"001001010",
  44323=>"111010011",
  44324=>"101001100",
  44325=>"111110110",
  44326=>"001111111",
  44327=>"010111110",
  44328=>"110100101",
  44329=>"111110110",
  44330=>"100000100",
  44331=>"010001101",
  44332=>"101110110",
  44333=>"111101000",
  44334=>"110001000",
  44335=>"101101101",
  44336=>"011010110",
  44337=>"101110001",
  44338=>"000000111",
  44339=>"001111010",
  44340=>"110110110",
  44341=>"110110011",
  44342=>"011010111",
  44343=>"101110101",
  44344=>"001001100",
  44345=>"010011111",
  44346=>"100101001",
  44347=>"000001010",
  44348=>"011010000",
  44349=>"111011111",
  44350=>"111001000",
  44351=>"111111111",
  44352=>"111110110",
  44353=>"010000010",
  44354=>"111011110",
  44355=>"101001101",
  44356=>"111100111",
  44357=>"111111010",
  44358=>"011100000",
  44359=>"010010001",
  44360=>"011010111",
  44361=>"011100111",
  44362=>"101001110",
  44363=>"010000111",
  44364=>"000011100",
  44365=>"010110100",
  44366=>"110000000",
  44367=>"011110111",
  44368=>"110010011",
  44369=>"011111111",
  44370=>"011001010",
  44371=>"010010011",
  44372=>"001011001",
  44373=>"101000111",
  44374=>"011101001",
  44375=>"000011000",
  44376=>"100001011",
  44377=>"001001101",
  44378=>"010011000",
  44379=>"001011101",
  44380=>"000001000",
  44381=>"100111111",
  44382=>"001010011",
  44383=>"110011101",
  44384=>"101110010",
  44385=>"011000001",
  44386=>"011000001",
  44387=>"101011111",
  44388=>"100100110",
  44389=>"011010110",
  44390=>"101100001",
  44391=>"101111110",
  44392=>"110011101",
  44393=>"110011000",
  44394=>"001001000",
  44395=>"110010100",
  44396=>"010110010",
  44397=>"000001000",
  44398=>"000110000",
  44399=>"110100001",
  44400=>"010001110",
  44401=>"111101110",
  44402=>"000011110",
  44403=>"100111101",
  44404=>"110101001",
  44405=>"000001111",
  44406=>"110100110",
  44407=>"000100011",
  44408=>"101001110",
  44409=>"001110001",
  44410=>"100100000",
  44411=>"111001010",
  44412=>"000000000",
  44413=>"101011000",
  44414=>"100001100",
  44415=>"111011000",
  44416=>"100001000",
  44417=>"111110000",
  44418=>"001110101",
  44419=>"010111111",
  44420=>"011110101",
  44421=>"110010100",
  44422=>"000010011",
  44423=>"101010101",
  44424=>"110101111",
  44425=>"001100001",
  44426=>"010001001",
  44427=>"000101011",
  44428=>"010100111",
  44429=>"110001111",
  44430=>"101001101",
  44431=>"011111101",
  44432=>"011100000",
  44433=>"100100011",
  44434=>"010011110",
  44435=>"111110011",
  44436=>"010011000",
  44437=>"110111110",
  44438=>"110100010",
  44439=>"111111100",
  44440=>"001001100",
  44441=>"010000010",
  44442=>"101111101",
  44443=>"000111000",
  44444=>"001110111",
  44445=>"111111111",
  44446=>"000010000",
  44447=>"011011100",
  44448=>"000110110",
  44449=>"111010011",
  44450=>"100101001",
  44451=>"100100001",
  44452=>"011100001",
  44453=>"111111001",
  44454=>"010000000",
  44455=>"000001000",
  44456=>"011000110",
  44457=>"101110101",
  44458=>"111100111",
  44459=>"111001100",
  44460=>"000010001",
  44461=>"001011111",
  44462=>"000000000",
  44463=>"101001001",
  44464=>"111010010",
  44465=>"110001101",
  44466=>"000110100",
  44467=>"111011110",
  44468=>"010001111",
  44469=>"111110101",
  44470=>"001110110",
  44471=>"111001000",
  44472=>"010101101",
  44473=>"100101110",
  44474=>"000100100",
  44475=>"101000000",
  44476=>"000111011",
  44477=>"101101001",
  44478=>"001110010",
  44479=>"111101010",
  44480=>"100001100",
  44481=>"010001000",
  44482=>"111101001",
  44483=>"111101101",
  44484=>"100100111",
  44485=>"011000011",
  44486=>"011111111",
  44487=>"111000101",
  44488=>"111010001",
  44489=>"111111110",
  44490=>"010101100",
  44491=>"110111011",
  44492=>"010101101",
  44493=>"000100101",
  44494=>"101101110",
  44495=>"010001010",
  44496=>"000010101",
  44497=>"000000000",
  44498=>"101101101",
  44499=>"110011000",
  44500=>"001001011",
  44501=>"110110100",
  44502=>"111000100",
  44503=>"100000001",
  44504=>"110001100",
  44505=>"001011110",
  44506=>"111101011",
  44507=>"110101011",
  44508=>"110000101",
  44509=>"101101011",
  44510=>"000001000",
  44511=>"010000000",
  44512=>"011001100",
  44513=>"011110101",
  44514=>"101000100",
  44515=>"111001100",
  44516=>"100110100",
  44517=>"100000001",
  44518=>"101010100",
  44519=>"111010111",
  44520=>"100100100",
  44521=>"000011011",
  44522=>"011101100",
  44523=>"000010010",
  44524=>"000110110",
  44525=>"011111110",
  44526=>"010110110",
  44527=>"011100000",
  44528=>"101110101",
  44529=>"011100110",
  44530=>"011001010",
  44531=>"101010101",
  44532=>"111101001",
  44533=>"001100011",
  44534=>"000101000",
  44535=>"011011010",
  44536=>"100100101",
  44537=>"111100110",
  44538=>"111010010",
  44539=>"011000001",
  44540=>"111010001",
  44541=>"001110001",
  44542=>"001100000",
  44543=>"111010001",
  44544=>"100110000",
  44545=>"010010100",
  44546=>"111100010",
  44547=>"100111110",
  44548=>"111100100",
  44549=>"100000001",
  44550=>"110100110",
  44551=>"001111001",
  44552=>"110110001",
  44553=>"100011100",
  44554=>"001111000",
  44555=>"011100100",
  44556=>"011001000",
  44557=>"001101010",
  44558=>"111000111",
  44559=>"001100100",
  44560=>"011101010",
  44561=>"000111000",
  44562=>"111111100",
  44563=>"111011101",
  44564=>"010010100",
  44565=>"111011101",
  44566=>"001110000",
  44567=>"010101010",
  44568=>"000110001",
  44569=>"010100111",
  44570=>"110100000",
  44571=>"101011101",
  44572=>"111101011",
  44573=>"010100000",
  44574=>"111110101",
  44575=>"110010010",
  44576=>"010100110",
  44577=>"101111110",
  44578=>"110001111",
  44579=>"000100100",
  44580=>"000011110",
  44581=>"000010001",
  44582=>"111011111",
  44583=>"101010100",
  44584=>"101101111",
  44585=>"000100001",
  44586=>"110100111",
  44587=>"010010101",
  44588=>"000010101",
  44589=>"000000001",
  44590=>"011011111",
  44591=>"001001000",
  44592=>"111000111",
  44593=>"100110001",
  44594=>"111111111",
  44595=>"010111110",
  44596=>"010000011",
  44597=>"001011001",
  44598=>"100000100",
  44599=>"001100111",
  44600=>"111001000",
  44601=>"011001110",
  44602=>"001000011",
  44603=>"110011101",
  44604=>"010111011",
  44605=>"001000000",
  44606=>"110000001",
  44607=>"001010000",
  44608=>"111110111",
  44609=>"110111011",
  44610=>"010101101",
  44611=>"101111110",
  44612=>"110111100",
  44613=>"001011001",
  44614=>"001110111",
  44615=>"011011001",
  44616=>"110011100",
  44617=>"011111101",
  44618=>"011000100",
  44619=>"100001001",
  44620=>"001000001",
  44621=>"101001111",
  44622=>"001010000",
  44623=>"011010000",
  44624=>"101110000",
  44625=>"001101111",
  44626=>"101110110",
  44627=>"000101110",
  44628=>"101001110",
  44629=>"001010000",
  44630=>"100110011",
  44631=>"110000110",
  44632=>"100001001",
  44633=>"110001000",
  44634=>"110001111",
  44635=>"001000111",
  44636=>"111010111",
  44637=>"011000111",
  44638=>"000001000",
  44639=>"101111000",
  44640=>"010110111",
  44641=>"101100011",
  44642=>"111110100",
  44643=>"000011110",
  44644=>"100001111",
  44645=>"111011110",
  44646=>"001100011",
  44647=>"100000010",
  44648=>"000000111",
  44649=>"000010000",
  44650=>"010011111",
  44651=>"001100000",
  44652=>"010001010",
  44653=>"011000001",
  44654=>"100101001",
  44655=>"000110110",
  44656=>"001101100",
  44657=>"101000110",
  44658=>"001010001",
  44659=>"101111100",
  44660=>"110101001",
  44661=>"111000111",
  44662=>"100111000",
  44663=>"000010111",
  44664=>"101011011",
  44665=>"111011100",
  44666=>"011010111",
  44667=>"100001000",
  44668=>"110001010",
  44669=>"111110101",
  44670=>"111100000",
  44671=>"000111111",
  44672=>"110100111",
  44673=>"001001000",
  44674=>"111011101",
  44675=>"010001010",
  44676=>"100000011",
  44677=>"110000011",
  44678=>"001101101",
  44679=>"010100101",
  44680=>"011111000",
  44681=>"111010100",
  44682=>"001011101",
  44683=>"000010110",
  44684=>"010000001",
  44685=>"110100100",
  44686=>"111111011",
  44687=>"110110101",
  44688=>"100111111",
  44689=>"001001011",
  44690=>"110100101",
  44691=>"010100110",
  44692=>"001010000",
  44693=>"001101010",
  44694=>"111110001",
  44695=>"101000000",
  44696=>"010000110",
  44697=>"101110001",
  44698=>"010011011",
  44699=>"010110100",
  44700=>"111110111",
  44701=>"000111010",
  44702=>"110100110",
  44703=>"100110111",
  44704=>"111111000",
  44705=>"110111111",
  44706=>"111111011",
  44707=>"001000101",
  44708=>"100010101",
  44709=>"011001111",
  44710=>"110100011",
  44711=>"001000011",
  44712=>"000011001",
  44713=>"111111101",
  44714=>"011100101",
  44715=>"010001000",
  44716=>"000101111",
  44717=>"001000101",
  44718=>"100001111",
  44719=>"010100010",
  44720=>"110010111",
  44721=>"010011011",
  44722=>"010000010",
  44723=>"000001101",
  44724=>"011100011",
  44725=>"011010110",
  44726=>"111101011",
  44727=>"000000111",
  44728=>"010000110",
  44729=>"011011110",
  44730=>"001100001",
  44731=>"000101000",
  44732=>"111010100",
  44733=>"001101000",
  44734=>"111010110",
  44735=>"001011001",
  44736=>"011000000",
  44737=>"100100001",
  44738=>"100001110",
  44739=>"011101100",
  44740=>"000000111",
  44741=>"100110000",
  44742=>"000000000",
  44743=>"100111101",
  44744=>"111110000",
  44745=>"010100001",
  44746=>"011001111",
  44747=>"111011010",
  44748=>"011001011",
  44749=>"110000001",
  44750=>"001110100",
  44751=>"001111011",
  44752=>"001110000",
  44753=>"101100001",
  44754=>"011010001",
  44755=>"101101001",
  44756=>"101100011",
  44757=>"011001010",
  44758=>"010111110",
  44759=>"010000011",
  44760=>"000001001",
  44761=>"111010000",
  44762=>"001000111",
  44763=>"001110010",
  44764=>"111100010",
  44765=>"111011110",
  44766=>"000010111",
  44767=>"011010001",
  44768=>"110010110",
  44769=>"101010111",
  44770=>"110111011",
  44771=>"111111111",
  44772=>"101111101",
  44773=>"101100110",
  44774=>"111100111",
  44775=>"111100110",
  44776=>"110111001",
  44777=>"111000101",
  44778=>"100101100",
  44779=>"101111101",
  44780=>"000100101",
  44781=>"001101011",
  44782=>"010010000",
  44783=>"001010101",
  44784=>"011101101",
  44785=>"000000111",
  44786=>"011100001",
  44787=>"011001000",
  44788=>"110001110",
  44789=>"111010000",
  44790=>"010010111",
  44791=>"111101100",
  44792=>"011011001",
  44793=>"100011011",
  44794=>"010101101",
  44795=>"010000001",
  44796=>"101100101",
  44797=>"111000101",
  44798=>"111001110",
  44799=>"010011001",
  44800=>"000010001",
  44801=>"111001101",
  44802=>"111110000",
  44803=>"100110000",
  44804=>"101011001",
  44805=>"111110000",
  44806=>"000010111",
  44807=>"111010111",
  44808=>"001111110",
  44809=>"010001001",
  44810=>"111010011",
  44811=>"111111111",
  44812=>"100010000",
  44813=>"011101011",
  44814=>"011010001",
  44815=>"000100001",
  44816=>"110010001",
  44817=>"110000100",
  44818=>"111110010",
  44819=>"001110110",
  44820=>"001001001",
  44821=>"110111001",
  44822=>"111010110",
  44823=>"000011001",
  44824=>"111101100",
  44825=>"011100010",
  44826=>"000101111",
  44827=>"000110110",
  44828=>"110001111",
  44829=>"010011100",
  44830=>"111101101",
  44831=>"000000111",
  44832=>"000010101",
  44833=>"000000010",
  44834=>"111101000",
  44835=>"111100101",
  44836=>"001001010",
  44837=>"000101010",
  44838=>"101100110",
  44839=>"011110101",
  44840=>"111111111",
  44841=>"110011110",
  44842=>"011111010",
  44843=>"111100010",
  44844=>"011001011",
  44845=>"010011001",
  44846=>"111110100",
  44847=>"100011110",
  44848=>"001010110",
  44849=>"101011010",
  44850=>"000100000",
  44851=>"100110101",
  44852=>"011001010",
  44853=>"101110110",
  44854=>"110110010",
  44855=>"110011100",
  44856=>"100111110",
  44857=>"101101100",
  44858=>"010011000",
  44859=>"011001000",
  44860=>"111001110",
  44861=>"010011000",
  44862=>"111001110",
  44863=>"000101101",
  44864=>"101111001",
  44865=>"101000001",
  44866=>"101111111",
  44867=>"010110111",
  44868=>"001100100",
  44869=>"101000001",
  44870=>"111100101",
  44871=>"110011010",
  44872=>"011000010",
  44873=>"011011100",
  44874=>"010011000",
  44875=>"000001001",
  44876=>"001100011",
  44877=>"110110101",
  44878=>"110010101",
  44879=>"001010101",
  44880=>"111000000",
  44881=>"100101111",
  44882=>"110101000",
  44883=>"101000111",
  44884=>"000010101",
  44885=>"100101110",
  44886=>"000100011",
  44887=>"001011001",
  44888=>"010110111",
  44889=>"000111011",
  44890=>"101011000",
  44891=>"110010001",
  44892=>"100111001",
  44893=>"010001011",
  44894=>"111110111",
  44895=>"000001001",
  44896=>"000010111",
  44897=>"100001100",
  44898=>"110111101",
  44899=>"011101000",
  44900=>"101100001",
  44901=>"010111111",
  44902=>"111001110",
  44903=>"001110000",
  44904=>"110010000",
  44905=>"100010010",
  44906=>"110100111",
  44907=>"100100111",
  44908=>"101101011",
  44909=>"111111101",
  44910=>"110101011",
  44911=>"010010100",
  44912=>"010010110",
  44913=>"100001000",
  44914=>"101010010",
  44915=>"101100100",
  44916=>"011000111",
  44917=>"101111000",
  44918=>"000000000",
  44919=>"100101111",
  44920=>"111001001",
  44921=>"110110100",
  44922=>"111001011",
  44923=>"001100011",
  44924=>"011000101",
  44925=>"001100001",
  44926=>"100001000",
  44927=>"011001101",
  44928=>"000100110",
  44929=>"010111000",
  44930=>"110100111",
  44931=>"001001001",
  44932=>"010100011",
  44933=>"101101001",
  44934=>"101101110",
  44935=>"111100000",
  44936=>"000111111",
  44937=>"000111000",
  44938=>"000110011",
  44939=>"010110110",
  44940=>"000110000",
  44941=>"010000010",
  44942=>"101101111",
  44943=>"000101000",
  44944=>"101011010",
  44945=>"010110011",
  44946=>"001100101",
  44947=>"111100100",
  44948=>"101111100",
  44949=>"011010011",
  44950=>"100111110",
  44951=>"110001101",
  44952=>"111100100",
  44953=>"010000000",
  44954=>"000000101",
  44955=>"101111101",
  44956=>"010000111",
  44957=>"101100000",
  44958=>"101011010",
  44959=>"001100001",
  44960=>"000110010",
  44961=>"001110000",
  44962=>"110010101",
  44963=>"000100100",
  44964=>"111011010",
  44965=>"011111101",
  44966=>"000101010",
  44967=>"010001011",
  44968=>"010110110",
  44969=>"011011111",
  44970=>"011010111",
  44971=>"000100000",
  44972=>"011100000",
  44973=>"111111000",
  44974=>"111111110",
  44975=>"110101100",
  44976=>"000000001",
  44977=>"010011010",
  44978=>"100001000",
  44979=>"000000111",
  44980=>"010010001",
  44981=>"001100101",
  44982=>"000010100",
  44983=>"111001111",
  44984=>"101001100",
  44985=>"010111110",
  44986=>"101000000",
  44987=>"000110001",
  44988=>"101101001",
  44989=>"111011001",
  44990=>"111101101",
  44991=>"010000100",
  44992=>"101100110",
  44993=>"110111000",
  44994=>"000110010",
  44995=>"111101111",
  44996=>"100110010",
  44997=>"010111010",
  44998=>"010101000",
  44999=>"101001001",
  45000=>"000011001",
  45001=>"011111101",
  45002=>"111100110",
  45003=>"011101110",
  45004=>"001011100",
  45005=>"100111011",
  45006=>"011100010",
  45007=>"100001010",
  45008=>"100000100",
  45009=>"101111111",
  45010=>"000100001",
  45011=>"100000000",
  45012=>"110111000",
  45013=>"011100000",
  45014=>"001000101",
  45015=>"111110010",
  45016=>"101100101",
  45017=>"101010110",
  45018=>"000100011",
  45019=>"010011011",
  45020=>"100011100",
  45021=>"110010111",
  45022=>"101101110",
  45023=>"011000011",
  45024=>"110111011",
  45025=>"100001001",
  45026=>"011101100",
  45027=>"111100110",
  45028=>"100000000",
  45029=>"110000110",
  45030=>"000000011",
  45031=>"110001001",
  45032=>"000011101",
  45033=>"001010001",
  45034=>"101000101",
  45035=>"110101111",
  45036=>"101000011",
  45037=>"111001110",
  45038=>"011101111",
  45039=>"111111010",
  45040=>"011101111",
  45041=>"000010000",
  45042=>"000110000",
  45043=>"000001001",
  45044=>"111010001",
  45045=>"010100011",
  45046=>"101100111",
  45047=>"100101010",
  45048=>"001011011",
  45049=>"011100000",
  45050=>"111111111",
  45051=>"000111110",
  45052=>"100000001",
  45053=>"111111100",
  45054=>"011100011",
  45055=>"110101110",
  45056=>"100011011",
  45057=>"000000000",
  45058=>"010111000",
  45059=>"110010001",
  45060=>"011111100",
  45061=>"101000011",
  45062=>"000100101",
  45063=>"101100001",
  45064=>"000100110",
  45065=>"111101011",
  45066=>"011100101",
  45067=>"010001001",
  45068=>"010010011",
  45069=>"010111110",
  45070=>"011111101",
  45071=>"000111001",
  45072=>"000101100",
  45073=>"100101011",
  45074=>"111100001",
  45075=>"100000101",
  45076=>"010100100",
  45077=>"101000000",
  45078=>"000011000",
  45079=>"100101110",
  45080=>"010101011",
  45081=>"101001011",
  45082=>"001001011",
  45083=>"001010111",
  45084=>"011001100",
  45085=>"110110010",
  45086=>"100001011",
  45087=>"001001001",
  45088=>"000100110",
  45089=>"101011100",
  45090=>"000110101",
  45091=>"011000010",
  45092=>"100110000",
  45093=>"010001111",
  45094=>"000110110",
  45095=>"101011001",
  45096=>"111101011",
  45097=>"011110011",
  45098=>"011011010",
  45099=>"110000000",
  45100=>"000001111",
  45101=>"001000111",
  45102=>"010000111",
  45103=>"101001111",
  45104=>"111011110",
  45105=>"111111100",
  45106=>"011100010",
  45107=>"100110110",
  45108=>"110101100",
  45109=>"100000001",
  45110=>"001100111",
  45111=>"011000100",
  45112=>"010100011",
  45113=>"001000100",
  45114=>"110101110",
  45115=>"010000011",
  45116=>"100000011",
  45117=>"100101010",
  45118=>"100001000",
  45119=>"010110001",
  45120=>"100100111",
  45121=>"110011000",
  45122=>"011011010",
  45123=>"001000100",
  45124=>"011011111",
  45125=>"001011111",
  45126=>"100011111",
  45127=>"110011111",
  45128=>"101010000",
  45129=>"110010111",
  45130=>"011010011",
  45131=>"011100110",
  45132=>"110010111",
  45133=>"111111000",
  45134=>"101101101",
  45135=>"101111100",
  45136=>"110111101",
  45137=>"011101100",
  45138=>"001001110",
  45139=>"000101100",
  45140=>"101000001",
  45141=>"011000000",
  45142=>"110001010",
  45143=>"010101000",
  45144=>"110110101",
  45145=>"111001001",
  45146=>"111001100",
  45147=>"001100001",
  45148=>"001100000",
  45149=>"011011100",
  45150=>"100010011",
  45151=>"111100101",
  45152=>"111100001",
  45153=>"000111001",
  45154=>"110011010",
  45155=>"000010110",
  45156=>"001111001",
  45157=>"110000000",
  45158=>"000010000",
  45159=>"100000101",
  45160=>"100011011",
  45161=>"100001001",
  45162=>"111001110",
  45163=>"100110101",
  45164=>"111100110",
  45165=>"000000110",
  45166=>"101100110",
  45167=>"010011101",
  45168=>"010100000",
  45169=>"101100110",
  45170=>"110111010",
  45171=>"111110101",
  45172=>"000110001",
  45173=>"011110110",
  45174=>"111001100",
  45175=>"110101110",
  45176=>"010100110",
  45177=>"110100101",
  45178=>"000000110",
  45179=>"001011111",
  45180=>"000000111",
  45181=>"110010100",
  45182=>"000100011",
  45183=>"111111001",
  45184=>"101010000",
  45185=>"111001000",
  45186=>"111011101",
  45187=>"101000101",
  45188=>"010010111",
  45189=>"111100111",
  45190=>"011100111",
  45191=>"101101000",
  45192=>"000111110",
  45193=>"100111000",
  45194=>"100000101",
  45195=>"101110101",
  45196=>"100010001",
  45197=>"010010111",
  45198=>"000001000",
  45199=>"100010101",
  45200=>"010011100",
  45201=>"111010100",
  45202=>"101010010",
  45203=>"001000001",
  45204=>"111001101",
  45205=>"100000101",
  45206=>"011111110",
  45207=>"111110011",
  45208=>"010111011",
  45209=>"101010111",
  45210=>"111011101",
  45211=>"011100101",
  45212=>"001110101",
  45213=>"101000000",
  45214=>"000100000",
  45215=>"101001001",
  45216=>"010101000",
  45217=>"010001001",
  45218=>"111000110",
  45219=>"111101000",
  45220=>"001011011",
  45221=>"000101100",
  45222=>"100000001",
  45223=>"100100101",
  45224=>"011011110",
  45225=>"110111100",
  45226=>"100000111",
  45227=>"110100001",
  45228=>"011001100",
  45229=>"111100100",
  45230=>"000101011",
  45231=>"000001110",
  45232=>"101000011",
  45233=>"001010010",
  45234=>"110100101",
  45235=>"100011100",
  45236=>"101000000",
  45237=>"110111100",
  45238=>"010100010",
  45239=>"000000011",
  45240=>"100111100",
  45241=>"100100001",
  45242=>"010011100",
  45243=>"000110110",
  45244=>"011111100",
  45245=>"101110000",
  45246=>"010011111",
  45247=>"000110001",
  45248=>"001010110",
  45249=>"110100001",
  45250=>"101010101",
  45251=>"100000100",
  45252=>"001101011",
  45253=>"011011111",
  45254=>"111100010",
  45255=>"101110110",
  45256=>"000010011",
  45257=>"001100101",
  45258=>"100010110",
  45259=>"001010000",
  45260=>"001110101",
  45261=>"101110011",
  45262=>"010110100",
  45263=>"000111111",
  45264=>"100100011",
  45265=>"111011110",
  45266=>"000011110",
  45267=>"111011001",
  45268=>"011001110",
  45269=>"011110100",
  45270=>"010010110",
  45271=>"101111110",
  45272=>"000011000",
  45273=>"101101110",
  45274=>"000100101",
  45275=>"000110101",
  45276=>"100011101",
  45277=>"101110100",
  45278=>"010101011",
  45279=>"011001011",
  45280=>"111100001",
  45281=>"011010001",
  45282=>"010100111",
  45283=>"100000000",
  45284=>"011100110",
  45285=>"101001101",
  45286=>"110110000",
  45287=>"000001100",
  45288=>"001111010",
  45289=>"110111101",
  45290=>"111100101",
  45291=>"100101010",
  45292=>"000011100",
  45293=>"101000000",
  45294=>"111001011",
  45295=>"101111000",
  45296=>"010101011",
  45297=>"101101110",
  45298=>"111000111",
  45299=>"011011100",
  45300=>"100000011",
  45301=>"110010111",
  45302=>"001100111",
  45303=>"110100001",
  45304=>"000000101",
  45305=>"000111000",
  45306=>"101110110",
  45307=>"000111001",
  45308=>"000100111",
  45309=>"001000010",
  45310=>"000110101",
  45311=>"001001000",
  45312=>"110010001",
  45313=>"100101110",
  45314=>"110101111",
  45315=>"110111111",
  45316=>"001110101",
  45317=>"101100111",
  45318=>"000000010",
  45319=>"110010010",
  45320=>"111011111",
  45321=>"001110010",
  45322=>"110110001",
  45323=>"101111001",
  45324=>"111110011",
  45325=>"101010010",
  45326=>"010001111",
  45327=>"111111011",
  45328=>"011011010",
  45329=>"100101010",
  45330=>"011111100",
  45331=>"101111010",
  45332=>"111110111",
  45333=>"100000000",
  45334=>"101011100",
  45335=>"000000011",
  45336=>"011101011",
  45337=>"101101001",
  45338=>"011010001",
  45339=>"010000100",
  45340=>"110100010",
  45341=>"001100110",
  45342=>"111100010",
  45343=>"000100110",
  45344=>"011101010",
  45345=>"001001111",
  45346=>"000001101",
  45347=>"011001011",
  45348=>"000001111",
  45349=>"011011000",
  45350=>"100100000",
  45351=>"100010011",
  45352=>"011100110",
  45353=>"010010101",
  45354=>"011100110",
  45355=>"111011001",
  45356=>"111100001",
  45357=>"110001010",
  45358=>"110100111",
  45359=>"011010101",
  45360=>"010001000",
  45361=>"010000010",
  45362=>"100111010",
  45363=>"111010010",
  45364=>"000001001",
  45365=>"011110101",
  45366=>"101010100",
  45367=>"100110011",
  45368=>"001101000",
  45369=>"100101001",
  45370=>"101001000",
  45371=>"000100101",
  45372=>"000110010",
  45373=>"111110000",
  45374=>"010001010",
  45375=>"111101001",
  45376=>"100101110",
  45377=>"011111001",
  45378=>"011010011",
  45379=>"101010110",
  45380=>"001111001",
  45381=>"011101111",
  45382=>"100110101",
  45383=>"110001001",
  45384=>"101101100",
  45385=>"010010000",
  45386=>"100110000",
  45387=>"001101010",
  45388=>"000011010",
  45389=>"101101111",
  45390=>"111010110",
  45391=>"100100011",
  45392=>"101010100",
  45393=>"001101101",
  45394=>"100010111",
  45395=>"111011010",
  45396=>"111111000",
  45397=>"110110111",
  45398=>"101100011",
  45399=>"001111000",
  45400=>"000000111",
  45401=>"101110000",
  45402=>"110111000",
  45403=>"011000011",
  45404=>"011011011",
  45405=>"000110111",
  45406=>"010110101",
  45407=>"101110000",
  45408=>"101101011",
  45409=>"010000101",
  45410=>"110110001",
  45411=>"000000001",
  45412=>"101100101",
  45413=>"010100101",
  45414=>"010001001",
  45415=>"010010100",
  45416=>"101000100",
  45417=>"001101111",
  45418=>"111111101",
  45419=>"010111011",
  45420=>"110111010",
  45421=>"110101101",
  45422=>"011000001",
  45423=>"111011010",
  45424=>"010001101",
  45425=>"100100101",
  45426=>"010000111",
  45427=>"000000101",
  45428=>"100101111",
  45429=>"100001101",
  45430=>"101011001",
  45431=>"100111101",
  45432=>"000111100",
  45433=>"010010110",
  45434=>"010010101",
  45435=>"010010100",
  45436=>"100010011",
  45437=>"111111001",
  45438=>"011001000",
  45439=>"101110101",
  45440=>"000111111",
  45441=>"011001101",
  45442=>"111111100",
  45443=>"111001111",
  45444=>"111010110",
  45445=>"011001100",
  45446=>"100000110",
  45447=>"100011100",
  45448=>"100011111",
  45449=>"110101001",
  45450=>"001010000",
  45451=>"011111100",
  45452=>"001110010",
  45453=>"111111100",
  45454=>"010110110",
  45455=>"100100001",
  45456=>"100011111",
  45457=>"001110011",
  45458=>"000010011",
  45459=>"011011111",
  45460=>"010011111",
  45461=>"111110101",
  45462=>"000110011",
  45463=>"000110010",
  45464=>"111111100",
  45465=>"110001100",
  45466=>"110111011",
  45467=>"001010101",
  45468=>"011011100",
  45469=>"010101001",
  45470=>"001101011",
  45471=>"011000001",
  45472=>"001010000",
  45473=>"111101000",
  45474=>"000110000",
  45475=>"111111111",
  45476=>"111100010",
  45477=>"101000100",
  45478=>"110001100",
  45479=>"010100000",
  45480=>"010100011",
  45481=>"110101000",
  45482=>"100000100",
  45483=>"111001000",
  45484=>"110001100",
  45485=>"000101010",
  45486=>"011100100",
  45487=>"111100111",
  45488=>"001010000",
  45489=>"110111010",
  45490=>"110000110",
  45491=>"001111101",
  45492=>"001100101",
  45493=>"111100011",
  45494=>"000001001",
  45495=>"010101111",
  45496=>"111100111",
  45497=>"110000101",
  45498=>"110100100",
  45499=>"111110111",
  45500=>"101001111",
  45501=>"010010000",
  45502=>"101111100",
  45503=>"011110100",
  45504=>"100101110",
  45505=>"001110100",
  45506=>"000100101",
  45507=>"110010000",
  45508=>"010111110",
  45509=>"011011100",
  45510=>"101110101",
  45511=>"110010010",
  45512=>"111110101",
  45513=>"110100010",
  45514=>"010010111",
  45515=>"011111011",
  45516=>"001011101",
  45517=>"111010100",
  45518=>"110110100",
  45519=>"011101001",
  45520=>"101101000",
  45521=>"110000110",
  45522=>"000001000",
  45523=>"010111101",
  45524=>"011011111",
  45525=>"101110001",
  45526=>"001000111",
  45527=>"000100111",
  45528=>"001000001",
  45529=>"001101011",
  45530=>"011011110",
  45531=>"001010000",
  45532=>"101001110",
  45533=>"110111000",
  45534=>"000000000",
  45535=>"110000110",
  45536=>"111000000",
  45537=>"001010100",
  45538=>"100000001",
  45539=>"100010000",
  45540=>"100001000",
  45541=>"000001110",
  45542=>"000101000",
  45543=>"010100011",
  45544=>"001100111",
  45545=>"111101000",
  45546=>"100010111",
  45547=>"100101111",
  45548=>"111111001",
  45549=>"010001100",
  45550=>"100000011",
  45551=>"001100111",
  45552=>"100010011",
  45553=>"010100111",
  45554=>"000001101",
  45555=>"101110101",
  45556=>"011110010",
  45557=>"000110011",
  45558=>"111101110",
  45559=>"010110110",
  45560=>"101010000",
  45561=>"110011111",
  45562=>"101111000",
  45563=>"000010101",
  45564=>"010011011",
  45565=>"110100111",
  45566=>"100000110",
  45567=>"001001110",
  45568=>"110010000",
  45569=>"110000111",
  45570=>"110010101",
  45571=>"110100001",
  45572=>"001110101",
  45573=>"111000000",
  45574=>"111110010",
  45575=>"010111101",
  45576=>"000110001",
  45577=>"111100011",
  45578=>"010101101",
  45579=>"110010110",
  45580=>"100010010",
  45581=>"010100010",
  45582=>"110100010",
  45583=>"001101001",
  45584=>"010110111",
  45585=>"011110001",
  45586=>"111111111",
  45587=>"110101101",
  45588=>"010100011",
  45589=>"110000100",
  45590=>"001011100",
  45591=>"000000101",
  45592=>"000001000",
  45593=>"101011100",
  45594=>"111000000",
  45595=>"110001001",
  45596=>"010101000",
  45597=>"100000100",
  45598=>"110001111",
  45599=>"101100011",
  45600=>"101010010",
  45601=>"111110100",
  45602=>"011010010",
  45603=>"110000000",
  45604=>"011111000",
  45605=>"100110011",
  45606=>"000110000",
  45607=>"001111100",
  45608=>"000110100",
  45609=>"011000101",
  45610=>"100010100",
  45611=>"101111001",
  45612=>"000101110",
  45613=>"100100100",
  45614=>"000111111",
  45615=>"111001010",
  45616=>"101000110",
  45617=>"011111100",
  45618=>"100110001",
  45619=>"010101111",
  45620=>"011100011",
  45621=>"010100100",
  45622=>"010000101",
  45623=>"101111001",
  45624=>"000011010",
  45625=>"001110011",
  45626=>"000000111",
  45627=>"011100001",
  45628=>"000001110",
  45629=>"010101010",
  45630=>"001010011",
  45631=>"011110111",
  45632=>"100101000",
  45633=>"001010101",
  45634=>"000010000",
  45635=>"100010000",
  45636=>"011000101",
  45637=>"100110010",
  45638=>"000101000",
  45639=>"011111001",
  45640=>"010010011",
  45641=>"101000100",
  45642=>"001111100",
  45643=>"010000010",
  45644=>"001000101",
  45645=>"100011010",
  45646=>"111111101",
  45647=>"100110101",
  45648=>"111010100",
  45649=>"001110010",
  45650=>"000011001",
  45651=>"001101110",
  45652=>"010011000",
  45653=>"100100110",
  45654=>"001000001",
  45655=>"100000110",
  45656=>"111110011",
  45657=>"110100111",
  45658=>"110000111",
  45659=>"000010011",
  45660=>"010101100",
  45661=>"011010001",
  45662=>"010001100",
  45663=>"010111110",
  45664=>"101110100",
  45665=>"000110000",
  45666=>"001100111",
  45667=>"110101000",
  45668=>"101101001",
  45669=>"111111010",
  45670=>"010101000",
  45671=>"000101001",
  45672=>"001010001",
  45673=>"110110110",
  45674=>"101101011",
  45675=>"100010000",
  45676=>"100110111",
  45677=>"111001100",
  45678=>"000010000",
  45679=>"110100010",
  45680=>"010011010",
  45681=>"000011010",
  45682=>"111111101",
  45683=>"001100010",
  45684=>"110010101",
  45685=>"001101010",
  45686=>"111101101",
  45687=>"100000001",
  45688=>"010000110",
  45689=>"000101010",
  45690=>"110000100",
  45691=>"001101001",
  45692=>"001111101",
  45693=>"101101110",
  45694=>"001100010",
  45695=>"000101011",
  45696=>"000101100",
  45697=>"111101111",
  45698=>"100100000",
  45699=>"110111010",
  45700=>"110000100",
  45701=>"010001111",
  45702=>"010110010",
  45703=>"010111101",
  45704=>"111000101",
  45705=>"010101011",
  45706=>"000110100",
  45707=>"010111100",
  45708=>"011100110",
  45709=>"111001010",
  45710=>"101101100",
  45711=>"000110011",
  45712=>"111000101",
  45713=>"011101001",
  45714=>"111001100",
  45715=>"000111110",
  45716=>"011111001",
  45717=>"111111111",
  45718=>"110110110",
  45719=>"100010110",
  45720=>"111111111",
  45721=>"000010001",
  45722=>"111100011",
  45723=>"110110111",
  45724=>"100001110",
  45725=>"011010001",
  45726=>"001001001",
  45727=>"110000100",
  45728=>"111001110",
  45729=>"010100100",
  45730=>"100010101",
  45731=>"001011010",
  45732=>"111101011",
  45733=>"111101100",
  45734=>"101001011",
  45735=>"010000000",
  45736=>"110101000",
  45737=>"101101111",
  45738=>"010101000",
  45739=>"100110101",
  45740=>"011000100",
  45741=>"111001101",
  45742=>"100010000",
  45743=>"101011010",
  45744=>"010000111",
  45745=>"011011011",
  45746=>"100100110",
  45747=>"010010101",
  45748=>"011100001",
  45749=>"011011000",
  45750=>"001111101",
  45751=>"010100010",
  45752=>"101011110",
  45753=>"011011001",
  45754=>"101101101",
  45755=>"101000100",
  45756=>"111111001",
  45757=>"010110001",
  45758=>"100111101",
  45759=>"100011101",
  45760=>"101010100",
  45761=>"010010000",
  45762=>"100101100",
  45763=>"101010101",
  45764=>"010001001",
  45765=>"110000100",
  45766=>"001111010",
  45767=>"010000000",
  45768=>"011010001",
  45769=>"101011101",
  45770=>"101100010",
  45771=>"100000000",
  45772=>"011101000",
  45773=>"000011010",
  45774=>"000100011",
  45775=>"110111000",
  45776=>"101001000",
  45777=>"010001001",
  45778=>"100011001",
  45779=>"110110101",
  45780=>"000010111",
  45781=>"001010101",
  45782=>"011001010",
  45783=>"000011010",
  45784=>"100011010",
  45785=>"001000011",
  45786=>"010001011",
  45787=>"100100001",
  45788=>"111101010",
  45789=>"110001100",
  45790=>"110001101",
  45791=>"110110101",
  45792=>"000100000",
  45793=>"001101000",
  45794=>"100011110",
  45795=>"101001101",
  45796=>"110001101",
  45797=>"110100010",
  45798=>"001000111",
  45799=>"100110001",
  45800=>"010111101",
  45801=>"011001010",
  45802=>"011010000",
  45803=>"110010011",
  45804=>"100101010",
  45805=>"010000011",
  45806=>"110100001",
  45807=>"011010111",
  45808=>"011001111",
  45809=>"100110010",
  45810=>"011001101",
  45811=>"010111001",
  45812=>"011111011",
  45813=>"011001111",
  45814=>"011110110",
  45815=>"000000001",
  45816=>"100101011",
  45817=>"101100110",
  45818=>"000011101",
  45819=>"101100010",
  45820=>"101000010",
  45821=>"100001011",
  45822=>"101110100",
  45823=>"010101111",
  45824=>"110001000",
  45825=>"111011000",
  45826=>"011100001",
  45827=>"110001110",
  45828=>"110101011",
  45829=>"011101110",
  45830=>"100010011",
  45831=>"011100111",
  45832=>"101000011",
  45833=>"001001100",
  45834=>"110101010",
  45835=>"001011100",
  45836=>"100000111",
  45837=>"001101111",
  45838=>"110100110",
  45839=>"000011010",
  45840=>"110010000",
  45841=>"001111001",
  45842=>"110101100",
  45843=>"011110100",
  45844=>"100011010",
  45845=>"111101000",
  45846=>"100011001",
  45847=>"011001110",
  45848=>"000110100",
  45849=>"001000101",
  45850=>"101111101",
  45851=>"101100101",
  45852=>"010001110",
  45853=>"011011010",
  45854=>"111110010",
  45855=>"100010010",
  45856=>"000111110",
  45857=>"011110000",
  45858=>"001100100",
  45859=>"011000100",
  45860=>"111101001",
  45861=>"001000010",
  45862=>"111111010",
  45863=>"000110000",
  45864=>"001100111",
  45865=>"001101101",
  45866=>"101110001",
  45867=>"111001100",
  45868=>"011100111",
  45869=>"000101101",
  45870=>"101001100",
  45871=>"100001001",
  45872=>"110110100",
  45873=>"101111101",
  45874=>"000111101",
  45875=>"011011011",
  45876=>"010100000",
  45877=>"100010000",
  45878=>"000010001",
  45879=>"101010111",
  45880=>"111111011",
  45881=>"011110101",
  45882=>"011000011",
  45883=>"000101000",
  45884=>"000110110",
  45885=>"111110111",
  45886=>"111111101",
  45887=>"101010101",
  45888=>"010010001",
  45889=>"010011100",
  45890=>"001010001",
  45891=>"010110001",
  45892=>"000010111",
  45893=>"100010101",
  45894=>"100111101",
  45895=>"100110110",
  45896=>"110101100",
  45897=>"101111100",
  45898=>"101001111",
  45899=>"011101110",
  45900=>"110010100",
  45901=>"001111000",
  45902=>"001100011",
  45903=>"111010101",
  45904=>"010010010",
  45905=>"011011011",
  45906=>"001100010",
  45907=>"010011111",
  45908=>"010001001",
  45909=>"110110001",
  45910=>"111100100",
  45911=>"101000001",
  45912=>"011110000",
  45913=>"111110000",
  45914=>"001011111",
  45915=>"000100101",
  45916=>"000010101",
  45917=>"110010101",
  45918=>"101111100",
  45919=>"110100101",
  45920=>"100101101",
  45921=>"101111100",
  45922=>"100101011",
  45923=>"110110100",
  45924=>"110011011",
  45925=>"100000001",
  45926=>"111100101",
  45927=>"001011011",
  45928=>"110011101",
  45929=>"001100011",
  45930=>"001011001",
  45931=>"101001111",
  45932=>"011010011",
  45933=>"100101000",
  45934=>"010001110",
  45935=>"000111100",
  45936=>"101000110",
  45937=>"001010110",
  45938=>"010101110",
  45939=>"001100010",
  45940=>"100001110",
  45941=>"000000000",
  45942=>"001110011",
  45943=>"101100011",
  45944=>"110001011",
  45945=>"000010001",
  45946=>"001010100",
  45947=>"110101101",
  45948=>"011000000",
  45949=>"011011110",
  45950=>"111010101",
  45951=>"001011100",
  45952=>"011010010",
  45953=>"110010111",
  45954=>"000100010",
  45955=>"000111001",
  45956=>"101000010",
  45957=>"001010101",
  45958=>"001110111",
  45959=>"100000101",
  45960=>"010001010",
  45961=>"001000011",
  45962=>"000011011",
  45963=>"110011011",
  45964=>"100010111",
  45965=>"101101101",
  45966=>"011001010",
  45967=>"000000001",
  45968=>"101101000",
  45969=>"011110110",
  45970=>"010111110",
  45971=>"001101100",
  45972=>"110110011",
  45973=>"111111000",
  45974=>"010011010",
  45975=>"010001101",
  45976=>"110101101",
  45977=>"001110000",
  45978=>"001001010",
  45979=>"011101000",
  45980=>"010101001",
  45981=>"111111110",
  45982=>"001000100",
  45983=>"000010010",
  45984=>"011100000",
  45985=>"111110000",
  45986=>"111110000",
  45987=>"100010001",
  45988=>"000001101",
  45989=>"101001111",
  45990=>"001000111",
  45991=>"010001011",
  45992=>"101010000",
  45993=>"110011100",
  45994=>"100100110",
  45995=>"100010010",
  45996=>"000010000",
  45997=>"010010111",
  45998=>"000111100",
  45999=>"010100001",
  46000=>"111111001",
  46001=>"110101010",
  46002=>"101100001",
  46003=>"000011111",
  46004=>"111011001",
  46005=>"100000100",
  46006=>"000001001",
  46007=>"100000001",
  46008=>"010101011",
  46009=>"101011010",
  46010=>"101011100",
  46011=>"110100111",
  46012=>"100100101",
  46013=>"001111101",
  46014=>"110000100",
  46015=>"010100000",
  46016=>"011100011",
  46017=>"001100111",
  46018=>"001011010",
  46019=>"100110000",
  46020=>"110010100",
  46021=>"000101111",
  46022=>"110110000",
  46023=>"110111110",
  46024=>"000101000",
  46025=>"011111110",
  46026=>"001000101",
  46027=>"000000100",
  46028=>"100100110",
  46029=>"011001110",
  46030=>"100000111",
  46031=>"111010100",
  46032=>"110010110",
  46033=>"011101010",
  46034=>"101001000",
  46035=>"010111111",
  46036=>"011000111",
  46037=>"101010000",
  46038=>"101110000",
  46039=>"010111000",
  46040=>"111010011",
  46041=>"010111111",
  46042=>"011011101",
  46043=>"011111101",
  46044=>"101111110",
  46045=>"101001010",
  46046=>"101111111",
  46047=>"001011101",
  46048=>"000010010",
  46049=>"110010100",
  46050=>"101001110",
  46051=>"101101110",
  46052=>"100010011",
  46053=>"110100001",
  46054=>"100001111",
  46055=>"001101100",
  46056=>"000000010",
  46057=>"101110000",
  46058=>"110100000",
  46059=>"001100000",
  46060=>"011101101",
  46061=>"100011010",
  46062=>"110100010",
  46063=>"010110111",
  46064=>"011011011",
  46065=>"010101110",
  46066=>"001001001",
  46067=>"100011100",
  46068=>"111001011",
  46069=>"011010001",
  46070=>"111100100",
  46071=>"101011011",
  46072=>"111110110",
  46073=>"000110110",
  46074=>"110100101",
  46075=>"111110011",
  46076=>"000000100",
  46077=>"100110011",
  46078=>"110111000",
  46079=>"000011000",
  46080=>"111101101",
  46081=>"100001011",
  46082=>"000011101",
  46083=>"100111101",
  46084=>"011011001",
  46085=>"010111101",
  46086=>"010001001",
  46087=>"111001000",
  46088=>"101110110",
  46089=>"001110101",
  46090=>"100011000",
  46091=>"110000001",
  46092=>"010001011",
  46093=>"011100000",
  46094=>"000001110",
  46095=>"010000111",
  46096=>"101001001",
  46097=>"000000010",
  46098=>"000110001",
  46099=>"000010000",
  46100=>"100110011",
  46101=>"000110111",
  46102=>"011100110",
  46103=>"110000011",
  46104=>"110101110",
  46105=>"011110100",
  46106=>"001010011",
  46107=>"101111101",
  46108=>"000101000",
  46109=>"101001101",
  46110=>"110000100",
  46111=>"101011101",
  46112=>"010100000",
  46113=>"001111111",
  46114=>"001101011",
  46115=>"101100001",
  46116=>"110010101",
  46117=>"001101000",
  46118=>"001010111",
  46119=>"011000000",
  46120=>"100110001",
  46121=>"010001000",
  46122=>"101010010",
  46123=>"001010101",
  46124=>"001110111",
  46125=>"101101010",
  46126=>"110000011",
  46127=>"001110111",
  46128=>"101011110",
  46129=>"101111101",
  46130=>"011100101",
  46131=>"110111010",
  46132=>"011000001",
  46133=>"000100100",
  46134=>"111111100",
  46135=>"100110011",
  46136=>"001000101",
  46137=>"011111000",
  46138=>"111101011",
  46139=>"000110101",
  46140=>"000000111",
  46141=>"110011110",
  46142=>"111001001",
  46143=>"101101100",
  46144=>"001101001",
  46145=>"100110101",
  46146=>"101001001",
  46147=>"000000000",
  46148=>"101001100",
  46149=>"110010111",
  46150=>"011011100",
  46151=>"000001000",
  46152=>"000111000",
  46153=>"001111001",
  46154=>"010110000",
  46155=>"011001101",
  46156=>"001000001",
  46157=>"000011011",
  46158=>"110111001",
  46159=>"101100111",
  46160=>"101101111",
  46161=>"111100110",
  46162=>"100001110",
  46163=>"101100101",
  46164=>"000101110",
  46165=>"001010010",
  46166=>"110111101",
  46167=>"110000010",
  46168=>"011110110",
  46169=>"110101101",
  46170=>"001011000",
  46171=>"110001111",
  46172=>"011100101",
  46173=>"000011000",
  46174=>"111001001",
  46175=>"001001110",
  46176=>"001001001",
  46177=>"101000000",
  46178=>"110011010",
  46179=>"101010101",
  46180=>"101001011",
  46181=>"000010111",
  46182=>"001101000",
  46183=>"000001010",
  46184=>"111111101",
  46185=>"001011101",
  46186=>"000010101",
  46187=>"000100001",
  46188=>"010100001",
  46189=>"011110010",
  46190=>"100011101",
  46191=>"111101010",
  46192=>"101011111",
  46193=>"110101010",
  46194=>"111001111",
  46195=>"111010001",
  46196=>"101001001",
  46197=>"101010011",
  46198=>"110000010",
  46199=>"111110110",
  46200=>"000001000",
  46201=>"000100010",
  46202=>"010101111",
  46203=>"010101011",
  46204=>"110000000",
  46205=>"001111111",
  46206=>"101010111",
  46207=>"010111110",
  46208=>"000101000",
  46209=>"000111111",
  46210=>"100010011",
  46211=>"111010100",
  46212=>"010010101",
  46213=>"111110001",
  46214=>"101010101",
  46215=>"110110101",
  46216=>"110110110",
  46217=>"100111001",
  46218=>"011000110",
  46219=>"100000101",
  46220=>"001011010",
  46221=>"000110011",
  46222=>"101110000",
  46223=>"001101111",
  46224=>"111111011",
  46225=>"110011100",
  46226=>"100110011",
  46227=>"000001100",
  46228=>"111000010",
  46229=>"111111100",
  46230=>"111100000",
  46231=>"101011000",
  46232=>"100001111",
  46233=>"001001111",
  46234=>"101010000",
  46235=>"010000111",
  46236=>"001010010",
  46237=>"110010000",
  46238=>"001111100",
  46239=>"011101001",
  46240=>"101000111",
  46241=>"000111100",
  46242=>"111110011",
  46243=>"011100111",
  46244=>"110100000",
  46245=>"000110000",
  46246=>"000111011",
  46247=>"101001101",
  46248=>"000010111",
  46249=>"001110111",
  46250=>"001011001",
  46251=>"111000011",
  46252=>"111111000",
  46253=>"101100011",
  46254=>"110100110",
  46255=>"101100111",
  46256=>"000110111",
  46257=>"010110011",
  46258=>"010010100",
  46259=>"000110000",
  46260=>"111001000",
  46261=>"111110111",
  46262=>"010110010",
  46263=>"001010111",
  46264=>"111000111",
  46265=>"011001000",
  46266=>"101011110",
  46267=>"111001011",
  46268=>"001010011",
  46269=>"101000101",
  46270=>"010011110",
  46271=>"011000111",
  46272=>"000011000",
  46273=>"010110011",
  46274=>"111110100",
  46275=>"011100000",
  46276=>"100110111",
  46277=>"111110000",
  46278=>"100011000",
  46279=>"001110010",
  46280=>"001111100",
  46281=>"101100000",
  46282=>"011001111",
  46283=>"110100100",
  46284=>"010101001",
  46285=>"000101010",
  46286=>"101101101",
  46287=>"111100011",
  46288=>"100111011",
  46289=>"010011011",
  46290=>"101001011",
  46291=>"010010000",
  46292=>"111111001",
  46293=>"000011101",
  46294=>"101010101",
  46295=>"011110110",
  46296=>"010000101",
  46297=>"100110000",
  46298=>"111100011",
  46299=>"000010011",
  46300=>"011001010",
  46301=>"100010100",
  46302=>"001001010",
  46303=>"010001010",
  46304=>"100000011",
  46305=>"101100111",
  46306=>"000100010",
  46307=>"010010011",
  46308=>"000110111",
  46309=>"000100000",
  46310=>"000101000",
  46311=>"110010010",
  46312=>"111101110",
  46313=>"000111101",
  46314=>"000111111",
  46315=>"000000111",
  46316=>"110111110",
  46317=>"110001000",
  46318=>"011101111",
  46319=>"100011111",
  46320=>"011001110",
  46321=>"010000110",
  46322=>"001011101",
  46323=>"111010001",
  46324=>"010011001",
  46325=>"101110110",
  46326=>"000010000",
  46327=>"100001110",
  46328=>"101111010",
  46329=>"100111111",
  46330=>"011010001",
  46331=>"110000010",
  46332=>"000011111",
  46333=>"111111111",
  46334=>"110110100",
  46335=>"010111101",
  46336=>"010101001",
  46337=>"010110000",
  46338=>"001100001",
  46339=>"111111001",
  46340=>"001111111",
  46341=>"111010111",
  46342=>"101101100",
  46343=>"000001011",
  46344=>"000111111",
  46345=>"100011111",
  46346=>"000010000",
  46347=>"011110010",
  46348=>"100110000",
  46349=>"011010000",
  46350=>"000111001",
  46351=>"110100100",
  46352=>"010010000",
  46353=>"100101000",
  46354=>"001000010",
  46355=>"111011001",
  46356=>"111101000",
  46357=>"100011010",
  46358=>"000001100",
  46359=>"000001100",
  46360=>"100011111",
  46361=>"010111111",
  46362=>"011100001",
  46363=>"001111111",
  46364=>"101001100",
  46365=>"000011011",
  46366=>"110100011",
  46367=>"011101010",
  46368=>"011011000",
  46369=>"101101010",
  46370=>"001000001",
  46371=>"111010010",
  46372=>"000101100",
  46373=>"001110010",
  46374=>"100100001",
  46375=>"011000110",
  46376=>"000110000",
  46377=>"110010110",
  46378=>"111101101",
  46379=>"101111001",
  46380=>"110101011",
  46381=>"110100000",
  46382=>"011000001",
  46383=>"110001001",
  46384=>"100011101",
  46385=>"111001101",
  46386=>"010111100",
  46387=>"101001111",
  46388=>"000011110",
  46389=>"000101101",
  46390=>"101111000",
  46391=>"111110101",
  46392=>"000111100",
  46393=>"111001101",
  46394=>"001001011",
  46395=>"001010010",
  46396=>"010100010",
  46397=>"100000001",
  46398=>"101011101",
  46399=>"111111001",
  46400=>"101111100",
  46401=>"000001100",
  46402=>"100011111",
  46403=>"101110010",
  46404=>"110001001",
  46405=>"000111000",
  46406=>"100100010",
  46407=>"001010100",
  46408=>"111011010",
  46409=>"111110101",
  46410=>"000110000",
  46411=>"110100111",
  46412=>"010111101",
  46413=>"101000111",
  46414=>"000110111",
  46415=>"101101000",
  46416=>"011111000",
  46417=>"111101111",
  46418=>"010111111",
  46419=>"011101000",
  46420=>"000000010",
  46421=>"010111110",
  46422=>"111011111",
  46423=>"111100000",
  46424=>"000111101",
  46425=>"001110000",
  46426=>"001001101",
  46427=>"000111100",
  46428=>"010001010",
  46429=>"100101101",
  46430=>"000111000",
  46431=>"101100010",
  46432=>"110110100",
  46433=>"001001100",
  46434=>"100010101",
  46435=>"001101011",
  46436=>"011100000",
  46437=>"010010111",
  46438=>"010000010",
  46439=>"100000000",
  46440=>"011010101",
  46441=>"111100010",
  46442=>"110110001",
  46443=>"001100111",
  46444=>"001101110",
  46445=>"100000101",
  46446=>"101110000",
  46447=>"100101101",
  46448=>"000101101",
  46449=>"100111110",
  46450=>"110011011",
  46451=>"011000100",
  46452=>"011011111",
  46453=>"000110010",
  46454=>"000010101",
  46455=>"001001011",
  46456=>"000110000",
  46457=>"101101101",
  46458=>"000010101",
  46459=>"100001111",
  46460=>"111100010",
  46461=>"111111001",
  46462=>"101010101",
  46463=>"010000000",
  46464=>"111000111",
  46465=>"101101000",
  46466=>"101011111",
  46467=>"100011010",
  46468=>"001110000",
  46469=>"010000110",
  46470=>"010000000",
  46471=>"010010011",
  46472=>"010001000",
  46473=>"111010001",
  46474=>"101100111",
  46475=>"110101010",
  46476=>"111110110",
  46477=>"101011010",
  46478=>"110010110",
  46479=>"111111000",
  46480=>"111111001",
  46481=>"000110100",
  46482=>"111001010",
  46483=>"100110110",
  46484=>"100000101",
  46485=>"011111111",
  46486=>"111111111",
  46487=>"000000111",
  46488=>"111111001",
  46489=>"000000101",
  46490=>"100000110",
  46491=>"001011000",
  46492=>"110010101",
  46493=>"011000010",
  46494=>"101100101",
  46495=>"010110100",
  46496=>"110111010",
  46497=>"100000110",
  46498=>"101111111",
  46499=>"010001000",
  46500=>"011111110",
  46501=>"011010111",
  46502=>"011100111",
  46503=>"100100001",
  46504=>"011000000",
  46505=>"001011001",
  46506=>"100000010",
  46507=>"100001010",
  46508=>"011100001",
  46509=>"010001111",
  46510=>"101111001",
  46511=>"101010010",
  46512=>"001101011",
  46513=>"010001100",
  46514=>"000010100",
  46515=>"000000011",
  46516=>"010100010",
  46517=>"100111101",
  46518=>"101001011",
  46519=>"101101101",
  46520=>"000110000",
  46521=>"000100001",
  46522=>"001001110",
  46523=>"111001011",
  46524=>"010111001",
  46525=>"111001010",
  46526=>"011111000",
  46527=>"111000101",
  46528=>"010101010",
  46529=>"011000011",
  46530=>"010011100",
  46531=>"110110111",
  46532=>"111110100",
  46533=>"010011011",
  46534=>"111101100",
  46535=>"111000110",
  46536=>"000001000",
  46537=>"010101111",
  46538=>"000101110",
  46539=>"110111000",
  46540=>"101110111",
  46541=>"111011111",
  46542=>"001100101",
  46543=>"011100010",
  46544=>"110000111",
  46545=>"110111011",
  46546=>"111101001",
  46547=>"101000001",
  46548=>"101010000",
  46549=>"011001101",
  46550=>"110011111",
  46551=>"010010110",
  46552=>"101111110",
  46553=>"010001001",
  46554=>"100000001",
  46555=>"011010011",
  46556=>"000010110",
  46557=>"101011101",
  46558=>"111011101",
  46559=>"010111000",
  46560=>"000010100",
  46561=>"010000010",
  46562=>"110011001",
  46563=>"010010100",
  46564=>"000110111",
  46565=>"000001010",
  46566=>"001001010",
  46567=>"011001111",
  46568=>"110111111",
  46569=>"100010011",
  46570=>"011000101",
  46571=>"000101011",
  46572=>"010001000",
  46573=>"110101001",
  46574=>"110001001",
  46575=>"000010010",
  46576=>"001110110",
  46577=>"110101111",
  46578=>"000011111",
  46579=>"100010100",
  46580=>"011001011",
  46581=>"000010001",
  46582=>"110011010",
  46583=>"010111101",
  46584=>"000010100",
  46585=>"000000111",
  46586=>"011001001",
  46587=>"001000110",
  46588=>"010111000",
  46589=>"011001110",
  46590=>"011000111",
  46591=>"010011101",
  46592=>"110011010",
  46593=>"000110110",
  46594=>"111010100",
  46595=>"101001001",
  46596=>"000101001",
  46597=>"011111010",
  46598=>"011000110",
  46599=>"101011100",
  46600=>"101010101",
  46601=>"011110101",
  46602=>"111111100",
  46603=>"011100001",
  46604=>"101001001",
  46605=>"011000000",
  46606=>"010101010",
  46607=>"000110101",
  46608=>"001111000",
  46609=>"110110001",
  46610=>"101101001",
  46611=>"111100100",
  46612=>"000101101",
  46613=>"001000100",
  46614=>"100001010",
  46615=>"000011101",
  46616=>"100011010",
  46617=>"000011100",
  46618=>"111110101",
  46619=>"001011000",
  46620=>"001000110",
  46621=>"000001010",
  46622=>"010010000",
  46623=>"010000001",
  46624=>"010100110",
  46625=>"100011001",
  46626=>"101001111",
  46627=>"001111101",
  46628=>"011001010",
  46629=>"001110101",
  46630=>"101101010",
  46631=>"000001110",
  46632=>"110010111",
  46633=>"110000110",
  46634=>"010000111",
  46635=>"101110111",
  46636=>"011000010",
  46637=>"110010001",
  46638=>"011011100",
  46639=>"001000111",
  46640=>"100111111",
  46641=>"010000010",
  46642=>"011001010",
  46643=>"001000001",
  46644=>"001001011",
  46645=>"001101000",
  46646=>"010100101",
  46647=>"111111010",
  46648=>"110100101",
  46649=>"111111011",
  46650=>"001100011",
  46651=>"111111111",
  46652=>"110111100",
  46653=>"001110000",
  46654=>"111110000",
  46655=>"011011011",
  46656=>"111010111",
  46657=>"010001001",
  46658=>"100000110",
  46659=>"000001000",
  46660=>"001001010",
  46661=>"100001100",
  46662=>"010010011",
  46663=>"111001001",
  46664=>"101101011",
  46665=>"011011000",
  46666=>"000100001",
  46667=>"011100100",
  46668=>"000011001",
  46669=>"101010010",
  46670=>"101000000",
  46671=>"110101100",
  46672=>"100000000",
  46673=>"101011100",
  46674=>"010111110",
  46675=>"100001111",
  46676=>"010100000",
  46677=>"000000010",
  46678=>"011010100",
  46679=>"000111010",
  46680=>"111111110",
  46681=>"111110000",
  46682=>"100001111",
  46683=>"010100001",
  46684=>"001110010",
  46685=>"000101100",
  46686=>"001011110",
  46687=>"111101001",
  46688=>"001010111",
  46689=>"100100111",
  46690=>"000100110",
  46691=>"110111000",
  46692=>"111000010",
  46693=>"011010010",
  46694=>"001100000",
  46695=>"000010010",
  46696=>"110001101",
  46697=>"000000101",
  46698=>"011000101",
  46699=>"111011110",
  46700=>"110011111",
  46701=>"011110110",
  46702=>"110110111",
  46703=>"101110101",
  46704=>"001000000",
  46705=>"111000111",
  46706=>"111111001",
  46707=>"000010111",
  46708=>"001000001",
  46709=>"111111110",
  46710=>"101111111",
  46711=>"100111101",
  46712=>"010000010",
  46713=>"011100100",
  46714=>"111010111",
  46715=>"001100001",
  46716=>"101010110",
  46717=>"000000000",
  46718=>"001111111",
  46719=>"010100000",
  46720=>"100111011",
  46721=>"111001110",
  46722=>"111011010",
  46723=>"100111111",
  46724=>"111001111",
  46725=>"001000110",
  46726=>"111111111",
  46727=>"111000101",
  46728=>"000100111",
  46729=>"101001000",
  46730=>"001100100",
  46731=>"011101111",
  46732=>"001101000",
  46733=>"110111011",
  46734=>"001101001",
  46735=>"011010111",
  46736=>"100110100",
  46737=>"111010110",
  46738=>"110000000",
  46739=>"110011100",
  46740=>"001010110",
  46741=>"111011111",
  46742=>"101110100",
  46743=>"001101011",
  46744=>"000000011",
  46745=>"111001001",
  46746=>"111111110",
  46747=>"101011000",
  46748=>"100000101",
  46749=>"110001101",
  46750=>"010101000",
  46751=>"010001011",
  46752=>"000101111",
  46753=>"110000111",
  46754=>"001001111",
  46755=>"101010001",
  46756=>"000011001",
  46757=>"011100111",
  46758=>"010001010",
  46759=>"001100100",
  46760=>"111101101",
  46761=>"100010110",
  46762=>"100000001",
  46763=>"010111000",
  46764=>"111110101",
  46765=>"111011110",
  46766=>"010100011",
  46767=>"101011010",
  46768=>"111100100",
  46769=>"111111111",
  46770=>"011111100",
  46771=>"111010101",
  46772=>"011001001",
  46773=>"001000100",
  46774=>"100010100",
  46775=>"111101110",
  46776=>"001000110",
  46777=>"001100000",
  46778=>"000100011",
  46779=>"010001100",
  46780=>"111101001",
  46781=>"100101000",
  46782=>"110011111",
  46783=>"011011000",
  46784=>"110111010",
  46785=>"011000001",
  46786=>"101111011",
  46787=>"111101100",
  46788=>"010111000",
  46789=>"001000000",
  46790=>"011101000",
  46791=>"101110000",
  46792=>"111010001",
  46793=>"001111110",
  46794=>"000100001",
  46795=>"110111010",
  46796=>"101111110",
  46797=>"001010101",
  46798=>"100101000",
  46799=>"100011010",
  46800=>"110010001",
  46801=>"011110111",
  46802=>"110001101",
  46803=>"101010011",
  46804=>"010111111",
  46805=>"000101010",
  46806=>"101111011",
  46807=>"010000010",
  46808=>"011110100",
  46809=>"100101111",
  46810=>"010010100",
  46811=>"100101010",
  46812=>"010100011",
  46813=>"000110100",
  46814=>"110010011",
  46815=>"101111111",
  46816=>"110010110",
  46817=>"100100000",
  46818=>"111010101",
  46819=>"010100010",
  46820=>"011111001",
  46821=>"010110010",
  46822=>"101111110",
  46823=>"000111110",
  46824=>"011000010",
  46825=>"001100011",
  46826=>"010011011",
  46827=>"000110010",
  46828=>"000100111",
  46829=>"001100010",
  46830=>"111110101",
  46831=>"010001101",
  46832=>"110110011",
  46833=>"010011001",
  46834=>"000000111",
  46835=>"011010000",
  46836=>"100011111",
  46837=>"100000110",
  46838=>"000101010",
  46839=>"101010001",
  46840=>"001111000",
  46841=>"101100111",
  46842=>"000100100",
  46843=>"101001000",
  46844=>"101011111",
  46845=>"011100000",
  46846=>"011101011",
  46847=>"011110010",
  46848=>"111100111",
  46849=>"110000111",
  46850=>"000010000",
  46851=>"001001001",
  46852=>"111010111",
  46853=>"111001100",
  46854=>"000010100",
  46855=>"100110011",
  46856=>"111010101",
  46857=>"110001001",
  46858=>"001010110",
  46859=>"110101010",
  46860=>"110111101",
  46861=>"001101111",
  46862=>"111011010",
  46863=>"101001110",
  46864=>"100111001",
  46865=>"111111110",
  46866=>"011010100",
  46867=>"001010101",
  46868=>"011111101",
  46869=>"110110100",
  46870=>"111101110",
  46871=>"111000000",
  46872=>"000110100",
  46873=>"010011110",
  46874=>"000000110",
  46875=>"011011110",
  46876=>"000010011",
  46877=>"011011010",
  46878=>"010010000",
  46879=>"001000111",
  46880=>"110110000",
  46881=>"011010110",
  46882=>"001101010",
  46883=>"001100010",
  46884=>"100010011",
  46885=>"111101010",
  46886=>"110101011",
  46887=>"100001110",
  46888=>"111110111",
  46889=>"010100110",
  46890=>"000101001",
  46891=>"111010001",
  46892=>"111001000",
  46893=>"010000111",
  46894=>"011111010",
  46895=>"001110110",
  46896=>"101111101",
  46897=>"001101111",
  46898=>"000111110",
  46899=>"010101110",
  46900=>"001001101",
  46901=>"110101001",
  46902=>"111000101",
  46903=>"010011111",
  46904=>"110001100",
  46905=>"110100000",
  46906=>"110010000",
  46907=>"010011001",
  46908=>"010010101",
  46909=>"101001111",
  46910=>"100101101",
  46911=>"111011000",
  46912=>"110101010",
  46913=>"000100111",
  46914=>"010000111",
  46915=>"101101011",
  46916=>"110111011",
  46917=>"001010001",
  46918=>"100111011",
  46919=>"110110010",
  46920=>"101000110",
  46921=>"000110101",
  46922=>"111011110",
  46923=>"110100111",
  46924=>"111111101",
  46925=>"000011100",
  46926=>"011110111",
  46927=>"001000110",
  46928=>"111000000",
  46929=>"000100001",
  46930=>"000001101",
  46931=>"001001011",
  46932=>"000000100",
  46933=>"110100001",
  46934=>"110101001",
  46935=>"011011000",
  46936=>"101100011",
  46937=>"111011001",
  46938=>"111100000",
  46939=>"111001100",
  46940=>"000100100",
  46941=>"001000110",
  46942=>"101110001",
  46943=>"011100011",
  46944=>"010111010",
  46945=>"100000001",
  46946=>"000101100",
  46947=>"001111110",
  46948=>"101001011",
  46949=>"000011010",
  46950=>"101100110",
  46951=>"010011010",
  46952=>"111110110",
  46953=>"011010011",
  46954=>"011101110",
  46955=>"110011100",
  46956=>"000010010",
  46957=>"010001011",
  46958=>"110010010",
  46959=>"101001110",
  46960=>"010010101",
  46961=>"000011010",
  46962=>"101110000",
  46963=>"001100010",
  46964=>"000101111",
  46965=>"101101111",
  46966=>"101001000",
  46967=>"101010101",
  46968=>"100010111",
  46969=>"000000010",
  46970=>"010010011",
  46971=>"111111111",
  46972=>"010111110",
  46973=>"011011100",
  46974=>"000100100",
  46975=>"101001010",
  46976=>"010000011",
  46977=>"000101101",
  46978=>"010000010",
  46979=>"100000010",
  46980=>"000000001",
  46981=>"011010000",
  46982=>"101111110",
  46983=>"001000011",
  46984=>"011000101",
  46985=>"001001001",
  46986=>"101011110",
  46987=>"010101000",
  46988=>"000110101",
  46989=>"111001010",
  46990=>"101000001",
  46991=>"011101001",
  46992=>"010011111",
  46993=>"110111100",
  46994=>"111111101",
  46995=>"110001010",
  46996=>"011101000",
  46997=>"001011000",
  46998=>"110011000",
  46999=>"011111111",
  47000=>"001101011",
  47001=>"000100010",
  47002=>"101010001",
  47003=>"100001001",
  47004=>"010111011",
  47005=>"110011000",
  47006=>"111001110",
  47007=>"000100101",
  47008=>"011011101",
  47009=>"100011110",
  47010=>"101101000",
  47011=>"011000000",
  47012=>"000010010",
  47013=>"111110111",
  47014=>"101111100",
  47015=>"000110011",
  47016=>"111111101",
  47017=>"000111010",
  47018=>"100111110",
  47019=>"110101001",
  47020=>"000000110",
  47021=>"011000110",
  47022=>"001100101",
  47023=>"111000010",
  47024=>"100111010",
  47025=>"100101000",
  47026=>"101011011",
  47027=>"001111100",
  47028=>"111000001",
  47029=>"110010110",
  47030=>"001010011",
  47031=>"110000101",
  47032=>"010000000",
  47033=>"100111011",
  47034=>"101010100",
  47035=>"001100000",
  47036=>"010100111",
  47037=>"001011011",
  47038=>"001001000",
  47039=>"111111110",
  47040=>"001110110",
  47041=>"010011110",
  47042=>"101000100",
  47043=>"001101010",
  47044=>"000110011",
  47045=>"011011011",
  47046=>"111100110",
  47047=>"100011000",
  47048=>"101000010",
  47049=>"100111110",
  47050=>"101111001",
  47051=>"101000010",
  47052=>"010110001",
  47053=>"110100111",
  47054=>"110011000",
  47055=>"000110001",
  47056=>"100000001",
  47057=>"110000111",
  47058=>"110100001",
  47059=>"010011111",
  47060=>"101101010",
  47061=>"000011011",
  47062=>"010010111",
  47063=>"101100100",
  47064=>"001110111",
  47065=>"100000010",
  47066=>"000000001",
  47067=>"011000000",
  47068=>"000010101",
  47069=>"011011101",
  47070=>"001101110",
  47071=>"000010011",
  47072=>"010001111",
  47073=>"001001100",
  47074=>"101101111",
  47075=>"010000000",
  47076=>"010111011",
  47077=>"011001000",
  47078=>"001000100",
  47079=>"010110110",
  47080=>"000011100",
  47081=>"111111001",
  47082=>"011000110",
  47083=>"010001000",
  47084=>"011110101",
  47085=>"001101101",
  47086=>"001100100",
  47087=>"000110101",
  47088=>"110010010",
  47089=>"110100000",
  47090=>"011100101",
  47091=>"010001011",
  47092=>"101101110",
  47093=>"000000101",
  47094=>"101101101",
  47095=>"111100111",
  47096=>"011010100",
  47097=>"100000111",
  47098=>"011000000",
  47099=>"010100110",
  47100=>"100110010",
  47101=>"011101111",
  47102=>"110001101",
  47103=>"000011010",
  47104=>"100111111",
  47105=>"110010000",
  47106=>"011000101",
  47107=>"010101100",
  47108=>"101011100",
  47109=>"100010010",
  47110=>"111010001",
  47111=>"100010000",
  47112=>"111010110",
  47113=>"001101100",
  47114=>"001000111",
  47115=>"010100011",
  47116=>"111110000",
  47117=>"001100111",
  47118=>"110110100",
  47119=>"111100101",
  47120=>"110111010",
  47121=>"101111010",
  47122=>"000001000",
  47123=>"110111001",
  47124=>"000000000",
  47125=>"001101011",
  47126=>"100101111",
  47127=>"000011010",
  47128=>"111001001",
  47129=>"101000100",
  47130=>"001111101",
  47131=>"111111010",
  47132=>"110101110",
  47133=>"100111101",
  47134=>"001011110",
  47135=>"100100011",
  47136=>"100101010",
  47137=>"101011001",
  47138=>"100011011",
  47139=>"111011011",
  47140=>"111000100",
  47141=>"010001010",
  47142=>"100110100",
  47143=>"101100001",
  47144=>"000111100",
  47145=>"000010000",
  47146=>"110011101",
  47147=>"010100011",
  47148=>"011101101",
  47149=>"010011111",
  47150=>"000011011",
  47151=>"111010110",
  47152=>"101010010",
  47153=>"110001000",
  47154=>"011001101",
  47155=>"100001100",
  47156=>"111101100",
  47157=>"010110110",
  47158=>"010111111",
  47159=>"001010001",
  47160=>"000011001",
  47161=>"011100110",
  47162=>"100010000",
  47163=>"101100101",
  47164=>"100000100",
  47165=>"101010011",
  47166=>"000001010",
  47167=>"011011101",
  47168=>"111011001",
  47169=>"000010001",
  47170=>"011011000",
  47171=>"011110000",
  47172=>"001101010",
  47173=>"000001011",
  47174=>"101010000",
  47175=>"110000001",
  47176=>"100111110",
  47177=>"110111000",
  47178=>"000000100",
  47179=>"011000101",
  47180=>"011101100",
  47181=>"011111001",
  47182=>"000011110",
  47183=>"100110000",
  47184=>"101011101",
  47185=>"111110011",
  47186=>"111100011",
  47187=>"000100001",
  47188=>"010101000",
  47189=>"110101100",
  47190=>"100010000",
  47191=>"111100110",
  47192=>"001110110",
  47193=>"001101111",
  47194=>"000110110",
  47195=>"101000001",
  47196=>"000010110",
  47197=>"101010000",
  47198=>"011011001",
  47199=>"011001111",
  47200=>"100111110",
  47201=>"111001001",
  47202=>"010100100",
  47203=>"001101000",
  47204=>"100000000",
  47205=>"011001001",
  47206=>"011100101",
  47207=>"100010000",
  47208=>"001001000",
  47209=>"110000011",
  47210=>"111100101",
  47211=>"010000011",
  47212=>"110110010",
  47213=>"110000000",
  47214=>"011101001",
  47215=>"110001000",
  47216=>"000101000",
  47217=>"100011110",
  47218=>"111000011",
  47219=>"000100000",
  47220=>"100101100",
  47221=>"101011111",
  47222=>"001100001",
  47223=>"010111110",
  47224=>"000100100",
  47225=>"000000101",
  47226=>"010011111",
  47227=>"001100010",
  47228=>"001100101",
  47229=>"001101110",
  47230=>"100101011",
  47231=>"111000100",
  47232=>"101001011",
  47233=>"111101101",
  47234=>"010000101",
  47235=>"000000010",
  47236=>"100101000",
  47237=>"100111000",
  47238=>"100001010",
  47239=>"100111011",
  47240=>"110111000",
  47241=>"111000110",
  47242=>"000000100",
  47243=>"101001111",
  47244=>"101001101",
  47245=>"101000000",
  47246=>"101010110",
  47247=>"110000000",
  47248=>"111111000",
  47249=>"110110110",
  47250=>"001001111",
  47251=>"100101000",
  47252=>"011000000",
  47253=>"001010001",
  47254=>"110011110",
  47255=>"100000010",
  47256=>"010111011",
  47257=>"111011110",
  47258=>"010100011",
  47259=>"111001000",
  47260=>"010100111",
  47261=>"001010011",
  47262=>"111110010",
  47263=>"000101100",
  47264=>"011110011",
  47265=>"110110101",
  47266=>"001011100",
  47267=>"111111100",
  47268=>"111110111",
  47269=>"000011111",
  47270=>"100011110",
  47271=>"001010111",
  47272=>"011010010",
  47273=>"011000101",
  47274=>"001101011",
  47275=>"010011100",
  47276=>"100010110",
  47277=>"001000100",
  47278=>"110011110",
  47279=>"110011110",
  47280=>"111011010",
  47281=>"010101111",
  47282=>"001000111",
  47283=>"000100000",
  47284=>"000001111",
  47285=>"100000111",
  47286=>"100111001",
  47287=>"011100110",
  47288=>"000000001",
  47289=>"110111100",
  47290=>"001111101",
  47291=>"110101001",
  47292=>"010001101",
  47293=>"011000001",
  47294=>"110001010",
  47295=>"110101100",
  47296=>"110010001",
  47297=>"001001000",
  47298=>"101100110",
  47299=>"101110000",
  47300=>"111010101",
  47301=>"111100110",
  47302=>"011000001",
  47303=>"010111001",
  47304=>"001111111",
  47305=>"101001110",
  47306=>"001111001",
  47307=>"111111111",
  47308=>"000000001",
  47309=>"101011110",
  47310=>"011000100",
  47311=>"111100111",
  47312=>"010010111",
  47313=>"100111111",
  47314=>"001001011",
  47315=>"010010001",
  47316=>"011001100",
  47317=>"010001100",
  47318=>"110001101",
  47319=>"101011001",
  47320=>"011111011",
  47321=>"010000010",
  47322=>"000100010",
  47323=>"110101111",
  47324=>"001001011",
  47325=>"101001111",
  47326=>"100000010",
  47327=>"110011111",
  47328=>"000001000",
  47329=>"010011111",
  47330=>"001110111",
  47331=>"001110110",
  47332=>"110010011",
  47333=>"101001010",
  47334=>"001010010",
  47335=>"110111010",
  47336=>"000010101",
  47337=>"101010010",
  47338=>"000100101",
  47339=>"101001011",
  47340=>"111000111",
  47341=>"010001001",
  47342=>"100110111",
  47343=>"110001011",
  47344=>"111011111",
  47345=>"001011011",
  47346=>"000110101",
  47347=>"001010010",
  47348=>"111111010",
  47349=>"110000100",
  47350=>"010000010",
  47351=>"000100011",
  47352=>"111010001",
  47353=>"011101001",
  47354=>"010110100",
  47355=>"010010100",
  47356=>"000000100",
  47357=>"001010111",
  47358=>"110001100",
  47359=>"001010110",
  47360=>"111011011",
  47361=>"000001101",
  47362=>"000101110",
  47363=>"100001100",
  47364=>"010101011",
  47365=>"101110100",
  47366=>"101110110",
  47367=>"000000111",
  47368=>"011111101",
  47369=>"100000111",
  47370=>"011011000",
  47371=>"111101000",
  47372=>"000111111",
  47373=>"011010100",
  47374=>"000100110",
  47375=>"001001111",
  47376=>"011110000",
  47377=>"100101011",
  47378=>"011110000",
  47379=>"000100010",
  47380=>"110101011",
  47381=>"111100110",
  47382=>"100001011",
  47383=>"111101000",
  47384=>"101101000",
  47385=>"100110001",
  47386=>"101001000",
  47387=>"001001000",
  47388=>"001010010",
  47389=>"100101111",
  47390=>"101100000",
  47391=>"001000010",
  47392=>"001101101",
  47393=>"010001001",
  47394=>"010000000",
  47395=>"000011011",
  47396=>"101010111",
  47397=>"000000000",
  47398=>"001110111",
  47399=>"001111011",
  47400=>"010000001",
  47401=>"100111110",
  47402=>"010001110",
  47403=>"110001101",
  47404=>"010100000",
  47405=>"100000001",
  47406=>"001111101",
  47407=>"110100101",
  47408=>"100001000",
  47409=>"011100100",
  47410=>"001011001",
  47411=>"011010110",
  47412=>"001001001",
  47413=>"010010110",
  47414=>"001111000",
  47415=>"100101111",
  47416=>"011100010",
  47417=>"110010100",
  47418=>"100010110",
  47419=>"111010111",
  47420=>"011010010",
  47421=>"011100010",
  47422=>"001010000",
  47423=>"001111011",
  47424=>"101100011",
  47425=>"110100110",
  47426=>"000000011",
  47427=>"000001000",
  47428=>"010111101",
  47429=>"010110100",
  47430=>"100101011",
  47431=>"011001001",
  47432=>"100011100",
  47433=>"101011010",
  47434=>"110111110",
  47435=>"000000000",
  47436=>"010000100",
  47437=>"111110100",
  47438=>"110100010",
  47439=>"110000100",
  47440=>"101000111",
  47441=>"010101000",
  47442=>"001101001",
  47443=>"000001001",
  47444=>"111000011",
  47445=>"010100101",
  47446=>"000011101",
  47447=>"101111000",
  47448=>"101111100",
  47449=>"110011110",
  47450=>"110111101",
  47451=>"011010010",
  47452=>"110000001",
  47453=>"111111000",
  47454=>"110000110",
  47455=>"011010111",
  47456=>"101010011",
  47457=>"111001111",
  47458=>"100110110",
  47459=>"110000101",
  47460=>"110100110",
  47461=>"001010111",
  47462=>"000000111",
  47463=>"000101000",
  47464=>"011111011",
  47465=>"111110001",
  47466=>"010001000",
  47467=>"000011001",
  47468=>"011010101",
  47469=>"000110010",
  47470=>"101000011",
  47471=>"001001000",
  47472=>"001000011",
  47473=>"101101110",
  47474=>"110100111",
  47475=>"011101110",
  47476=>"100000100",
  47477=>"111111011",
  47478=>"000110100",
  47479=>"000100101",
  47480=>"100010110",
  47481=>"010100001",
  47482=>"101010000",
  47483=>"111101001",
  47484=>"000000101",
  47485=>"011000111",
  47486=>"010110011",
  47487=>"111100010",
  47488=>"000010011",
  47489=>"011101010",
  47490=>"110010111",
  47491=>"010001000",
  47492=>"101010011",
  47493=>"010101101",
  47494=>"100001011",
  47495=>"010100010",
  47496=>"000011000",
  47497=>"010011001",
  47498=>"011011011",
  47499=>"101110111",
  47500=>"101111010",
  47501=>"100100110",
  47502=>"011001110",
  47503=>"000001110",
  47504=>"100110111",
  47505=>"100101101",
  47506=>"001010110",
  47507=>"010100100",
  47508=>"001100100",
  47509=>"001000010",
  47510=>"010001010",
  47511=>"110111110",
  47512=>"110010010",
  47513=>"001101011",
  47514=>"001000000",
  47515=>"011010100",
  47516=>"011011010",
  47517=>"110100011",
  47518=>"001100010",
  47519=>"101111000",
  47520=>"000100110",
  47521=>"001111000",
  47522=>"111101000",
  47523=>"101011110",
  47524=>"101101100",
  47525=>"001110001",
  47526=>"000111011",
  47527=>"110101100",
  47528=>"110001110",
  47529=>"001000010",
  47530=>"110111000",
  47531=>"000001011",
  47532=>"100001100",
  47533=>"001000010",
  47534=>"011010010",
  47535=>"100101001",
  47536=>"000000111",
  47537=>"011000001",
  47538=>"001101100",
  47539=>"111110100",
  47540=>"010101111",
  47541=>"110100101",
  47542=>"100111001",
  47543=>"001101100",
  47544=>"101101110",
  47545=>"000000000",
  47546=>"001010100",
  47547=>"111101111",
  47548=>"011111011",
  47549=>"100000011",
  47550=>"011111010",
  47551=>"000011000",
  47552=>"110101000",
  47553=>"011110111",
  47554=>"001111110",
  47555=>"001110001",
  47556=>"100101011",
  47557=>"010001111",
  47558=>"101111110",
  47559=>"011101001",
  47560=>"101110001",
  47561=>"000111011",
  47562=>"000100000",
  47563=>"001001111",
  47564=>"111111101",
  47565=>"010000010",
  47566=>"100011111",
  47567=>"010101110",
  47568=>"111101111",
  47569=>"000001000",
  47570=>"000111011",
  47571=>"001110000",
  47572=>"011001111",
  47573=>"011000011",
  47574=>"001001111",
  47575=>"011111111",
  47576=>"000010010",
  47577=>"110010111",
  47578=>"010000100",
  47579=>"101111010",
  47580=>"100111110",
  47581=>"010101000",
  47582=>"100110111",
  47583=>"001111110",
  47584=>"000011001",
  47585=>"011000001",
  47586=>"111001010",
  47587=>"010111000",
  47588=>"101010011",
  47589=>"000000010",
  47590=>"000000010",
  47591=>"010101011",
  47592=>"001010110",
  47593=>"101111010",
  47594=>"010011110",
  47595=>"111101011",
  47596=>"000000011",
  47597=>"001000000",
  47598=>"011010001",
  47599=>"000101110",
  47600=>"100100111",
  47601=>"011100010",
  47602=>"110111000",
  47603=>"100010000",
  47604=>"101001010",
  47605=>"001101011",
  47606=>"110111110",
  47607=>"001001010",
  47608=>"001010110",
  47609=>"111111010",
  47610=>"110010001",
  47611=>"101100110",
  47612=>"111101111",
  47613=>"000101100",
  47614=>"000001011",
  47615=>"111101101",
  47616=>"010101111",
  47617=>"110111000",
  47618=>"110101001",
  47619=>"111001010",
  47620=>"111100110",
  47621=>"101100101",
  47622=>"001001000",
  47623=>"001010001",
  47624=>"101111000",
  47625=>"010101101",
  47626=>"100111111",
  47627=>"011100000",
  47628=>"001111111",
  47629=>"111001111",
  47630=>"000010000",
  47631=>"000101010",
  47632=>"111000000",
  47633=>"110101001",
  47634=>"100100101",
  47635=>"001000010",
  47636=>"011111111",
  47637=>"110011100",
  47638=>"000100111",
  47639=>"110000011",
  47640=>"111110110",
  47641=>"000010111",
  47642=>"010101011",
  47643=>"011000011",
  47644=>"101100010",
  47645=>"100001100",
  47646=>"101101000",
  47647=>"110111111",
  47648=>"000011100",
  47649=>"001010000",
  47650=>"000011001",
  47651=>"000000111",
  47652=>"100010001",
  47653=>"011100100",
  47654=>"111011110",
  47655=>"001000000",
  47656=>"001011000",
  47657=>"011001001",
  47658=>"100111111",
  47659=>"010001011",
  47660=>"101010101",
  47661=>"100000101",
  47662=>"111001010",
  47663=>"010010100",
  47664=>"010101010",
  47665=>"010011101",
  47666=>"111101000",
  47667=>"100110001",
  47668=>"001010110",
  47669=>"110111000",
  47670=>"110001100",
  47671=>"101111001",
  47672=>"010010101",
  47673=>"001010010",
  47674=>"011110001",
  47675=>"101011100",
  47676=>"011100111",
  47677=>"011100100",
  47678=>"100001010",
  47679=>"110010101",
  47680=>"000100111",
  47681=>"011000000",
  47682=>"010001110",
  47683=>"111011110",
  47684=>"101100011",
  47685=>"000101100",
  47686=>"000101100",
  47687=>"100110100",
  47688=>"001111001",
  47689=>"100010000",
  47690=>"001101111",
  47691=>"010010010",
  47692=>"000100010",
  47693=>"111110010",
  47694=>"100011101",
  47695=>"001011100",
  47696=>"000100110",
  47697=>"111001110",
  47698=>"000000010",
  47699=>"000101111",
  47700=>"111010110",
  47701=>"001111100",
  47702=>"011110100",
  47703=>"110011110",
  47704=>"101010101",
  47705=>"100101100",
  47706=>"011100100",
  47707=>"010011010",
  47708=>"011101000",
  47709=>"110100010",
  47710=>"100010100",
  47711=>"100001100",
  47712=>"101010011",
  47713=>"100000001",
  47714=>"000000101",
  47715=>"101111111",
  47716=>"001101001",
  47717=>"011010000",
  47718=>"011101000",
  47719=>"010110000",
  47720=>"001101100",
  47721=>"011010100",
  47722=>"110110110",
  47723=>"011110000",
  47724=>"011110001",
  47725=>"000010111",
  47726=>"100010111",
  47727=>"111011001",
  47728=>"010000100",
  47729=>"001000100",
  47730=>"101110110",
  47731=>"010100110",
  47732=>"001110001",
  47733=>"111110101",
  47734=>"111101111",
  47735=>"100010100",
  47736=>"011101100",
  47737=>"111111111",
  47738=>"101010111",
  47739=>"000111010",
  47740=>"101010010",
  47741=>"101000111",
  47742=>"000100010",
  47743=>"110010001",
  47744=>"000000010",
  47745=>"000011101",
  47746=>"000000100",
  47747=>"001001001",
  47748=>"010100001",
  47749=>"100011110",
  47750=>"010110111",
  47751=>"110101010",
  47752=>"011110010",
  47753=>"011000010",
  47754=>"111011001",
  47755=>"001000010",
  47756=>"010101110",
  47757=>"100101110",
  47758=>"010010000",
  47759=>"111101111",
  47760=>"100111110",
  47761=>"111001010",
  47762=>"111000100",
  47763=>"000110110",
  47764=>"110101101",
  47765=>"011110111",
  47766=>"110000011",
  47767=>"110100100",
  47768=>"010000001",
  47769=>"001011111",
  47770=>"011011011",
  47771=>"000010101",
  47772=>"001110000",
  47773=>"111101010",
  47774=>"110101100",
  47775=>"011110011",
  47776=>"001000010",
  47777=>"101111010",
  47778=>"010110110",
  47779=>"011001111",
  47780=>"011001000",
  47781=>"011010100",
  47782=>"000010011",
  47783=>"000010101",
  47784=>"011100011",
  47785=>"011000100",
  47786=>"110111011",
  47787=>"001010001",
  47788=>"001011011",
  47789=>"100101111",
  47790=>"110000001",
  47791=>"010001010",
  47792=>"111000111",
  47793=>"100010110",
  47794=>"011000011",
  47795=>"110011101",
  47796=>"010101110",
  47797=>"100010111",
  47798=>"000110110",
  47799=>"110100010",
  47800=>"011110100",
  47801=>"011101011",
  47802=>"111111111",
  47803=>"101000010",
  47804=>"110100010",
  47805=>"000110001",
  47806=>"000101000",
  47807=>"100110000",
  47808=>"010010001",
  47809=>"111110000",
  47810=>"010011001",
  47811=>"001110101",
  47812=>"111111000",
  47813=>"011010010",
  47814=>"001100011",
  47815=>"001000101",
  47816=>"010000100",
  47817=>"101010000",
  47818=>"111100110",
  47819=>"001010001",
  47820=>"010110101",
  47821=>"010100011",
  47822=>"000110011",
  47823=>"101111011",
  47824=>"001000001",
  47825=>"011101010",
  47826=>"011011010",
  47827=>"000110101",
  47828=>"010011111",
  47829=>"001011001",
  47830=>"100100100",
  47831=>"010110000",
  47832=>"110101000",
  47833=>"010111100",
  47834=>"100101001",
  47835=>"001101000",
  47836=>"111010101",
  47837=>"000010011",
  47838=>"011001000",
  47839=>"000011101",
  47840=>"000110000",
  47841=>"000011100",
  47842=>"100101001",
  47843=>"101000000",
  47844=>"100011010",
  47845=>"011011100",
  47846=>"001001101",
  47847=>"000001010",
  47848=>"010111000",
  47849=>"000011111",
  47850=>"000010111",
  47851=>"101001000",
  47852=>"000101000",
  47853=>"000110010",
  47854=>"010010111",
  47855=>"001101100",
  47856=>"001101100",
  47857=>"000010010",
  47858=>"110110101",
  47859=>"111111001",
  47860=>"010010100",
  47861=>"010001110",
  47862=>"110111000",
  47863=>"101101001",
  47864=>"001101111",
  47865=>"011001100",
  47866=>"101001000",
  47867=>"101011000",
  47868=>"100101000",
  47869=>"011011000",
  47870=>"000011100",
  47871=>"111101110",
  47872=>"000100111",
  47873=>"001100001",
  47874=>"110011101",
  47875=>"111001100",
  47876=>"101011000",
  47877=>"101101111",
  47878=>"011100111",
  47879=>"011010010",
  47880=>"101010000",
  47881=>"100111010",
  47882=>"101011110",
  47883=>"010011111",
  47884=>"001010001",
  47885=>"101011101",
  47886=>"000100011",
  47887=>"011011101",
  47888=>"011110000",
  47889=>"100000001",
  47890=>"111000010",
  47891=>"110011011",
  47892=>"101001100",
  47893=>"000010101",
  47894=>"001001100",
  47895=>"100010111",
  47896=>"110110110",
  47897=>"000100111",
  47898=>"010110110",
  47899=>"010011100",
  47900=>"111011110",
  47901=>"010010011",
  47902=>"000011000",
  47903=>"111111000",
  47904=>"000000100",
  47905=>"111110110",
  47906=>"010111011",
  47907=>"110010110",
  47908=>"101110011",
  47909=>"000100100",
  47910=>"100000110",
  47911=>"000010110",
  47912=>"000010100",
  47913=>"010001111",
  47914=>"110110010",
  47915=>"110010001",
  47916=>"110101101",
  47917=>"010000100",
  47918=>"110101101",
  47919=>"101101111",
  47920=>"110000011",
  47921=>"010111011",
  47922=>"001001111",
  47923=>"111100100",
  47924=>"111110111",
  47925=>"110000000",
  47926=>"001110000",
  47927=>"001101010",
  47928=>"010100000",
  47929=>"010001111",
  47930=>"000111111",
  47931=>"010111011",
  47932=>"011100000",
  47933=>"000110001",
  47934=>"110001100",
  47935=>"000110010",
  47936=>"001001000",
  47937=>"000100100",
  47938=>"111001000",
  47939=>"100100011",
  47940=>"011101001",
  47941=>"001111111",
  47942=>"000010001",
  47943=>"110000010",
  47944=>"111101000",
  47945=>"110100010",
  47946=>"001100011",
  47947=>"010010001",
  47948=>"010000101",
  47949=>"010111101",
  47950=>"001011000",
  47951=>"011111001",
  47952=>"001000011",
  47953=>"000010000",
  47954=>"000110110",
  47955=>"000110001",
  47956=>"110111001",
  47957=>"111110010",
  47958=>"101110100",
  47959=>"110010111",
  47960=>"001000010",
  47961=>"000011001",
  47962=>"110101011",
  47963=>"000100100",
  47964=>"000101011",
  47965=>"111101111",
  47966=>"010101010",
  47967=>"001111111",
  47968=>"010101110",
  47969=>"011011111",
  47970=>"111110000",
  47971=>"001001001",
  47972=>"011010000",
  47973=>"011110000",
  47974=>"100000001",
  47975=>"111101001",
  47976=>"010010010",
  47977=>"101100111",
  47978=>"010101110",
  47979=>"000110001",
  47980=>"101001101",
  47981=>"101010000",
  47982=>"010000000",
  47983=>"010100001",
  47984=>"111100010",
  47985=>"000000101",
  47986=>"001011000",
  47987=>"010000011",
  47988=>"000110000",
  47989=>"011001000",
  47990=>"111001111",
  47991=>"011011011",
  47992=>"101111010",
  47993=>"000110001",
  47994=>"110100001",
  47995=>"111011000",
  47996=>"000000100",
  47997=>"010110000",
  47998=>"001100001",
  47999=>"011101100",
  48000=>"111101000",
  48001=>"001111000",
  48002=>"100000011",
  48003=>"010000011",
  48004=>"110100011",
  48005=>"000000110",
  48006=>"000000000",
  48007=>"000010000",
  48008=>"010001000",
  48009=>"001010100",
  48010=>"100000111",
  48011=>"111111111",
  48012=>"000110111",
  48013=>"000000100",
  48014=>"011110100",
  48015=>"100011010",
  48016=>"010010000",
  48017=>"000101101",
  48018=>"001100000",
  48019=>"101001000",
  48020=>"010101010",
  48021=>"110111001",
  48022=>"011110011",
  48023=>"100001001",
  48024=>"001101111",
  48025=>"000000000",
  48026=>"010110011",
  48027=>"101110101",
  48028=>"001111010",
  48029=>"111001110",
  48030=>"110010001",
  48031=>"001000111",
  48032=>"010010000",
  48033=>"110100111",
  48034=>"010100111",
  48035=>"101001101",
  48036=>"001011110",
  48037=>"111111010",
  48038=>"111011011",
  48039=>"110101111",
  48040=>"000101011",
  48041=>"010101010",
  48042=>"100100010",
  48043=>"000010100",
  48044=>"100010101",
  48045=>"000100101",
  48046=>"110011000",
  48047=>"101011001",
  48048=>"111011000",
  48049=>"110011111",
  48050=>"000110000",
  48051=>"010101100",
  48052=>"001101110",
  48053=>"100010100",
  48054=>"010000111",
  48055=>"001111111",
  48056=>"001001100",
  48057=>"001101111",
  48058=>"100001000",
  48059=>"011100011",
  48060=>"100000111",
  48061=>"100000100",
  48062=>"000110111",
  48063=>"011010110",
  48064=>"011011000",
  48065=>"101010111",
  48066=>"000010000",
  48067=>"000100010",
  48068=>"000010000",
  48069=>"011010101",
  48070=>"010001011",
  48071=>"110001111",
  48072=>"011100110",
  48073=>"010010010",
  48074=>"101111000",
  48075=>"111100001",
  48076=>"011100100",
  48077=>"111001111",
  48078=>"000110010",
  48079=>"001101011",
  48080=>"101100101",
  48081=>"101101111",
  48082=>"100000001",
  48083=>"110011000",
  48084=>"111111111",
  48085=>"000100100",
  48086=>"000000011",
  48087=>"000100111",
  48088=>"011100110",
  48089=>"000001100",
  48090=>"011101001",
  48091=>"001000001",
  48092=>"001001110",
  48093=>"000101000",
  48094=>"010000011",
  48095=>"111001011",
  48096=>"000011011",
  48097=>"000001100",
  48098=>"011101100",
  48099=>"100111111",
  48100=>"100100101",
  48101=>"110100111",
  48102=>"000101011",
  48103=>"000110000",
  48104=>"110111100",
  48105=>"001100111",
  48106=>"100001010",
  48107=>"100010000",
  48108=>"001001000",
  48109=>"010010110",
  48110=>"000100000",
  48111=>"111110011",
  48112=>"111101010",
  48113=>"000011010",
  48114=>"111000001",
  48115=>"001001100",
  48116=>"101101011",
  48117=>"001000001",
  48118=>"001010010",
  48119=>"110100101",
  48120=>"000010100",
  48121=>"001110110",
  48122=>"010111100",
  48123=>"110001100",
  48124=>"110010110",
  48125=>"010011100",
  48126=>"011011101",
  48127=>"111001000",
  48128=>"001000010",
  48129=>"000110000",
  48130=>"101110011",
  48131=>"000111010",
  48132=>"000111001",
  48133=>"100100010",
  48134=>"010001111",
  48135=>"110001100",
  48136=>"100010000",
  48137=>"100010000",
  48138=>"001001100",
  48139=>"000011101",
  48140=>"011111110",
  48141=>"001011010",
  48142=>"111001111",
  48143=>"001000111",
  48144=>"010110001",
  48145=>"000000001",
  48146=>"010100101",
  48147=>"001100000",
  48148=>"110011101",
  48149=>"001111100",
  48150=>"001101101",
  48151=>"001110110",
  48152=>"011010100",
  48153=>"101101000",
  48154=>"000101010",
  48155=>"111010101",
  48156=>"100010011",
  48157=>"101001000",
  48158=>"011111110",
  48159=>"100110100",
  48160=>"001100100",
  48161=>"111110001",
  48162=>"100001110",
  48163=>"011011011",
  48164=>"010101011",
  48165=>"101001100",
  48166=>"011011000",
  48167=>"101111000",
  48168=>"111110010",
  48169=>"010000001",
  48170=>"101000011",
  48171=>"100110101",
  48172=>"111010101",
  48173=>"101101110",
  48174=>"110100001",
  48175=>"110110000",
  48176=>"110111000",
  48177=>"011011000",
  48178=>"010010100",
  48179=>"100100000",
  48180=>"011010000",
  48181=>"101111010",
  48182=>"100101111",
  48183=>"010100001",
  48184=>"110010110",
  48185=>"111100000",
  48186=>"000000010",
  48187=>"001000000",
  48188=>"001011010",
  48189=>"000100000",
  48190=>"010000110",
  48191=>"001001111",
  48192=>"110100010",
  48193=>"000100001",
  48194=>"100001100",
  48195=>"101010000",
  48196=>"010110010",
  48197=>"111100001",
  48198=>"001011011",
  48199=>"100111000",
  48200=>"010111100",
  48201=>"010010100",
  48202=>"101010110",
  48203=>"001100010",
  48204=>"111100000",
  48205=>"100111101",
  48206=>"111001001",
  48207=>"101101011",
  48208=>"001111011",
  48209=>"000100100",
  48210=>"001001011",
  48211=>"111001001",
  48212=>"000000011",
  48213=>"000100000",
  48214=>"010100111",
  48215=>"010110010",
  48216=>"110000011",
  48217=>"110001001",
  48218=>"110010111",
  48219=>"010101111",
  48220=>"001110101",
  48221=>"011000000",
  48222=>"101101100",
  48223=>"000000001",
  48224=>"010001100",
  48225=>"110111100",
  48226=>"010101111",
  48227=>"111101100",
  48228=>"101100000",
  48229=>"111100011",
  48230=>"100000111",
  48231=>"010110000",
  48232=>"100100000",
  48233=>"001100011",
  48234=>"101100111",
  48235=>"001110010",
  48236=>"011001000",
  48237=>"001110010",
  48238=>"110110000",
  48239=>"111011111",
  48240=>"101000110",
  48241=>"101011001",
  48242=>"110001111",
  48243=>"000010010",
  48244=>"101111100",
  48245=>"011110111",
  48246=>"110101010",
  48247=>"110110000",
  48248=>"111100111",
  48249=>"000111000",
  48250=>"101001000",
  48251=>"111011101",
  48252=>"101001000",
  48253=>"001100110",
  48254=>"000100001",
  48255=>"000110001",
  48256=>"011000010",
  48257=>"001110100",
  48258=>"101100100",
  48259=>"000101010",
  48260=>"001110101",
  48261=>"000000011",
  48262=>"011000111",
  48263=>"101111010",
  48264=>"111111111",
  48265=>"001011101",
  48266=>"010001110",
  48267=>"001010111",
  48268=>"001011010",
  48269=>"110000100",
  48270=>"010101101",
  48271=>"100111010",
  48272=>"011010110",
  48273=>"000110001",
  48274=>"010110001",
  48275=>"101001000",
  48276=>"110001011",
  48277=>"100010001",
  48278=>"100001000",
  48279=>"010010101",
  48280=>"000001111",
  48281=>"110111100",
  48282=>"110100000",
  48283=>"101111010",
  48284=>"110001100",
  48285=>"111111011",
  48286=>"110000100",
  48287=>"100111111",
  48288=>"100000111",
  48289=>"000000100",
  48290=>"101111101",
  48291=>"010011111",
  48292=>"111011111",
  48293=>"000000101",
  48294=>"010000111",
  48295=>"101011100",
  48296=>"110111111",
  48297=>"011001010",
  48298=>"111100110",
  48299=>"000101011",
  48300=>"111110011",
  48301=>"111100111",
  48302=>"000011010",
  48303=>"010110101",
  48304=>"111000100",
  48305=>"000110010",
  48306=>"000000111",
  48307=>"100100101",
  48308=>"100000001",
  48309=>"000111100",
  48310=>"111100100",
  48311=>"011011010",
  48312=>"111000110",
  48313=>"000001100",
  48314=>"110000101",
  48315=>"110001111",
  48316=>"001000001",
  48317=>"011011011",
  48318=>"000000001",
  48319=>"000010010",
  48320=>"001011000",
  48321=>"101010010",
  48322=>"000101110",
  48323=>"111000001",
  48324=>"100111000",
  48325=>"110010111",
  48326=>"010010110",
  48327=>"100111111",
  48328=>"001101001",
  48329=>"111001110",
  48330=>"101011111",
  48331=>"001110110",
  48332=>"110000101",
  48333=>"100010111",
  48334=>"000110100",
  48335=>"101111001",
  48336=>"100010000",
  48337=>"110001100",
  48338=>"001011000",
  48339=>"110001000",
  48340=>"111001011",
  48341=>"100000110",
  48342=>"101110001",
  48343=>"010111110",
  48344=>"111010011",
  48345=>"111101101",
  48346=>"110001110",
  48347=>"110100100",
  48348=>"100101101",
  48349=>"100001011",
  48350=>"001101001",
  48351=>"011010001",
  48352=>"001001011",
  48353=>"001011001",
  48354=>"111111100",
  48355=>"011100100",
  48356=>"010010111",
  48357=>"001010111",
  48358=>"001101100",
  48359=>"100010011",
  48360=>"011001001",
  48361=>"111101100",
  48362=>"111111010",
  48363=>"010011001",
  48364=>"001111110",
  48365=>"000101101",
  48366=>"000011111",
  48367=>"011010011",
  48368=>"110011000",
  48369=>"010011100",
  48370=>"100101111",
  48371=>"011000110",
  48372=>"000110110",
  48373=>"011100111",
  48374=>"100010011",
  48375=>"000011101",
  48376=>"000011101",
  48377=>"011001110",
  48378=>"111100011",
  48379=>"110010011",
  48380=>"011011010",
  48381=>"111101111",
  48382=>"110110101",
  48383=>"011100111",
  48384=>"011111101",
  48385=>"001011111",
  48386=>"101011111",
  48387=>"001001100",
  48388=>"111111111",
  48389=>"111101010",
  48390=>"010011110",
  48391=>"010111000",
  48392=>"111110111",
  48393=>"110010010",
  48394=>"010000111",
  48395=>"101010100",
  48396=>"101011100",
  48397=>"000010100",
  48398=>"100110010",
  48399=>"100101101",
  48400=>"001110111",
  48401=>"010100111",
  48402=>"011100010",
  48403=>"111000010",
  48404=>"010111000",
  48405=>"000101011",
  48406=>"001000010",
  48407=>"010110011",
  48408=>"100010000",
  48409=>"101000001",
  48410=>"011110010",
  48411=>"011011010",
  48412=>"000111000",
  48413=>"111010010",
  48414=>"011001000",
  48415=>"000010011",
  48416=>"100011110",
  48417=>"111111101",
  48418=>"011110110",
  48419=>"111111011",
  48420=>"110001101",
  48421=>"111000010",
  48422=>"111110000",
  48423=>"011110111",
  48424=>"010000110",
  48425=>"101010001",
  48426=>"000010010",
  48427=>"101100101",
  48428=>"101111000",
  48429=>"010010100",
  48430=>"011000100",
  48431=>"001011010",
  48432=>"001000110",
  48433=>"001010110",
  48434=>"111010111",
  48435=>"100100010",
  48436=>"111010010",
  48437=>"001000000",
  48438=>"001011100",
  48439=>"010011011",
  48440=>"010011011",
  48441=>"100011110",
  48442=>"101000110",
  48443=>"111100011",
  48444=>"101011100",
  48445=>"001000100",
  48446=>"010101100",
  48447=>"101111001",
  48448=>"000111111",
  48449=>"111011111",
  48450=>"001001011",
  48451=>"100110101",
  48452=>"111010110",
  48453=>"100011111",
  48454=>"111111100",
  48455=>"011000000",
  48456=>"101110111",
  48457=>"011110000",
  48458=>"001110011",
  48459=>"011001000",
  48460=>"000100001",
  48461=>"110001000",
  48462=>"100010000",
  48463=>"101001100",
  48464=>"101010101",
  48465=>"001000100",
  48466=>"100000001",
  48467=>"001111001",
  48468=>"111001011",
  48469=>"010111101",
  48470=>"000010100",
  48471=>"000110000",
  48472=>"000010001",
  48473=>"101110111",
  48474=>"011010100",
  48475=>"000111000",
  48476=>"111110001",
  48477=>"101001001",
  48478=>"011000001",
  48479=>"111010001",
  48480=>"000110001",
  48481=>"011001010",
  48482=>"010000111",
  48483=>"011010010",
  48484=>"100000010",
  48485=>"010001100",
  48486=>"101100000",
  48487=>"010001111",
  48488=>"001000010",
  48489=>"001111000",
  48490=>"011110000",
  48491=>"000000111",
  48492=>"010011010",
  48493=>"001111001",
  48494=>"011110101",
  48495=>"001110000",
  48496=>"001110001",
  48497=>"100011011",
  48498=>"110010011",
  48499=>"001000010",
  48500=>"000001101",
  48501=>"110011011",
  48502=>"010000011",
  48503=>"101110000",
  48504=>"101000110",
  48505=>"001011100",
  48506=>"111000100",
  48507=>"100001110",
  48508=>"001001011",
  48509=>"101100101",
  48510=>"001000100",
  48511=>"011001000",
  48512=>"101001001",
  48513=>"110101111",
  48514=>"101101111",
  48515=>"000000101",
  48516=>"001001111",
  48517=>"000110110",
  48518=>"101100101",
  48519=>"000100110",
  48520=>"001001101",
  48521=>"110010101",
  48522=>"100110110",
  48523=>"000000001",
  48524=>"110010111",
  48525=>"000010111",
  48526=>"010100011",
  48527=>"101001111",
  48528=>"101010011",
  48529=>"000111010",
  48530=>"010001011",
  48531=>"100111110",
  48532=>"001111000",
  48533=>"000001001",
  48534=>"000101010",
  48535=>"111101010",
  48536=>"001100110",
  48537=>"001000001",
  48538=>"101011101",
  48539=>"111111100",
  48540=>"101011111",
  48541=>"000010101",
  48542=>"101110101",
  48543=>"110110111",
  48544=>"011011111",
  48545=>"110000011",
  48546=>"101111111",
  48547=>"101000011",
  48548=>"001001010",
  48549=>"101110111",
  48550=>"010010101",
  48551=>"101110110",
  48552=>"101101011",
  48553=>"110011011",
  48554=>"110000010",
  48555=>"100111101",
  48556=>"011000110",
  48557=>"010011000",
  48558=>"100010110",
  48559=>"001011010",
  48560=>"111111010",
  48561=>"010101110",
  48562=>"000110111",
  48563=>"101110010",
  48564=>"100001010",
  48565=>"010101001",
  48566=>"010011101",
  48567=>"110100001",
  48568=>"001101001",
  48569=>"101011110",
  48570=>"000000000",
  48571=>"000100000",
  48572=>"101110001",
  48573=>"101110001",
  48574=>"011110011",
  48575=>"001101111",
  48576=>"110010000",
  48577=>"000001101",
  48578=>"000001111",
  48579=>"100011000",
  48580=>"101100001",
  48581=>"001101110",
  48582=>"010101000",
  48583=>"000110010",
  48584=>"111000011",
  48585=>"100010010",
  48586=>"111101001",
  48587=>"011101111",
  48588=>"011010101",
  48589=>"101001101",
  48590=>"110110011",
  48591=>"101111011",
  48592=>"011000100",
  48593=>"100111111",
  48594=>"000011110",
  48595=>"010111010",
  48596=>"111101000",
  48597=>"000100000",
  48598=>"011001101",
  48599=>"110001000",
  48600=>"001111111",
  48601=>"010011010",
  48602=>"100100100",
  48603=>"111010101",
  48604=>"110010000",
  48605=>"011110000",
  48606=>"001101010",
  48607=>"011000100",
  48608=>"111100111",
  48609=>"111100000",
  48610=>"101010111",
  48611=>"010000100",
  48612=>"110100100",
  48613=>"111011111",
  48614=>"010001000",
  48615=>"000100111",
  48616=>"000000000",
  48617=>"100011010",
  48618=>"111001010",
  48619=>"111110110",
  48620=>"010011000",
  48621=>"001001000",
  48622=>"010011101",
  48623=>"000011110",
  48624=>"000001011",
  48625=>"000000101",
  48626=>"101100111",
  48627=>"101001000",
  48628=>"000010101",
  48629=>"111110010",
  48630=>"010101100",
  48631=>"100111001",
  48632=>"110001100",
  48633=>"000010011",
  48634=>"100110011",
  48635=>"011101100",
  48636=>"110000100",
  48637=>"101010011",
  48638=>"100101111",
  48639=>"010000010",
  48640=>"011001011",
  48641=>"010000000",
  48642=>"010110101",
  48643=>"111011000",
  48644=>"101010010",
  48645=>"100010000",
  48646=>"010000110",
  48647=>"111111111",
  48648=>"000001010",
  48649=>"101110011",
  48650=>"000110110",
  48651=>"101000001",
  48652=>"001011010",
  48653=>"001111001",
  48654=>"000011000",
  48655=>"111111001",
  48656=>"000000100",
  48657=>"100111001",
  48658=>"101100010",
  48659=>"100000101",
  48660=>"000001010",
  48661=>"010111001",
  48662=>"101111101",
  48663=>"000001001",
  48664=>"111011010",
  48665=>"001101011",
  48666=>"010100000",
  48667=>"111111001",
  48668=>"100000101",
  48669=>"101100100",
  48670=>"000110111",
  48671=>"010110010",
  48672=>"010001101",
  48673=>"011110111",
  48674=>"101100100",
  48675=>"000101000",
  48676=>"101101101",
  48677=>"110110011",
  48678=>"110001010",
  48679=>"011111000",
  48680=>"100010010",
  48681=>"111011110",
  48682=>"111101111",
  48683=>"110110010",
  48684=>"000000000",
  48685=>"111111111",
  48686=>"000000011",
  48687=>"001001110",
  48688=>"011011010",
  48689=>"101010010",
  48690=>"110010001",
  48691=>"011101110",
  48692=>"011101111",
  48693=>"110000010",
  48694=>"100100011",
  48695=>"110101010",
  48696=>"001100111",
  48697=>"111111000",
  48698=>"001000010",
  48699=>"100001101",
  48700=>"110100101",
  48701=>"111110000",
  48702=>"100000001",
  48703=>"111010101",
  48704=>"110001101",
  48705=>"011101110",
  48706=>"100000011",
  48707=>"000010101",
  48708=>"000111110",
  48709=>"111100010",
  48710=>"011001111",
  48711=>"000111100",
  48712=>"010101101",
  48713=>"111110100",
  48714=>"001000001",
  48715=>"010000101",
  48716=>"000000100",
  48717=>"111000000",
  48718=>"001000110",
  48719=>"100101001",
  48720=>"001001101",
  48721=>"000111101",
  48722=>"010000101",
  48723=>"110010001",
  48724=>"111100001",
  48725=>"111110010",
  48726=>"110000110",
  48727=>"110010001",
  48728=>"001100111",
  48729=>"111101001",
  48730=>"001111100",
  48731=>"100001101",
  48732=>"001010011",
  48733=>"110000100",
  48734=>"110111100",
  48735=>"010001101",
  48736=>"000111001",
  48737=>"010110000",
  48738=>"110001101",
  48739=>"000000000",
  48740=>"001011010",
  48741=>"111110110",
  48742=>"001111110",
  48743=>"000001000",
  48744=>"001001010",
  48745=>"001100010",
  48746=>"111111110",
  48747=>"010101100",
  48748=>"000001001",
  48749=>"111101010",
  48750=>"000010111",
  48751=>"100000010",
  48752=>"101110000",
  48753=>"011100011",
  48754=>"101101101",
  48755=>"111001100",
  48756=>"001001001",
  48757=>"101111000",
  48758=>"000111000",
  48759=>"110001010",
  48760=>"001111001",
  48761=>"010000100",
  48762=>"111001001",
  48763=>"000111010",
  48764=>"110100011",
  48765=>"110010110",
  48766=>"000110010",
  48767=>"110110010",
  48768=>"010101100",
  48769=>"110111111",
  48770=>"010000100",
  48771=>"001000011",
  48772=>"000110100",
  48773=>"101010101",
  48774=>"101000101",
  48775=>"111101011",
  48776=>"111100101",
  48777=>"000000000",
  48778=>"010011101",
  48779=>"101110010",
  48780=>"110011111",
  48781=>"011101000",
  48782=>"101101001",
  48783=>"110001000",
  48784=>"111000111",
  48785=>"100001001",
  48786=>"000101001",
  48787=>"100010010",
  48788=>"111111111",
  48789=>"011010110",
  48790=>"011010111",
  48791=>"101111000",
  48792=>"111101111",
  48793=>"001110110",
  48794=>"000000111",
  48795=>"000000000",
  48796=>"000101000",
  48797=>"100001111",
  48798=>"110101110",
  48799=>"010000011",
  48800=>"000001110",
  48801=>"001110011",
  48802=>"010010100",
  48803=>"010011001",
  48804=>"100011001",
  48805=>"110010101",
  48806=>"111011100",
  48807=>"001000110",
  48808=>"011100010",
  48809=>"000001011",
  48810=>"111010110",
  48811=>"001011111",
  48812=>"110001011",
  48813=>"001001001",
  48814=>"001100000",
  48815=>"011111011",
  48816=>"101000000",
  48817=>"010010100",
  48818=>"011011111",
  48819=>"001011100",
  48820=>"001011110",
  48821=>"001101010",
  48822=>"011101101",
  48823=>"011100001",
  48824=>"100001011",
  48825=>"100101101",
  48826=>"110100010",
  48827=>"101101001",
  48828=>"000011110",
  48829=>"111110101",
  48830=>"111110010",
  48831=>"100111101",
  48832=>"010110111",
  48833=>"000010111",
  48834=>"101010010",
  48835=>"000100011",
  48836=>"010010100",
  48837=>"111011011",
  48838=>"101101101",
  48839=>"100111101",
  48840=>"011001101",
  48841=>"100011100",
  48842=>"101011110",
  48843=>"110011001",
  48844=>"000010100",
  48845=>"000110011",
  48846=>"100010101",
  48847=>"110000000",
  48848=>"110101011",
  48849=>"000110001",
  48850=>"010101011",
  48851=>"000011010",
  48852=>"101110001",
  48853=>"001001001",
  48854=>"000011001",
  48855=>"001000011",
  48856=>"010101100",
  48857=>"110111010",
  48858=>"100000100",
  48859=>"100100000",
  48860=>"101111101",
  48861=>"100111100",
  48862=>"001001010",
  48863=>"000100011",
  48864=>"100110000",
  48865=>"001001100",
  48866=>"101110000",
  48867=>"001000010",
  48868=>"101101011",
  48869=>"011101100",
  48870=>"100011100",
  48871=>"011001001",
  48872=>"110101011",
  48873=>"111100000",
  48874=>"100111101",
  48875=>"101011001",
  48876=>"010110100",
  48877=>"001000111",
  48878=>"111111111",
  48879=>"100111011",
  48880=>"010111101",
  48881=>"100010000",
  48882=>"010100000",
  48883=>"000001101",
  48884=>"111000111",
  48885=>"110011010",
  48886=>"011011100",
  48887=>"010001000",
  48888=>"011110000",
  48889=>"110011001",
  48890=>"010000000",
  48891=>"001101101",
  48892=>"111000010",
  48893=>"100000100",
  48894=>"101011010",
  48895=>"001100000",
  48896=>"110100011",
  48897=>"000010110",
  48898=>"101100110",
  48899=>"101001101",
  48900=>"100001000",
  48901=>"100100100",
  48902=>"111001100",
  48903=>"110110000",
  48904=>"011100000",
  48905=>"001111000",
  48906=>"101111000",
  48907=>"000010010",
  48908=>"111101011",
  48909=>"010110011",
  48910=>"111000110",
  48911=>"101101101",
  48912=>"100010001",
  48913=>"000010000",
  48914=>"110101101",
  48915=>"111000111",
  48916=>"000110000",
  48917=>"010100101",
  48918=>"011001110",
  48919=>"011010000",
  48920=>"010000010",
  48921=>"100110111",
  48922=>"010100100",
  48923=>"111101011",
  48924=>"001000110",
  48925=>"010000110",
  48926=>"000011110",
  48927=>"011110110",
  48928=>"110001001",
  48929=>"011011100",
  48930=>"111010111",
  48931=>"001001111",
  48932=>"011001111",
  48933=>"111101110",
  48934=>"011001110",
  48935=>"001001010",
  48936=>"011000101",
  48937=>"100001000",
  48938=>"001110100",
  48939=>"011010011",
  48940=>"111101001",
  48941=>"110000111",
  48942=>"001100010",
  48943=>"100000101",
  48944=>"000000000",
  48945=>"000000011",
  48946=>"000111010",
  48947=>"000100100",
  48948=>"111011011",
  48949=>"011000100",
  48950=>"110111111",
  48951=>"010110011",
  48952=>"100100111",
  48953=>"100100101",
  48954=>"111011100",
  48955=>"000100101",
  48956=>"000100011",
  48957=>"110000011",
  48958=>"110111100",
  48959=>"100110001",
  48960=>"001100111",
  48961=>"011010101",
  48962=>"000010000",
  48963=>"111111001",
  48964=>"111011110",
  48965=>"101101111",
  48966=>"101111000",
  48967=>"001011100",
  48968=>"010011101",
  48969=>"001101110",
  48970=>"000001001",
  48971=>"101000010",
  48972=>"001111001",
  48973=>"111111010",
  48974=>"100101000",
  48975=>"101010111",
  48976=>"111101000",
  48977=>"100100010",
  48978=>"010011011",
  48979=>"000001000",
  48980=>"110111011",
  48981=>"010100001",
  48982=>"001001011",
  48983=>"011000101",
  48984=>"000010010",
  48985=>"101111010",
  48986=>"101111011",
  48987=>"000000100",
  48988=>"001100011",
  48989=>"110010100",
  48990=>"010000111",
  48991=>"111010000",
  48992=>"011110010",
  48993=>"111101100",
  48994=>"010011001",
  48995=>"000001000",
  48996=>"110001101",
  48997=>"000010101",
  48998=>"000000001",
  48999=>"010101100",
  49000=>"001010011",
  49001=>"010010011",
  49002=>"101110101",
  49003=>"101101100",
  49004=>"110101111",
  49005=>"101110001",
  49006=>"101011010",
  49007=>"001101010",
  49008=>"111000001",
  49009=>"010110111",
  49010=>"101111110",
  49011=>"110011000",
  49012=>"011110010",
  49013=>"000010111",
  49014=>"011111110",
  49015=>"111110001",
  49016=>"011000100",
  49017=>"111001000",
  49018=>"110000110",
  49019=>"101101110",
  49020=>"101111111",
  49021=>"010100011",
  49022=>"000000101",
  49023=>"010000110",
  49024=>"110011010",
  49025=>"001010011",
  49026=>"111001110",
  49027=>"000000110",
  49028=>"001010010",
  49029=>"000111100",
  49030=>"110001111",
  49031=>"000010000",
  49032=>"101110101",
  49033=>"001001010",
  49034=>"101000011",
  49035=>"111111100",
  49036=>"101011010",
  49037=>"000011111",
  49038=>"001000010",
  49039=>"100010100",
  49040=>"100010010",
  49041=>"101000000",
  49042=>"100010110",
  49043=>"110011010",
  49044=>"111111100",
  49045=>"110011010",
  49046=>"000101101",
  49047=>"110000001",
  49048=>"110110010",
  49049=>"001100100",
  49050=>"100010000",
  49051=>"101111100",
  49052=>"010001000",
  49053=>"000010100",
  49054=>"010110000",
  49055=>"001100000",
  49056=>"010110110",
  49057=>"000110101",
  49058=>"011001110",
  49059=>"101010101",
  49060=>"101110001",
  49061=>"100000010",
  49062=>"011011111",
  49063=>"001100001",
  49064=>"110100111",
  49065=>"110100101",
  49066=>"111010000",
  49067=>"111000100",
  49068=>"010110010",
  49069=>"111000111",
  49070=>"001011101",
  49071=>"111011000",
  49072=>"010001001",
  49073=>"001101000",
  49074=>"111101111",
  49075=>"110000000",
  49076=>"011111101",
  49077=>"010111011",
  49078=>"101010101",
  49079=>"110111011",
  49080=>"101001000",
  49081=>"001000100",
  49082=>"000111100",
  49083=>"011001110",
  49084=>"100101110",
  49085=>"111111100",
  49086=>"101100011",
  49087=>"011100101",
  49088=>"011010011",
  49089=>"100100111",
  49090=>"010111001",
  49091=>"110001010",
  49092=>"010011111",
  49093=>"000100001",
  49094=>"010001010",
  49095=>"010100111",
  49096=>"000100101",
  49097=>"010011000",
  49098=>"000001100",
  49099=>"110001110",
  49100=>"011010010",
  49101=>"010101111",
  49102=>"101111001",
  49103=>"100100011",
  49104=>"101100100",
  49105=>"010000000",
  49106=>"101100000",
  49107=>"111001110",
  49108=>"111001000",
  49109=>"111011001",
  49110=>"111110101",
  49111=>"111110010",
  49112=>"011000110",
  49113=>"110011011",
  49114=>"100111110",
  49115=>"011110101",
  49116=>"111001010",
  49117=>"001100010",
  49118=>"111111000",
  49119=>"101100100",
  49120=>"000100000",
  49121=>"100111000",
  49122=>"111011011",
  49123=>"101000001",
  49124=>"110011000",
  49125=>"110110101",
  49126=>"101101000",
  49127=>"110101100",
  49128=>"001010010",
  49129=>"110100010",
  49130=>"101100000",
  49131=>"101010101",
  49132=>"011110111",
  49133=>"010001101",
  49134=>"000100100",
  49135=>"101111010",
  49136=>"111010111",
  49137=>"000010111",
  49138=>"011000101",
  49139=>"010100011",
  49140=>"100111100",
  49141=>"000100100",
  49142=>"101110101",
  49143=>"101101111",
  49144=>"011101000",
  49145=>"011111110",
  49146=>"000001111",
  49147=>"101010000",
  49148=>"101001101",
  49149=>"000101101",
  49150=>"000011000",
  49151=>"110010011",
  49152=>"110000111",
  49153=>"011110011",
  49154=>"110011010",
  49155=>"010001010",
  49156=>"001100101",
  49157=>"101101110",
  49158=>"100110111",
  49159=>"001000001",
  49160=>"101101111",
  49161=>"111101010",
  49162=>"011001011",
  49163=>"001110100",
  49164=>"010001100",
  49165=>"101111101",
  49166=>"101000001",
  49167=>"010000001",
  49168=>"011010001",
  49169=>"101101100",
  49170=>"100000010",
  49171=>"111010101",
  49172=>"100110110",
  49173=>"011101010",
  49174=>"001101001",
  49175=>"011111101",
  49176=>"000100111",
  49177=>"110011011",
  49178=>"010110111",
  49179=>"111110100",
  49180=>"100001101",
  49181=>"100101101",
  49182=>"101100011",
  49183=>"100000101",
  49184=>"001010001",
  49185=>"011010100",
  49186=>"110111111",
  49187=>"000110011",
  49188=>"100110111",
  49189=>"100000111",
  49190=>"111100111",
  49191=>"011000010",
  49192=>"000010100",
  49193=>"110011101",
  49194=>"111101100",
  49195=>"001010010",
  49196=>"100011010",
  49197=>"010000000",
  49198=>"110101100",
  49199=>"111000011",
  49200=>"011001000",
  49201=>"010100101",
  49202=>"111110101",
  49203=>"110110000",
  49204=>"011000111",
  49205=>"011101001",
  49206=>"100010100",
  49207=>"011111001",
  49208=>"110100010",
  49209=>"001101111",
  49210=>"110011111",
  49211=>"111010101",
  49212=>"111101000",
  49213=>"111111111",
  49214=>"100000101",
  49215=>"000000110",
  49216=>"111110101",
  49217=>"110001110",
  49218=>"011011000",
  49219=>"011101110",
  49220=>"010110000",
  49221=>"100111011",
  49222=>"111010111",
  49223=>"100101101",
  49224=>"111010001",
  49225=>"001100000",
  49226=>"101011000",
  49227=>"000000101",
  49228=>"010011010",
  49229=>"011011011",
  49230=>"100010111",
  49231=>"111111111",
  49232=>"010100001",
  49233=>"000000100",
  49234=>"101001110",
  49235=>"111101111",
  49236=>"110111010",
  49237=>"111000000",
  49238=>"111000110",
  49239=>"110111001",
  49240=>"010011011",
  49241=>"111111110",
  49242=>"000101111",
  49243=>"101011100",
  49244=>"000100101",
  49245=>"100101100",
  49246=>"111110000",
  49247=>"010000100",
  49248=>"000000110",
  49249=>"111101111",
  49250=>"000010110",
  49251=>"101010100",
  49252=>"101010010",
  49253=>"010011000",
  49254=>"110110010",
  49255=>"000000010",
  49256=>"100001010",
  49257=>"110000011",
  49258=>"001101011",
  49259=>"101110111",
  49260=>"000101001",
  49261=>"001000010",
  49262=>"110001101",
  49263=>"000100101",
  49264=>"100111101",
  49265=>"111001111",
  49266=>"001101000",
  49267=>"010111101",
  49268=>"001000000",
  49269=>"111100101",
  49270=>"011101111",
  49271=>"000110101",
  49272=>"000110100",
  49273=>"110101010",
  49274=>"001111010",
  49275=>"100011110",
  49276=>"000100011",
  49277=>"000011110",
  49278=>"010001111",
  49279=>"000000001",
  49280=>"101001001",
  49281=>"111111101",
  49282=>"101011000",
  49283=>"101100000",
  49284=>"101101010",
  49285=>"010000010",
  49286=>"100001110",
  49287=>"110001111",
  49288=>"010000010",
  49289=>"011011111",
  49290=>"111101010",
  49291=>"101011100",
  49292=>"100010000",
  49293=>"001001101",
  49294=>"000001001",
  49295=>"001111001",
  49296=>"001010010",
  49297=>"100111000",
  49298=>"100011001",
  49299=>"101010001",
  49300=>"100001101",
  49301=>"100101011",
  49302=>"010111101",
  49303=>"111110011",
  49304=>"011001001",
  49305=>"111011110",
  49306=>"011100011",
  49307=>"110000000",
  49308=>"001000110",
  49309=>"001110000",
  49310=>"000000010",
  49311=>"010110111",
  49312=>"000011110",
  49313=>"001010010",
  49314=>"000011000",
  49315=>"000001001",
  49316=>"011110011",
  49317=>"001100111",
  49318=>"101010110",
  49319=>"100001000",
  49320=>"000010011",
  49321=>"000011100",
  49322=>"100001000",
  49323=>"000001111",
  49324=>"010111011",
  49325=>"111011111",
  49326=>"100000111",
  49327=>"110010011",
  49328=>"011110110",
  49329=>"011111110",
  49330=>"110101000",
  49331=>"000000101",
  49332=>"011001000",
  49333=>"010001101",
  49334=>"000100100",
  49335=>"101111001",
  49336=>"101000011",
  49337=>"111100111",
  49338=>"101010001",
  49339=>"101100100",
  49340=>"100101010",
  49341=>"101101100",
  49342=>"111100110",
  49343=>"101000010",
  49344=>"011000100",
  49345=>"111010110",
  49346=>"000101001",
  49347=>"001100100",
  49348=>"100010111",
  49349=>"011101111",
  49350=>"001010111",
  49351=>"111010111",
  49352=>"111110000",
  49353=>"110101000",
  49354=>"110011000",
  49355=>"010000111",
  49356=>"010110100",
  49357=>"011000100",
  49358=>"011010110",
  49359=>"110010101",
  49360=>"111111000",
  49361=>"111010110",
  49362=>"010101110",
  49363=>"101010010",
  49364=>"111011111",
  49365=>"000100111",
  49366=>"111001111",
  49367=>"001000000",
  49368=>"110011101",
  49369=>"001011000",
  49370=>"010000111",
  49371=>"101000001",
  49372=>"100110010",
  49373=>"000111110",
  49374=>"101100101",
  49375=>"111100111",
  49376=>"111111100",
  49377=>"000001001",
  49378=>"110001110",
  49379=>"000101001",
  49380=>"101010011",
  49381=>"000001100",
  49382=>"101100101",
  49383=>"001100011",
  49384=>"001111100",
  49385=>"000010000",
  49386=>"100001010",
  49387=>"101011010",
  49388=>"001011000",
  49389=>"011100111",
  49390=>"000000000",
  49391=>"001100000",
  49392=>"001110100",
  49393=>"100010100",
  49394=>"010010010",
  49395=>"010101101",
  49396=>"111011000",
  49397=>"111100100",
  49398=>"011000001",
  49399=>"111101001",
  49400=>"011001001",
  49401=>"101101111",
  49402=>"110001000",
  49403=>"101000101",
  49404=>"001101100",
  49405=>"011000010",
  49406=>"010011000",
  49407=>"110001001",
  49408=>"001011011",
  49409=>"101101010",
  49410=>"111100000",
  49411=>"101111110",
  49412=>"010000100",
  49413=>"100011010",
  49414=>"110011010",
  49415=>"001001001",
  49416=>"100100111",
  49417=>"101000010",
  49418=>"001101011",
  49419=>"000100011",
  49420=>"011111110",
  49421=>"101000110",
  49422=>"001000100",
  49423=>"100100000",
  49424=>"111110111",
  49425=>"111001011",
  49426=>"000000111",
  49427=>"111010010",
  49428=>"011110111",
  49429=>"001011011",
  49430=>"000100110",
  49431=>"110111111",
  49432=>"011011111",
  49433=>"010111010",
  49434=>"100101001",
  49435=>"001100000",
  49436=>"110001111",
  49437=>"101011000",
  49438=>"010110001",
  49439=>"000100010",
  49440=>"010100011",
  49441=>"001001110",
  49442=>"100111000",
  49443=>"010111110",
  49444=>"111101001",
  49445=>"011001100",
  49446=>"100000001",
  49447=>"000010100",
  49448=>"011001110",
  49449=>"111001010",
  49450=>"111001101",
  49451=>"010100100",
  49452=>"111110001",
  49453=>"110010110",
  49454=>"010001011",
  49455=>"110110000",
  49456=>"111101110",
  49457=>"101011011",
  49458=>"111100010",
  49459=>"000010000",
  49460=>"111110111",
  49461=>"111010111",
  49462=>"010111000",
  49463=>"101000110",
  49464=>"011100000",
  49465=>"101011110",
  49466=>"101111101",
  49467=>"001000110",
  49468=>"001001000",
  49469=>"100001100",
  49470=>"110111101",
  49471=>"001100000",
  49472=>"111101110",
  49473=>"010000000",
  49474=>"101111001",
  49475=>"110101110",
  49476=>"101100011",
  49477=>"010110001",
  49478=>"110001100",
  49479=>"011000000",
  49480=>"110000111",
  49481=>"110101011",
  49482=>"100000111",
  49483=>"110001110",
  49484=>"101001000",
  49485=>"001000000",
  49486=>"110010001",
  49487=>"110000110",
  49488=>"101000011",
  49489=>"011101100",
  49490=>"100001000",
  49491=>"101101110",
  49492=>"011111101",
  49493=>"100001110",
  49494=>"000001100",
  49495=>"000101111",
  49496=>"111110100",
  49497=>"011010000",
  49498=>"100101000",
  49499=>"010100000",
  49500=>"101010101",
  49501=>"100001111",
  49502=>"101010100",
  49503=>"001110101",
  49504=>"101100000",
  49505=>"000000111",
  49506=>"000000000",
  49507=>"111011111",
  49508=>"111000111",
  49509=>"111110100",
  49510=>"001110011",
  49511=>"110011110",
  49512=>"100011010",
  49513=>"000111001",
  49514=>"110100101",
  49515=>"100001011",
  49516=>"010101010",
  49517=>"101111111",
  49518=>"101010110",
  49519=>"011000000",
  49520=>"111001001",
  49521=>"000111100",
  49522=>"110110101",
  49523=>"010100010",
  49524=>"011101011",
  49525=>"101001100",
  49526=>"011110011",
  49527=>"101101100",
  49528=>"000001001",
  49529=>"100001101",
  49530=>"000010111",
  49531=>"000100001",
  49532=>"110100101",
  49533=>"100001100",
  49534=>"101010101",
  49535=>"101110111",
  49536=>"010100010",
  49537=>"011001000",
  49538=>"110010100",
  49539=>"111011110",
  49540=>"001101101",
  49541=>"111100101",
  49542=>"000011011",
  49543=>"100110111",
  49544=>"101001101",
  49545=>"000001000",
  49546=>"011101100",
  49547=>"001011000",
  49548=>"101101001",
  49549=>"010001010",
  49550=>"111110111",
  49551=>"010110000",
  49552=>"101001101",
  49553=>"101110100",
  49554=>"111101111",
  49555=>"110000011",
  49556=>"001111111",
  49557=>"000100100",
  49558=>"011111111",
  49559=>"000000000",
  49560=>"001100101",
  49561=>"111011101",
  49562=>"001010111",
  49563=>"010000011",
  49564=>"011000000",
  49565=>"011111101",
  49566=>"010110000",
  49567=>"100111110",
  49568=>"001000110",
  49569=>"100001000",
  49570=>"011011101",
  49571=>"010011010",
  49572=>"110101001",
  49573=>"100001110",
  49574=>"101001111",
  49575=>"110110100",
  49576=>"011000100",
  49577=>"101011010",
  49578=>"101001110",
  49579=>"010101110",
  49580=>"100111100",
  49581=>"000001000",
  49582=>"000001111",
  49583=>"100111111",
  49584=>"111111001",
  49585=>"100001011",
  49586=>"100110110",
  49587=>"001110101",
  49588=>"101100100",
  49589=>"000100110",
  49590=>"111101100",
  49591=>"111001011",
  49592=>"011110100",
  49593=>"000000111",
  49594=>"101001000",
  49595=>"111000010",
  49596=>"110010011",
  49597=>"111010000",
  49598=>"111100111",
  49599=>"011110110",
  49600=>"001011010",
  49601=>"010010011",
  49602=>"110010101",
  49603=>"000010010",
  49604=>"110011100",
  49605=>"010101101",
  49606=>"010110011",
  49607=>"101101110",
  49608=>"001101110",
  49609=>"111110111",
  49610=>"001010110",
  49611=>"000100101",
  49612=>"110000001",
  49613=>"001001011",
  49614=>"000011110",
  49615=>"000101000",
  49616=>"010010100",
  49617=>"100011110",
  49618=>"001010110",
  49619=>"110100101",
  49620=>"000111100",
  49621=>"010101110",
  49622=>"100100011",
  49623=>"111011111",
  49624=>"001011110",
  49625=>"001101011",
  49626=>"001100110",
  49627=>"000111101",
  49628=>"010001101",
  49629=>"101111010",
  49630=>"101110011",
  49631=>"011110001",
  49632=>"100010001",
  49633=>"110101101",
  49634=>"110111111",
  49635=>"011011100",
  49636=>"101100011",
  49637=>"011111110",
  49638=>"101011011",
  49639=>"010011001",
  49640=>"111111000",
  49641=>"101000111",
  49642=>"110000110",
  49643=>"010011001",
  49644=>"111010110",
  49645=>"111101001",
  49646=>"010000110",
  49647=>"101100001",
  49648=>"001000111",
  49649=>"001011000",
  49650=>"001000110",
  49651=>"101111110",
  49652=>"110100110",
  49653=>"001001110",
  49654=>"100100000",
  49655=>"111111101",
  49656=>"110100111",
  49657=>"000001001",
  49658=>"110000110",
  49659=>"010001010",
  49660=>"110101011",
  49661=>"101111101",
  49662=>"101100100",
  49663=>"111110101",
  49664=>"000100101",
  49665=>"001111000",
  49666=>"011000101",
  49667=>"010101111",
  49668=>"110111110",
  49669=>"000100000",
  49670=>"100100100",
  49671=>"101110110",
  49672=>"001011011",
  49673=>"001111110",
  49674=>"010101011",
  49675=>"010010000",
  49676=>"101011011",
  49677=>"000110001",
  49678=>"100000101",
  49679=>"011000110",
  49680=>"100111010",
  49681=>"001011111",
  49682=>"101000000",
  49683=>"000111001",
  49684=>"110001101",
  49685=>"111010110",
  49686=>"001011000",
  49687=>"101100010",
  49688=>"101001000",
  49689=>"000100111",
  49690=>"110010111",
  49691=>"000101011",
  49692=>"010000001",
  49693=>"001000000",
  49694=>"110000110",
  49695=>"110111100",
  49696=>"101111010",
  49697=>"110110100",
  49698=>"001111111",
  49699=>"101010101",
  49700=>"101100111",
  49701=>"000010001",
  49702=>"100010010",
  49703=>"000001010",
  49704=>"111110100",
  49705=>"110111100",
  49706=>"100110010",
  49707=>"100000101",
  49708=>"000001111",
  49709=>"010000111",
  49710=>"001101101",
  49711=>"110100000",
  49712=>"011101011",
  49713=>"001000100",
  49714=>"000100010",
  49715=>"001101011",
  49716=>"010011111",
  49717=>"010010110",
  49718=>"010100001",
  49719=>"110110111",
  49720=>"111111101",
  49721=>"100100010",
  49722=>"101000010",
  49723=>"001011001",
  49724=>"111001100",
  49725=>"000010010",
  49726=>"000111100",
  49727=>"001100010",
  49728=>"111111101",
  49729=>"100111110",
  49730=>"001111010",
  49731=>"101010111",
  49732=>"101010101",
  49733=>"101111010",
  49734=>"001011010",
  49735=>"001011000",
  49736=>"111001110",
  49737=>"000000011",
  49738=>"100001101",
  49739=>"101011111",
  49740=>"101111000",
  49741=>"010000001",
  49742=>"001000101",
  49743=>"000101000",
  49744=>"001000001",
  49745=>"010001001",
  49746=>"000100001",
  49747=>"010010001",
  49748=>"110001010",
  49749=>"110100101",
  49750=>"110101011",
  49751=>"101011001",
  49752=>"011100000",
  49753=>"001011100",
  49754=>"000101100",
  49755=>"011000110",
  49756=>"001111000",
  49757=>"010010100",
  49758=>"001000011",
  49759=>"101011001",
  49760=>"001110000",
  49761=>"010000000",
  49762=>"010010011",
  49763=>"100101010",
  49764=>"001100111",
  49765=>"111001111",
  49766=>"011011000",
  49767=>"110110101",
  49768=>"101110111",
  49769=>"001101001",
  49770=>"001101101",
  49771=>"111001111",
  49772=>"111011110",
  49773=>"100000011",
  49774=>"011100000",
  49775=>"010111111",
  49776=>"111101110",
  49777=>"010010110",
  49778=>"010100101",
  49779=>"000010101",
  49780=>"100110010",
  49781=>"011011000",
  49782=>"110000110",
  49783=>"110000101",
  49784=>"101100110",
  49785=>"000010111",
  49786=>"001000011",
  49787=>"101110010",
  49788=>"001101010",
  49789=>"100101001",
  49790=>"110001010",
  49791=>"000010011",
  49792=>"010001111",
  49793=>"001010111",
  49794=>"011011001",
  49795=>"010001001",
  49796=>"111101000",
  49797=>"100010110",
  49798=>"010001010",
  49799=>"110110110",
  49800=>"001111011",
  49801=>"000010101",
  49802=>"000010110",
  49803=>"100010110",
  49804=>"111000100",
  49805=>"001111011",
  49806=>"100101111",
  49807=>"011000010",
  49808=>"111011110",
  49809=>"010111001",
  49810=>"100000110",
  49811=>"010101001",
  49812=>"100000011",
  49813=>"100111001",
  49814=>"000010001",
  49815=>"000000110",
  49816=>"110110000",
  49817=>"011000101",
  49818=>"100111110",
  49819=>"111011101",
  49820=>"100011101",
  49821=>"111010010",
  49822=>"000010111",
  49823=>"000100100",
  49824=>"000000110",
  49825=>"010011000",
  49826=>"111011110",
  49827=>"111000000",
  49828=>"001101001",
  49829=>"101000100",
  49830=>"110011101",
  49831=>"110000000",
  49832=>"110000110",
  49833=>"110111011",
  49834=>"100101100",
  49835=>"011000001",
  49836=>"111000001",
  49837=>"000100111",
  49838=>"110111001",
  49839=>"111111111",
  49840=>"010000001",
  49841=>"101001110",
  49842=>"110001110",
  49843=>"001010101",
  49844=>"001101010",
  49845=>"100000001",
  49846=>"000011101",
  49847=>"011110110",
  49848=>"100100001",
  49849=>"110011100",
  49850=>"011000000",
  49851=>"110111001",
  49852=>"110001111",
  49853=>"001110101",
  49854=>"111101000",
  49855=>"001110100",
  49856=>"111000111",
  49857=>"011110011",
  49858=>"001101000",
  49859=>"101010010",
  49860=>"010111111",
  49861=>"111011110",
  49862=>"100010011",
  49863=>"011000010",
  49864=>"010001101",
  49865=>"100101000",
  49866=>"010010110",
  49867=>"010000000",
  49868=>"011110010",
  49869=>"111010010",
  49870=>"010101101",
  49871=>"110011011",
  49872=>"010111111",
  49873=>"010000001",
  49874=>"010011001",
  49875=>"000010011",
  49876=>"001101011",
  49877=>"111001110",
  49878=>"000111010",
  49879=>"001001110",
  49880=>"111011101",
  49881=>"000111011",
  49882=>"000000010",
  49883=>"010010111",
  49884=>"011000100",
  49885=>"010110011",
  49886=>"111000011",
  49887=>"001110111",
  49888=>"110011011",
  49889=>"000010010",
  49890=>"111101000",
  49891=>"010011010",
  49892=>"110111110",
  49893=>"110000110",
  49894=>"010000101",
  49895=>"000001101",
  49896=>"011010110",
  49897=>"110001111",
  49898=>"100101110",
  49899=>"110010011",
  49900=>"100000010",
  49901=>"100101010",
  49902=>"100111001",
  49903=>"011101100",
  49904=>"011000001",
  49905=>"010101111",
  49906=>"001101001",
  49907=>"010001010",
  49908=>"111110100",
  49909=>"000110101",
  49910=>"111111111",
  49911=>"000001110",
  49912=>"011001111",
  49913=>"110111000",
  49914=>"110000001",
  49915=>"100000010",
  49916=>"010010000",
  49917=>"100011101",
  49918=>"101100011",
  49919=>"000010111",
  49920=>"111110010",
  49921=>"010111001",
  49922=>"001110001",
  49923=>"111010011",
  49924=>"011011100",
  49925=>"110010000",
  49926=>"010100111",
  49927=>"010101111",
  49928=>"001010011",
  49929=>"011101001",
  49930=>"111101111",
  49931=>"111111010",
  49932=>"010110101",
  49933=>"000010100",
  49934=>"000111000",
  49935=>"000111000",
  49936=>"000100000",
  49937=>"101100001",
  49938=>"101110001",
  49939=>"110001000",
  49940=>"011111111",
  49941=>"110101000",
  49942=>"110100000",
  49943=>"111101010",
  49944=>"000001010",
  49945=>"101001110",
  49946=>"110010011",
  49947=>"110011001",
  49948=>"001001011",
  49949=>"111100010",
  49950=>"111100110",
  49951=>"110001000",
  49952=>"111110111",
  49953=>"101001100",
  49954=>"100010100",
  49955=>"111111111",
  49956=>"110110010",
  49957=>"001100011",
  49958=>"100110101",
  49959=>"010111111",
  49960=>"110001111",
  49961=>"101100000",
  49962=>"010100100",
  49963=>"110010100",
  49964=>"001000100",
  49965=>"101111011",
  49966=>"010110111",
  49967=>"100000110",
  49968=>"010101000",
  49969=>"110111110",
  49970=>"101100001",
  49971=>"100111100",
  49972=>"101001001",
  49973=>"100100100",
  49974=>"101111001",
  49975=>"001110111",
  49976=>"010100100",
  49977=>"011000101",
  49978=>"011000101",
  49979=>"011011010",
  49980=>"101010000",
  49981=>"110101111",
  49982=>"101010010",
  49983=>"100111100",
  49984=>"110110111",
  49985=>"001110101",
  49986=>"011101100",
  49987=>"111110110",
  49988=>"101011111",
  49989=>"000111001",
  49990=>"100011000",
  49991=>"110111010",
  49992=>"011110001",
  49993=>"110111101",
  49994=>"110000011",
  49995=>"100001100",
  49996=>"001011100",
  49997=>"000001011",
  49998=>"111011011",
  49999=>"011000000",
  50000=>"110000111",
  50001=>"111111010",
  50002=>"100000010",
  50003=>"100100001",
  50004=>"100110000",
  50005=>"100000101",
  50006=>"110011001",
  50007=>"110110101",
  50008=>"110011100",
  50009=>"110110011",
  50010=>"100000111",
  50011=>"101100010",
  50012=>"100001011",
  50013=>"111111100",
  50014=>"111010001",
  50015=>"110111011",
  50016=>"011101010",
  50017=>"010010111",
  50018=>"000110011",
  50019=>"111111011",
  50020=>"111110001",
  50021=>"111101011",
  50022=>"011001010",
  50023=>"100010000",
  50024=>"110010000",
  50025=>"101101010",
  50026=>"110010001",
  50027=>"100100001",
  50028=>"111100101",
  50029=>"110110111",
  50030=>"111100010",
  50031=>"111100101",
  50032=>"110001111",
  50033=>"100001000",
  50034=>"110001001",
  50035=>"010011011",
  50036=>"111101110",
  50037=>"000110001",
  50038=>"101111111",
  50039=>"100111100",
  50040=>"101011111",
  50041=>"010100001",
  50042=>"001111000",
  50043=>"001001000",
  50044=>"000101110",
  50045=>"000110000",
  50046=>"100000010",
  50047=>"101001010",
  50048=>"011000111",
  50049=>"000000101",
  50050=>"011111111",
  50051=>"111111101",
  50052=>"111101010",
  50053=>"011000101",
  50054=>"110110000",
  50055=>"010110100",
  50056=>"110111011",
  50057=>"011101010",
  50058=>"001000111",
  50059=>"100011000",
  50060=>"000111100",
  50061=>"111101000",
  50062=>"111110111",
  50063=>"101001001",
  50064=>"100111101",
  50065=>"110110100",
  50066=>"100000010",
  50067=>"001001101",
  50068=>"110000101",
  50069=>"111001011",
  50070=>"001101101",
  50071=>"111011010",
  50072=>"011010111",
  50073=>"000010111",
  50074=>"000100101",
  50075=>"110101000",
  50076=>"011110010",
  50077=>"100100000",
  50078=>"011101001",
  50079=>"011011010",
  50080=>"100000011",
  50081=>"101101111",
  50082=>"010101100",
  50083=>"010100010",
  50084=>"100010100",
  50085=>"010100100",
  50086=>"011111010",
  50087=>"011111111",
  50088=>"011110111",
  50089=>"000000000",
  50090=>"110111101",
  50091=>"100001111",
  50092=>"011110011",
  50093=>"111011011",
  50094=>"010100111",
  50095=>"110111100",
  50096=>"110010001",
  50097=>"000001010",
  50098=>"110111010",
  50099=>"101110101",
  50100=>"000100001",
  50101=>"111001000",
  50102=>"000101000",
  50103=>"000000011",
  50104=>"110111000",
  50105=>"110111011",
  50106=>"111011111",
  50107=>"001111100",
  50108=>"100100000",
  50109=>"100001001",
  50110=>"010011111",
  50111=>"110001111",
  50112=>"101010000",
  50113=>"111011111",
  50114=>"110101101",
  50115=>"111011010",
  50116=>"000110100",
  50117=>"011110000",
  50118=>"100001000",
  50119=>"110011011",
  50120=>"001111011",
  50121=>"011110000",
  50122=>"001000100",
  50123=>"100111101",
  50124=>"000110000",
  50125=>"010100100",
  50126=>"111100111",
  50127=>"101010100",
  50128=>"010000100",
  50129=>"101010110",
  50130=>"100100100",
  50131=>"101110001",
  50132=>"110011010",
  50133=>"011100100",
  50134=>"011110011",
  50135=>"101101100",
  50136=>"001100001",
  50137=>"010101000",
  50138=>"000000010",
  50139=>"110101100",
  50140=>"010000000",
  50141=>"000111110",
  50142=>"110110111",
  50143=>"001110001",
  50144=>"011110001",
  50145=>"001000000",
  50146=>"000010101",
  50147=>"110010010",
  50148=>"111101111",
  50149=>"011000110",
  50150=>"111100010",
  50151=>"011011000",
  50152=>"011000010",
  50153=>"011100000",
  50154=>"111111100",
  50155=>"111110011",
  50156=>"111100010",
  50157=>"100011011",
  50158=>"110001110",
  50159=>"110111001",
  50160=>"101010000",
  50161=>"101110100",
  50162=>"011101100",
  50163=>"111101111",
  50164=>"111111111",
  50165=>"101011110",
  50166=>"111101100",
  50167=>"111101000",
  50168=>"011101101",
  50169=>"100011110",
  50170=>"110101010",
  50171=>"000101011",
  50172=>"000000000",
  50173=>"001011001",
  50174=>"011011001",
  50175=>"001111010",
  50176=>"010010010",
  50177=>"001000111",
  50178=>"100001000",
  50179=>"001011000",
  50180=>"100011110",
  50181=>"001011101",
  50182=>"000000101",
  50183=>"001110011",
  50184=>"010111000",
  50185=>"011010000",
  50186=>"111111101",
  50187=>"100000100",
  50188=>"010100110",
  50189=>"110010000",
  50190=>"100101000",
  50191=>"000111011",
  50192=>"000100101",
  50193=>"100001111",
  50194=>"100110000",
  50195=>"011101011",
  50196=>"100000010",
  50197=>"010100001",
  50198=>"110110000",
  50199=>"011001010",
  50200=>"100010010",
  50201=>"111100111",
  50202=>"100001100",
  50203=>"110001100",
  50204=>"111001111",
  50205=>"011111000",
  50206=>"011000010",
  50207=>"100110111",
  50208=>"011000010",
  50209=>"000101110",
  50210=>"011000101",
  50211=>"101011110",
  50212=>"100001011",
  50213=>"010110111",
  50214=>"110010010",
  50215=>"111011011",
  50216=>"000101000",
  50217=>"010100011",
  50218=>"011100011",
  50219=>"001001110",
  50220=>"000111010",
  50221=>"111111000",
  50222=>"111100000",
  50223=>"000000101",
  50224=>"111111101",
  50225=>"111011001",
  50226=>"010001011",
  50227=>"110011101",
  50228=>"011111110",
  50229=>"110100101",
  50230=>"110100110",
  50231=>"111111010",
  50232=>"000000110",
  50233=>"011100011",
  50234=>"001101111",
  50235=>"101110110",
  50236=>"111111101",
  50237=>"111111000",
  50238=>"011110011",
  50239=>"011111110",
  50240=>"001010101",
  50241=>"100111111",
  50242=>"101101001",
  50243=>"110001000",
  50244=>"010101111",
  50245=>"100000111",
  50246=>"111111001",
  50247=>"000011101",
  50248=>"101000000",
  50249=>"100010000",
  50250=>"100101110",
  50251=>"110101101",
  50252=>"000111110",
  50253=>"101011010",
  50254=>"010011101",
  50255=>"010000010",
  50256=>"110010010",
  50257=>"100101100",
  50258=>"101111101",
  50259=>"011101101",
  50260=>"000001010",
  50261=>"011111101",
  50262=>"010001010",
  50263=>"001110111",
  50264=>"000000110",
  50265=>"111000110",
  50266=>"100101111",
  50267=>"000010000",
  50268=>"000111000",
  50269=>"111011100",
  50270=>"111001110",
  50271=>"110110110",
  50272=>"010010011",
  50273=>"011001001",
  50274=>"110111001",
  50275=>"000000110",
  50276=>"000101101",
  50277=>"011001000",
  50278=>"101011101",
  50279=>"001001110",
  50280=>"011100100",
  50281=>"010000110",
  50282=>"011001011",
  50283=>"001000100",
  50284=>"011011001",
  50285=>"101100010",
  50286=>"101000110",
  50287=>"111111010",
  50288=>"100110111",
  50289=>"111010100",
  50290=>"001100001",
  50291=>"001101111",
  50292=>"011111111",
  50293=>"111001111",
  50294=>"011100011",
  50295=>"001001001",
  50296=>"001111001",
  50297=>"100101111",
  50298=>"000001010",
  50299=>"101101011",
  50300=>"110000101",
  50301=>"001000111",
  50302=>"110100000",
  50303=>"010100001",
  50304=>"110000011",
  50305=>"100101001",
  50306=>"110111011",
  50307=>"110000110",
  50308=>"101110110",
  50309=>"011000101",
  50310=>"000011100",
  50311=>"010111110",
  50312=>"011101101",
  50313=>"101100110",
  50314=>"100100010",
  50315=>"001110001",
  50316=>"001000100",
  50317=>"110000000",
  50318=>"111110101",
  50319=>"011101001",
  50320=>"111010011",
  50321=>"011110001",
  50322=>"000001111",
  50323=>"100010011",
  50324=>"001101000",
  50325=>"101111100",
  50326=>"111100101",
  50327=>"101101100",
  50328=>"100100111",
  50329=>"110111111",
  50330=>"110111000",
  50331=>"001110000",
  50332=>"000010001",
  50333=>"000111110",
  50334=>"001110101",
  50335=>"110100001",
  50336=>"000100000",
  50337=>"011111001",
  50338=>"011000001",
  50339=>"001001000",
  50340=>"100101111",
  50341=>"001011001",
  50342=>"000110111",
  50343=>"001010010",
  50344=>"011101111",
  50345=>"111010011",
  50346=>"100011011",
  50347=>"001100001",
  50348=>"100111111",
  50349=>"101101111",
  50350=>"110110010",
  50351=>"111011000",
  50352=>"110001111",
  50353=>"110011001",
  50354=>"110001100",
  50355=>"111110011",
  50356=>"100100100",
  50357=>"111000101",
  50358=>"000111000",
  50359=>"101000000",
  50360=>"100010110",
  50361=>"010110110",
  50362=>"100111100",
  50363=>"100101000",
  50364=>"000101000",
  50365=>"100110010",
  50366=>"000000000",
  50367=>"100000111",
  50368=>"000110001",
  50369=>"101101110",
  50370=>"110011011",
  50371=>"101100100",
  50372=>"111101010",
  50373=>"100011000",
  50374=>"000100011",
  50375=>"100011010",
  50376=>"111010010",
  50377=>"010011111",
  50378=>"000110010",
  50379=>"011010000",
  50380=>"011111101",
  50381=>"001001000",
  50382=>"100000010",
  50383=>"110100110",
  50384=>"001111011",
  50385=>"001100111",
  50386=>"010110001",
  50387=>"010011110",
  50388=>"000101111",
  50389=>"110011100",
  50390=>"000111111",
  50391=>"111001100",
  50392=>"010101011",
  50393=>"111010101",
  50394=>"001011111",
  50395=>"101000001",
  50396=>"001100001",
  50397=>"110000101",
  50398=>"110100001",
  50399=>"111110000",
  50400=>"111000101",
  50401=>"100100011",
  50402=>"110010001",
  50403=>"101110100",
  50404=>"111111100",
  50405=>"001111101",
  50406=>"100110001",
  50407=>"010111000",
  50408=>"110010011",
  50409=>"101000101",
  50410=>"100010001",
  50411=>"101111111",
  50412=>"000011100",
  50413=>"001010111",
  50414=>"110000011",
  50415=>"011111111",
  50416=>"110100000",
  50417=>"011000100",
  50418=>"100101101",
  50419=>"111001110",
  50420=>"101100111",
  50421=>"001000101",
  50422=>"111101001",
  50423=>"011010110",
  50424=>"000101101",
  50425=>"010110101",
  50426=>"111011001",
  50427=>"010111110",
  50428=>"010110111",
  50429=>"101011000",
  50430=>"101011100",
  50431=>"110101011",
  50432=>"000111110",
  50433=>"010111000",
  50434=>"011110111",
  50435=>"110010111",
  50436=>"001111100",
  50437=>"111110001",
  50438=>"100000111",
  50439=>"000111100",
  50440=>"111100001",
  50441=>"100010000",
  50442=>"000101001",
  50443=>"010101001",
  50444=>"101000100",
  50445=>"000111110",
  50446=>"000100010",
  50447=>"100100100",
  50448=>"111010101",
  50449=>"110101101",
  50450=>"101001100",
  50451=>"011010111",
  50452=>"001011111",
  50453=>"001010111",
  50454=>"111010100",
  50455=>"101000000",
  50456=>"111011001",
  50457=>"111011110",
  50458=>"000010001",
  50459=>"001101111",
  50460=>"001111000",
  50461=>"101001011",
  50462=>"001110100",
  50463=>"010000000",
  50464=>"100111110",
  50465=>"110010000",
  50466=>"101010001",
  50467=>"111101000",
  50468=>"011000010",
  50469=>"101111001",
  50470=>"100110011",
  50471=>"101100101",
  50472=>"011001101",
  50473=>"101101111",
  50474=>"001111011",
  50475=>"100110010",
  50476=>"011110000",
  50477=>"010010110",
  50478=>"111110001",
  50479=>"011101010",
  50480=>"000010010",
  50481=>"111100100",
  50482=>"001100100",
  50483=>"111100011",
  50484=>"001011110",
  50485=>"000001100",
  50486=>"000101001",
  50487=>"101101111",
  50488=>"100101010",
  50489=>"011001110",
  50490=>"000010001",
  50491=>"011111000",
  50492=>"110010100",
  50493=>"000000101",
  50494=>"010101010",
  50495=>"010111011",
  50496=>"010010111",
  50497=>"101101111",
  50498=>"101001010",
  50499=>"000001000",
  50500=>"011101111",
  50501=>"011101010",
  50502=>"100000000",
  50503=>"111010011",
  50504=>"101100000",
  50505=>"000100000",
  50506=>"111110100",
  50507=>"001101011",
  50508=>"101110001",
  50509=>"000011011",
  50510=>"101101011",
  50511=>"101111110",
  50512=>"010111001",
  50513=>"000110010",
  50514=>"010001101",
  50515=>"100101001",
  50516=>"010111101",
  50517=>"100011110",
  50518=>"111101001",
  50519=>"011011001",
  50520=>"111110101",
  50521=>"111101101",
  50522=>"001010111",
  50523=>"010110101",
  50524=>"000011110",
  50525=>"110011111",
  50526=>"100101101",
  50527=>"000000000",
  50528=>"101110011",
  50529=>"111011001",
  50530=>"000000010",
  50531=>"101101101",
  50532=>"010110110",
  50533=>"000010011",
  50534=>"110101100",
  50535=>"100001100",
  50536=>"110101000",
  50537=>"111001100",
  50538=>"110000111",
  50539=>"011010110",
  50540=>"101110111",
  50541=>"010000011",
  50542=>"000100110",
  50543=>"111101111",
  50544=>"000000001",
  50545=>"110011111",
  50546=>"111111101",
  50547=>"100000101",
  50548=>"101001111",
  50549=>"010010000",
  50550=>"100010000",
  50551=>"100010000",
  50552=>"000110011",
  50553=>"010011011",
  50554=>"000001111",
  50555=>"111011100",
  50556=>"110100101",
  50557=>"111010100",
  50558=>"111010001",
  50559=>"001100111",
  50560=>"111100101",
  50561=>"000110001",
  50562=>"100010000",
  50563=>"000111001",
  50564=>"110000010",
  50565=>"110110101",
  50566=>"000110001",
  50567=>"110100010",
  50568=>"101111000",
  50569=>"111011010",
  50570=>"011010110",
  50571=>"000000001",
  50572=>"110011100",
  50573=>"101111000",
  50574=>"101100101",
  50575=>"111110110",
  50576=>"010101101",
  50577=>"010100000",
  50578=>"111001100",
  50579=>"100111000",
  50580=>"111000000",
  50581=>"111100111",
  50582=>"101100011",
  50583=>"111011101",
  50584=>"010001000",
  50585=>"010000000",
  50586=>"010100110",
  50587=>"010111100",
  50588=>"001010111",
  50589=>"000101000",
  50590=>"111111001",
  50591=>"110000111",
  50592=>"001111010",
  50593=>"110011000",
  50594=>"111111111",
  50595=>"100101100",
  50596=>"100100001",
  50597=>"111011100",
  50598=>"011000100",
  50599=>"000111100",
  50600=>"011110010",
  50601=>"011000000",
  50602=>"001001000",
  50603=>"000011010",
  50604=>"111111101",
  50605=>"110010110",
  50606=>"101000011",
  50607=>"110101101",
  50608=>"001000000",
  50609=>"011011110",
  50610=>"000110000",
  50611=>"101000011",
  50612=>"100101011",
  50613=>"001111100",
  50614=>"101000111",
  50615=>"001101010",
  50616=>"101001110",
  50617=>"001100101",
  50618=>"111011000",
  50619=>"101101110",
  50620=>"101010101",
  50621=>"010111000",
  50622=>"101101000",
  50623=>"010100001",
  50624=>"100001010",
  50625=>"001111000",
  50626=>"010001000",
  50627=>"110110100",
  50628=>"111111001",
  50629=>"001000000",
  50630=>"010000101",
  50631=>"101010100",
  50632=>"100000011",
  50633=>"110000011",
  50634=>"001000111",
  50635=>"000011000",
  50636=>"100111001",
  50637=>"000111111",
  50638=>"110111000",
  50639=>"110111100",
  50640=>"100101111",
  50641=>"010011001",
  50642=>"101010001",
  50643=>"000000110",
  50644=>"110000101",
  50645=>"101001100",
  50646=>"001000010",
  50647=>"010001000",
  50648=>"100110010",
  50649=>"010000000",
  50650=>"101110110",
  50651=>"101101011",
  50652=>"000000010",
  50653=>"010001010",
  50654=>"011111010",
  50655=>"001011010",
  50656=>"111100000",
  50657=>"100110001",
  50658=>"010001000",
  50659=>"011001001",
  50660=>"110101010",
  50661=>"000100010",
  50662=>"110011011",
  50663=>"100100100",
  50664=>"000000111",
  50665=>"011001110",
  50666=>"010011001",
  50667=>"101001010",
  50668=>"011000100",
  50669=>"010011100",
  50670=>"000001110",
  50671=>"110110100",
  50672=>"000001011",
  50673=>"010111111",
  50674=>"010011010",
  50675=>"001001110",
  50676=>"001010000",
  50677=>"010110101",
  50678=>"000100011",
  50679=>"011010001",
  50680=>"110110010",
  50681=>"010001010",
  50682=>"111111011",
  50683=>"101011110",
  50684=>"010001101",
  50685=>"111010011",
  50686=>"011101011",
  50687=>"010110100",
  50688=>"111111000",
  50689=>"111011010",
  50690=>"010111001",
  50691=>"111100111",
  50692=>"000000010",
  50693=>"001100001",
  50694=>"011101010",
  50695=>"110010101",
  50696=>"000000001",
  50697=>"011011001",
  50698=>"111010010",
  50699=>"100000000",
  50700=>"100010001",
  50701=>"100100000",
  50702=>"001110000",
  50703=>"001100000",
  50704=>"010000011",
  50705=>"111001111",
  50706=>"111000101",
  50707=>"101110011",
  50708=>"001011111",
  50709=>"111010011",
  50710=>"001100111",
  50711=>"001010111",
  50712=>"011001110",
  50713=>"010011011",
  50714=>"000001000",
  50715=>"000101100",
  50716=>"111100001",
  50717=>"100100111",
  50718=>"110110011",
  50719=>"011001001",
  50720=>"100100111",
  50721=>"111101101",
  50722=>"000010001",
  50723=>"101110110",
  50724=>"011001101",
  50725=>"101110011",
  50726=>"011010010",
  50727=>"011100100",
  50728=>"001100101",
  50729=>"101011011",
  50730=>"000000000",
  50731=>"011011010",
  50732=>"000000100",
  50733=>"110010101",
  50734=>"001110000",
  50735=>"000111101",
  50736=>"100111100",
  50737=>"011101000",
  50738=>"111101011",
  50739=>"111001111",
  50740=>"011111011",
  50741=>"111001001",
  50742=>"011001110",
  50743=>"101011001",
  50744=>"110110111",
  50745=>"110011000",
  50746=>"100111100",
  50747=>"101111111",
  50748=>"001110010",
  50749=>"010010111",
  50750=>"010000110",
  50751=>"011010111",
  50752=>"111111111",
  50753=>"010011011",
  50754=>"101111110",
  50755=>"100000111",
  50756=>"010110101",
  50757=>"000011010",
  50758=>"101000010",
  50759=>"010001011",
  50760=>"000010000",
  50761=>"101101001",
  50762=>"101111110",
  50763=>"100111111",
  50764=>"011010000",
  50765=>"110101100",
  50766=>"101111111",
  50767=>"111111000",
  50768=>"110010110",
  50769=>"100000100",
  50770=>"000011001",
  50771=>"000001101",
  50772=>"110001111",
  50773=>"001001111",
  50774=>"100000100",
  50775=>"000110101",
  50776=>"110011000",
  50777=>"010110000",
  50778=>"011001111",
  50779=>"111100110",
  50780=>"101111000",
  50781=>"010101010",
  50782=>"001001111",
  50783=>"001001100",
  50784=>"000101100",
  50785=>"111000100",
  50786=>"010101011",
  50787=>"111001011",
  50788=>"001010010",
  50789=>"001110111",
  50790=>"010111111",
  50791=>"101011100",
  50792=>"000111000",
  50793=>"001001001",
  50794=>"000011110",
  50795=>"010011110",
  50796=>"010001001",
  50797=>"110100000",
  50798=>"101011101",
  50799=>"010001101",
  50800=>"010011100",
  50801=>"101001101",
  50802=>"101011011",
  50803=>"110000111",
  50804=>"100100100",
  50805=>"000111111",
  50806=>"111111001",
  50807=>"010011011",
  50808=>"011101011",
  50809=>"010100001",
  50810=>"100010111",
  50811=>"011000100",
  50812=>"100111100",
  50813=>"101001110",
  50814=>"110110011",
  50815=>"111110111",
  50816=>"111110111",
  50817=>"100111010",
  50818=>"111000011",
  50819=>"111100011",
  50820=>"011011011",
  50821=>"110100101",
  50822=>"101110011",
  50823=>"011100110",
  50824=>"111010101",
  50825=>"001011000",
  50826=>"010110011",
  50827=>"111110011",
  50828=>"110000100",
  50829=>"111010110",
  50830=>"111001100",
  50831=>"101111101",
  50832=>"011011011",
  50833=>"010100010",
  50834=>"101000111",
  50835=>"110101101",
  50836=>"011110100",
  50837=>"111010111",
  50838=>"111100110",
  50839=>"101000100",
  50840=>"101000000",
  50841=>"111011100",
  50842=>"011110011",
  50843=>"110010100",
  50844=>"001010011",
  50845=>"110110101",
  50846=>"011111110",
  50847=>"111011101",
  50848=>"111100101",
  50849=>"100101001",
  50850=>"001000000",
  50851=>"010111111",
  50852=>"110110101",
  50853=>"010010100",
  50854=>"011011110",
  50855=>"100011000",
  50856=>"101000110",
  50857=>"111010101",
  50858=>"010101100",
  50859=>"011101110",
  50860=>"010000111",
  50861=>"011111000",
  50862=>"100010001",
  50863=>"001100011",
  50864=>"011010010",
  50865=>"101110001",
  50866=>"010110001",
  50867=>"110011000",
  50868=>"010100100",
  50869=>"101110000",
  50870=>"101010101",
  50871=>"110010111",
  50872=>"101111101",
  50873=>"100000110",
  50874=>"001100101",
  50875=>"110001100",
  50876=>"111010110",
  50877=>"010110011",
  50878=>"001000011",
  50879=>"011011010",
  50880=>"010111100",
  50881=>"010110011",
  50882=>"101000111",
  50883=>"011100100",
  50884=>"101001000",
  50885=>"001110101",
  50886=>"010001100",
  50887=>"001110011",
  50888=>"101000000",
  50889=>"010101100",
  50890=>"100010100",
  50891=>"110100011",
  50892=>"010001100",
  50893=>"101110000",
  50894=>"100000001",
  50895=>"101100011",
  50896=>"101011011",
  50897=>"101101001",
  50898=>"010011111",
  50899=>"000100110",
  50900=>"011000000",
  50901=>"000000110",
  50902=>"101100101",
  50903=>"011001010",
  50904=>"010000100",
  50905=>"011010000",
  50906=>"001001011",
  50907=>"110110100",
  50908=>"101001011",
  50909=>"010100001",
  50910=>"110101001",
  50911=>"111110101",
  50912=>"101011101",
  50913=>"010001000",
  50914=>"010100111",
  50915=>"011100010",
  50916=>"100110111",
  50917=>"100101001",
  50918=>"011011011",
  50919=>"100111110",
  50920=>"000110110",
  50921=>"111001000",
  50922=>"100010110",
  50923=>"110011001",
  50924=>"100000110",
  50925=>"011110100",
  50926=>"101110001",
  50927=>"101101110",
  50928=>"100010101",
  50929=>"100110110",
  50930=>"100001110",
  50931=>"001101100",
  50932=>"011111011",
  50933=>"010001101",
  50934=>"111101000",
  50935=>"000100110",
  50936=>"010000111",
  50937=>"110101000",
  50938=>"000010100",
  50939=>"110000001",
  50940=>"110000010",
  50941=>"011010001",
  50942=>"111101011",
  50943=>"100010111",
  50944=>"110010100",
  50945=>"100000001",
  50946=>"011001000",
  50947=>"010000011",
  50948=>"000101010",
  50949=>"010011110",
  50950=>"010100010",
  50951=>"000001000",
  50952=>"101010111",
  50953=>"011000111",
  50954=>"101000001",
  50955=>"000001101",
  50956=>"011000100",
  50957=>"000111001",
  50958=>"111111110",
  50959=>"011010101",
  50960=>"101100000",
  50961=>"110001101",
  50962=>"100101001",
  50963=>"001101100",
  50964=>"101010010",
  50965=>"011101011",
  50966=>"110100101",
  50967=>"111110110",
  50968=>"000110011",
  50969=>"111101110",
  50970=>"000010010",
  50971=>"001000010",
  50972=>"010110110",
  50973=>"010011101",
  50974=>"101110100",
  50975=>"010010110",
  50976=>"001110100",
  50977=>"110011000",
  50978=>"000000011",
  50979=>"110000000",
  50980=>"100111000",
  50981=>"100001100",
  50982=>"111100111",
  50983=>"001011011",
  50984=>"110011111",
  50985=>"000001101",
  50986=>"001100111",
  50987=>"111110111",
  50988=>"011000101",
  50989=>"000011101",
  50990=>"000110001",
  50991=>"111101011",
  50992=>"010001001",
  50993=>"000101000",
  50994=>"001101110",
  50995=>"111101111",
  50996=>"001000101",
  50997=>"111110111",
  50998=>"100111000",
  50999=>"110010000",
  51000=>"001010111",
  51001=>"000101111",
  51002=>"100011001",
  51003=>"001110011",
  51004=>"110011010",
  51005=>"100011111",
  51006=>"101101000",
  51007=>"000110000",
  51008=>"011001001",
  51009=>"011111000",
  51010=>"100111101",
  51011=>"011010111",
  51012=>"100110101",
  51013=>"001100111",
  51014=>"100111011",
  51015=>"010100001",
  51016=>"011000011",
  51017=>"111101111",
  51018=>"010100100",
  51019=>"011100110",
  51020=>"010101011",
  51021=>"101010101",
  51022=>"100000101",
  51023=>"010110111",
  51024=>"010010000",
  51025=>"111001111",
  51026=>"011101111",
  51027=>"110010101",
  51028=>"101001110",
  51029=>"010010011",
  51030=>"111110000",
  51031=>"010011010",
  51032=>"101010010",
  51033=>"100011110",
  51034=>"110100101",
  51035=>"101101111",
  51036=>"000100000",
  51037=>"110001101",
  51038=>"000011111",
  51039=>"001011110",
  51040=>"011111000",
  51041=>"110110110",
  51042=>"110001011",
  51043=>"000010110",
  51044=>"010110100",
  51045=>"100101010",
  51046=>"111100000",
  51047=>"101111000",
  51048=>"001000100",
  51049=>"111111101",
  51050=>"100110100",
  51051=>"000111011",
  51052=>"100100101",
  51053=>"110101100",
  51054=>"001011001",
  51055=>"110101001",
  51056=>"001010001",
  51057=>"110110010",
  51058=>"000101100",
  51059=>"100010110",
  51060=>"000111011",
  51061=>"010111011",
  51062=>"110000000",
  51063=>"101001011",
  51064=>"000100110",
  51065=>"011011111",
  51066=>"100100000",
  51067=>"000010110",
  51068=>"000110010",
  51069=>"101110110",
  51070=>"100011010",
  51071=>"110000001",
  51072=>"001001011",
  51073=>"110100001",
  51074=>"110100100",
  51075=>"111100000",
  51076=>"110001110",
  51077=>"101010101",
  51078=>"110010101",
  51079=>"111000100",
  51080=>"110110100",
  51081=>"001101001",
  51082=>"000110101",
  51083=>"111001001",
  51084=>"011011111",
  51085=>"010100000",
  51086=>"110010011",
  51087=>"101011011",
  51088=>"110111010",
  51089=>"100111111",
  51090=>"100000001",
  51091=>"011111100",
  51092=>"001110101",
  51093=>"111011001",
  51094=>"110111100",
  51095=>"101010001",
  51096=>"001101101",
  51097=>"010011101",
  51098=>"010110010",
  51099=>"010001011",
  51100=>"001111110",
  51101=>"111110110",
  51102=>"010000110",
  51103=>"010001010",
  51104=>"100001111",
  51105=>"010010011",
  51106=>"000110100",
  51107=>"000001100",
  51108=>"011110100",
  51109=>"011100010",
  51110=>"000000010",
  51111=>"010000010",
  51112=>"010011011",
  51113=>"011011010",
  51114=>"011110001",
  51115=>"001101001",
  51116=>"110100101",
  51117=>"000010110",
  51118=>"110101001",
  51119=>"101011111",
  51120=>"100110010",
  51121=>"011101110",
  51122=>"110100110",
  51123=>"001010011",
  51124=>"111101110",
  51125=>"011010001",
  51126=>"110100110",
  51127=>"110111110",
  51128=>"000000101",
  51129=>"101011001",
  51130=>"110010101",
  51131=>"110110100",
  51132=>"000100001",
  51133=>"000000110",
  51134=>"101111101",
  51135=>"011111100",
  51136=>"001000111",
  51137=>"010010101",
  51138=>"100000101",
  51139=>"100100111",
  51140=>"011111100",
  51141=>"101011010",
  51142=>"111101101",
  51143=>"010100111",
  51144=>"001010100",
  51145=>"110111000",
  51146=>"100100100",
  51147=>"011110010",
  51148=>"110100100",
  51149=>"110001000",
  51150=>"101001111",
  51151=>"000011000",
  51152=>"110101111",
  51153=>"101000100",
  51154=>"000000100",
  51155=>"010010111",
  51156=>"101010010",
  51157=>"000101111",
  51158=>"010100001",
  51159=>"000100010",
  51160=>"010101001",
  51161=>"110100110",
  51162=>"111110000",
  51163=>"001011100",
  51164=>"100000110",
  51165=>"111110100",
  51166=>"110000000",
  51167=>"110000010",
  51168=>"001100000",
  51169=>"111101110",
  51170=>"011010111",
  51171=>"001111001",
  51172=>"011001110",
  51173=>"101111000",
  51174=>"100000101",
  51175=>"100011011",
  51176=>"011000010",
  51177=>"011101010",
  51178=>"010000011",
  51179=>"101101001",
  51180=>"110100101",
  51181=>"001110111",
  51182=>"010100100",
  51183=>"101100000",
  51184=>"010100010",
  51185=>"011011000",
  51186=>"010111111",
  51187=>"111101011",
  51188=>"111010011",
  51189=>"100010000",
  51190=>"111101001",
  51191=>"111100011",
  51192=>"111001110",
  51193=>"111010110",
  51194=>"010011100",
  51195=>"111100000",
  51196=>"001001101",
  51197=>"000001111",
  51198=>"000001011",
  51199=>"101100110",
  51200=>"111011000",
  51201=>"011000010",
  51202=>"111110100",
  51203=>"110100111",
  51204=>"010101100",
  51205=>"101101110",
  51206=>"100010100",
  51207=>"001111100",
  51208=>"110111001",
  51209=>"111111110",
  51210=>"101100111",
  51211=>"101111010",
  51212=>"100111000",
  51213=>"111000100",
  51214=>"101110001",
  51215=>"000101111",
  51216=>"011111011",
  51217=>"001100111",
  51218=>"100011001",
  51219=>"101011000",
  51220=>"101000111",
  51221=>"111000011",
  51222=>"110111101",
  51223=>"001100111",
  51224=>"010001110",
  51225=>"111111010",
  51226=>"011100110",
  51227=>"011111110",
  51228=>"101101111",
  51229=>"001100000",
  51230=>"111011000",
  51231=>"111101110",
  51232=>"001011101",
  51233=>"011001010",
  51234=>"010010010",
  51235=>"001010011",
  51236=>"110111101",
  51237=>"011111010",
  51238=>"010000010",
  51239=>"110011011",
  51240=>"101111111",
  51241=>"010100100",
  51242=>"010001011",
  51243=>"010111110",
  51244=>"000111011",
  51245=>"100100111",
  51246=>"100000101",
  51247=>"110001000",
  51248=>"101110011",
  51249=>"101001110",
  51250=>"110000100",
  51251=>"111010011",
  51252=>"010001111",
  51253=>"001010001",
  51254=>"110111111",
  51255=>"110001110",
  51256=>"011100001",
  51257=>"110110111",
  51258=>"100010101",
  51259=>"111101100",
  51260=>"111111100",
  51261=>"111101000",
  51262=>"010101111",
  51263=>"100110101",
  51264=>"001000111",
  51265=>"100101000",
  51266=>"000101000",
  51267=>"011010100",
  51268=>"000010011",
  51269=>"110111111",
  51270=>"011100100",
  51271=>"001110010",
  51272=>"101111001",
  51273=>"110010100",
  51274=>"000101010",
  51275=>"010010010",
  51276=>"010100001",
  51277=>"100110001",
  51278=>"110001011",
  51279=>"100101001",
  51280=>"100111100",
  51281=>"110000000",
  51282=>"011100100",
  51283=>"100001110",
  51284=>"001000110",
  51285=>"111000000",
  51286=>"000111001",
  51287=>"100101110",
  51288=>"111011111",
  51289=>"000110101",
  51290=>"100000001",
  51291=>"010010111",
  51292=>"000011011",
  51293=>"010001001",
  51294=>"111001000",
  51295=>"101011011",
  51296=>"000110000",
  51297=>"111101101",
  51298=>"011010011",
  51299=>"011011011",
  51300=>"111001101",
  51301=>"000010001",
  51302=>"000100000",
  51303=>"000011011",
  51304=>"111001101",
  51305=>"010111010",
  51306=>"111111101",
  51307=>"100010100",
  51308=>"001100100",
  51309=>"101111001",
  51310=>"011110010",
  51311=>"000111111",
  51312=>"101111001",
  51313=>"111001110",
  51314=>"100100001",
  51315=>"010000010",
  51316=>"011110000",
  51317=>"010110101",
  51318=>"000100000",
  51319=>"101100001",
  51320=>"000111000",
  51321=>"001010000",
  51322=>"011000000",
  51323=>"101100111",
  51324=>"110001100",
  51325=>"011101010",
  51326=>"010101001",
  51327=>"111000011",
  51328=>"100011100",
  51329=>"001001100",
  51330=>"110100101",
  51331=>"000100001",
  51332=>"110010101",
  51333=>"001101010",
  51334=>"100011111",
  51335=>"100100110",
  51336=>"011101101",
  51337=>"011001111",
  51338=>"100001001",
  51339=>"110001110",
  51340=>"000011100",
  51341=>"111001010",
  51342=>"100110000",
  51343=>"011000111",
  51344=>"101101010",
  51345=>"001001111",
  51346=>"100010000",
  51347=>"010011001",
  51348=>"111011001",
  51349=>"011011011",
  51350=>"011101100",
  51351=>"101000100",
  51352=>"110011010",
  51353=>"110100010",
  51354=>"000011101",
  51355=>"000011001",
  51356=>"000100010",
  51357=>"001000110",
  51358=>"011010100",
  51359=>"110011110",
  51360=>"111010101",
  51361=>"011101000",
  51362=>"101011111",
  51363=>"000100101",
  51364=>"100011001",
  51365=>"110000011",
  51366=>"111000101",
  51367=>"111110101",
  51368=>"100001000",
  51369=>"100011001",
  51370=>"100010010",
  51371=>"000101101",
  51372=>"100011011",
  51373=>"000110000",
  51374=>"001100100",
  51375=>"001000100",
  51376=>"001011000",
  51377=>"111111000",
  51378=>"110001001",
  51379=>"001010100",
  51380=>"111001100",
  51381=>"001100110",
  51382=>"111010000",
  51383=>"000110110",
  51384=>"111000110",
  51385=>"110001001",
  51386=>"111100001",
  51387=>"101010111",
  51388=>"100000010",
  51389=>"001110111",
  51390=>"101110111",
  51391=>"111100111",
  51392=>"101001101",
  51393=>"111011000",
  51394=>"010010001",
  51395=>"100111001",
  51396=>"101011110",
  51397=>"100000011",
  51398=>"110010100",
  51399=>"010000011",
  51400=>"111101000",
  51401=>"111011110",
  51402=>"100010111",
  51403=>"111100001",
  51404=>"111001110",
  51405=>"011100101",
  51406=>"011111101",
  51407=>"010111110",
  51408=>"111110001",
  51409=>"101101100",
  51410=>"011011001",
  51411=>"001111001",
  51412=>"011010011",
  51413=>"111010010",
  51414=>"001110101",
  51415=>"100111111",
  51416=>"100110100",
  51417=>"110010000",
  51418=>"000010011",
  51419=>"011101101",
  51420=>"011010011",
  51421=>"101101101",
  51422=>"110110010",
  51423=>"000110110",
  51424=>"011001001",
  51425=>"011111000",
  51426=>"011110000",
  51427=>"001101110",
  51428=>"000100101",
  51429=>"011110010",
  51430=>"100000000",
  51431=>"100011111",
  51432=>"111110000",
  51433=>"011011010",
  51434=>"110110101",
  51435=>"011010111",
  51436=>"101101100",
  51437=>"011001100",
  51438=>"010011110",
  51439=>"101000010",
  51440=>"001010011",
  51441=>"111010100",
  51442=>"010111100",
  51443=>"111010101",
  51444=>"101000000",
  51445=>"000100110",
  51446=>"100101100",
  51447=>"101111001",
  51448=>"100110011",
  51449=>"100100101",
  51450=>"111011101",
  51451=>"111000100",
  51452=>"011100011",
  51453=>"111010010",
  51454=>"011111110",
  51455=>"100001110",
  51456=>"001101100",
  51457=>"101000000",
  51458=>"010010111",
  51459=>"111100110",
  51460=>"000001000",
  51461=>"010001111",
  51462=>"001001001",
  51463=>"111101100",
  51464=>"111111101",
  51465=>"111000011",
  51466=>"111011001",
  51467=>"001110100",
  51468=>"000111000",
  51469=>"000101101",
  51470=>"011001010",
  51471=>"001010001",
  51472=>"010000100",
  51473=>"110000010",
  51474=>"010101000",
  51475=>"001110001",
  51476=>"010011100",
  51477=>"110111101",
  51478=>"100111000",
  51479=>"100100111",
  51480=>"100111011",
  51481=>"111100011",
  51482=>"101110100",
  51483=>"001111011",
  51484=>"110011001",
  51485=>"011001100",
  51486=>"000100001",
  51487=>"100110001",
  51488=>"110111110",
  51489=>"110011001",
  51490=>"001001111",
  51491=>"101000010",
  51492=>"011101101",
  51493=>"100010010",
  51494=>"101110100",
  51495=>"011001011",
  51496=>"101000001",
  51497=>"111001101",
  51498=>"010111100",
  51499=>"000100000",
  51500=>"111100011",
  51501=>"011011000",
  51502=>"001000100",
  51503=>"011001100",
  51504=>"111110000",
  51505=>"111000011",
  51506=>"111111011",
  51507=>"110011001",
  51508=>"111100101",
  51509=>"000100000",
  51510=>"010111011",
  51511=>"111001001",
  51512=>"100001000",
  51513=>"010010111",
  51514=>"110000110",
  51515=>"111111100",
  51516=>"110110001",
  51517=>"001100001",
  51518=>"000100010",
  51519=>"010101011",
  51520=>"000000101",
  51521=>"000101001",
  51522=>"101111101",
  51523=>"101000011",
  51524=>"101000011",
  51525=>"101110111",
  51526=>"001001110",
  51527=>"101110010",
  51528=>"010110010",
  51529=>"001100100",
  51530=>"100000111",
  51531=>"010000000",
  51532=>"101000101",
  51533=>"001110101",
  51534=>"110100100",
  51535=>"011011000",
  51536=>"001001011",
  51537=>"101001111",
  51538=>"000000011",
  51539=>"110110000",
  51540=>"000110100",
  51541=>"100001010",
  51542=>"101001111",
  51543=>"000000000",
  51544=>"100011010",
  51545=>"001011001",
  51546=>"000101000",
  51547=>"011000011",
  51548=>"101000001",
  51549=>"011011111",
  51550=>"011011000",
  51551=>"001001001",
  51552=>"010011001",
  51553=>"110001011",
  51554=>"110101111",
  51555=>"011000100",
  51556=>"110000110",
  51557=>"111011100",
  51558=>"011000010",
  51559=>"101110011",
  51560=>"010001011",
  51561=>"101101000",
  51562=>"101111111",
  51563=>"110000100",
  51564=>"111010100",
  51565=>"101100010",
  51566=>"001011100",
  51567=>"111010000",
  51568=>"001111001",
  51569=>"111101000",
  51570=>"011010110",
  51571=>"011000111",
  51572=>"101110011",
  51573=>"100000111",
  51574=>"010000100",
  51575=>"110101011",
  51576=>"100110111",
  51577=>"101000011",
  51578=>"010011000",
  51579=>"010110001",
  51580=>"101010101",
  51581=>"110011000",
  51582=>"001011000",
  51583=>"101001001",
  51584=>"000111111",
  51585=>"101000111",
  51586=>"100011101",
  51587=>"100100010",
  51588=>"110010111",
  51589=>"110101100",
  51590=>"000000011",
  51591=>"101111110",
  51592=>"111110001",
  51593=>"100011011",
  51594=>"111001000",
  51595=>"100110111",
  51596=>"010010010",
  51597=>"110111000",
  51598=>"001110001",
  51599=>"000000010",
  51600=>"010010110",
  51601=>"111111111",
  51602=>"110000100",
  51603=>"100101011",
  51604=>"010111010",
  51605=>"101111111",
  51606=>"100001000",
  51607=>"000111000",
  51608=>"100100101",
  51609=>"001010000",
  51610=>"111000001",
  51611=>"000000101",
  51612=>"110110000",
  51613=>"100000010",
  51614=>"010010000",
  51615=>"111101110",
  51616=>"000000101",
  51617=>"110110010",
  51618=>"111001011",
  51619=>"001001110",
  51620=>"001110011",
  51621=>"010010101",
  51622=>"000011100",
  51623=>"011110010",
  51624=>"011001100",
  51625=>"001101000",
  51626=>"000010000",
  51627=>"011011011",
  51628=>"110000101",
  51629=>"110110000",
  51630=>"000110001",
  51631=>"001100011",
  51632=>"010000011",
  51633=>"110100100",
  51634=>"010010111",
  51635=>"010001000",
  51636=>"001011000",
  51637=>"101110010",
  51638=>"100111110",
  51639=>"101110100",
  51640=>"100101000",
  51641=>"110001010",
  51642=>"010010111",
  51643=>"111100001",
  51644=>"111110101",
  51645=>"001111110",
  51646=>"010001001",
  51647=>"010011011",
  51648=>"110001010",
  51649=>"110011010",
  51650=>"111100000",
  51651=>"101111001",
  51652=>"111000101",
  51653=>"111101101",
  51654=>"100010010",
  51655=>"111011110",
  51656=>"100001001",
  51657=>"011010011",
  51658=>"111111110",
  51659=>"001010101",
  51660=>"000110110",
  51661=>"100100000",
  51662=>"101101111",
  51663=>"111110111",
  51664=>"101001110",
  51665=>"111011000",
  51666=>"000111110",
  51667=>"101110000",
  51668=>"011011000",
  51669=>"001000101",
  51670=>"010010000",
  51671=>"101000010",
  51672=>"110010100",
  51673=>"110110101",
  51674=>"111101011",
  51675=>"110110110",
  51676=>"010101111",
  51677=>"011001111",
  51678=>"010000011",
  51679=>"011110100",
  51680=>"100101111",
  51681=>"111010010",
  51682=>"100011101",
  51683=>"101010111",
  51684=>"000011010",
  51685=>"100010100",
  51686=>"110010001",
  51687=>"011111011",
  51688=>"101000011",
  51689=>"111111001",
  51690=>"100111001",
  51691=>"100101001",
  51692=>"010001001",
  51693=>"111110101",
  51694=>"001110000",
  51695=>"111010111",
  51696=>"110011010",
  51697=>"010010110",
  51698=>"011101010",
  51699=>"111001110",
  51700=>"111100000",
  51701=>"100001010",
  51702=>"010001111",
  51703=>"000000000",
  51704=>"100010010",
  51705=>"010010011",
  51706=>"001110000",
  51707=>"000100100",
  51708=>"110010001",
  51709=>"110011110",
  51710=>"101001000",
  51711=>"111011011",
  51712=>"011100000",
  51713=>"111011111",
  51714=>"111110010",
  51715=>"000101101",
  51716=>"000001001",
  51717=>"110110000",
  51718=>"111100100",
  51719=>"101101111",
  51720=>"110100101",
  51721=>"001011010",
  51722=>"011001001",
  51723=>"110110001",
  51724=>"011010001",
  51725=>"000000111",
  51726=>"111111000",
  51727=>"110100000",
  51728=>"010010100",
  51729=>"110011101",
  51730=>"110100011",
  51731=>"100111010",
  51732=>"110100000",
  51733=>"000111110",
  51734=>"110100101",
  51735=>"001110011",
  51736=>"000111000",
  51737=>"000001010",
  51738=>"000000001",
  51739=>"111000000",
  51740=>"101101011",
  51741=>"110111000",
  51742=>"011000101",
  51743=>"111111010",
  51744=>"111111010",
  51745=>"011000011",
  51746=>"001010100",
  51747=>"111101111",
  51748=>"010111000",
  51749=>"001111111",
  51750=>"110111101",
  51751=>"001001000",
  51752=>"001011100",
  51753=>"110110111",
  51754=>"100011010",
  51755=>"100000010",
  51756=>"110110100",
  51757=>"110101011",
  51758=>"101101010",
  51759=>"101100010",
  51760=>"110110001",
  51761=>"001101001",
  51762=>"000000001",
  51763=>"100100001",
  51764=>"010011111",
  51765=>"001000100",
  51766=>"101100001",
  51767=>"001010011",
  51768=>"011001111",
  51769=>"010111000",
  51770=>"000111011",
  51771=>"001010011",
  51772=>"111110110",
  51773=>"100111110",
  51774=>"000011100",
  51775=>"100111011",
  51776=>"111001100",
  51777=>"010101000",
  51778=>"110010000",
  51779=>"101110001",
  51780=>"101000100",
  51781=>"001000001",
  51782=>"100001011",
  51783=>"001101110",
  51784=>"000001101",
  51785=>"010010001",
  51786=>"101001101",
  51787=>"010110001",
  51788=>"100110110",
  51789=>"010110010",
  51790=>"011101010",
  51791=>"011110011",
  51792=>"101001000",
  51793=>"110011100",
  51794=>"011011010",
  51795=>"011001100",
  51796=>"010001100",
  51797=>"111110011",
  51798=>"011100001",
  51799=>"001001100",
  51800=>"101111001",
  51801=>"011000111",
  51802=>"000110100",
  51803=>"001000001",
  51804=>"100110010",
  51805=>"001010010",
  51806=>"000001001",
  51807=>"000010000",
  51808=>"011100000",
  51809=>"000101100",
  51810=>"000010000",
  51811=>"111001011",
  51812=>"011101000",
  51813=>"001001111",
  51814=>"000101101",
  51815=>"000110000",
  51816=>"010110001",
  51817=>"011011010",
  51818=>"101101111",
  51819=>"111101110",
  51820=>"010000100",
  51821=>"011100010",
  51822=>"001111101",
  51823=>"010101001",
  51824=>"101100111",
  51825=>"100110100",
  51826=>"100010000",
  51827=>"111001010",
  51828=>"101000000",
  51829=>"001111100",
  51830=>"001110110",
  51831=>"100111110",
  51832=>"110100010",
  51833=>"010110111",
  51834=>"111101111",
  51835=>"100001100",
  51836=>"001010010",
  51837=>"100100010",
  51838=>"100110000",
  51839=>"011000100",
  51840=>"010111110",
  51841=>"111100100",
  51842=>"000000010",
  51843=>"000001100",
  51844=>"011001000",
  51845=>"011010101",
  51846=>"100110001",
  51847=>"001101010",
  51848=>"110001111",
  51849=>"110000000",
  51850=>"010110101",
  51851=>"001001001",
  51852=>"011100101",
  51853=>"101101100",
  51854=>"111001100",
  51855=>"000010001",
  51856=>"111010010",
  51857=>"111011111",
  51858=>"111010011",
  51859=>"110101101",
  51860=>"000100001",
  51861=>"101000101",
  51862=>"001001011",
  51863=>"001001100",
  51864=>"111100010",
  51865=>"111110100",
  51866=>"010001101",
  51867=>"111100101",
  51868=>"101100000",
  51869=>"111111001",
  51870=>"010101110",
  51871=>"011001100",
  51872=>"010000101",
  51873=>"100101101",
  51874=>"101010111",
  51875=>"111111001",
  51876=>"011011001",
  51877=>"111110111",
  51878=>"110100001",
  51879=>"101110000",
  51880=>"000100011",
  51881=>"101000110",
  51882=>"101000011",
  51883=>"111100010",
  51884=>"000111011",
  51885=>"111001010",
  51886=>"011010010",
  51887=>"110000110",
  51888=>"000001111",
  51889=>"111101110",
  51890=>"000110110",
  51891=>"000111110",
  51892=>"011011010",
  51893=>"101011001",
  51894=>"000101100",
  51895=>"110101111",
  51896=>"010001000",
  51897=>"100000111",
  51898=>"011110101",
  51899=>"010001111",
  51900=>"010001011",
  51901=>"111110001",
  51902=>"010100100",
  51903=>"111111010",
  51904=>"000101010",
  51905=>"101100110",
  51906=>"111101001",
  51907=>"111011001",
  51908=>"000011111",
  51909=>"001100010",
  51910=>"011010110",
  51911=>"111101001",
  51912=>"000101011",
  51913=>"110101101",
  51914=>"100001010",
  51915=>"001101001",
  51916=>"001010010",
  51917=>"011100100",
  51918=>"010010111",
  51919=>"111000100",
  51920=>"011110010",
  51921=>"101111101",
  51922=>"100111110",
  51923=>"110010111",
  51924=>"011000001",
  51925=>"010110111",
  51926=>"111101000",
  51927=>"000000010",
  51928=>"100000010",
  51929=>"111110000",
  51930=>"101001000",
  51931=>"111110101",
  51932=>"100100111",
  51933=>"100010111",
  51934=>"000000011",
  51935=>"111000001",
  51936=>"011111010",
  51937=>"100110101",
  51938=>"100011000",
  51939=>"111001100",
  51940=>"001101110",
  51941=>"000101011",
  51942=>"000011001",
  51943=>"111101010",
  51944=>"100011111",
  51945=>"111101111",
  51946=>"011101001",
  51947=>"010100001",
  51948=>"001000111",
  51949=>"111101110",
  51950=>"001010101",
  51951=>"010100000",
  51952=>"000100111",
  51953=>"111111001",
  51954=>"101000100",
  51955=>"001011110",
  51956=>"011110000",
  51957=>"000100001",
  51958=>"001111110",
  51959=>"110111110",
  51960=>"110010111",
  51961=>"000101110",
  51962=>"110001111",
  51963=>"101000101",
  51964=>"010010111",
  51965=>"101101000",
  51966=>"111101011",
  51967=>"000010111",
  51968=>"000111010",
  51969=>"011011001",
  51970=>"111101011",
  51971=>"000011111",
  51972=>"101110000",
  51973=>"000011111",
  51974=>"111010110",
  51975=>"110000111",
  51976=>"011001001",
  51977=>"000101011",
  51978=>"001110100",
  51979=>"111100001",
  51980=>"000001011",
  51981=>"010000110",
  51982=>"100110110",
  51983=>"000010011",
  51984=>"101111111",
  51985=>"000001001",
  51986=>"110010001",
  51987=>"101000101",
  51988=>"001000110",
  51989=>"010101011",
  51990=>"011110010",
  51991=>"111001100",
  51992=>"101000001",
  51993=>"001011001",
  51994=>"000000100",
  51995=>"100000000",
  51996=>"110101001",
  51997=>"110100000",
  51998=>"111000100",
  51999=>"011111011",
  52000=>"011101001",
  52001=>"011110000",
  52002=>"000101011",
  52003=>"010001000",
  52004=>"100011110",
  52005=>"000100100",
  52006=>"110010110",
  52007=>"010100101",
  52008=>"101111110",
  52009=>"111101011",
  52010=>"010101110",
  52011=>"000001010",
  52012=>"101110110",
  52013=>"011101010",
  52014=>"011000100",
  52015=>"001000000",
  52016=>"011100111",
  52017=>"101110111",
  52018=>"001100001",
  52019=>"100111011",
  52020=>"001100001",
  52021=>"100100110",
  52022=>"100110110",
  52023=>"101110110",
  52024=>"001101011",
  52025=>"101101000",
  52026=>"111111101",
  52027=>"100010100",
  52028=>"010100010",
  52029=>"000110010",
  52030=>"001100001",
  52031=>"111111101",
  52032=>"011111011",
  52033=>"100000111",
  52034=>"111100111",
  52035=>"010000110",
  52036=>"101000101",
  52037=>"000110000",
  52038=>"101001101",
  52039=>"101100110",
  52040=>"001101001",
  52041=>"000011011",
  52042=>"000101100",
  52043=>"011110011",
  52044=>"011000001",
  52045=>"111110010",
  52046=>"111010100",
  52047=>"010111110",
  52048=>"000100111",
  52049=>"101010101",
  52050=>"010101101",
  52051=>"101100001",
  52052=>"011010101",
  52053=>"111101101",
  52054=>"011111001",
  52055=>"011001110",
  52056=>"000100011",
  52057=>"110000010",
  52058=>"111111110",
  52059=>"001000100",
  52060=>"000111001",
  52061=>"101101110",
  52062=>"001010101",
  52063=>"111010000",
  52064=>"000101111",
  52065=>"111100001",
  52066=>"101001111",
  52067=>"111010110",
  52068=>"011000010",
  52069=>"000001011",
  52070=>"110110010",
  52071=>"000111111",
  52072=>"101001001",
  52073=>"110110111",
  52074=>"010101111",
  52075=>"000010011",
  52076=>"100111000",
  52077=>"101001001",
  52078=>"110001111",
  52079=>"011011010",
  52080=>"011101110",
  52081=>"010011110",
  52082=>"000011111",
  52083=>"100011010",
  52084=>"010010001",
  52085=>"111100100",
  52086=>"101110010",
  52087=>"001101110",
  52088=>"010100110",
  52089=>"110110011",
  52090=>"101011110",
  52091=>"010111001",
  52092=>"011000010",
  52093=>"100101000",
  52094=>"001110101",
  52095=>"110110011",
  52096=>"000001010",
  52097=>"111011000",
  52098=>"001000101",
  52099=>"100001111",
  52100=>"101110001",
  52101=>"001110000",
  52102=>"111110010",
  52103=>"000000010",
  52104=>"000101110",
  52105=>"111100101",
  52106=>"111000000",
  52107=>"000000100",
  52108=>"010011100",
  52109=>"110011111",
  52110=>"000011101",
  52111=>"110000100",
  52112=>"011111110",
  52113=>"110111110",
  52114=>"100000000",
  52115=>"001111000",
  52116=>"011011101",
  52117=>"010110010",
  52118=>"101000001",
  52119=>"110110001",
  52120=>"001111110",
  52121=>"110010011",
  52122=>"111110100",
  52123=>"110010010",
  52124=>"000000011",
  52125=>"101110001",
  52126=>"100111001",
  52127=>"110111000",
  52128=>"001000101",
  52129=>"010010110",
  52130=>"000000110",
  52131=>"101100111",
  52132=>"111110110",
  52133=>"100001110",
  52134=>"010110001",
  52135=>"000111111",
  52136=>"101001100",
  52137=>"101000011",
  52138=>"010100100",
  52139=>"111001010",
  52140=>"011011010",
  52141=>"110110110",
  52142=>"000010110",
  52143=>"100000011",
  52144=>"000001111",
  52145=>"110101100",
  52146=>"101001100",
  52147=>"110111101",
  52148=>"111100110",
  52149=>"011110010",
  52150=>"001000111",
  52151=>"011100011",
  52152=>"111100111",
  52153=>"101100110",
  52154=>"100111110",
  52155=>"010111001",
  52156=>"101011111",
  52157=>"101111101",
  52158=>"110000000",
  52159=>"111101100",
  52160=>"000001000",
  52161=>"110010110",
  52162=>"000010110",
  52163=>"001100001",
  52164=>"110110011",
  52165=>"001101011",
  52166=>"000110001",
  52167=>"110011000",
  52168=>"000000001",
  52169=>"000110000",
  52170=>"010000001",
  52171=>"010101111",
  52172=>"111110010",
  52173=>"111100001",
  52174=>"010011001",
  52175=>"111110111",
  52176=>"011000100",
  52177=>"011110110",
  52178=>"100110011",
  52179=>"000011100",
  52180=>"100001110",
  52181=>"010000010",
  52182=>"110001001",
  52183=>"011001011",
  52184=>"111011111",
  52185=>"001000100",
  52186=>"010010111",
  52187=>"100101010",
  52188=>"000101011",
  52189=>"111001100",
  52190=>"100011101",
  52191=>"010110111",
  52192=>"001010010",
  52193=>"101001010",
  52194=>"101111001",
  52195=>"110000000",
  52196=>"101010100",
  52197=>"110111000",
  52198=>"000110000",
  52199=>"001110100",
  52200=>"110000111",
  52201=>"011010111",
  52202=>"011010010",
  52203=>"000110100",
  52204=>"000011000",
  52205=>"011011101",
  52206=>"110000010",
  52207=>"001010001",
  52208=>"101001000",
  52209=>"001001101",
  52210=>"000101101",
  52211=>"001101100",
  52212=>"011101010",
  52213=>"111011100",
  52214=>"010101000",
  52215=>"011011000",
  52216=>"110001010",
  52217=>"001010101",
  52218=>"111001101",
  52219=>"100111011",
  52220=>"100101110",
  52221=>"010100110",
  52222=>"001000001",
  52223=>"100010111",
  52224=>"110010111",
  52225=>"110001100",
  52226=>"000101111",
  52227=>"011100011",
  52228=>"000100000",
  52229=>"001000110",
  52230=>"110111010",
  52231=>"111000100",
  52232=>"110010100",
  52233=>"100010001",
  52234=>"111011111",
  52235=>"110001010",
  52236=>"100101111",
  52237=>"111101010",
  52238=>"000001000",
  52239=>"111110000",
  52240=>"101100111",
  52241=>"000111110",
  52242=>"110000000",
  52243=>"001101100",
  52244=>"011100010",
  52245=>"110011110",
  52246=>"000011011",
  52247=>"000001001",
  52248=>"101000000",
  52249=>"001101110",
  52250=>"101100101",
  52251=>"111000010",
  52252=>"111110100",
  52253=>"100000000",
  52254=>"000111100",
  52255=>"111000011",
  52256=>"011100101",
  52257=>"011101110",
  52258=>"111100010",
  52259=>"110001110",
  52260=>"111000010",
  52261=>"110000110",
  52262=>"101011011",
  52263=>"011011001",
  52264=>"101011011",
  52265=>"001101100",
  52266=>"111100111",
  52267=>"001011011",
  52268=>"101010011",
  52269=>"010100010",
  52270=>"000010110",
  52271=>"100010000",
  52272=>"010101001",
  52273=>"001010100",
  52274=>"010010011",
  52275=>"000000101",
  52276=>"000001101",
  52277=>"011000100",
  52278=>"000100000",
  52279=>"111100101",
  52280=>"101001101",
  52281=>"110111111",
  52282=>"000110010",
  52283=>"000101000",
  52284=>"000110110",
  52285=>"011010001",
  52286=>"110011011",
  52287=>"100010000",
  52288=>"000011001",
  52289=>"000000100",
  52290=>"010010010",
  52291=>"001111000",
  52292=>"010110100",
  52293=>"001101110",
  52294=>"000101000",
  52295=>"100000110",
  52296=>"111011010",
  52297=>"101010010",
  52298=>"111111001",
  52299=>"011111001",
  52300=>"000010000",
  52301=>"011111011",
  52302=>"111101111",
  52303=>"001101011",
  52304=>"100011001",
  52305=>"000101100",
  52306=>"110010101",
  52307=>"111110101",
  52308=>"100001001",
  52309=>"010101001",
  52310=>"001101000",
  52311=>"111101111",
  52312=>"100001111",
  52313=>"111011110",
  52314=>"100010111",
  52315=>"000010001",
  52316=>"001100001",
  52317=>"001011010",
  52318=>"101010101",
  52319=>"110111011",
  52320=>"100100000",
  52321=>"100001101",
  52322=>"011111010",
  52323=>"000110110",
  52324=>"011000000",
  52325=>"101001000",
  52326=>"000000000",
  52327=>"111111111",
  52328=>"000011100",
  52329=>"010100110",
  52330=>"000110010",
  52331=>"110110000",
  52332=>"110100001",
  52333=>"000101000",
  52334=>"010001001",
  52335=>"001101010",
  52336=>"110010001",
  52337=>"011100101",
  52338=>"110100110",
  52339=>"111101111",
  52340=>"000001110",
  52341=>"000011000",
  52342=>"011110001",
  52343=>"000101101",
  52344=>"110111010",
  52345=>"001110000",
  52346=>"110011110",
  52347=>"011000001",
  52348=>"110001110",
  52349=>"101100010",
  52350=>"011010110",
  52351=>"100001011",
  52352=>"100011111",
  52353=>"010101001",
  52354=>"010010000",
  52355=>"101001100",
  52356=>"000000100",
  52357=>"100010110",
  52358=>"110011110",
  52359=>"000000011",
  52360=>"001010100",
  52361=>"011011011",
  52362=>"010000001",
  52363=>"011111001",
  52364=>"101101111",
  52365=>"100001011",
  52366=>"100000010",
  52367=>"011011101",
  52368=>"010111110",
  52369=>"100010000",
  52370=>"110001000",
  52371=>"000110011",
  52372=>"001010000",
  52373=>"000100100",
  52374=>"010011111",
  52375=>"100101000",
  52376=>"110101111",
  52377=>"100111101",
  52378=>"010000100",
  52379=>"001010100",
  52380=>"000001010",
  52381=>"100001001",
  52382=>"101000001",
  52383=>"000010010",
  52384=>"111011001",
  52385=>"011111101",
  52386=>"000011001",
  52387=>"100000000",
  52388=>"111100000",
  52389=>"100111101",
  52390=>"011110011",
  52391=>"110110010",
  52392=>"110111000",
  52393=>"101000001",
  52394=>"011001001",
  52395=>"011101111",
  52396=>"001100000",
  52397=>"111000001",
  52398=>"101000011",
  52399=>"110111101",
  52400=>"101001101",
  52401=>"011110100",
  52402=>"010111001",
  52403=>"011010010",
  52404=>"101011010",
  52405=>"001011101",
  52406=>"110001101",
  52407=>"010101010",
  52408=>"010001011",
  52409=>"000101100",
  52410=>"000000110",
  52411=>"000100010",
  52412=>"111101111",
  52413=>"110010110",
  52414=>"100010011",
  52415=>"110110100",
  52416=>"100001101",
  52417=>"111110101",
  52418=>"111100101",
  52419=>"100010110",
  52420=>"111100110",
  52421=>"100001100",
  52422=>"000010001",
  52423=>"111110011",
  52424=>"100111001",
  52425=>"010000101",
  52426=>"010000000",
  52427=>"010111010",
  52428=>"111001001",
  52429=>"000001000",
  52430=>"111011110",
  52431=>"110110000",
  52432=>"100010001",
  52433=>"000100010",
  52434=>"001111110",
  52435=>"101100011",
  52436=>"101000101",
  52437=>"010011001",
  52438=>"001110000",
  52439=>"111011000",
  52440=>"111101101",
  52441=>"110100111",
  52442=>"100000110",
  52443=>"010010000",
  52444=>"101011011",
  52445=>"001000100",
  52446=>"001111010",
  52447=>"000110100",
  52448=>"010101110",
  52449=>"000111000",
  52450=>"010100100",
  52451=>"110111111",
  52452=>"110001101",
  52453=>"110101011",
  52454=>"011001111",
  52455=>"111000110",
  52456=>"011101111",
  52457=>"111101111",
  52458=>"001111001",
  52459=>"101110000",
  52460=>"101111010",
  52461=>"100111010",
  52462=>"000111000",
  52463=>"011010000",
  52464=>"011010111",
  52465=>"000111010",
  52466=>"011101010",
  52467=>"100111001",
  52468=>"111001110",
  52469=>"001011001",
  52470=>"101000011",
  52471=>"000011001",
  52472=>"011111100",
  52473=>"001010000",
  52474=>"011000000",
  52475=>"000111111",
  52476=>"011001101",
  52477=>"101011110",
  52478=>"001001000",
  52479=>"011101100",
  52480=>"101001001",
  52481=>"100101111",
  52482=>"001011110",
  52483=>"101011111",
  52484=>"100001110",
  52485=>"001100111",
  52486=>"010000110",
  52487=>"100110100",
  52488=>"011010011",
  52489=>"000111001",
  52490=>"100101110",
  52491=>"110000011",
  52492=>"011100000",
  52493=>"001010100",
  52494=>"000101001",
  52495=>"000010100",
  52496=>"000000000",
  52497=>"011100100",
  52498=>"101000111",
  52499=>"111011000",
  52500=>"101010111",
  52501=>"010000111",
  52502=>"010010011",
  52503=>"000011111",
  52504=>"010010000",
  52505=>"000000000",
  52506=>"100100000",
  52507=>"100010101",
  52508=>"000100001",
  52509=>"100100111",
  52510=>"001010000",
  52511=>"000001010",
  52512=>"100101100",
  52513=>"000000101",
  52514=>"010000111",
  52515=>"000001010",
  52516=>"010000000",
  52517=>"001000100",
  52518=>"111101110",
  52519=>"111111111",
  52520=>"001110011",
  52521=>"101001111",
  52522=>"111000111",
  52523=>"111011000",
  52524=>"101011110",
  52525=>"111111011",
  52526=>"111000010",
  52527=>"010100001",
  52528=>"101101111",
  52529=>"001011100",
  52530=>"111101100",
  52531=>"001000001",
  52532=>"101101111",
  52533=>"010000000",
  52534=>"111110100",
  52535=>"001111111",
  52536=>"000010000",
  52537=>"110000100",
  52538=>"000010000",
  52539=>"011100100",
  52540=>"100010001",
  52541=>"000100111",
  52542=>"010000011",
  52543=>"101101001",
  52544=>"010000010",
  52545=>"100100010",
  52546=>"011110111",
  52547=>"100111101",
  52548=>"111010011",
  52549=>"010110011",
  52550=>"100010001",
  52551=>"011011110",
  52552=>"011101011",
  52553=>"110101110",
  52554=>"011100110",
  52555=>"000100101",
  52556=>"001110011",
  52557=>"100000100",
  52558=>"001011111",
  52559=>"111011111",
  52560=>"000110110",
  52561=>"011111010",
  52562=>"010101111",
  52563=>"100001001",
  52564=>"010101000",
  52565=>"010110000",
  52566=>"100100011",
  52567=>"001111011",
  52568=>"011101010",
  52569=>"011110101",
  52570=>"111101000",
  52571=>"001001101",
  52572=>"011110111",
  52573=>"110001100",
  52574=>"010101100",
  52575=>"001000100",
  52576=>"011101011",
  52577=>"000010001",
  52578=>"100000111",
  52579=>"101101101",
  52580=>"001010011",
  52581=>"000110101",
  52582=>"010101100",
  52583=>"000011011",
  52584=>"110101111",
  52585=>"010100001",
  52586=>"010010100",
  52587=>"000101011",
  52588=>"111011011",
  52589=>"001011011",
  52590=>"111100101",
  52591=>"111010000",
  52592=>"000011010",
  52593=>"111010001",
  52594=>"000011101",
  52595=>"111000101",
  52596=>"000000101",
  52597=>"000010000",
  52598=>"011110111",
  52599=>"011000110",
  52600=>"101110010",
  52601=>"110011100",
  52602=>"011101111",
  52603=>"110011111",
  52604=>"000010010",
  52605=>"011111011",
  52606=>"000000110",
  52607=>"100000101",
  52608=>"111010100",
  52609=>"010010111",
  52610=>"011101110",
  52611=>"100111100",
  52612=>"011001111",
  52613=>"110100010",
  52614=>"011111111",
  52615=>"101001011",
  52616=>"111110100",
  52617=>"010011010",
  52618=>"011001110",
  52619=>"011010000",
  52620=>"100001011",
  52621=>"000001011",
  52622=>"000011100",
  52623=>"001011110",
  52624=>"100000110",
  52625=>"000011001",
  52626=>"111101010",
  52627=>"000101011",
  52628=>"110010101",
  52629=>"001001111",
  52630=>"011100111",
  52631=>"001100000",
  52632=>"010000110",
  52633=>"000110011",
  52634=>"000001101",
  52635=>"100111010",
  52636=>"111110010",
  52637=>"010110011",
  52638=>"101011010",
  52639=>"001100000",
  52640=>"111100011",
  52641=>"010000100",
  52642=>"010100111",
  52643=>"100010100",
  52644=>"110000001",
  52645=>"111101011",
  52646=>"000000110",
  52647=>"001000010",
  52648=>"101010010",
  52649=>"110001110",
  52650=>"111111000",
  52651=>"010010010",
  52652=>"000110100",
  52653=>"111110100",
  52654=>"010010101",
  52655=>"101111000",
  52656=>"100000111",
  52657=>"010010000",
  52658=>"111010111",
  52659=>"101111111",
  52660=>"111110000",
  52661=>"010001100",
  52662=>"111111010",
  52663=>"100101001",
  52664=>"101100111",
  52665=>"001010100",
  52666=>"110011001",
  52667=>"000110101",
  52668=>"001100101",
  52669=>"000011101",
  52670=>"011011011",
  52671=>"110111111",
  52672=>"001000101",
  52673=>"001100110",
  52674=>"100001111",
  52675=>"011111110",
  52676=>"100010010",
  52677=>"110000001",
  52678=>"001001001",
  52679=>"001011000",
  52680=>"010011001",
  52681=>"110100101",
  52682=>"000011010",
  52683=>"101001110",
  52684=>"010100000",
  52685=>"111100001",
  52686=>"010110111",
  52687=>"000011110",
  52688=>"001011011",
  52689=>"011100001",
  52690=>"101100110",
  52691=>"011010000",
  52692=>"101100101",
  52693=>"010000100",
  52694=>"000000011",
  52695=>"010010101",
  52696=>"000001010",
  52697=>"011110001",
  52698=>"001001010",
  52699=>"011011110",
  52700=>"111100000",
  52701=>"100000001",
  52702=>"111000111",
  52703=>"000100110",
  52704=>"111111100",
  52705=>"001000101",
  52706=>"100111011",
  52707=>"100010101",
  52708=>"110100000",
  52709=>"101000010",
  52710=>"011011111",
  52711=>"100111001",
  52712=>"010111111",
  52713=>"000010111",
  52714=>"001001001",
  52715=>"101110111",
  52716=>"001010011",
  52717=>"101111000",
  52718=>"000011100",
  52719=>"101000000",
  52720=>"011010111",
  52721=>"101010110",
  52722=>"001111101",
  52723=>"000010110",
  52724=>"101100101",
  52725=>"001101111",
  52726=>"111011110",
  52727=>"111010110",
  52728=>"001110000",
  52729=>"000111000",
  52730=>"010010010",
  52731=>"111010111",
  52732=>"001001001",
  52733=>"001000110",
  52734=>"000010101",
  52735=>"011010101",
  52736=>"101010100",
  52737=>"000101111",
  52738=>"111111110",
  52739=>"010010111",
  52740=>"110000111",
  52741=>"000001010",
  52742=>"000011110",
  52743=>"010001010",
  52744=>"111000010",
  52745=>"010110100",
  52746=>"111001010",
  52747=>"001001000",
  52748=>"010101010",
  52749=>"110110110",
  52750=>"000101000",
  52751=>"010110100",
  52752=>"010111111",
  52753=>"110000111",
  52754=>"000111101",
  52755=>"011011101",
  52756=>"000000011",
  52757=>"010111110",
  52758=>"110010000",
  52759=>"011110010",
  52760=>"111101100",
  52761=>"100111001",
  52762=>"110110111",
  52763=>"110010101",
  52764=>"001100001",
  52765=>"110101101",
  52766=>"110110100",
  52767=>"010101000",
  52768=>"001010111",
  52769=>"001001011",
  52770=>"111110001",
  52771=>"011101011",
  52772=>"101010100",
  52773=>"110000101",
  52774=>"010010000",
  52775=>"111101111",
  52776=>"000100001",
  52777=>"000011111",
  52778=>"110011101",
  52779=>"101011100",
  52780=>"010101000",
  52781=>"000110111",
  52782=>"111101000",
  52783=>"001000000",
  52784=>"101001001",
  52785=>"001010111",
  52786=>"110011111",
  52787=>"001000010",
  52788=>"010001000",
  52789=>"001001000",
  52790=>"100000010",
  52791=>"010110000",
  52792=>"110101101",
  52793=>"010100110",
  52794=>"111001011",
  52795=>"110001000",
  52796=>"100100100",
  52797=>"110010100",
  52798=>"100010101",
  52799=>"111100001",
  52800=>"011111110",
  52801=>"011101111",
  52802=>"110101100",
  52803=>"111010011",
  52804=>"011110101",
  52805=>"101000010",
  52806=>"000001011",
  52807=>"111000010",
  52808=>"100010100",
  52809=>"010000111",
  52810=>"100110000",
  52811=>"110101111",
  52812=>"000000111",
  52813=>"011111011",
  52814=>"011000001",
  52815=>"110001010",
  52816=>"101001101",
  52817=>"000100001",
  52818=>"011101100",
  52819=>"001011010",
  52820=>"000110000",
  52821=>"100001010",
  52822=>"111101011",
  52823=>"000111111",
  52824=>"110101011",
  52825=>"111101101",
  52826=>"011101010",
  52827=>"001001110",
  52828=>"001010111",
  52829=>"111101001",
  52830=>"010011010",
  52831=>"000010010",
  52832=>"010001011",
  52833=>"100101000",
  52834=>"010101010",
  52835=>"000101000",
  52836=>"100110100",
  52837=>"101011110",
  52838=>"011100110",
  52839=>"100010011",
  52840=>"100001101",
  52841=>"110100010",
  52842=>"110111000",
  52843=>"011000010",
  52844=>"000100110",
  52845=>"000110100",
  52846=>"000010001",
  52847=>"010011101",
  52848=>"101000111",
  52849=>"100100010",
  52850=>"011010001",
  52851=>"110011010",
  52852=>"011000001",
  52853=>"100010100",
  52854=>"011011110",
  52855=>"010011111",
  52856=>"001111001",
  52857=>"000000000",
  52858=>"110011011",
  52859=>"011101011",
  52860=>"010010101",
  52861=>"101111010",
  52862=>"000000000",
  52863=>"011111010",
  52864=>"000100000",
  52865=>"111011010",
  52866=>"010011011",
  52867=>"011000110",
  52868=>"100001100",
  52869=>"101111100",
  52870=>"110110001",
  52871=>"111101001",
  52872=>"000110000",
  52873=>"101000000",
  52874=>"110000011",
  52875=>"100101111",
  52876=>"100110001",
  52877=>"010011000",
  52878=>"100100000",
  52879=>"011111100",
  52880=>"001100110",
  52881=>"111110000",
  52882=>"110010001",
  52883=>"101001110",
  52884=>"010001100",
  52885=>"101011110",
  52886=>"101101000",
  52887=>"010111100",
  52888=>"100001000",
  52889=>"000111011",
  52890=>"101101101",
  52891=>"011110100",
  52892=>"000011001",
  52893=>"100100011",
  52894=>"011101010",
  52895=>"111001100",
  52896=>"111010100",
  52897=>"010111001",
  52898=>"001110001",
  52899=>"111011110",
  52900=>"111010001",
  52901=>"110111011",
  52902=>"111000000",
  52903=>"001000001",
  52904=>"000001111",
  52905=>"000100010",
  52906=>"111000101",
  52907=>"001010000",
  52908=>"010000000",
  52909=>"000100100",
  52910=>"001110110",
  52911=>"100000111",
  52912=>"010100100",
  52913=>"000010000",
  52914=>"001000100",
  52915=>"111011110",
  52916=>"110011100",
  52917=>"101111101",
  52918=>"110010101",
  52919=>"011110001",
  52920=>"000100001",
  52921=>"001001000",
  52922=>"011000101",
  52923=>"011010010",
  52924=>"001001000",
  52925=>"111011001",
  52926=>"100111111",
  52927=>"000110100",
  52928=>"101111000",
  52929=>"111101001",
  52930=>"110001011",
  52931=>"110000000",
  52932=>"100000111",
  52933=>"111011001",
  52934=>"111100011",
  52935=>"001110000",
  52936=>"000110001",
  52937=>"001000101",
  52938=>"001110110",
  52939=>"111011001",
  52940=>"000101010",
  52941=>"101110011",
  52942=>"100000100",
  52943=>"011001010",
  52944=>"001010101",
  52945=>"100100000",
  52946=>"011000010",
  52947=>"111011101",
  52948=>"000101010",
  52949=>"000111111",
  52950=>"111010010",
  52951=>"110110010",
  52952=>"010001111",
  52953=>"011010110",
  52954=>"010011110",
  52955=>"010010110",
  52956=>"111111100",
  52957=>"010011011",
  52958=>"010111111",
  52959=>"100001001",
  52960=>"101101101",
  52961=>"111011001",
  52962=>"000101110",
  52963=>"101101101",
  52964=>"000001101",
  52965=>"010010011",
  52966=>"100101000",
  52967=>"110100100",
  52968=>"101010110",
  52969=>"001110101",
  52970=>"111110001",
  52971=>"100000001",
  52972=>"011011010",
  52973=>"010110111",
  52974=>"010101110",
  52975=>"010011111",
  52976=>"111100101",
  52977=>"110111110",
  52978=>"010110111",
  52979=>"011011101",
  52980=>"010111001",
  52981=>"000000100",
  52982=>"100001001",
  52983=>"100100001",
  52984=>"100100011",
  52985=>"101100110",
  52986=>"111011011",
  52987=>"011010010",
  52988=>"110011101",
  52989=>"010110011",
  52990=>"101110100",
  52991=>"110110001",
  52992=>"111010001",
  52993=>"111110100",
  52994=>"110101011",
  52995=>"011001010",
  52996=>"101100001",
  52997=>"101100100",
  52998=>"110100011",
  52999=>"010101100",
  53000=>"010101100",
  53001=>"011110101",
  53002=>"111110001",
  53003=>"110011010",
  53004=>"000000111",
  53005=>"100001110",
  53006=>"011010010",
  53007=>"100000001",
  53008=>"001110010",
  53009=>"010011101",
  53010=>"001000000",
  53011=>"011111111",
  53012=>"011100100",
  53013=>"010001100",
  53014=>"111010111",
  53015=>"000011101",
  53016=>"110000000",
  53017=>"010100010",
  53018=>"001100001",
  53019=>"110111100",
  53020=>"011000100",
  53021=>"011110010",
  53022=>"010010000",
  53023=>"000101001",
  53024=>"101100001",
  53025=>"001011110",
  53026=>"100001001",
  53027=>"000110001",
  53028=>"011001111",
  53029=>"000001000",
  53030=>"010010011",
  53031=>"010110100",
  53032=>"101010100",
  53033=>"001011010",
  53034=>"000010110",
  53035=>"100010111",
  53036=>"010010010",
  53037=>"100110101",
  53038=>"000101100",
  53039=>"000101100",
  53040=>"011001000",
  53041=>"100000110",
  53042=>"001011111",
  53043=>"000010110",
  53044=>"001110000",
  53045=>"101010110",
  53046=>"101110011",
  53047=>"001000011",
  53048=>"011000011",
  53049=>"000101001",
  53050=>"101000010",
  53051=>"110001000",
  53052=>"010000000",
  53053=>"010010101",
  53054=>"000001001",
  53055=>"000111010",
  53056=>"100001000",
  53057=>"100011001",
  53058=>"110111011",
  53059=>"000001101",
  53060=>"100010011",
  53061=>"010010111",
  53062=>"000001110",
  53063=>"111010011",
  53064=>"100100011",
  53065=>"001101010",
  53066=>"111001010",
  53067=>"001110010",
  53068=>"010010011",
  53069=>"111111111",
  53070=>"010111001",
  53071=>"110000000",
  53072=>"101101100",
  53073=>"000111001",
  53074=>"000010110",
  53075=>"001000001",
  53076=>"110010010",
  53077=>"001001111",
  53078=>"001111000",
  53079=>"100101010",
  53080=>"100010111",
  53081=>"100111000",
  53082=>"011111100",
  53083=>"111111010",
  53084=>"110010101",
  53085=>"000110010",
  53086=>"101101000",
  53087=>"001001110",
  53088=>"110110000",
  53089=>"111110001",
  53090=>"110100110",
  53091=>"001001101",
  53092=>"001010111",
  53093=>"100001001",
  53094=>"011000010",
  53095=>"100011111",
  53096=>"000101100",
  53097=>"110100100",
  53098=>"100101000",
  53099=>"110001101",
  53100=>"001001111",
  53101=>"100010000",
  53102=>"011001001",
  53103=>"101000010",
  53104=>"101000110",
  53105=>"001000010",
  53106=>"000100111",
  53107=>"011011010",
  53108=>"011100010",
  53109=>"000100101",
  53110=>"101001100",
  53111=>"100100100",
  53112=>"110000011",
  53113=>"101000111",
  53114=>"011101001",
  53115=>"100011000",
  53116=>"101011000",
  53117=>"001101000",
  53118=>"111100100",
  53119=>"011101011",
  53120=>"010000011",
  53121=>"100101011",
  53122=>"110101110",
  53123=>"011111110",
  53124=>"000110011",
  53125=>"111010100",
  53126=>"001111100",
  53127=>"000010110",
  53128=>"010001111",
  53129=>"000001010",
  53130=>"001010101",
  53131=>"010100000",
  53132=>"100001001",
  53133=>"011011001",
  53134=>"011101011",
  53135=>"000111000",
  53136=>"000001100",
  53137=>"101000000",
  53138=>"000000000",
  53139=>"001011100",
  53140=>"110010110",
  53141=>"001110101",
  53142=>"110110101",
  53143=>"001101100",
  53144=>"101101110",
  53145=>"110011101",
  53146=>"100101111",
  53147=>"001011000",
  53148=>"000111111",
  53149=>"101100010",
  53150=>"100100010",
  53151=>"111100100",
  53152=>"101010010",
  53153=>"010010111",
  53154=>"111101010",
  53155=>"110000010",
  53156=>"011001001",
  53157=>"110101000",
  53158=>"110111100",
  53159=>"001011011",
  53160=>"100000010",
  53161=>"101111110",
  53162=>"111111110",
  53163=>"001110010",
  53164=>"000110101",
  53165=>"001110111",
  53166=>"011011011",
  53167=>"111001011",
  53168=>"111011100",
  53169=>"001011100",
  53170=>"100111111",
  53171=>"001100010",
  53172=>"011110011",
  53173=>"110010000",
  53174=>"000110101",
  53175=>"011101011",
  53176=>"001000100",
  53177=>"000000110",
  53178=>"101100111",
  53179=>"000110000",
  53180=>"011000001",
  53181=>"111010000",
  53182=>"000111010",
  53183=>"000000100",
  53184=>"111001010",
  53185=>"001110001",
  53186=>"100000100",
  53187=>"111110001",
  53188=>"010001010",
  53189=>"101000110",
  53190=>"111010010",
  53191=>"001000110",
  53192=>"000110111",
  53193=>"111011101",
  53194=>"100000111",
  53195=>"101011010",
  53196=>"100101101",
  53197=>"100000010",
  53198=>"111110011",
  53199=>"010001001",
  53200=>"001011110",
  53201=>"000010111",
  53202=>"101100011",
  53203=>"100000001",
  53204=>"000000010",
  53205=>"100000110",
  53206=>"001011000",
  53207=>"100000101",
  53208=>"010001110",
  53209=>"100010011",
  53210=>"100000011",
  53211=>"000001110",
  53212=>"011010010",
  53213=>"011011010",
  53214=>"100110101",
  53215=>"111000011",
  53216=>"101100110",
  53217=>"000000000",
  53218=>"110110010",
  53219=>"101111100",
  53220=>"100011000",
  53221=>"010110101",
  53222=>"111011001",
  53223=>"000001100",
  53224=>"111110101",
  53225=>"100101100",
  53226=>"110011100",
  53227=>"000010001",
  53228=>"100010010",
  53229=>"010001000",
  53230=>"101011101",
  53231=>"101111001",
  53232=>"011010000",
  53233=>"110010010",
  53234=>"001100001",
  53235=>"001010111",
  53236=>"010110001",
  53237=>"000101100",
  53238=>"100010000",
  53239=>"011000100",
  53240=>"100010110",
  53241=>"110000111",
  53242=>"101101100",
  53243=>"111111001",
  53244=>"110011100",
  53245=>"001001100",
  53246=>"000100001",
  53247=>"111001101",
  53248=>"101110001",
  53249=>"011000111",
  53250=>"010111101",
  53251=>"011101011",
  53252=>"001000011",
  53253=>"000100101",
  53254=>"110011010",
  53255=>"100110011",
  53256=>"110001111",
  53257=>"111111110",
  53258=>"100100101",
  53259=>"000100010",
  53260=>"100100111",
  53261=>"110101100",
  53262=>"110101010",
  53263=>"011110100",
  53264=>"111111001",
  53265=>"001001101",
  53266=>"001100100",
  53267=>"101000011",
  53268=>"101101010",
  53269=>"000010010",
  53270=>"110111111",
  53271=>"010000111",
  53272=>"101111111",
  53273=>"010000101",
  53274=>"101000100",
  53275=>"100110011",
  53276=>"101111000",
  53277=>"001111010",
  53278=>"011101111",
  53279=>"010101110",
  53280=>"001001000",
  53281=>"110011011",
  53282=>"000100100",
  53283=>"110000111",
  53284=>"011111011",
  53285=>"100100011",
  53286=>"000101100",
  53287=>"000011011",
  53288=>"111001000",
  53289=>"101010001",
  53290=>"000110110",
  53291=>"101110000",
  53292=>"000001000",
  53293=>"101011101",
  53294=>"101111101",
  53295=>"001010000",
  53296=>"000100101",
  53297=>"010000100",
  53298=>"101010011",
  53299=>"001010111",
  53300=>"101110011",
  53301=>"010000101",
  53302=>"111101111",
  53303=>"100001110",
  53304=>"011000011",
  53305=>"100001110",
  53306=>"101110000",
  53307=>"100101100",
  53308=>"011101110",
  53309=>"111011011",
  53310=>"011001100",
  53311=>"001001000",
  53312=>"000010100",
  53313=>"001000001",
  53314=>"010000111",
  53315=>"010110110",
  53316=>"100100100",
  53317=>"011010000",
  53318=>"001110000",
  53319=>"100101011",
  53320=>"010110011",
  53321=>"010000001",
  53322=>"001100110",
  53323=>"000000100",
  53324=>"110100111",
  53325=>"110111100",
  53326=>"100110101",
  53327=>"010011100",
  53328=>"011011000",
  53329=>"111000001",
  53330=>"011001101",
  53331=>"000100111",
  53332=>"111001110",
  53333=>"000100100",
  53334=>"101011111",
  53335=>"101010011",
  53336=>"111001010",
  53337=>"110010010",
  53338=>"111101011",
  53339=>"100110010",
  53340=>"000000111",
  53341=>"111100111",
  53342=>"000110101",
  53343=>"110011100",
  53344=>"101100110",
  53345=>"001011010",
  53346=>"101001000",
  53347=>"001001110",
  53348=>"111110101",
  53349=>"101001011",
  53350=>"110010110",
  53351=>"010001001",
  53352=>"101100000",
  53353=>"101100101",
  53354=>"011001111",
  53355=>"000000010",
  53356=>"011010010",
  53357=>"000000010",
  53358=>"001111111",
  53359=>"001100010",
  53360=>"000011111",
  53361=>"101000011",
  53362=>"100111110",
  53363=>"101110111",
  53364=>"010111101",
  53365=>"101111010",
  53366=>"111100101",
  53367=>"111001110",
  53368=>"000000010",
  53369=>"111011000",
  53370=>"010000010",
  53371=>"100111111",
  53372=>"001010001",
  53373=>"000001011",
  53374=>"010100101",
  53375=>"011101111",
  53376=>"111011000",
  53377=>"001111101",
  53378=>"100101001",
  53379=>"110000110",
  53380=>"001110100",
  53381=>"001001011",
  53382=>"001001110",
  53383=>"100100110",
  53384=>"111111001",
  53385=>"111111111",
  53386=>"100100100",
  53387=>"010011111",
  53388=>"001100100",
  53389=>"000111111",
  53390=>"000100111",
  53391=>"110010001",
  53392=>"100011010",
  53393=>"011000010",
  53394=>"110101010",
  53395=>"111000111",
  53396=>"011110100",
  53397=>"010000011",
  53398=>"110000111",
  53399=>"100110010",
  53400=>"100001100",
  53401=>"101001101",
  53402=>"101010000",
  53403=>"011011110",
  53404=>"000101100",
  53405=>"010011110",
  53406=>"001011001",
  53407=>"011001111",
  53408=>"000000101",
  53409=>"000001010",
  53410=>"011110000",
  53411=>"111101110",
  53412=>"000100111",
  53413=>"100010101",
  53414=>"101011001",
  53415=>"010000000",
  53416=>"001010001",
  53417=>"011010000",
  53418=>"101000101",
  53419=>"110101000",
  53420=>"111010000",
  53421=>"000101110",
  53422=>"010000000",
  53423=>"111100010",
  53424=>"100101000",
  53425=>"111100000",
  53426=>"100111110",
  53427=>"000110011",
  53428=>"001011010",
  53429=>"101010001",
  53430=>"001010110",
  53431=>"101101101",
  53432=>"001100101",
  53433=>"100100110",
  53434=>"101101100",
  53435=>"000010010",
  53436=>"010001100",
  53437=>"010111111",
  53438=>"001110000",
  53439=>"001010111",
  53440=>"111101010",
  53441=>"101001100",
  53442=>"101111110",
  53443=>"100110110",
  53444=>"011011101",
  53445=>"111100011",
  53446=>"000101011",
  53447=>"000001000",
  53448=>"000111010",
  53449=>"100011111",
  53450=>"011101011",
  53451=>"110011100",
  53452=>"110100011",
  53453=>"001011111",
  53454=>"110011001",
  53455=>"111110111",
  53456=>"010101000",
  53457=>"101001110",
  53458=>"110110101",
  53459=>"000011001",
  53460=>"010010101",
  53461=>"010000101",
  53462=>"110101101",
  53463=>"011011100",
  53464=>"000000100",
  53465=>"011011101",
  53466=>"010101111",
  53467=>"111111110",
  53468=>"110110011",
  53469=>"101000101",
  53470=>"001100111",
  53471=>"011011100",
  53472=>"101101000",
  53473=>"000000001",
  53474=>"011001110",
  53475=>"110001111",
  53476=>"100010101",
  53477=>"001101110",
  53478=>"001010110",
  53479=>"110110101",
  53480=>"011000010",
  53481=>"110110110",
  53482=>"011011101",
  53483=>"001001011",
  53484=>"001100101",
  53485=>"111101110",
  53486=>"110000001",
  53487=>"100101001",
  53488=>"110110110",
  53489=>"001001111",
  53490=>"010111001",
  53491=>"111100100",
  53492=>"011010000",
  53493=>"101100000",
  53494=>"001101000",
  53495=>"110001101",
  53496=>"000000000",
  53497=>"001111000",
  53498=>"100100100",
  53499=>"101100111",
  53500=>"101100011",
  53501=>"001010111",
  53502=>"110110000",
  53503=>"011101000",
  53504=>"001010011",
  53505=>"101011000",
  53506=>"100001111",
  53507=>"100010000",
  53508=>"000001110",
  53509=>"001010010",
  53510=>"001001010",
  53511=>"111101100",
  53512=>"101111111",
  53513=>"100111011",
  53514=>"010000000",
  53515=>"001011111",
  53516=>"101000010",
  53517=>"000101010",
  53518=>"111001100",
  53519=>"000110111",
  53520=>"100001001",
  53521=>"010100000",
  53522=>"011011111",
  53523=>"101101000",
  53524=>"110001011",
  53525=>"100101011",
  53526=>"000111111",
  53527=>"000000000",
  53528=>"011001001",
  53529=>"010101011",
  53530=>"100111011",
  53531=>"000010011",
  53532=>"111111011",
  53533=>"111000001",
  53534=>"001010011",
  53535=>"010110001",
  53536=>"110010101",
  53537=>"011110111",
  53538=>"111100101",
  53539=>"010000011",
  53540=>"000101100",
  53541=>"100110000",
  53542=>"010000111",
  53543=>"001001001",
  53544=>"110010010",
  53545=>"010100011",
  53546=>"111011011",
  53547=>"000110100",
  53548=>"101011100",
  53549=>"101101111",
  53550=>"110010100",
  53551=>"101000001",
  53552=>"111010110",
  53553=>"110101011",
  53554=>"110001001",
  53555=>"111110111",
  53556=>"111001001",
  53557=>"001000001",
  53558=>"000110011",
  53559=>"001000101",
  53560=>"111110011",
  53561=>"100101011",
  53562=>"110101001",
  53563=>"100011001",
  53564=>"001000101",
  53565=>"100111110",
  53566=>"110100110",
  53567=>"100101110",
  53568=>"100101111",
  53569=>"100101010",
  53570=>"011110100",
  53571=>"111010100",
  53572=>"011000000",
  53573=>"000010001",
  53574=>"000111100",
  53575=>"110100101",
  53576=>"100000110",
  53577=>"111101100",
  53578=>"001110000",
  53579=>"000011000",
  53580=>"111010101",
  53581=>"000001100",
  53582=>"011001101",
  53583=>"111101000",
  53584=>"100010010",
  53585=>"111010100",
  53586=>"100010001",
  53587=>"110000110",
  53588=>"000001000",
  53589=>"011001010",
  53590=>"001100100",
  53591=>"000001010",
  53592=>"010000010",
  53593=>"110110000",
  53594=>"100000011",
  53595=>"001001111",
  53596=>"110001001",
  53597=>"010100111",
  53598=>"010011011",
  53599=>"111100111",
  53600=>"110111110",
  53601=>"100010100",
  53602=>"111001110",
  53603=>"111000100",
  53604=>"111101001",
  53605=>"001000001",
  53606=>"010010111",
  53607=>"011000101",
  53608=>"111001010",
  53609=>"100000010",
  53610=>"000000010",
  53611=>"110000010",
  53612=>"000110111",
  53613=>"011000111",
  53614=>"111111101",
  53615=>"001011101",
  53616=>"000111110",
  53617=>"111111110",
  53618=>"010001110",
  53619=>"001001000",
  53620=>"011001011",
  53621=>"101100011",
  53622=>"100011111",
  53623=>"101010001",
  53624=>"001110110",
  53625=>"011100011",
  53626=>"111100000",
  53627=>"000000010",
  53628=>"001000000",
  53629=>"100111011",
  53630=>"100110101",
  53631=>"100110001",
  53632=>"000010001",
  53633=>"111111101",
  53634=>"001111001",
  53635=>"001011011",
  53636=>"010010001",
  53637=>"010101000",
  53638=>"010111110",
  53639=>"111001100",
  53640=>"111111100",
  53641=>"010000101",
  53642=>"010000010",
  53643=>"011101011",
  53644=>"101001110",
  53645=>"100000101",
  53646=>"111011111",
  53647=>"011101100",
  53648=>"010111000",
  53649=>"111010111",
  53650=>"110011111",
  53651=>"110001001",
  53652=>"011001110",
  53653=>"100111101",
  53654=>"101110000",
  53655=>"111110110",
  53656=>"010111001",
  53657=>"101110010",
  53658=>"000111010",
  53659=>"000100011",
  53660=>"110010001",
  53661=>"101110101",
  53662=>"100010110",
  53663=>"111111111",
  53664=>"010100111",
  53665=>"011100011",
  53666=>"100110010",
  53667=>"000001001",
  53668=>"100100101",
  53669=>"100111000",
  53670=>"011100000",
  53671=>"011100100",
  53672=>"100000001",
  53673=>"100010000",
  53674=>"011100100",
  53675=>"111000111",
  53676=>"101100001",
  53677=>"010011110",
  53678=>"010101101",
  53679=>"110101000",
  53680=>"101110110",
  53681=>"011110011",
  53682=>"010111100",
  53683=>"111101010",
  53684=>"001101111",
  53685=>"001100101",
  53686=>"000111101",
  53687=>"111100101",
  53688=>"111111110",
  53689=>"100101110",
  53690=>"111101100",
  53691=>"010011011",
  53692=>"000101011",
  53693=>"001010001",
  53694=>"011010110",
  53695=>"000110011",
  53696=>"001100111",
  53697=>"101001110",
  53698=>"000011111",
  53699=>"010110010",
  53700=>"101000010",
  53701=>"010110000",
  53702=>"110011011",
  53703=>"101100111",
  53704=>"100101101",
  53705=>"101110100",
  53706=>"111101000",
  53707=>"100011000",
  53708=>"010100110",
  53709=>"100100111",
  53710=>"100110011",
  53711=>"100111000",
  53712=>"010011011",
  53713=>"111011010",
  53714=>"110011110",
  53715=>"101111101",
  53716=>"001011111",
  53717=>"101110011",
  53718=>"100010100",
  53719=>"010010001",
  53720=>"111001100",
  53721=>"100000110",
  53722=>"000000100",
  53723=>"010000010",
  53724=>"111000001",
  53725=>"101100010",
  53726=>"011100111",
  53727=>"110011110",
  53728=>"001101000",
  53729=>"000110100",
  53730=>"001101000",
  53731=>"000101001",
  53732=>"101110001",
  53733=>"000001000",
  53734=>"000111100",
  53735=>"101001001",
  53736=>"001011110",
  53737=>"101110011",
  53738=>"011000110",
  53739=>"111011010",
  53740=>"100010101",
  53741=>"111111000",
  53742=>"110000110",
  53743=>"111010101",
  53744=>"110110111",
  53745=>"001111110",
  53746=>"111001000",
  53747=>"000000110",
  53748=>"101000001",
  53749=>"011010111",
  53750=>"011110000",
  53751=>"010100101",
  53752=>"101111110",
  53753=>"101010010",
  53754=>"010001101",
  53755=>"011111110",
  53756=>"000000010",
  53757=>"011011111",
  53758=>"100000111",
  53759=>"111000010",
  53760=>"110101111",
  53761=>"000000000",
  53762=>"111110111",
  53763=>"110100000",
  53764=>"001010100",
  53765=>"110000111",
  53766=>"000110011",
  53767=>"011010011",
  53768=>"011000001",
  53769=>"100011100",
  53770=>"110011011",
  53771=>"011000000",
  53772=>"111000110",
  53773=>"101101101",
  53774=>"111000000",
  53775=>"001110101",
  53776=>"100111011",
  53777=>"010101011",
  53778=>"010100010",
  53779=>"101001110",
  53780=>"001100101",
  53781=>"000000000",
  53782=>"100111011",
  53783=>"000100101",
  53784=>"111001010",
  53785=>"100011100",
  53786=>"010101100",
  53787=>"010010011",
  53788=>"111001010",
  53789=>"011110100",
  53790=>"001011000",
  53791=>"100111000",
  53792=>"010111000",
  53793=>"011100101",
  53794=>"011010000",
  53795=>"000011111",
  53796=>"011101101",
  53797=>"110110100",
  53798=>"110111011",
  53799=>"010110110",
  53800=>"011000100",
  53801=>"000011111",
  53802=>"001100010",
  53803=>"001110001",
  53804=>"001100000",
  53805=>"011110010",
  53806=>"111101010",
  53807=>"110000011",
  53808=>"101000000",
  53809=>"110100110",
  53810=>"011011101",
  53811=>"001000111",
  53812=>"001100001",
  53813=>"010100101",
  53814=>"001010111",
  53815=>"111000001",
  53816=>"111011011",
  53817=>"000001001",
  53818=>"101101111",
  53819=>"010111111",
  53820=>"000011110",
  53821=>"010001100",
  53822=>"001001000",
  53823=>"010000000",
  53824=>"000010111",
  53825=>"111110110",
  53826=>"001100100",
  53827=>"111010001",
  53828=>"111101100",
  53829=>"001011110",
  53830=>"000101001",
  53831=>"011011000",
  53832=>"000111001",
  53833=>"010001111",
  53834=>"100011000",
  53835=>"001001011",
  53836=>"011000111",
  53837=>"101011000",
  53838=>"010011000",
  53839=>"011101101",
  53840=>"001001101",
  53841=>"111001111",
  53842=>"100101101",
  53843=>"000100011",
  53844=>"100000011",
  53845=>"010100101",
  53846=>"110100110",
  53847=>"011110011",
  53848=>"000101110",
  53849=>"011100100",
  53850=>"101000001",
  53851=>"111001011",
  53852=>"011111101",
  53853=>"101000100",
  53854=>"100110100",
  53855=>"101110010",
  53856=>"101101101",
  53857=>"101110110",
  53858=>"110100111",
  53859=>"011011100",
  53860=>"110001101",
  53861=>"110100000",
  53862=>"011001010",
  53863=>"010000010",
  53864=>"000110011",
  53865=>"011001100",
  53866=>"001100011",
  53867=>"101101101",
  53868=>"100110000",
  53869=>"010000111",
  53870=>"000110011",
  53871=>"100010000",
  53872=>"110110000",
  53873=>"100000000",
  53874=>"110101101",
  53875=>"000000010",
  53876=>"100100101",
  53877=>"111010001",
  53878=>"101001111",
  53879=>"100111111",
  53880=>"011100001",
  53881=>"101000110",
  53882=>"000110000",
  53883=>"101101111",
  53884=>"000111101",
  53885=>"111001011",
  53886=>"110100101",
  53887=>"000001001",
  53888=>"101101111",
  53889=>"011101010",
  53890=>"000001111",
  53891=>"001100100",
  53892=>"001011010",
  53893=>"111011010",
  53894=>"111100101",
  53895=>"111101000",
  53896=>"010000101",
  53897=>"011010100",
  53898=>"011100110",
  53899=>"001010011",
  53900=>"110011001",
  53901=>"101000000",
  53902=>"100010111",
  53903=>"001110100",
  53904=>"100000001",
  53905=>"110100001",
  53906=>"001001101",
  53907=>"111010000",
  53908=>"100011110",
  53909=>"100101011",
  53910=>"000100001",
  53911=>"111110100",
  53912=>"111111010",
  53913=>"100101010",
  53914=>"000110100",
  53915=>"000010010",
  53916=>"111010110",
  53917=>"010000100",
  53918=>"110001000",
  53919=>"000100110",
  53920=>"111011110",
  53921=>"100000100",
  53922=>"111000011",
  53923=>"111000001",
  53924=>"010010011",
  53925=>"111100111",
  53926=>"001100101",
  53927=>"101011100",
  53928=>"010010000",
  53929=>"000000101",
  53930=>"111011010",
  53931=>"100110011",
  53932=>"010101011",
  53933=>"000101100",
  53934=>"101101010",
  53935=>"000001000",
  53936=>"101110110",
  53937=>"000001001",
  53938=>"111100110",
  53939=>"111000001",
  53940=>"010001111",
  53941=>"001000000",
  53942=>"001111101",
  53943=>"100100000",
  53944=>"110001011",
  53945=>"011001011",
  53946=>"001100110",
  53947=>"111011000",
  53948=>"001101111",
  53949=>"010011001",
  53950=>"011101000",
  53951=>"110011111",
  53952=>"101010101",
  53953=>"100101011",
  53954=>"111010010",
  53955=>"110101001",
  53956=>"101111000",
  53957=>"111100100",
  53958=>"011110100",
  53959=>"111000010",
  53960=>"111101000",
  53961=>"100100101",
  53962=>"100011000",
  53963=>"000010111",
  53964=>"100100101",
  53965=>"111101011",
  53966=>"011011101",
  53967=>"110001001",
  53968=>"111111010",
  53969=>"001000110",
  53970=>"000000101",
  53971=>"000101111",
  53972=>"001011111",
  53973=>"011101101",
  53974=>"010100111",
  53975=>"110100001",
  53976=>"001010100",
  53977=>"001000000",
  53978=>"111010100",
  53979=>"101111011",
  53980=>"001101010",
  53981=>"000110001",
  53982=>"001100010",
  53983=>"101100001",
  53984=>"111011001",
  53985=>"101011001",
  53986=>"001100010",
  53987=>"110011011",
  53988=>"101110101",
  53989=>"001110101",
  53990=>"110101111",
  53991=>"111011101",
  53992=>"100101101",
  53993=>"111001000",
  53994=>"001011010",
  53995=>"010111000",
  53996=>"011111101",
  53997=>"010001011",
  53998=>"101111000",
  53999=>"010111110",
  54000=>"001111111",
  54001=>"010010101",
  54002=>"111110100",
  54003=>"001101000",
  54004=>"101011110",
  54005=>"011100110",
  54006=>"101101010",
  54007=>"001011111",
  54008=>"001100001",
  54009=>"110011101",
  54010=>"111001001",
  54011=>"001111000",
  54012=>"110001111",
  54013=>"111001100",
  54014=>"111011000",
  54015=>"011010101",
  54016=>"010001010",
  54017=>"111000001",
  54018=>"010110100",
  54019=>"110000111",
  54020=>"000101000",
  54021=>"011000110",
  54022=>"100011000",
  54023=>"001011000",
  54024=>"001001011",
  54025=>"101001001",
  54026=>"001010101",
  54027=>"100001000",
  54028=>"101101001",
  54029=>"010111100",
  54030=>"111111100",
  54031=>"011001100",
  54032=>"110111111",
  54033=>"001101011",
  54034=>"011010100",
  54035=>"110111101",
  54036=>"110001010",
  54037=>"000101011",
  54038=>"111101110",
  54039=>"111010100",
  54040=>"101101101",
  54041=>"111100100",
  54042=>"010011100",
  54043=>"010101000",
  54044=>"110111001",
  54045=>"110111101",
  54046=>"111101011",
  54047=>"101111011",
  54048=>"111101100",
  54049=>"100000100",
  54050=>"000000000",
  54051=>"001101101",
  54052=>"011000111",
  54053=>"100011100",
  54054=>"011010010",
  54055=>"111110101",
  54056=>"110110110",
  54057=>"100110000",
  54058=>"101001101",
  54059=>"101101110",
  54060=>"100010010",
  54061=>"111111101",
  54062=>"011110100",
  54063=>"111111111",
  54064=>"111101011",
  54065=>"001110100",
  54066=>"110100010",
  54067=>"010010111",
  54068=>"010001111",
  54069=>"011001110",
  54070=>"000010011",
  54071=>"100010110",
  54072=>"110011001",
  54073=>"011011000",
  54074=>"101000001",
  54075=>"000110100",
  54076=>"000000011",
  54077=>"000000000",
  54078=>"111001011",
  54079=>"011000111",
  54080=>"101101111",
  54081=>"000010001",
  54082=>"011110111",
  54083=>"111101001",
  54084=>"111100001",
  54085=>"010001010",
  54086=>"111010101",
  54087=>"101001111",
  54088=>"000010010",
  54089=>"000101100",
  54090=>"001111111",
  54091=>"011011010",
  54092=>"010101101",
  54093=>"110110011",
  54094=>"111000000",
  54095=>"111001110",
  54096=>"000110100",
  54097=>"011101111",
  54098=>"101111101",
  54099=>"001000100",
  54100=>"101101100",
  54101=>"111000000",
  54102=>"111110001",
  54103=>"100010011",
  54104=>"111010011",
  54105=>"100111011",
  54106=>"100100100",
  54107=>"111111110",
  54108=>"100110111",
  54109=>"000011001",
  54110=>"100111001",
  54111=>"110100010",
  54112=>"000000000",
  54113=>"110001100",
  54114=>"001110101",
  54115=>"011110100",
  54116=>"101011100",
  54117=>"010101000",
  54118=>"110001111",
  54119=>"000100101",
  54120=>"010011110",
  54121=>"000010001",
  54122=>"100111100",
  54123=>"110010000",
  54124=>"101100110",
  54125=>"110001000",
  54126=>"100000111",
  54127=>"010000001",
  54128=>"100100001",
  54129=>"101110010",
  54130=>"010011100",
  54131=>"011101010",
  54132=>"010110000",
  54133=>"111001111",
  54134=>"101101001",
  54135=>"000001000",
  54136=>"101100001",
  54137=>"010100101",
  54138=>"001001100",
  54139=>"110101100",
  54140=>"001101100",
  54141=>"000101111",
  54142=>"100111010",
  54143=>"010011010",
  54144=>"101011011",
  54145=>"000101101",
  54146=>"101000010",
  54147=>"010111001",
  54148=>"000100010",
  54149=>"010111110",
  54150=>"000110101",
  54151=>"010011111",
  54152=>"110000001",
  54153=>"011001111",
  54154=>"101111110",
  54155=>"001011111",
  54156=>"000101010",
  54157=>"111000011",
  54158=>"110101111",
  54159=>"111010011",
  54160=>"001010011",
  54161=>"011100001",
  54162=>"011000101",
  54163=>"110100000",
  54164=>"100000101",
  54165=>"011001100",
  54166=>"100000010",
  54167=>"001110101",
  54168=>"100010010",
  54169=>"000010001",
  54170=>"111001001",
  54171=>"100111100",
  54172=>"100011110",
  54173=>"001000100",
  54174=>"111100111",
  54175=>"110101100",
  54176=>"001111011",
  54177=>"010111100",
  54178=>"101110111",
  54179=>"011011001",
  54180=>"111100101",
  54181=>"010110110",
  54182=>"101000010",
  54183=>"001110000",
  54184=>"001001101",
  54185=>"011111111",
  54186=>"111101110",
  54187=>"011101010",
  54188=>"100000001",
  54189=>"011101001",
  54190=>"110010101",
  54191=>"011111000",
  54192=>"100001000",
  54193=>"000010101",
  54194=>"110000001",
  54195=>"010000111",
  54196=>"101111011",
  54197=>"000101111",
  54198=>"011000011",
  54199=>"101000111",
  54200=>"100011000",
  54201=>"011101100",
  54202=>"101110010",
  54203=>"010100011",
  54204=>"010110110",
  54205=>"000101010",
  54206=>"100111111",
  54207=>"111100111",
  54208=>"111010011",
  54209=>"110001010",
  54210=>"111101001",
  54211=>"011010010",
  54212=>"001101100",
  54213=>"000111010",
  54214=>"110100100",
  54215=>"000010010",
  54216=>"000011001",
  54217=>"010010000",
  54218=>"101101111",
  54219=>"000101111",
  54220=>"100001111",
  54221=>"110011111",
  54222=>"101001111",
  54223=>"000101111",
  54224=>"100100001",
  54225=>"100110011",
  54226=>"111110010",
  54227=>"111000100",
  54228=>"100110011",
  54229=>"111110100",
  54230=>"100001000",
  54231=>"101101111",
  54232=>"000000101",
  54233=>"011110110",
  54234=>"111001100",
  54235=>"100100000",
  54236=>"000010001",
  54237=>"011101101",
  54238=>"101110110",
  54239=>"110011100",
  54240=>"000001101",
  54241=>"010111101",
  54242=>"010011101",
  54243=>"111001000",
  54244=>"010000011",
  54245=>"101001111",
  54246=>"011001001",
  54247=>"111001110",
  54248=>"111111000",
  54249=>"010110000",
  54250=>"101000000",
  54251=>"010011000",
  54252=>"010111101",
  54253=>"110000011",
  54254=>"001101101",
  54255=>"010100011",
  54256=>"001000011",
  54257=>"110001011",
  54258=>"000100110",
  54259=>"001100011",
  54260=>"101100011",
  54261=>"100101001",
  54262=>"101100001",
  54263=>"001101001",
  54264=>"101001110",
  54265=>"100000011",
  54266=>"000100001",
  54267=>"111110100",
  54268=>"010000011",
  54269=>"100001110",
  54270=>"001111110",
  54271=>"100010011",
  54272=>"101001111",
  54273=>"111001101",
  54274=>"011011101",
  54275=>"001000100",
  54276=>"110110111",
  54277=>"101000000",
  54278=>"010101010",
  54279=>"001101011",
  54280=>"110101011",
  54281=>"111010101",
  54282=>"000001000",
  54283=>"101011100",
  54284=>"111000111",
  54285=>"010100101",
  54286=>"111000001",
  54287=>"001101010",
  54288=>"011010111",
  54289=>"110101101",
  54290=>"110001001",
  54291=>"000011101",
  54292=>"010111100",
  54293=>"100001101",
  54294=>"110011111",
  54295=>"111111111",
  54296=>"100100010",
  54297=>"010101011",
  54298=>"001101110",
  54299=>"011011111",
  54300=>"011110110",
  54301=>"101111111",
  54302=>"001111010",
  54303=>"101101000",
  54304=>"000110111",
  54305=>"011101001",
  54306=>"000111110",
  54307=>"000100011",
  54308=>"110111100",
  54309=>"110000001",
  54310=>"100101011",
  54311=>"101010001",
  54312=>"100111001",
  54313=>"000010110",
  54314=>"000010110",
  54315=>"100100100",
  54316=>"101111001",
  54317=>"010100110",
  54318=>"001000010",
  54319=>"110111000",
  54320=>"101111101",
  54321=>"000001011",
  54322=>"101101100",
  54323=>"100011110",
  54324=>"010010000",
  54325=>"000110111",
  54326=>"111010111",
  54327=>"010000100",
  54328=>"100000100",
  54329=>"011000000",
  54330=>"001011111",
  54331=>"000000111",
  54332=>"111000001",
  54333=>"000000010",
  54334=>"101100111",
  54335=>"000101000",
  54336=>"111111110",
  54337=>"101100110",
  54338=>"110010100",
  54339=>"000111000",
  54340=>"010000001",
  54341=>"011011100",
  54342=>"110010101",
  54343=>"000000101",
  54344=>"000010100",
  54345=>"011011011",
  54346=>"001000110",
  54347=>"111001101",
  54348=>"101000100",
  54349=>"101101010",
  54350=>"110111111",
  54351=>"100000000",
  54352=>"110101100",
  54353=>"111101111",
  54354=>"100011001",
  54355=>"000011110",
  54356=>"100011101",
  54357=>"101111101",
  54358=>"001011111",
  54359=>"111111011",
  54360=>"011000111",
  54361=>"011110101",
  54362=>"111001100",
  54363=>"111010010",
  54364=>"000111110",
  54365=>"001001011",
  54366=>"001010011",
  54367=>"111110011",
  54368=>"010000010",
  54369=>"101001011",
  54370=>"110000000",
  54371=>"000011100",
  54372=>"101111000",
  54373=>"011100010",
  54374=>"000110000",
  54375=>"111011111",
  54376=>"111100010",
  54377=>"000011000",
  54378=>"010010010",
  54379=>"010010100",
  54380=>"111001001",
  54381=>"101011011",
  54382=>"000111010",
  54383=>"011100001",
  54384=>"111010011",
  54385=>"010111101",
  54386=>"111101011",
  54387=>"100111100",
  54388=>"110001100",
  54389=>"111000110",
  54390=>"000110110",
  54391=>"000101110",
  54392=>"010100100",
  54393=>"001001101",
  54394=>"110101011",
  54395=>"100010010",
  54396=>"111110101",
  54397=>"111111110",
  54398=>"111010000",
  54399=>"010101000",
  54400=>"101010100",
  54401=>"001001011",
  54402=>"110101110",
  54403=>"101001111",
  54404=>"010110000",
  54405=>"000001000",
  54406=>"001111110",
  54407=>"000011010",
  54408=>"000101110",
  54409=>"100000110",
  54410=>"111010010",
  54411=>"010101000",
  54412=>"001110110",
  54413=>"010011110",
  54414=>"101001111",
  54415=>"000100100",
  54416=>"110001000",
  54417=>"100001011",
  54418=>"111101110",
  54419=>"011000010",
  54420=>"011110111",
  54421=>"010011111",
  54422=>"111011111",
  54423=>"110011100",
  54424=>"100010001",
  54425=>"100111010",
  54426=>"101111111",
  54427=>"011011111",
  54428=>"101110011",
  54429=>"001010001",
  54430=>"011111010",
  54431=>"001000010",
  54432=>"001101111",
  54433=>"100111000",
  54434=>"000010010",
  54435=>"010011101",
  54436=>"101110101",
  54437=>"111010010",
  54438=>"100100000",
  54439=>"000001010",
  54440=>"011000101",
  54441=>"011001011",
  54442=>"100111111",
  54443=>"101010111",
  54444=>"101000101",
  54445=>"110001100",
  54446=>"010110111",
  54447=>"111001111",
  54448=>"010101110",
  54449=>"001000100",
  54450=>"011001101",
  54451=>"101111111",
  54452=>"100000001",
  54453=>"110101000",
  54454=>"000111000",
  54455=>"101000111",
  54456=>"011111001",
  54457=>"111011110",
  54458=>"101101100",
  54459=>"100101001",
  54460=>"000000001",
  54461=>"101000110",
  54462=>"111111101",
  54463=>"010000000",
  54464=>"110101010",
  54465=>"111101000",
  54466=>"100111111",
  54467=>"000010011",
  54468=>"010001110",
  54469=>"111110011",
  54470=>"111110110",
  54471=>"111011101",
  54472=>"010100000",
  54473=>"011010011",
  54474=>"111101100",
  54475=>"011100010",
  54476=>"101110111",
  54477=>"101000101",
  54478=>"011110011",
  54479=>"010000100",
  54480=>"010100111",
  54481=>"001111000",
  54482=>"101011110",
  54483=>"101100101",
  54484=>"001100001",
  54485=>"010010000",
  54486=>"101011110",
  54487=>"101111000",
  54488=>"010010001",
  54489=>"101101111",
  54490=>"000111000",
  54491=>"111101111",
  54492=>"111000011",
  54493=>"000110010",
  54494=>"101011011",
  54495=>"100011011",
  54496=>"010110111",
  54497=>"111111111",
  54498=>"000110001",
  54499=>"111110000",
  54500=>"101000101",
  54501=>"011010010",
  54502=>"111011101",
  54503=>"111110100",
  54504=>"110100100",
  54505=>"011001000",
  54506=>"010111111",
  54507=>"101010011",
  54508=>"110111111",
  54509=>"111101010",
  54510=>"011111011",
  54511=>"001000000",
  54512=>"111000011",
  54513=>"101000000",
  54514=>"011010111",
  54515=>"111111101",
  54516=>"001101010",
  54517=>"110111111",
  54518=>"011111110",
  54519=>"100011001",
  54520=>"010001011",
  54521=>"001000100",
  54522=>"001010101",
  54523=>"000100011",
  54524=>"011100101",
  54525=>"011000011",
  54526=>"001001000",
  54527=>"001101101",
  54528=>"100110110",
  54529=>"011000100",
  54530=>"111011010",
  54531=>"000011010",
  54532=>"100010010",
  54533=>"010110000",
  54534=>"001110011",
  54535=>"100000000",
  54536=>"001111101",
  54537=>"000001101",
  54538=>"000100100",
  54539=>"111100011",
  54540=>"011110010",
  54541=>"110011000",
  54542=>"111111011",
  54543=>"101000000",
  54544=>"100111111",
  54545=>"110011110",
  54546=>"100110001",
  54547=>"110100101",
  54548=>"111111111",
  54549=>"011110001",
  54550=>"100100101",
  54551=>"101111100",
  54552=>"100100011",
  54553=>"100001101",
  54554=>"001100011",
  54555=>"100101001",
  54556=>"011000010",
  54557=>"101001001",
  54558=>"001010110",
  54559=>"000001011",
  54560=>"010001001",
  54561=>"011000101",
  54562=>"101011011",
  54563=>"000001110",
  54564=>"100000000",
  54565=>"001000101",
  54566=>"110001000",
  54567=>"000111001",
  54568=>"000001001",
  54569=>"001001101",
  54570=>"011101001",
  54571=>"001011100",
  54572=>"000111111",
  54573=>"101011010",
  54574=>"010110111",
  54575=>"110111101",
  54576=>"000101101",
  54577=>"011010000",
  54578=>"110101111",
  54579=>"000010001",
  54580=>"000111011",
  54581=>"001001100",
  54582=>"000001000",
  54583=>"111101010",
  54584=>"000111100",
  54585=>"111001000",
  54586=>"010010010",
  54587=>"010000100",
  54588=>"110110100",
  54589=>"110010011",
  54590=>"001000010",
  54591=>"110100111",
  54592=>"100000000",
  54593=>"000000111",
  54594=>"101111100",
  54595=>"100100100",
  54596=>"111111110",
  54597=>"101010111",
  54598=>"110111101",
  54599=>"000110101",
  54600=>"000100011",
  54601=>"001000001",
  54602=>"101110010",
  54603=>"011101100",
  54604=>"010001111",
  54605=>"110010011",
  54606=>"000000000",
  54607=>"100011110",
  54608=>"000010000",
  54609=>"100110111",
  54610=>"110001010",
  54611=>"001001001",
  54612=>"100001010",
  54613=>"101000111",
  54614=>"011001110",
  54615=>"101101000",
  54616=>"101100111",
  54617=>"000000111",
  54618=>"011101001",
  54619=>"101011111",
  54620=>"010110011",
  54621=>"100001110",
  54622=>"001000100",
  54623=>"101101000",
  54624=>"110100010",
  54625=>"101010100",
  54626=>"111001111",
  54627=>"000111010",
  54628=>"001000010",
  54629=>"011110010",
  54630=>"010000000",
  54631=>"011010000",
  54632=>"111100110",
  54633=>"111001011",
  54634=>"101000110",
  54635=>"000000010",
  54636=>"101000101",
  54637=>"111001001",
  54638=>"101001110",
  54639=>"100110100",
  54640=>"010001110",
  54641=>"010000111",
  54642=>"111001011",
  54643=>"001101000",
  54644=>"111001000",
  54645=>"111001100",
  54646=>"000001000",
  54647=>"101011000",
  54648=>"100000011",
  54649=>"110101110",
  54650=>"110110110",
  54651=>"110111000",
  54652=>"001111111",
  54653=>"101010010",
  54654=>"110011001",
  54655=>"011011011",
  54656=>"111011000",
  54657=>"001100100",
  54658=>"110111100",
  54659=>"001011111",
  54660=>"101010011",
  54661=>"101101010",
  54662=>"110000000",
  54663=>"110011110",
  54664=>"010111011",
  54665=>"100000111",
  54666=>"011011010",
  54667=>"010010001",
  54668=>"000011100",
  54669=>"001101111",
  54670=>"100010001",
  54671=>"100110100",
  54672=>"101100101",
  54673=>"101111111",
  54674=>"111100111",
  54675=>"011000011",
  54676=>"011011000",
  54677=>"010000001",
  54678=>"001100100",
  54679=>"110000001",
  54680=>"100000111",
  54681=>"110000010",
  54682=>"111001100",
  54683=>"111111100",
  54684=>"111011001",
  54685=>"111100111",
  54686=>"010011101",
  54687=>"111111101",
  54688=>"000101011",
  54689=>"000010001",
  54690=>"000010111",
  54691=>"111000010",
  54692=>"001101001",
  54693=>"011100110",
  54694=>"001001011",
  54695=>"111000010",
  54696=>"111010011",
  54697=>"101111000",
  54698=>"000000110",
  54699=>"110110101",
  54700=>"110011111",
  54701=>"111100011",
  54702=>"111100000",
  54703=>"010010010",
  54704=>"011110101",
  54705=>"110100100",
  54706=>"001000101",
  54707=>"111010001",
  54708=>"100001111",
  54709=>"011101110",
  54710=>"001000100",
  54711=>"110111111",
  54712=>"001001111",
  54713=>"111011111",
  54714=>"001111100",
  54715=>"011010011",
  54716=>"110110010",
  54717=>"110101010",
  54718=>"110001111",
  54719=>"011110010",
  54720=>"101110010",
  54721=>"111110010",
  54722=>"010110010",
  54723=>"010100100",
  54724=>"100000111",
  54725=>"101101010",
  54726=>"000101100",
  54727=>"100101001",
  54728=>"000001101",
  54729=>"011110010",
  54730=>"111100010",
  54731=>"100110011",
  54732=>"010001000",
  54733=>"000010111",
  54734=>"010010100",
  54735=>"001101100",
  54736=>"010100110",
  54737=>"010101011",
  54738=>"111111100",
  54739=>"101111101",
  54740=>"100011000",
  54741=>"010011001",
  54742=>"010000010",
  54743=>"101000111",
  54744=>"110001000",
  54745=>"000010101",
  54746=>"110011001",
  54747=>"001011001",
  54748=>"010011110",
  54749=>"111001000",
  54750=>"111111010",
  54751=>"100100111",
  54752=>"000111101",
  54753=>"000101010",
  54754=>"111001001",
  54755=>"010100000",
  54756=>"110110001",
  54757=>"111001111",
  54758=>"111011010",
  54759=>"111111010",
  54760=>"111010111",
  54761=>"010111011",
  54762=>"101101010",
  54763=>"100010100",
  54764=>"000010001",
  54765=>"011000000",
  54766=>"010000000",
  54767=>"000000110",
  54768=>"110000000",
  54769=>"011110101",
  54770=>"011010010",
  54771=>"101100011",
  54772=>"011111100",
  54773=>"100100101",
  54774=>"101000100",
  54775=>"000101101",
  54776=>"011011111",
  54777=>"101110101",
  54778=>"011111110",
  54779=>"001000111",
  54780=>"000001100",
  54781=>"011010010",
  54782=>"001010111",
  54783=>"000110011",
  54784=>"100010110",
  54785=>"101001000",
  54786=>"001100001",
  54787=>"000101000",
  54788=>"110110000",
  54789=>"011010011",
  54790=>"111100001",
  54791=>"110001101",
  54792=>"010101111",
  54793=>"110000101",
  54794=>"001001001",
  54795=>"000100110",
  54796=>"101011101",
  54797=>"000101101",
  54798=>"101001110",
  54799=>"111101010",
  54800=>"011111111",
  54801=>"011100111",
  54802=>"100111110",
  54803=>"000101101",
  54804=>"010001000",
  54805=>"101111011",
  54806=>"100000000",
  54807=>"010100001",
  54808=>"001010111",
  54809=>"011010001",
  54810=>"010110000",
  54811=>"101000000",
  54812=>"001111011",
  54813=>"001010111",
  54814=>"001100110",
  54815=>"111110111",
  54816=>"001011000",
  54817=>"110010011",
  54818=>"001100010",
  54819=>"010001111",
  54820=>"010100110",
  54821=>"110111111",
  54822=>"111001011",
  54823=>"101010001",
  54824=>"000010010",
  54825=>"001101110",
  54826=>"011010101",
  54827=>"101111001",
  54828=>"000101000",
  54829=>"101111100",
  54830=>"000010011",
  54831=>"111100111",
  54832=>"101010111",
  54833=>"111111111",
  54834=>"110111100",
  54835=>"101101001",
  54836=>"001010101",
  54837=>"101001111",
  54838=>"001010010",
  54839=>"010001000",
  54840=>"000010110",
  54841=>"101000010",
  54842=>"011010110",
  54843=>"111011010",
  54844=>"110010110",
  54845=>"111111100",
  54846=>"011110010",
  54847=>"001010111",
  54848=>"111000001",
  54849=>"101111110",
  54850=>"100101110",
  54851=>"000110111",
  54852=>"011000100",
  54853=>"110000001",
  54854=>"101011100",
  54855=>"001101100",
  54856=>"100001000",
  54857=>"110011101",
  54858=>"101101000",
  54859=>"011010010",
  54860=>"000010101",
  54861=>"101100011",
  54862=>"011111010",
  54863=>"000100010",
  54864=>"010101111",
  54865=>"101010000",
  54866=>"111010010",
  54867=>"001000011",
  54868=>"100001010",
  54869=>"111111101",
  54870=>"000110101",
  54871=>"010100010",
  54872=>"000010101",
  54873=>"010000000",
  54874=>"000000101",
  54875=>"000111110",
  54876=>"011101110",
  54877=>"111101100",
  54878=>"010111011",
  54879=>"110001100",
  54880=>"110111010",
  54881=>"001111011",
  54882=>"111111110",
  54883=>"111000000",
  54884=>"011010000",
  54885=>"100000011",
  54886=>"111100011",
  54887=>"011110000",
  54888=>"101101001",
  54889=>"111101000",
  54890=>"111001011",
  54891=>"101000101",
  54892=>"001000011",
  54893=>"110011011",
  54894=>"111001011",
  54895=>"111111111",
  54896=>"110010111",
  54897=>"011010101",
  54898=>"100110101",
  54899=>"101101010",
  54900=>"000011100",
  54901=>"000111110",
  54902=>"000100111",
  54903=>"000111001",
  54904=>"000100100",
  54905=>"111111110",
  54906=>"111010001",
  54907=>"000011001",
  54908=>"010100000",
  54909=>"010011011",
  54910=>"100000101",
  54911=>"011001010",
  54912=>"101001000",
  54913=>"011100011",
  54914=>"000000000",
  54915=>"110010110",
  54916=>"000101101",
  54917=>"100110001",
  54918=>"000111011",
  54919=>"110000100",
  54920=>"111110111",
  54921=>"110000000",
  54922=>"100001100",
  54923=>"110000011",
  54924=>"010010000",
  54925=>"000100111",
  54926=>"100101000",
  54927=>"001010110",
  54928=>"100011101",
  54929=>"000011011",
  54930=>"110101100",
  54931=>"110010011",
  54932=>"010110110",
  54933=>"001001111",
  54934=>"110111011",
  54935=>"001010011",
  54936=>"001010000",
  54937=>"110111110",
  54938=>"111010101",
  54939=>"100111100",
  54940=>"111111100",
  54941=>"000011000",
  54942=>"011010111",
  54943=>"000110011",
  54944=>"010011101",
  54945=>"011101101",
  54946=>"110100110",
  54947=>"000001111",
  54948=>"011101101",
  54949=>"110001011",
  54950=>"011011010",
  54951=>"101011011",
  54952=>"011101101",
  54953=>"110100000",
  54954=>"110111111",
  54955=>"011000010",
  54956=>"010110000",
  54957=>"110110111",
  54958=>"000001011",
  54959=>"111011000",
  54960=>"000011001",
  54961=>"110011000",
  54962=>"001001010",
  54963=>"110100000",
  54964=>"010101011",
  54965=>"111101111",
  54966=>"001001101",
  54967=>"000100101",
  54968=>"110100100",
  54969=>"011100101",
  54970=>"101111100",
  54971=>"111111100",
  54972=>"111000001",
  54973=>"011000111",
  54974=>"101101010",
  54975=>"000000011",
  54976=>"111100111",
  54977=>"010111101",
  54978=>"000101011",
  54979=>"111011100",
  54980=>"001100001",
  54981=>"011000101",
  54982=>"110101110",
  54983=>"000111001",
  54984=>"001111001",
  54985=>"110101100",
  54986=>"100100001",
  54987=>"110101010",
  54988=>"101111011",
  54989=>"110000011",
  54990=>"010011100",
  54991=>"011110011",
  54992=>"111110011",
  54993=>"100010111",
  54994=>"110110111",
  54995=>"001100001",
  54996=>"101010100",
  54997=>"101000000",
  54998=>"110101011",
  54999=>"001010000",
  55000=>"010110011",
  55001=>"100011000",
  55002=>"000100000",
  55003=>"100111000",
  55004=>"001010101",
  55005=>"110111110",
  55006=>"010010101",
  55007=>"110101111",
  55008=>"100010101",
  55009=>"000010011",
  55010=>"010000100",
  55011=>"011000100",
  55012=>"001000001",
  55013=>"101110100",
  55014=>"111000000",
  55015=>"101101000",
  55016=>"111001011",
  55017=>"011100001",
  55018=>"010100111",
  55019=>"111011111",
  55020=>"101010000",
  55021=>"100111110",
  55022=>"001100001",
  55023=>"011101000",
  55024=>"111001100",
  55025=>"001100010",
  55026=>"101101101",
  55027=>"010100111",
  55028=>"101011011",
  55029=>"011111000",
  55030=>"000010000",
  55031=>"110011111",
  55032=>"100101011",
  55033=>"000011110",
  55034=>"101011110",
  55035=>"010010010",
  55036=>"010101011",
  55037=>"110101110",
  55038=>"010001001",
  55039=>"000100000",
  55040=>"111111011",
  55041=>"000100111",
  55042=>"101010111",
  55043=>"100001101",
  55044=>"101110001",
  55045=>"111100111",
  55046=>"101000011",
  55047=>"001000100",
  55048=>"000000000",
  55049=>"010011100",
  55050=>"000111111",
  55051=>"001001100",
  55052=>"100000111",
  55053=>"000000000",
  55054=>"100001011",
  55055=>"100101011",
  55056=>"001010111",
  55057=>"000010111",
  55058=>"110010110",
  55059=>"110101111",
  55060=>"101101011",
  55061=>"111110000",
  55062=>"010110111",
  55063=>"100000011",
  55064=>"110000111",
  55065=>"001101110",
  55066=>"111010000",
  55067=>"000100000",
  55068=>"011011000",
  55069=>"001001010",
  55070=>"110101011",
  55071=>"000011011",
  55072=>"110111101",
  55073=>"111000111",
  55074=>"110001000",
  55075=>"101001101",
  55076=>"000001100",
  55077=>"111010110",
  55078=>"010011000",
  55079=>"011101101",
  55080=>"000100111",
  55081=>"000110100",
  55082=>"111011111",
  55083=>"000010111",
  55084=>"100100000",
  55085=>"000110000",
  55086=>"011101011",
  55087=>"101001110",
  55088=>"111011111",
  55089=>"001101101",
  55090=>"001011111",
  55091=>"101001110",
  55092=>"101100010",
  55093=>"100101000",
  55094=>"001111100",
  55095=>"111100100",
  55096=>"110110001",
  55097=>"010110010",
  55098=>"001111111",
  55099=>"100010111",
  55100=>"100100100",
  55101=>"001110000",
  55102=>"111100100",
  55103=>"011100001",
  55104=>"101110001",
  55105=>"111011101",
  55106=>"001000101",
  55107=>"010100011",
  55108=>"100101101",
  55109=>"001100101",
  55110=>"011101011",
  55111=>"101011010",
  55112=>"000100100",
  55113=>"010110110",
  55114=>"011100100",
  55115=>"111101110",
  55116=>"010011110",
  55117=>"100101100",
  55118=>"000010100",
  55119=>"100101101",
  55120=>"111011010",
  55121=>"011011010",
  55122=>"111100100",
  55123=>"101010000",
  55124=>"111011111",
  55125=>"001110111",
  55126=>"000100111",
  55127=>"011010111",
  55128=>"111111011",
  55129=>"100011101",
  55130=>"001101101",
  55131=>"100001101",
  55132=>"110101110",
  55133=>"001010100",
  55134=>"011111110",
  55135=>"100001101",
  55136=>"010110110",
  55137=>"111011010",
  55138=>"001000110",
  55139=>"010000100",
  55140=>"000111011",
  55141=>"000011010",
  55142=>"100011110",
  55143=>"000110100",
  55144=>"110100000",
  55145=>"111000001",
  55146=>"000011100",
  55147=>"010011010",
  55148=>"011011000",
  55149=>"011010101",
  55150=>"111100101",
  55151=>"010011011",
  55152=>"110101101",
  55153=>"101101111",
  55154=>"000110110",
  55155=>"110110111",
  55156=>"000001100",
  55157=>"101100100",
  55158=>"100000011",
  55159=>"101010011",
  55160=>"110000001",
  55161=>"011011110",
  55162=>"001001001",
  55163=>"000000011",
  55164=>"001010100",
  55165=>"110101110",
  55166=>"111000100",
  55167=>"111100101",
  55168=>"010111011",
  55169=>"000010100",
  55170=>"010010100",
  55171=>"010010000",
  55172=>"111111111",
  55173=>"001010000",
  55174=>"010111000",
  55175=>"001010001",
  55176=>"000011101",
  55177=>"101111101",
  55178=>"000000000",
  55179=>"100101000",
  55180=>"001011010",
  55181=>"100110001",
  55182=>"011001100",
  55183=>"111010100",
  55184=>"000101011",
  55185=>"001010001",
  55186=>"100011101",
  55187=>"001011111",
  55188=>"100011110",
  55189=>"011011001",
  55190=>"011100001",
  55191=>"001011010",
  55192=>"100110110",
  55193=>"010010000",
  55194=>"001001110",
  55195=>"100000101",
  55196=>"000000100",
  55197=>"010001001",
  55198=>"100011101",
  55199=>"110111000",
  55200=>"111110000",
  55201=>"111001111",
  55202=>"001001111",
  55203=>"101011101",
  55204=>"010100110",
  55205=>"101111110",
  55206=>"011000111",
  55207=>"000011010",
  55208=>"001000010",
  55209=>"011010010",
  55210=>"011110010",
  55211=>"011010000",
  55212=>"000101001",
  55213=>"101111111",
  55214=>"011010100",
  55215=>"100111101",
  55216=>"000010110",
  55217=>"001000000",
  55218=>"110111000",
  55219=>"010101101",
  55220=>"101100010",
  55221=>"111011001",
  55222=>"011011111",
  55223=>"110100101",
  55224=>"011101000",
  55225=>"000100001",
  55226=>"001110111",
  55227=>"001110000",
  55228=>"101111010",
  55229=>"101001111",
  55230=>"011110010",
  55231=>"010000101",
  55232=>"100110111",
  55233=>"010110101",
  55234=>"010000100",
  55235=>"100010110",
  55236=>"001100011",
  55237=>"011011111",
  55238=>"101011011",
  55239=>"001000000",
  55240=>"110001000",
  55241=>"000000010",
  55242=>"001100111",
  55243=>"111000100",
  55244=>"111111111",
  55245=>"001101101",
  55246=>"110111111",
  55247=>"010010001",
  55248=>"011101101",
  55249=>"001100100",
  55250=>"100101010",
  55251=>"011111101",
  55252=>"101011010",
  55253=>"111001011",
  55254=>"000110001",
  55255=>"010001000",
  55256=>"101000001",
  55257=>"001111000",
  55258=>"010011011",
  55259=>"100010010",
  55260=>"001000101",
  55261=>"001111010",
  55262=>"110110100",
  55263=>"001110011",
  55264=>"011001010",
  55265=>"101001011",
  55266=>"111111101",
  55267=>"000110110",
  55268=>"001011011",
  55269=>"101000101",
  55270=>"101010101",
  55271=>"001011101",
  55272=>"101111100",
  55273=>"100001000",
  55274=>"011100101",
  55275=>"101011111",
  55276=>"000110010",
  55277=>"011001011",
  55278=>"011001111",
  55279=>"110000101",
  55280=>"101001111",
  55281=>"111001101",
  55282=>"101011000",
  55283=>"000001100",
  55284=>"100011110",
  55285=>"000010100",
  55286=>"101011111",
  55287=>"010101110",
  55288=>"011100001",
  55289=>"100110100",
  55290=>"101011100",
  55291=>"010000110",
  55292=>"110101101",
  55293=>"011010001",
  55294=>"010101101",
  55295=>"101010000",
  55296=>"100000110",
  55297=>"000100111",
  55298=>"111010111",
  55299=>"111111000",
  55300=>"100000101",
  55301=>"100010011",
  55302=>"110000001",
  55303=>"011010110",
  55304=>"100000101",
  55305=>"111010111",
  55306=>"111010001",
  55307=>"001011101",
  55308=>"100100101",
  55309=>"001111101",
  55310=>"110100010",
  55311=>"011111001",
  55312=>"010101110",
  55313=>"001001001",
  55314=>"001010101",
  55315=>"000010100",
  55316=>"000111111",
  55317=>"110111000",
  55318=>"001010111",
  55319=>"100111110",
  55320=>"111101101",
  55321=>"011101010",
  55322=>"001010010",
  55323=>"001100001",
  55324=>"100001000",
  55325=>"101011010",
  55326=>"001110111",
  55327=>"000100001",
  55328=>"111110011",
  55329=>"001011001",
  55330=>"110000101",
  55331=>"100111111",
  55332=>"000000011",
  55333=>"100000100",
  55334=>"000100110",
  55335=>"100010101",
  55336=>"001001010",
  55337=>"111101011",
  55338=>"111011010",
  55339=>"100110011",
  55340=>"000010100",
  55341=>"000101011",
  55342=>"110001111",
  55343=>"100100101",
  55344=>"000011000",
  55345=>"011111100",
  55346=>"101001010",
  55347=>"011011111",
  55348=>"000000011",
  55349=>"010000001",
  55350=>"011010100",
  55351=>"101110000",
  55352=>"010001110",
  55353=>"100110000",
  55354=>"110100100",
  55355=>"100010000",
  55356=>"011010101",
  55357=>"000011010",
  55358=>"100100001",
  55359=>"000111010",
  55360=>"010000000",
  55361=>"011110110",
  55362=>"111101111",
  55363=>"101010100",
  55364=>"111001000",
  55365=>"001001111",
  55366=>"000001111",
  55367=>"000100111",
  55368=>"111110000",
  55369=>"101111010",
  55370=>"100111100",
  55371=>"111101100",
  55372=>"110110100",
  55373=>"101100011",
  55374=>"111011100",
  55375=>"100001011",
  55376=>"111101001",
  55377=>"000010000",
  55378=>"000001100",
  55379=>"010101100",
  55380=>"110110101",
  55381=>"010000111",
  55382=>"101100111",
  55383=>"111101001",
  55384=>"011110100",
  55385=>"000100000",
  55386=>"110011010",
  55387=>"000011011",
  55388=>"111010010",
  55389=>"100110101",
  55390=>"100011001",
  55391=>"001000010",
  55392=>"001010110",
  55393=>"110001111",
  55394=>"001010111",
  55395=>"010001000",
  55396=>"000010111",
  55397=>"100010001",
  55398=>"001001011",
  55399=>"001111101",
  55400=>"110111101",
  55401=>"001010101",
  55402=>"100111010",
  55403=>"010110010",
  55404=>"110010010",
  55405=>"010011101",
  55406=>"010111000",
  55407=>"000101111",
  55408=>"011111000",
  55409=>"010101111",
  55410=>"001000100",
  55411=>"001101100",
  55412=>"000000110",
  55413=>"111001110",
  55414=>"111101110",
  55415=>"000010110",
  55416=>"000000100",
  55417=>"000000010",
  55418=>"101000010",
  55419=>"111100011",
  55420=>"011111101",
  55421=>"101100101",
  55422=>"001010111",
  55423=>"000000010",
  55424=>"011011111",
  55425=>"010100000",
  55426=>"100010101",
  55427=>"101011111",
  55428=>"011011010",
  55429=>"110111000",
  55430=>"110111111",
  55431=>"000001101",
  55432=>"010000001",
  55433=>"011010101",
  55434=>"111111010",
  55435=>"111110101",
  55436=>"110111010",
  55437=>"100111010",
  55438=>"110111001",
  55439=>"100111111",
  55440=>"010011100",
  55441=>"000110000",
  55442=>"000110100",
  55443=>"101010100",
  55444=>"010100110",
  55445=>"011011111",
  55446=>"010101000",
  55447=>"110100010",
  55448=>"111111111",
  55449=>"101000111",
  55450=>"011011111",
  55451=>"110100101",
  55452=>"111110010",
  55453=>"110110001",
  55454=>"110010111",
  55455=>"101101010",
  55456=>"010011101",
  55457=>"111101011",
  55458=>"000101011",
  55459=>"011001110",
  55460=>"001100101",
  55461=>"100001101",
  55462=>"110010010",
  55463=>"110111111",
  55464=>"100000100",
  55465=>"110010000",
  55466=>"001100000",
  55467=>"111110111",
  55468=>"011111001",
  55469=>"000010010",
  55470=>"111110101",
  55471=>"001110110",
  55472=>"101100111",
  55473=>"001011110",
  55474=>"001001100",
  55475=>"000000101",
  55476=>"100100110",
  55477=>"010100001",
  55478=>"000001001",
  55479=>"100000010",
  55480=>"101000010",
  55481=>"001001101",
  55482=>"000100000",
  55483=>"110101111",
  55484=>"111100101",
  55485=>"101001011",
  55486=>"101010001",
  55487=>"111100010",
  55488=>"111011100",
  55489=>"110100011",
  55490=>"111110000",
  55491=>"010101111",
  55492=>"110111100",
  55493=>"011001101",
  55494=>"100000100",
  55495=>"111101101",
  55496=>"000001100",
  55497=>"000000111",
  55498=>"000101111",
  55499=>"101011101",
  55500=>"001100101",
  55501=>"010101101",
  55502=>"100001100",
  55503=>"001011111",
  55504=>"010110011",
  55505=>"110100011",
  55506=>"101000000",
  55507=>"100110011",
  55508=>"010111100",
  55509=>"000000011",
  55510=>"111011111",
  55511=>"110111101",
  55512=>"100110001",
  55513=>"110101000",
  55514=>"011111100",
  55515=>"101110111",
  55516=>"101000010",
  55517=>"000100101",
  55518=>"111101101",
  55519=>"110010100",
  55520=>"111011110",
  55521=>"010001011",
  55522=>"000111011",
  55523=>"000000110",
  55524=>"100111111",
  55525=>"101110111",
  55526=>"011011100",
  55527=>"001011001",
  55528=>"000001011",
  55529=>"001111110",
  55530=>"010110000",
  55531=>"010111011",
  55532=>"011000100",
  55533=>"010001110",
  55534=>"101101011",
  55535=>"011001101",
  55536=>"000000011",
  55537=>"101001100",
  55538=>"111001100",
  55539=>"010011101",
  55540=>"000101111",
  55541=>"001000011",
  55542=>"111100001",
  55543=>"110111011",
  55544=>"111000001",
  55545=>"111000100",
  55546=>"110111101",
  55547=>"000100011",
  55548=>"001010101",
  55549=>"110110111",
  55550=>"100011100",
  55551=>"000111000",
  55552=>"111111101",
  55553=>"101110100",
  55554=>"101000011",
  55555=>"100110111",
  55556=>"101000001",
  55557=>"000111011",
  55558=>"001110100",
  55559=>"101111011",
  55560=>"010011000",
  55561=>"011011001",
  55562=>"011010101",
  55563=>"101001110",
  55564=>"001100011",
  55565=>"011101100",
  55566=>"100101111",
  55567=>"001010100",
  55568=>"010101111",
  55569=>"010001011",
  55570=>"000011000",
  55571=>"101011101",
  55572=>"011000000",
  55573=>"000101001",
  55574=>"110110010",
  55575=>"000011111",
  55576=>"110010000",
  55577=>"111000100",
  55578=>"110001000",
  55579=>"100101100",
  55580=>"111001100",
  55581=>"000111101",
  55582=>"010110101",
  55583=>"111111010",
  55584=>"011011101",
  55585=>"011000111",
  55586=>"101001010",
  55587=>"100111101",
  55588=>"010000010",
  55589=>"001000000",
  55590=>"110101100",
  55591=>"111000111",
  55592=>"110101001",
  55593=>"110101111",
  55594=>"010100010",
  55595=>"100110000",
  55596=>"101010010",
  55597=>"010001000",
  55598=>"010100000",
  55599=>"000011101",
  55600=>"011010011",
  55601=>"001100101",
  55602=>"001001101",
  55603=>"101101011",
  55604=>"100001111",
  55605=>"011011000",
  55606=>"101111110",
  55607=>"000110001",
  55608=>"100000010",
  55609=>"010010100",
  55610=>"110010000",
  55611=>"000110000",
  55612=>"000000111",
  55613=>"010111111",
  55614=>"101110000",
  55615=>"111111111",
  55616=>"110110101",
  55617=>"111011000",
  55618=>"000111000",
  55619=>"111010101",
  55620=>"000000111",
  55621=>"110111001",
  55622=>"000101010",
  55623=>"000011000",
  55624=>"100010111",
  55625=>"001000000",
  55626=>"000011100",
  55627=>"111000010",
  55628=>"010000001",
  55629=>"101000111",
  55630=>"000111101",
  55631=>"101010010",
  55632=>"110001001",
  55633=>"011000111",
  55634=>"000100000",
  55635=>"010110000",
  55636=>"101111111",
  55637=>"101111111",
  55638=>"100010011",
  55639=>"011010001",
  55640=>"111001011",
  55641=>"100100000",
  55642=>"111111100",
  55643=>"111110001",
  55644=>"001100000",
  55645=>"011100011",
  55646=>"000001110",
  55647=>"111010010",
  55648=>"011100010",
  55649=>"000000010",
  55650=>"011101101",
  55651=>"110111000",
  55652=>"101110100",
  55653=>"100111111",
  55654=>"000111010",
  55655=>"001011011",
  55656=>"010100111",
  55657=>"000100100",
  55658=>"001101011",
  55659=>"111001011",
  55660=>"010101011",
  55661=>"010001000",
  55662=>"001111110",
  55663=>"001000001",
  55664=>"101011010",
  55665=>"110111110",
  55666=>"110110101",
  55667=>"011100101",
  55668=>"001011001",
  55669=>"001010100",
  55670=>"000100100",
  55671=>"110100011",
  55672=>"101000110",
  55673=>"110110011",
  55674=>"001001001",
  55675=>"110101110",
  55676=>"011001100",
  55677=>"001100110",
  55678=>"011000111",
  55679=>"010010000",
  55680=>"111111110",
  55681=>"101101110",
  55682=>"000101011",
  55683=>"010101000",
  55684=>"111010111",
  55685=>"100111000",
  55686=>"011100111",
  55687=>"110010011",
  55688=>"011100011",
  55689=>"111100000",
  55690=>"110100100",
  55691=>"101101000",
  55692=>"001110001",
  55693=>"010101110",
  55694=>"110001001",
  55695=>"101010001",
  55696=>"000001110",
  55697=>"001101100",
  55698=>"110001010",
  55699=>"011001000",
  55700=>"101110100",
  55701=>"001110111",
  55702=>"000101111",
  55703=>"110110011",
  55704=>"000110101",
  55705=>"101011110",
  55706=>"100100111",
  55707=>"000011001",
  55708=>"110111001",
  55709=>"010111101",
  55710=>"100000000",
  55711=>"110100011",
  55712=>"001101110",
  55713=>"101011111",
  55714=>"010010101",
  55715=>"111010001",
  55716=>"010100000",
  55717=>"111000001",
  55718=>"100000110",
  55719=>"001010000",
  55720=>"111001001",
  55721=>"101111100",
  55722=>"001010010",
  55723=>"101101101",
  55724=>"000000110",
  55725=>"111110101",
  55726=>"001110100",
  55727=>"010100000",
  55728=>"101011010",
  55729=>"111111110",
  55730=>"110110011",
  55731=>"101100110",
  55732=>"010001110",
  55733=>"001011111",
  55734=>"001101001",
  55735=>"110010011",
  55736=>"111001011",
  55737=>"001111000",
  55738=>"100001110",
  55739=>"110000000",
  55740=>"110110011",
  55741=>"011111101",
  55742=>"100010001",
  55743=>"111000000",
  55744=>"111101011",
  55745=>"111110010",
  55746=>"111111110",
  55747=>"101001011",
  55748=>"100000011",
  55749=>"111111101",
  55750=>"110010011",
  55751=>"100010101",
  55752=>"111101011",
  55753=>"111011000",
  55754=>"100111101",
  55755=>"011111010",
  55756=>"101011010",
  55757=>"100000110",
  55758=>"111110000",
  55759=>"111100111",
  55760=>"111010000",
  55761=>"110011000",
  55762=>"100100100",
  55763=>"001011111",
  55764=>"101001000",
  55765=>"110001101",
  55766=>"111011111",
  55767=>"110110011",
  55768=>"001000100",
  55769=>"101010011",
  55770=>"011100001",
  55771=>"011111100",
  55772=>"110000100",
  55773=>"101101000",
  55774=>"101110110",
  55775=>"000010100",
  55776=>"011000011",
  55777=>"100001110",
  55778=>"000010000",
  55779=>"010101100",
  55780=>"011010010",
  55781=>"110100111",
  55782=>"101011111",
  55783=>"100001010",
  55784=>"110110100",
  55785=>"011111101",
  55786=>"000010110",
  55787=>"011001110",
  55788=>"101001100",
  55789=>"101011001",
  55790=>"111100010",
  55791=>"000001100",
  55792=>"100011111",
  55793=>"001111111",
  55794=>"000011111",
  55795=>"110000000",
  55796=>"011101101",
  55797=>"000101010",
  55798=>"101100101",
  55799=>"011011011",
  55800=>"010101000",
  55801=>"000010000",
  55802=>"000100100",
  55803=>"101001101",
  55804=>"001111101",
  55805=>"100011110",
  55806=>"111110101",
  55807=>"101010101",
  55808=>"101101000",
  55809=>"001010110",
  55810=>"111111011",
  55811=>"000100101",
  55812=>"010010000",
  55813=>"010010100",
  55814=>"000001001",
  55815=>"010101101",
  55816=>"000011010",
  55817=>"011111000",
  55818=>"000110100",
  55819=>"001000001",
  55820=>"011000100",
  55821=>"100101010",
  55822=>"110100110",
  55823=>"111101001",
  55824=>"001100110",
  55825=>"000111011",
  55826=>"100000011",
  55827=>"101110000",
  55828=>"010101110",
  55829=>"111110111",
  55830=>"010010111",
  55831=>"101001001",
  55832=>"100010011",
  55833=>"001001110",
  55834=>"100100101",
  55835=>"010010110",
  55836=>"111101100",
  55837=>"011010010",
  55838=>"011100101",
  55839=>"010011110",
  55840=>"100110100",
  55841=>"011000110",
  55842=>"011100100",
  55843=>"100111010",
  55844=>"000000010",
  55845=>"111111111",
  55846=>"001001011",
  55847=>"100010111",
  55848=>"011100000",
  55849=>"011100100",
  55850=>"110010010",
  55851=>"001100011",
  55852=>"110000110",
  55853=>"011000001",
  55854=>"010111011",
  55855=>"110110110",
  55856=>"010011111",
  55857=>"001110000",
  55858=>"111111110",
  55859=>"111010100",
  55860=>"000000101",
  55861=>"000001100",
  55862=>"000001011",
  55863=>"101101111",
  55864=>"001100110",
  55865=>"100111111",
  55866=>"101001110",
  55867=>"001010010",
  55868=>"001001000",
  55869=>"011000010",
  55870=>"111000011",
  55871=>"001011010",
  55872=>"010000001",
  55873=>"001100001",
  55874=>"100011100",
  55875=>"110110100",
  55876=>"011111001",
  55877=>"110000100",
  55878=>"000001000",
  55879=>"101011111",
  55880=>"110110110",
  55881=>"001011100",
  55882=>"111111110",
  55883=>"111001000",
  55884=>"111111101",
  55885=>"011100001",
  55886=>"011000011",
  55887=>"101011111",
  55888=>"101011001",
  55889=>"101101111",
  55890=>"100000100",
  55891=>"101010100",
  55892=>"001001100",
  55893=>"000000000",
  55894=>"001011001",
  55895=>"010001001",
  55896=>"000001001",
  55897=>"010110000",
  55898=>"000000011",
  55899=>"111001000",
  55900=>"010100101",
  55901=>"011000100",
  55902=>"101011001",
  55903=>"010010011",
  55904=>"000001010",
  55905=>"000000010",
  55906=>"010110000",
  55907=>"001010000",
  55908=>"010001000",
  55909=>"000100000",
  55910=>"111101101",
  55911=>"100000001",
  55912=>"000000101",
  55913=>"110000000",
  55914=>"111110101",
  55915=>"010111000",
  55916=>"110011110",
  55917=>"100010010",
  55918=>"011111111",
  55919=>"000010100",
  55920=>"001001110",
  55921=>"111010000",
  55922=>"101000111",
  55923=>"100111001",
  55924=>"000111100",
  55925=>"001001110",
  55926=>"111100010",
  55927=>"101101111",
  55928=>"011110100",
  55929=>"001010010",
  55930=>"001111000",
  55931=>"101001100",
  55932=>"100011011",
  55933=>"110001011",
  55934=>"100110111",
  55935=>"011110011",
  55936=>"000111000",
  55937=>"100100111",
  55938=>"101111010",
  55939=>"000100110",
  55940=>"010111001",
  55941=>"000100111",
  55942=>"010001001",
  55943=>"110110100",
  55944=>"110010101",
  55945=>"101111101",
  55946=>"111001110",
  55947=>"110101011",
  55948=>"111110011",
  55949=>"110101011",
  55950=>"011111111",
  55951=>"111011010",
  55952=>"010011000",
  55953=>"110111000",
  55954=>"101100010",
  55955=>"111001011",
  55956=>"011110110",
  55957=>"011011001",
  55958=>"111101111",
  55959=>"101001011",
  55960=>"101111000",
  55961=>"000001101",
  55962=>"011011010",
  55963=>"101010100",
  55964=>"110101101",
  55965=>"011001011",
  55966=>"111111100",
  55967=>"100110010",
  55968=>"100110101",
  55969=>"011100001",
  55970=>"110110000",
  55971=>"011110000",
  55972=>"110001110",
  55973=>"000111111",
  55974=>"011001010",
  55975=>"011000110",
  55976=>"111111100",
  55977=>"001101111",
  55978=>"111100001",
  55979=>"001100001",
  55980=>"010101100",
  55981=>"000010010",
  55982=>"111001000",
  55983=>"000011111",
  55984=>"010000111",
  55985=>"010100010",
  55986=>"100101111",
  55987=>"100100110",
  55988=>"101100011",
  55989=>"011011010",
  55990=>"011111000",
  55991=>"010111011",
  55992=>"110010000",
  55993=>"111000101",
  55994=>"111101100",
  55995=>"011101011",
  55996=>"111110011",
  55997=>"110000000",
  55998=>"011100000",
  55999=>"000111110",
  56000=>"000111001",
  56001=>"011011100",
  56002=>"110011010",
  56003=>"010110011",
  56004=>"110101100",
  56005=>"001100011",
  56006=>"111000011",
  56007=>"110010000",
  56008=>"001111001",
  56009=>"000000000",
  56010=>"010001001",
  56011=>"100100011",
  56012=>"000011001",
  56013=>"000111111",
  56014=>"110010101",
  56015=>"110111100",
  56016=>"000010000",
  56017=>"011111110",
  56018=>"001100010",
  56019=>"110101001",
  56020=>"000110000",
  56021=>"100011101",
  56022=>"000011111",
  56023=>"010110000",
  56024=>"001000111",
  56025=>"001100011",
  56026=>"001011110",
  56027=>"101001110",
  56028=>"111110111",
  56029=>"000111011",
  56030=>"010001010",
  56031=>"100101110",
  56032=>"101111100",
  56033=>"100111100",
  56034=>"001101110",
  56035=>"111010101",
  56036=>"000101100",
  56037=>"000101111",
  56038=>"011100100",
  56039=>"110011101",
  56040=>"000110110",
  56041=>"110001110",
  56042=>"110100011",
  56043=>"111101010",
  56044=>"011011110",
  56045=>"000101001",
  56046=>"001001001",
  56047=>"101001010",
  56048=>"111000010",
  56049=>"010101100",
  56050=>"011101110",
  56051=>"110111101",
  56052=>"001101001",
  56053=>"000001100",
  56054=>"111101001",
  56055=>"101100111",
  56056=>"000000010",
  56057=>"111101100",
  56058=>"100110000",
  56059=>"101001001",
  56060=>"110101100",
  56061=>"000001010",
  56062=>"100010100",
  56063=>"001101000",
  56064=>"011000100",
  56065=>"111111101",
  56066=>"111000000",
  56067=>"100110100",
  56068=>"110100011",
  56069=>"011001111",
  56070=>"010011110",
  56071=>"100110011",
  56072=>"000010011",
  56073=>"110110100",
  56074=>"101110011",
  56075=>"100001110",
  56076=>"110001001",
  56077=>"100110110",
  56078=>"001011010",
  56079=>"000001010",
  56080=>"011110111",
  56081=>"100111010",
  56082=>"101100110",
  56083=>"110000110",
  56084=>"111110111",
  56085=>"101011110",
  56086=>"111111111",
  56087=>"001000101",
  56088=>"100101100",
  56089=>"110010110",
  56090=>"001010001",
  56091=>"001001010",
  56092=>"110101110",
  56093=>"100110100",
  56094=>"010110011",
  56095=>"100010011",
  56096=>"001111111",
  56097=>"100111001",
  56098=>"110101011",
  56099=>"000100001",
  56100=>"111010011",
  56101=>"011001000",
  56102=>"001000001",
  56103=>"101111010",
  56104=>"101011000",
  56105=>"101110100",
  56106=>"000001110",
  56107=>"001110011",
  56108=>"000100110",
  56109=>"010001101",
  56110=>"000101111",
  56111=>"001110000",
  56112=>"000001101",
  56113=>"000010111",
  56114=>"101001001",
  56115=>"001010000",
  56116=>"110001000",
  56117=>"110111000",
  56118=>"000001001",
  56119=>"011001000",
  56120=>"110110101",
  56121=>"001010100",
  56122=>"111000010",
  56123=>"000001011",
  56124=>"101000010",
  56125=>"000101010",
  56126=>"010010000",
  56127=>"001010101",
  56128=>"011000101",
  56129=>"000100110",
  56130=>"000111111",
  56131=>"110101000",
  56132=>"110001100",
  56133=>"000000000",
  56134=>"011111101",
  56135=>"010110101",
  56136=>"001100101",
  56137=>"110111101",
  56138=>"100001101",
  56139=>"111101000",
  56140=>"100110111",
  56141=>"010010001",
  56142=>"011111101",
  56143=>"110110100",
  56144=>"110100101",
  56145=>"111011010",
  56146=>"110000111",
  56147=>"111001110",
  56148=>"111110000",
  56149=>"101101010",
  56150=>"001000001",
  56151=>"101010101",
  56152=>"001100000",
  56153=>"101110100",
  56154=>"001100001",
  56155=>"100010001",
  56156=>"101101101",
  56157=>"001101100",
  56158=>"000001110",
  56159=>"001000000",
  56160=>"001100110",
  56161=>"100111000",
  56162=>"001101010",
  56163=>"001100101",
  56164=>"111011011",
  56165=>"010000011",
  56166=>"110000101",
  56167=>"001111011",
  56168=>"101111111",
  56169=>"011110111",
  56170=>"010110001",
  56171=>"101000011",
  56172=>"110000100",
  56173=>"011000000",
  56174=>"000001111",
  56175=>"011010000",
  56176=>"000101010",
  56177=>"111101100",
  56178=>"001001110",
  56179=>"011101000",
  56180=>"001111101",
  56181=>"001110110",
  56182=>"010010100",
  56183=>"100111111",
  56184=>"001110101",
  56185=>"011110100",
  56186=>"101111111",
  56187=>"100000001",
  56188=>"010001100",
  56189=>"011011101",
  56190=>"101001101",
  56191=>"101110111",
  56192=>"111001101",
  56193=>"101100110",
  56194=>"001100111",
  56195=>"111101001",
  56196=>"000101111",
  56197=>"000010110",
  56198=>"101100111",
  56199=>"100000001",
  56200=>"010011001",
  56201=>"100000010",
  56202=>"011001010",
  56203=>"100011111",
  56204=>"101000010",
  56205=>"110001100",
  56206=>"001100111",
  56207=>"100111101",
  56208=>"000101111",
  56209=>"100100111",
  56210=>"110011101",
  56211=>"001010000",
  56212=>"001011011",
  56213=>"101001010",
  56214=>"011101001",
  56215=>"100100110",
  56216=>"001000100",
  56217=>"110111101",
  56218=>"111000110",
  56219=>"111000001",
  56220=>"101111111",
  56221=>"101000100",
  56222=>"110011001",
  56223=>"111010011",
  56224=>"110101101",
  56225=>"100000001",
  56226=>"010101100",
  56227=>"100111111",
  56228=>"110000000",
  56229=>"011000000",
  56230=>"101001011",
  56231=>"110111100",
  56232=>"100000101",
  56233=>"111111001",
  56234=>"111000000",
  56235=>"110110001",
  56236=>"010110111",
  56237=>"000011100",
  56238=>"101000000",
  56239=>"000110110",
  56240=>"000110010",
  56241=>"010010111",
  56242=>"001110000",
  56243=>"011101100",
  56244=>"101100110",
  56245=>"010100011",
  56246=>"101101111",
  56247=>"001110010",
  56248=>"100101101",
  56249=>"000100000",
  56250=>"011101111",
  56251=>"100011000",
  56252=>"000101011",
  56253=>"000011000",
  56254=>"110100111",
  56255=>"000010111",
  56256=>"011000011",
  56257=>"010001001",
  56258=>"110001111",
  56259=>"000110110",
  56260=>"101000000",
  56261=>"000010110",
  56262=>"000011010",
  56263=>"111110110",
  56264=>"000010010",
  56265=>"001110111",
  56266=>"000010011",
  56267=>"111111110",
  56268=>"000100000",
  56269=>"111100110",
  56270=>"011100011",
  56271=>"011101110",
  56272=>"000000010",
  56273=>"001001001",
  56274=>"111111001",
  56275=>"001000010",
  56276=>"011100010",
  56277=>"111010010",
  56278=>"101101010",
  56279=>"100000001",
  56280=>"111111011",
  56281=>"011111000",
  56282=>"110010101",
  56283=>"110000010",
  56284=>"110001000",
  56285=>"001011011",
  56286=>"101110111",
  56287=>"100001101",
  56288=>"110110111",
  56289=>"000001100",
  56290=>"000001011",
  56291=>"000011100",
  56292=>"100001100",
  56293=>"001011001",
  56294=>"000111011",
  56295=>"110000011",
  56296=>"000101001",
  56297=>"101110010",
  56298=>"111110001",
  56299=>"010011111",
  56300=>"111110100",
  56301=>"011001100",
  56302=>"000110100",
  56303=>"101001010",
  56304=>"001101010",
  56305=>"011110001",
  56306=>"010011110",
  56307=>"000001001",
  56308=>"010110101",
  56309=>"100101100",
  56310=>"001101111",
  56311=>"101101000",
  56312=>"001111000",
  56313=>"001000110",
  56314=>"010011001",
  56315=>"001101011",
  56316=>"010110001",
  56317=>"000100010",
  56318=>"011110001",
  56319=>"010000010",
  56320=>"101000100",
  56321=>"010011000",
  56322=>"011110010",
  56323=>"100110110",
  56324=>"111010000",
  56325=>"000100001",
  56326=>"111101101",
  56327=>"010000101",
  56328=>"010010001",
  56329=>"010011000",
  56330=>"000001110",
  56331=>"010110101",
  56332=>"000011000",
  56333=>"000000110",
  56334=>"111110010",
  56335=>"111010001",
  56336=>"001110100",
  56337=>"011000000",
  56338=>"011110010",
  56339=>"000001000",
  56340=>"001100111",
  56341=>"011000001",
  56342=>"101100110",
  56343=>"001111110",
  56344=>"001101011",
  56345=>"101110100",
  56346=>"000000000",
  56347=>"001000001",
  56348=>"111101100",
  56349=>"010010010",
  56350=>"101111110",
  56351=>"100101111",
  56352=>"010010101",
  56353=>"010011100",
  56354=>"000111101",
  56355=>"111011101",
  56356=>"101101000",
  56357=>"011111001",
  56358=>"100110001",
  56359=>"110000011",
  56360=>"001001100",
  56361=>"101001101",
  56362=>"011011001",
  56363=>"101100101",
  56364=>"101011111",
  56365=>"000000010",
  56366=>"000001010",
  56367=>"010100000",
  56368=>"010101011",
  56369=>"111101000",
  56370=>"010001111",
  56371=>"001001000",
  56372=>"111101011",
  56373=>"000011010",
  56374=>"111100101",
  56375=>"001110100",
  56376=>"010010101",
  56377=>"101101110",
  56378=>"101010000",
  56379=>"111011000",
  56380=>"100110010",
  56381=>"000100110",
  56382=>"000000000",
  56383=>"010111111",
  56384=>"000001110",
  56385=>"000001110",
  56386=>"111101010",
  56387=>"011011110",
  56388=>"101110011",
  56389=>"101001101",
  56390=>"011101100",
  56391=>"101110011",
  56392=>"110011110",
  56393=>"000011010",
  56394=>"100010100",
  56395=>"011101011",
  56396=>"011100111",
  56397=>"111111011",
  56398=>"010110111",
  56399=>"000001100",
  56400=>"111111100",
  56401=>"000010010",
  56402=>"101010111",
  56403=>"011111010",
  56404=>"000011110",
  56405=>"101110101",
  56406=>"111011010",
  56407=>"011010101",
  56408=>"001111101",
  56409=>"011010100",
  56410=>"101101111",
  56411=>"100010001",
  56412=>"000100111",
  56413=>"010000101",
  56414=>"011000011",
  56415=>"000000001",
  56416=>"001001011",
  56417=>"111111111",
  56418=>"101111000",
  56419=>"100110101",
  56420=>"000101101",
  56421=>"001011111",
  56422=>"100111111",
  56423=>"001100011",
  56424=>"010110000",
  56425=>"010110001",
  56426=>"101001001",
  56427=>"111110110",
  56428=>"000000100",
  56429=>"101101010",
  56430=>"111000000",
  56431=>"011111000",
  56432=>"100110010",
  56433=>"000110000",
  56434=>"000100100",
  56435=>"001000111",
  56436=>"001101111",
  56437=>"010101001",
  56438=>"110001011",
  56439=>"001001111",
  56440=>"111010011",
  56441=>"101111101",
  56442=>"000001111",
  56443=>"001001101",
  56444=>"010111100",
  56445=>"000010011",
  56446=>"011010000",
  56447=>"101000111",
  56448=>"101111110",
  56449=>"001000110",
  56450=>"111011100",
  56451=>"100110100",
  56452=>"001100111",
  56453=>"000000000",
  56454=>"011011111",
  56455=>"001000011",
  56456=>"110001100",
  56457=>"010010100",
  56458=>"101000010",
  56459=>"000011101",
  56460=>"010001111",
  56461=>"101100110",
  56462=>"111111111",
  56463=>"011001001",
  56464=>"000000010",
  56465=>"110011111",
  56466=>"001001001",
  56467=>"111111101",
  56468=>"011110011",
  56469=>"011100100",
  56470=>"101000101",
  56471=>"000011111",
  56472=>"010011011",
  56473=>"110000011",
  56474=>"001010010",
  56475=>"011101001",
  56476=>"111100110",
  56477=>"011101101",
  56478=>"000110101",
  56479=>"110101010",
  56480=>"010011000",
  56481=>"010111110",
  56482=>"001010001",
  56483=>"001110100",
  56484=>"110110011",
  56485=>"100111111",
  56486=>"111100000",
  56487=>"111110000",
  56488=>"011010001",
  56489=>"010110111",
  56490=>"001001011",
  56491=>"111000000",
  56492=>"010101010",
  56493=>"010011101",
  56494=>"001111001",
  56495=>"100110111",
  56496=>"100001000",
  56497=>"000111111",
  56498=>"111000111",
  56499=>"100000000",
  56500=>"011011110",
  56501=>"111000000",
  56502=>"010011110",
  56503=>"101000010",
  56504=>"111000110",
  56505=>"010111100",
  56506=>"110110000",
  56507=>"000010111",
  56508=>"110111000",
  56509=>"000010110",
  56510=>"100010000",
  56511=>"100001000",
  56512=>"010010110",
  56513=>"001010000",
  56514=>"100001010",
  56515=>"000110001",
  56516=>"001101001",
  56517=>"111000111",
  56518=>"000000100",
  56519=>"100110001",
  56520=>"110011011",
  56521=>"000100101",
  56522=>"000110101",
  56523=>"000100111",
  56524=>"110001111",
  56525=>"110111101",
  56526=>"010001011",
  56527=>"010001111",
  56528=>"001101010",
  56529=>"110110110",
  56530=>"000111100",
  56531=>"101101100",
  56532=>"111001010",
  56533=>"010000110",
  56534=>"111110100",
  56535=>"001000001",
  56536=>"010110000",
  56537=>"110100101",
  56538=>"110001110",
  56539=>"001110000",
  56540=>"111100001",
  56541=>"010010110",
  56542=>"000000000",
  56543=>"111001111",
  56544=>"000000001",
  56545=>"010100111",
  56546=>"110010011",
  56547=>"101110111",
  56548=>"100001000",
  56549=>"100110000",
  56550=>"001110111",
  56551=>"000100111",
  56552=>"100100000",
  56553=>"000001000",
  56554=>"001000001",
  56555=>"101111110",
  56556=>"100010010",
  56557=>"101010001",
  56558=>"010000110",
  56559=>"111100101",
  56560=>"111111010",
  56561=>"001000011",
  56562=>"101111100",
  56563=>"110011000",
  56564=>"110000101",
  56565=>"010000010",
  56566=>"000010100",
  56567=>"010110010",
  56568=>"011000110",
  56569=>"001100001",
  56570=>"110100111",
  56571=>"100000110",
  56572=>"010010101",
  56573=>"101111110",
  56574=>"000000111",
  56575=>"101000111",
  56576=>"010111100",
  56577=>"000110100",
  56578=>"011100011",
  56579=>"010011100",
  56580=>"100010001",
  56581=>"101001001",
  56582=>"011000000",
  56583=>"011011101",
  56584=>"111100101",
  56585=>"001010110",
  56586=>"101101110",
  56587=>"010000010",
  56588=>"011110111",
  56589=>"011001000",
  56590=>"111000101",
  56591=>"100010110",
  56592=>"110110001",
  56593=>"001001010",
  56594=>"111100001",
  56595=>"001000101",
  56596=>"011110101",
  56597=>"111101000",
  56598=>"011001011",
  56599=>"011111101",
  56600=>"101110000",
  56601=>"001000110",
  56602=>"100101101",
  56603=>"010110001",
  56604=>"100010110",
  56605=>"010110110",
  56606=>"100000010",
  56607=>"100100001",
  56608=>"101011000",
  56609=>"000110000",
  56610=>"010010001",
  56611=>"011010011",
  56612=>"001101111",
  56613=>"110000011",
  56614=>"110101110",
  56615=>"111010001",
  56616=>"000100000",
  56617=>"010011000",
  56618=>"011111001",
  56619=>"100110101",
  56620=>"111110101",
  56621=>"000000001",
  56622=>"011100001",
  56623=>"010001101",
  56624=>"011000001",
  56625=>"011010111",
  56626=>"000111111",
  56627=>"111010010",
  56628=>"000100101",
  56629=>"001101001",
  56630=>"100010100",
  56631=>"101011010",
  56632=>"111111011",
  56633=>"011100010",
  56634=>"111100011",
  56635=>"001110000",
  56636=>"011100111",
  56637=>"101010001",
  56638=>"000001011",
  56639=>"110000110",
  56640=>"001000101",
  56641=>"011111101",
  56642=>"010101011",
  56643=>"001011010",
  56644=>"010100111",
  56645=>"001111001",
  56646=>"101100001",
  56647=>"111111011",
  56648=>"111010010",
  56649=>"010011110",
  56650=>"101011010",
  56651=>"100011001",
  56652=>"010100101",
  56653=>"110111101",
  56654=>"000101010",
  56655=>"111101111",
  56656=>"111111000",
  56657=>"110001100",
  56658=>"001001111",
  56659=>"111011000",
  56660=>"011001111",
  56661=>"111100000",
  56662=>"000011101",
  56663=>"111110000",
  56664=>"100011000",
  56665=>"111101000",
  56666=>"101010001",
  56667=>"111001011",
  56668=>"010000000",
  56669=>"000011111",
  56670=>"111000011",
  56671=>"010101110",
  56672=>"110000110",
  56673=>"111100101",
  56674=>"110011100",
  56675=>"001101110",
  56676=>"101111111",
  56677=>"110011001",
  56678=>"001000010",
  56679=>"101100110",
  56680=>"001000100",
  56681=>"110011001",
  56682=>"000101001",
  56683=>"011000010",
  56684=>"100100111",
  56685=>"000001110",
  56686=>"101010001",
  56687=>"101100000",
  56688=>"000011001",
  56689=>"001111100",
  56690=>"010001110",
  56691=>"000100100",
  56692=>"000010000",
  56693=>"101001110",
  56694=>"100000100",
  56695=>"111100100",
  56696=>"001100111",
  56697=>"110110110",
  56698=>"100011101",
  56699=>"010011010",
  56700=>"111001011",
  56701=>"010011000",
  56702=>"101100110",
  56703=>"011100110",
  56704=>"010010100",
  56705=>"100100101",
  56706=>"000011000",
  56707=>"101011101",
  56708=>"111000001",
  56709=>"101001010",
  56710=>"011100001",
  56711=>"010011100",
  56712=>"001111010",
  56713=>"000000000",
  56714=>"101001001",
  56715=>"001100001",
  56716=>"110110101",
  56717=>"010001011",
  56718=>"001111110",
  56719=>"110101100",
  56720=>"000100010",
  56721=>"101100001",
  56722=>"110110001",
  56723=>"101010111",
  56724=>"110111111",
  56725=>"101001111",
  56726=>"000101100",
  56727=>"011111101",
  56728=>"011111111",
  56729=>"101001001",
  56730=>"110111100",
  56731=>"000101100",
  56732=>"001011101",
  56733=>"001000010",
  56734=>"011110111",
  56735=>"001111010",
  56736=>"100101111",
  56737=>"001110100",
  56738=>"100001000",
  56739=>"001100001",
  56740=>"110101010",
  56741=>"111100110",
  56742=>"011001010",
  56743=>"101010100",
  56744=>"011101000",
  56745=>"111001110",
  56746=>"111111011",
  56747=>"010101010",
  56748=>"010100100",
  56749=>"001010011",
  56750=>"001101001",
  56751=>"001000110",
  56752=>"001101011",
  56753=>"110110011",
  56754=>"011100000",
  56755=>"101001111",
  56756=>"000010010",
  56757=>"100100000",
  56758=>"101011100",
  56759=>"011000001",
  56760=>"000011100",
  56761=>"111011011",
  56762=>"001000001",
  56763=>"010000000",
  56764=>"111110010",
  56765=>"001110000",
  56766=>"101110000",
  56767=>"000000011",
  56768=>"110011010",
  56769=>"100100111",
  56770=>"011000110",
  56771=>"110101010",
  56772=>"100010111",
  56773=>"111010001",
  56774=>"000000110",
  56775=>"010110010",
  56776=>"100111000",
  56777=>"001010100",
  56778=>"101011011",
  56779=>"100110101",
  56780=>"110001000",
  56781=>"001000010",
  56782=>"001111101",
  56783=>"000001011",
  56784=>"111101110",
  56785=>"011001011",
  56786=>"110100101",
  56787=>"100000110",
  56788=>"101111110",
  56789=>"011011111",
  56790=>"101010001",
  56791=>"100111110",
  56792=>"101111110",
  56793=>"001001011",
  56794=>"000010110",
  56795=>"001000011",
  56796=>"111000111",
  56797=>"100100110",
  56798=>"101100110",
  56799=>"110111010",
  56800=>"001000000",
  56801=>"110010110",
  56802=>"101101110",
  56803=>"100111110",
  56804=>"100000110",
  56805=>"101010111",
  56806=>"010101000",
  56807=>"100001111",
  56808=>"101111111",
  56809=>"110011100",
  56810=>"111001100",
  56811=>"011111000",
  56812=>"100110101",
  56813=>"100101000",
  56814=>"011011000",
  56815=>"111101001",
  56816=>"100010101",
  56817=>"111000110",
  56818=>"011010101",
  56819=>"000010001",
  56820=>"101000000",
  56821=>"111101000",
  56822=>"100111101",
  56823=>"101100011",
  56824=>"101011111",
  56825=>"100111100",
  56826=>"010111101",
  56827=>"011111001",
  56828=>"111111101",
  56829=>"010000101",
  56830=>"101110010",
  56831=>"100000111",
  56832=>"111011110",
  56833=>"000111101",
  56834=>"001100110",
  56835=>"010001001",
  56836=>"110001001",
  56837=>"010100110",
  56838=>"001110100",
  56839=>"101100001",
  56840=>"111011011",
  56841=>"000110111",
  56842=>"010000000",
  56843=>"111000000",
  56844=>"111010100",
  56845=>"101101111",
  56846=>"000000010",
  56847=>"110111111",
  56848=>"101001100",
  56849=>"001100010",
  56850=>"001101110",
  56851=>"110100001",
  56852=>"101111111",
  56853=>"101110110",
  56854=>"110001010",
  56855=>"111011011",
  56856=>"111001111",
  56857=>"100001000",
  56858=>"100111001",
  56859=>"001110001",
  56860=>"001101100",
  56861=>"101101100",
  56862=>"111110010",
  56863=>"101110000",
  56864=>"010010000",
  56865=>"101101011",
  56866=>"000101100",
  56867=>"000110001",
  56868=>"010101111",
  56869=>"001110001",
  56870=>"111100010",
  56871=>"100011100",
  56872=>"010010000",
  56873=>"111001101",
  56874=>"010001111",
  56875=>"111101011",
  56876=>"100111100",
  56877=>"011001101",
  56878=>"011101101",
  56879=>"001010010",
  56880=>"010100000",
  56881=>"100110010",
  56882=>"101111111",
  56883=>"100100110",
  56884=>"100001111",
  56885=>"101001110",
  56886=>"101011110",
  56887=>"100001001",
  56888=>"011110010",
  56889=>"101110101",
  56890=>"010110010",
  56891=>"101000001",
  56892=>"001010011",
  56893=>"001001110",
  56894=>"000000010",
  56895=>"101001011",
  56896=>"011000110",
  56897=>"110110001",
  56898=>"001111000",
  56899=>"100101111",
  56900=>"000001000",
  56901=>"101001000",
  56902=>"011100100",
  56903=>"001000010",
  56904=>"000100011",
  56905=>"010011000",
  56906=>"011100110",
  56907=>"100010000",
  56908=>"111111101",
  56909=>"000110101",
  56910=>"010011010",
  56911=>"001110000",
  56912=>"011101101",
  56913=>"011101110",
  56914=>"100000110",
  56915=>"100010001",
  56916=>"001111100",
  56917=>"001100110",
  56918=>"000001010",
  56919=>"111011000",
  56920=>"010000000",
  56921=>"011101101",
  56922=>"110100011",
  56923=>"000001111",
  56924=>"000100000",
  56925=>"011111001",
  56926=>"111011101",
  56927=>"101101001",
  56928=>"110000001",
  56929=>"100001111",
  56930=>"001001110",
  56931=>"111010101",
  56932=>"000011010",
  56933=>"001110110",
  56934=>"110110011",
  56935=>"001010011",
  56936=>"001100100",
  56937=>"111001010",
  56938=>"010101101",
  56939=>"111100010",
  56940=>"101000000",
  56941=>"101011011",
  56942=>"110010100",
  56943=>"111010110",
  56944=>"000010011",
  56945=>"111111111",
  56946=>"011001010",
  56947=>"010010100",
  56948=>"110101000",
  56949=>"000100000",
  56950=>"001110110",
  56951=>"010011111",
  56952=>"010000110",
  56953=>"100101010",
  56954=>"000010000",
  56955=>"011011011",
  56956=>"011111001",
  56957=>"000011101",
  56958=>"111010100",
  56959=>"110111010",
  56960=>"010111110",
  56961=>"011010110",
  56962=>"010111101",
  56963=>"001011000",
  56964=>"001011111",
  56965=>"001010101",
  56966=>"110001101",
  56967=>"010000101",
  56968=>"100111010",
  56969=>"110100100",
  56970=>"101001010",
  56971=>"110001000",
  56972=>"001110000",
  56973=>"000100011",
  56974=>"110000100",
  56975=>"011010001",
  56976=>"100011001",
  56977=>"100100010",
  56978=>"000110111",
  56979=>"100111000",
  56980=>"100011101",
  56981=>"100011111",
  56982=>"101001011",
  56983=>"111011001",
  56984=>"100101001",
  56985=>"101111111",
  56986=>"001100001",
  56987=>"010010110",
  56988=>"010011000",
  56989=>"010010111",
  56990=>"111110101",
  56991=>"100011110",
  56992=>"001011111",
  56993=>"010110000",
  56994=>"000000000",
  56995=>"111100011",
  56996=>"101010101",
  56997=>"110110100",
  56998=>"000000111",
  56999=>"110111101",
  57000=>"101010000",
  57001=>"101100001",
  57002=>"000100110",
  57003=>"101101010",
  57004=>"100010001",
  57005=>"111010101",
  57006=>"111101011",
  57007=>"100001000",
  57008=>"111111000",
  57009=>"111000111",
  57010=>"110011101",
  57011=>"111111100",
  57012=>"111001111",
  57013=>"010100110",
  57014=>"110000001",
  57015=>"001110011",
  57016=>"111110011",
  57017=>"000100001",
  57018=>"110011001",
  57019=>"111110000",
  57020=>"101110000",
  57021=>"110000111",
  57022=>"110010101",
  57023=>"110101110",
  57024=>"110100000",
  57025=>"111011111",
  57026=>"000001001",
  57027=>"111110010",
  57028=>"001100111",
  57029=>"011110000",
  57030=>"011011000",
  57031=>"110110000",
  57032=>"101101001",
  57033=>"000101101",
  57034=>"010001001",
  57035=>"110010101",
  57036=>"011000101",
  57037=>"110011000",
  57038=>"111001110",
  57039=>"000101000",
  57040=>"110000000",
  57041=>"010110001",
  57042=>"000001011",
  57043=>"100000101",
  57044=>"110100000",
  57045=>"111001100",
  57046=>"100101111",
  57047=>"000110011",
  57048=>"110010000",
  57049=>"110010001",
  57050=>"101101110",
  57051=>"000100001",
  57052=>"101101101",
  57053=>"011011111",
  57054=>"001111100",
  57055=>"101100111",
  57056=>"000111010",
  57057=>"010101111",
  57058=>"000101101",
  57059=>"110001000",
  57060=>"010010110",
  57061=>"101011110",
  57062=>"000100010",
  57063=>"000000010",
  57064=>"011000001",
  57065=>"111011110",
  57066=>"000100111",
  57067=>"001000011",
  57068=>"000001100",
  57069=>"000000100",
  57070=>"010110101",
  57071=>"111011101",
  57072=>"001111100",
  57073=>"000001101",
  57074=>"010110110",
  57075=>"111011011",
  57076=>"101111011",
  57077=>"011010001",
  57078=>"111110000",
  57079=>"111110011",
  57080=>"101101010",
  57081=>"111111000",
  57082=>"101100000",
  57083=>"101001110",
  57084=>"101011101",
  57085=>"111100100",
  57086=>"011000011",
  57087=>"000010010",
  57088=>"111000001",
  57089=>"101110001",
  57090=>"100100011",
  57091=>"111111011",
  57092=>"101011000",
  57093=>"101011010",
  57094=>"111111000",
  57095=>"000010101",
  57096=>"101011100",
  57097=>"110100001",
  57098=>"001000001",
  57099=>"101100011",
  57100=>"000011000",
  57101=>"110111111",
  57102=>"000010011",
  57103=>"100000010",
  57104=>"000011000",
  57105=>"110000010",
  57106=>"100000000",
  57107=>"111010001",
  57108=>"000000111",
  57109=>"001001001",
  57110=>"101000100",
  57111=>"011111001",
  57112=>"100001111",
  57113=>"100010110",
  57114=>"010011010",
  57115=>"101001111",
  57116=>"111001011",
  57117=>"010000011",
  57118=>"110011000",
  57119=>"100110011",
  57120=>"111010100",
  57121=>"100100011",
  57122=>"110010110",
  57123=>"101111011",
  57124=>"110111100",
  57125=>"111101110",
  57126=>"000000111",
  57127=>"001101000",
  57128=>"110110111",
  57129=>"111111010",
  57130=>"010100011",
  57131=>"111111011",
  57132=>"100110101",
  57133=>"100010010",
  57134=>"001001001",
  57135=>"000111000",
  57136=>"100001100",
  57137=>"100100100",
  57138=>"111011010",
  57139=>"001011001",
  57140=>"110111111",
  57141=>"011101101",
  57142=>"010011011",
  57143=>"101101101",
  57144=>"001100110",
  57145=>"000010010",
  57146=>"010010111",
  57147=>"111011110",
  57148=>"001000000",
  57149=>"111110110",
  57150=>"000011111",
  57151=>"101111001",
  57152=>"110000000",
  57153=>"100010110",
  57154=>"101000011",
  57155=>"100100011",
  57156=>"001101110",
  57157=>"001010101",
  57158=>"011111000",
  57159=>"000100101",
  57160=>"000101011",
  57161=>"110011000",
  57162=>"011010100",
  57163=>"111010011",
  57164=>"100011010",
  57165=>"001000101",
  57166=>"011110010",
  57167=>"100110110",
  57168=>"010110100",
  57169=>"101001000",
  57170=>"110000000",
  57171=>"111100100",
  57172=>"110110101",
  57173=>"010100011",
  57174=>"000110010",
  57175=>"001000111",
  57176=>"101100101",
  57177=>"001011101",
  57178=>"100010111",
  57179=>"001001000",
  57180=>"101100010",
  57181=>"001100101",
  57182=>"001110011",
  57183=>"010110010",
  57184=>"100100011",
  57185=>"010011110",
  57186=>"110011000",
  57187=>"010100100",
  57188=>"100001000",
  57189=>"011111011",
  57190=>"011111101",
  57191=>"010111101",
  57192=>"010110001",
  57193=>"010011011",
  57194=>"100101101",
  57195=>"111110110",
  57196=>"111110100",
  57197=>"111100101",
  57198=>"001000100",
  57199=>"010101011",
  57200=>"010011000",
  57201=>"111001100",
  57202=>"001110000",
  57203=>"000010101",
  57204=>"111111101",
  57205=>"010000110",
  57206=>"111000110",
  57207=>"101010011",
  57208=>"100101110",
  57209=>"001000100",
  57210=>"111100010",
  57211=>"011010000",
  57212=>"000010010",
  57213=>"101100111",
  57214=>"110100110",
  57215=>"111110011",
  57216=>"110001101",
  57217=>"010110011",
  57218=>"101001110",
  57219=>"010010110",
  57220=>"011111011",
  57221=>"100001001",
  57222=>"101001010",
  57223=>"000111101",
  57224=>"111011110",
  57225=>"011001100",
  57226=>"011110110",
  57227=>"011011101",
  57228=>"000101010",
  57229=>"001000110",
  57230=>"001000010",
  57231=>"110111110",
  57232=>"101100111",
  57233=>"100000011",
  57234=>"011111111",
  57235=>"000010011",
  57236=>"111010111",
  57237=>"111111000",
  57238=>"111010100",
  57239=>"010111101",
  57240=>"101000001",
  57241=>"000011001",
  57242=>"111110000",
  57243=>"100101010",
  57244=>"010111010",
  57245=>"111111011",
  57246=>"110100011",
  57247=>"011000000",
  57248=>"101110101",
  57249=>"111000101",
  57250=>"000110110",
  57251=>"010010110",
  57252=>"000110001",
  57253=>"011100001",
  57254=>"010000111",
  57255=>"100000001",
  57256=>"100110110",
  57257=>"010100000",
  57258=>"100110111",
  57259=>"111110100",
  57260=>"001001111",
  57261=>"101110100",
  57262=>"110011101",
  57263=>"000001110",
  57264=>"110010101",
  57265=>"010010111",
  57266=>"111011110",
  57267=>"111111100",
  57268=>"111100111",
  57269=>"001111011",
  57270=>"111101111",
  57271=>"111101101",
  57272=>"100101011",
  57273=>"101100001",
  57274=>"110000000",
  57275=>"011011101",
  57276=>"011011000",
  57277=>"000010000",
  57278=>"001111001",
  57279=>"010001100",
  57280=>"111110110",
  57281=>"100101001",
  57282=>"011001001",
  57283=>"110010000",
  57284=>"001000100",
  57285=>"101110010",
  57286=>"010010001",
  57287=>"110111101",
  57288=>"100011100",
  57289=>"011010110",
  57290=>"001010000",
  57291=>"101111011",
  57292=>"001000010",
  57293=>"110010010",
  57294=>"101010011",
  57295=>"101000001",
  57296=>"110010001",
  57297=>"011101111",
  57298=>"111111001",
  57299=>"010101000",
  57300=>"111010011",
  57301=>"110100111",
  57302=>"100001100",
  57303=>"011100000",
  57304=>"001110101",
  57305=>"100100101",
  57306=>"110100111",
  57307=>"110101111",
  57308=>"101001110",
  57309=>"010000111",
  57310=>"100010010",
  57311=>"000101011",
  57312=>"001111000",
  57313=>"011101110",
  57314=>"110010001",
  57315=>"101100100",
  57316=>"100101010",
  57317=>"111010000",
  57318=>"001101100",
  57319=>"000000001",
  57320=>"011001000",
  57321=>"111110110",
  57322=>"101001110",
  57323=>"001110100",
  57324=>"100001100",
  57325=>"110001100",
  57326=>"101000101",
  57327=>"011010010",
  57328=>"100100100",
  57329=>"000000000",
  57330=>"111000101",
  57331=>"110001001",
  57332=>"011101011",
  57333=>"000000000",
  57334=>"101101100",
  57335=>"010000010",
  57336=>"100001110",
  57337=>"110000111",
  57338=>"110100100",
  57339=>"100000100",
  57340=>"000111111",
  57341=>"011010100",
  57342=>"111100010",
  57343=>"011100101",
  57344=>"111000110",
  57345=>"101111010",
  57346=>"111010111",
  57347=>"001111101",
  57348=>"010000100",
  57349=>"110111000",
  57350=>"100101000",
  57351=>"100100101",
  57352=>"010101110",
  57353=>"101000111",
  57354=>"111101001",
  57355=>"100110111",
  57356=>"101111001",
  57357=>"010111000",
  57358=>"010001110",
  57359=>"100001001",
  57360=>"010000011",
  57361=>"000001000",
  57362=>"111101010",
  57363=>"001110010",
  57364=>"111001111",
  57365=>"011011000",
  57366=>"010111001",
  57367=>"110000000",
  57368=>"111011100",
  57369=>"110110110",
  57370=>"011111010",
  57371=>"111100110",
  57372=>"101110011",
  57373=>"110100101",
  57374=>"010100011",
  57375=>"011100010",
  57376=>"011001100",
  57377=>"010011110",
  57378=>"101011011",
  57379=>"000110000",
  57380=>"001001001",
  57381=>"010010000",
  57382=>"101001110",
  57383=>"101101010",
  57384=>"110100010",
  57385=>"000000010",
  57386=>"010111011",
  57387=>"100100010",
  57388=>"111111011",
  57389=>"000101010",
  57390=>"110111111",
  57391=>"011001111",
  57392=>"011100011",
  57393=>"011111100",
  57394=>"111000111",
  57395=>"010010010",
  57396=>"010000111",
  57397=>"000000110",
  57398=>"101000110",
  57399=>"100010110",
  57400=>"001001001",
  57401=>"001010100",
  57402=>"111111110",
  57403=>"101111010",
  57404=>"011110100",
  57405=>"100010100",
  57406=>"000010110",
  57407=>"100111001",
  57408=>"010110101",
  57409=>"110100111",
  57410=>"101101010",
  57411=>"010100100",
  57412=>"001100110",
  57413=>"111101001",
  57414=>"101110001",
  57415=>"101100000",
  57416=>"010111010",
  57417=>"011001101",
  57418=>"001000000",
  57419=>"000110011",
  57420=>"011010101",
  57421=>"100101111",
  57422=>"101010010",
  57423=>"010011001",
  57424=>"111101001",
  57425=>"111111011",
  57426=>"100010011",
  57427=>"001101100",
  57428=>"100001111",
  57429=>"000101000",
  57430=>"000101101",
  57431=>"000111001",
  57432=>"011100000",
  57433=>"001000101",
  57434=>"111110100",
  57435=>"010010111",
  57436=>"000011001",
  57437=>"000100111",
  57438=>"100011111",
  57439=>"111101111",
  57440=>"001000000",
  57441=>"111101110",
  57442=>"111110001",
  57443=>"110100110",
  57444=>"101010111",
  57445=>"000100001",
  57446=>"101001011",
  57447=>"101001101",
  57448=>"000110010",
  57449=>"101111000",
  57450=>"001010010",
  57451=>"011000011",
  57452=>"001001111",
  57453=>"100110010",
  57454=>"101011011",
  57455=>"111000000",
  57456=>"001011001",
  57457=>"110011001",
  57458=>"111000010",
  57459=>"001101111",
  57460=>"111011010",
  57461=>"110010100",
  57462=>"100010111",
  57463=>"000110010",
  57464=>"001011111",
  57465=>"111000010",
  57466=>"111101011",
  57467=>"001001111",
  57468=>"001000000",
  57469=>"101100001",
  57470=>"111110111",
  57471=>"010101100",
  57472=>"000011011",
  57473=>"110010101",
  57474=>"111110110",
  57475=>"100110000",
  57476=>"011101111",
  57477=>"101001000",
  57478=>"100111011",
  57479=>"111000110",
  57480=>"001101111",
  57481=>"000110110",
  57482=>"101001001",
  57483=>"001110101",
  57484=>"110101110",
  57485=>"010111101",
  57486=>"100100011",
  57487=>"010100010",
  57488=>"110000101",
  57489=>"010100110",
  57490=>"001000001",
  57491=>"110100010",
  57492=>"100100101",
  57493=>"000101000",
  57494=>"110001101",
  57495=>"000100111",
  57496=>"101101101",
  57497=>"110100000",
  57498=>"111000110",
  57499=>"111101010",
  57500=>"011000000",
  57501=>"110100000",
  57502=>"010010011",
  57503=>"110000100",
  57504=>"011110011",
  57505=>"011110000",
  57506=>"001101111",
  57507=>"100010000",
  57508=>"001100000",
  57509=>"101000000",
  57510=>"101100001",
  57511=>"010000000",
  57512=>"111000111",
  57513=>"111011101",
  57514=>"100100111",
  57515=>"100101100",
  57516=>"001011100",
  57517=>"111011010",
  57518=>"100001111",
  57519=>"001010010",
  57520=>"000001111",
  57521=>"110001111",
  57522=>"011011010",
  57523=>"010011011",
  57524=>"010110000",
  57525=>"010000111",
  57526=>"000110010",
  57527=>"101001100",
  57528=>"000010111",
  57529=>"100011110",
  57530=>"010010101",
  57531=>"100001100",
  57532=>"001010000",
  57533=>"010011110",
  57534=>"111001010",
  57535=>"111110110",
  57536=>"000001011",
  57537=>"010100101",
  57538=>"000001111",
  57539=>"011000010",
  57540=>"000110011",
  57541=>"101100110",
  57542=>"000010010",
  57543=>"001100011",
  57544=>"110100101",
  57545=>"101110101",
  57546=>"100000101",
  57547=>"001111111",
  57548=>"000111110",
  57549=>"101111010",
  57550=>"110111100",
  57551=>"101000000",
  57552=>"101011000",
  57553=>"111000010",
  57554=>"000011100",
  57555=>"011011111",
  57556=>"010011010",
  57557=>"101111011",
  57558=>"011010011",
  57559=>"111001011",
  57560=>"010000000",
  57561=>"100010000",
  57562=>"010001110",
  57563=>"101001010",
  57564=>"010010001",
  57565=>"000110001",
  57566=>"101111000",
  57567=>"000011101",
  57568=>"000110000",
  57569=>"010101001",
  57570=>"111010010",
  57571=>"000101110",
  57572=>"001011100",
  57573=>"101100001",
  57574=>"111111111",
  57575=>"011111100",
  57576=>"010011001",
  57577=>"110000000",
  57578=>"010111110",
  57579=>"000000100",
  57580=>"010000110",
  57581=>"001010010",
  57582=>"111000101",
  57583=>"101111000",
  57584=>"000000001",
  57585=>"111001011",
  57586=>"111010111",
  57587=>"010110100",
  57588=>"011000101",
  57589=>"010010011",
  57590=>"010001010",
  57591=>"101100010",
  57592=>"101010010",
  57593=>"100011101",
  57594=>"011100101",
  57595=>"111000011",
  57596=>"101110101",
  57597=>"110001000",
  57598=>"111111101",
  57599=>"100010010",
  57600=>"011001010",
  57601=>"000010001",
  57602=>"111110100",
  57603=>"101111010",
  57604=>"010000010",
  57605=>"110111101",
  57606=>"010010001",
  57607=>"111011011",
  57608=>"000110111",
  57609=>"000010111",
  57610=>"101101101",
  57611=>"000101001",
  57612=>"111000011",
  57613=>"101011011",
  57614=>"101101000",
  57615=>"000110001",
  57616=>"000001100",
  57617=>"010111111",
  57618=>"011110010",
  57619=>"001111011",
  57620=>"111110101",
  57621=>"101101101",
  57622=>"100101001",
  57623=>"111111100",
  57624=>"110011000",
  57625=>"110100001",
  57626=>"110001011",
  57627=>"100000111",
  57628=>"011011001",
  57629=>"101101111",
  57630=>"001011100",
  57631=>"100111111",
  57632=>"111010101",
  57633=>"011001001",
  57634=>"110111111",
  57635=>"010111001",
  57636=>"111100001",
  57637=>"010000000",
  57638=>"010110100",
  57639=>"110110000",
  57640=>"110100001",
  57641=>"011011111",
  57642=>"001000110",
  57643=>"100100010",
  57644=>"111000000",
  57645=>"101000111",
  57646=>"000011011",
  57647=>"001111111",
  57648=>"101000101",
  57649=>"000110010",
  57650=>"101110011",
  57651=>"101001001",
  57652=>"010110100",
  57653=>"111010000",
  57654=>"011101101",
  57655=>"111111101",
  57656=>"000100111",
  57657=>"110111111",
  57658=>"110101001",
  57659=>"000101011",
  57660=>"000001011",
  57661=>"100101001",
  57662=>"110110111",
  57663=>"011000000",
  57664=>"010111001",
  57665=>"000100011",
  57666=>"111010001",
  57667=>"111110011",
  57668=>"100101011",
  57669=>"000111101",
  57670=>"111011011",
  57671=>"110111101",
  57672=>"001101000",
  57673=>"111101111",
  57674=>"000110101",
  57675=>"101111001",
  57676=>"110011000",
  57677=>"010101110",
  57678=>"111001010",
  57679=>"111110110",
  57680=>"000100010",
  57681=>"111100000",
  57682=>"011111101",
  57683=>"010001111",
  57684=>"010101000",
  57685=>"011000001",
  57686=>"011000000",
  57687=>"100000101",
  57688=>"000110101",
  57689=>"100000000",
  57690=>"100000001",
  57691=>"111000000",
  57692=>"110110000",
  57693=>"111001001",
  57694=>"011001001",
  57695=>"111100101",
  57696=>"111100100",
  57697=>"011000000",
  57698=>"010000111",
  57699=>"111000111",
  57700=>"111001111",
  57701=>"101000111",
  57702=>"111110001",
  57703=>"111100110",
  57704=>"011100100",
  57705=>"010111101",
  57706=>"011100001",
  57707=>"010101111",
  57708=>"110000001",
  57709=>"001110001",
  57710=>"011110011",
  57711=>"100110110",
  57712=>"100001010",
  57713=>"111100000",
  57714=>"101000011",
  57715=>"111011000",
  57716=>"011111001",
  57717=>"101101101",
  57718=>"111111111",
  57719=>"111111001",
  57720=>"111000101",
  57721=>"111101100",
  57722=>"011101111",
  57723=>"000101000",
  57724=>"000101111",
  57725=>"111010011",
  57726=>"101101111",
  57727=>"110011011",
  57728=>"111110000",
  57729=>"001010001",
  57730=>"001101000",
  57731=>"001011001",
  57732=>"111100011",
  57733=>"100101101",
  57734=>"101000010",
  57735=>"100100010",
  57736=>"010010001",
  57737=>"111111110",
  57738=>"001011010",
  57739=>"100010111",
  57740=>"000001100",
  57741=>"110110000",
  57742=>"001000110",
  57743=>"111100000",
  57744=>"011101011",
  57745=>"101100111",
  57746=>"111000011",
  57747=>"100011110",
  57748=>"010110111",
  57749=>"101100101",
  57750=>"010001000",
  57751=>"101011010",
  57752=>"100000101",
  57753=>"101001100",
  57754=>"001100101",
  57755=>"111100101",
  57756=>"000101111",
  57757=>"001011010",
  57758=>"010101110",
  57759=>"011101001",
  57760=>"101101101",
  57761=>"000000100",
  57762=>"100100100",
  57763=>"100000010",
  57764=>"111000110",
  57765=>"001000100",
  57766=>"100011101",
  57767=>"111100100",
  57768=>"001000011",
  57769=>"000110011",
  57770=>"001001001",
  57771=>"010000101",
  57772=>"011101111",
  57773=>"111110100",
  57774=>"101101101",
  57775=>"100100001",
  57776=>"111110100",
  57777=>"100111111",
  57778=>"100111100",
  57779=>"000101000",
  57780=>"011111010",
  57781=>"111111001",
  57782=>"100100101",
  57783=>"110100011",
  57784=>"011111000",
  57785=>"000001110",
  57786=>"010001011",
  57787=>"011001100",
  57788=>"001110000",
  57789=>"100101000",
  57790=>"000010111",
  57791=>"110001011",
  57792=>"011110100",
  57793=>"011011010",
  57794=>"110101110",
  57795=>"111011000",
  57796=>"101111111",
  57797=>"000110000",
  57798=>"000000010",
  57799=>"011100110",
  57800=>"011101010",
  57801=>"001100011",
  57802=>"011010101",
  57803=>"011001111",
  57804=>"011100111",
  57805=>"010111000",
  57806=>"000101001",
  57807=>"001011011",
  57808=>"011001111",
  57809=>"111111110",
  57810=>"111100110",
  57811=>"000001101",
  57812=>"111101111",
  57813=>"110011101",
  57814=>"110010010",
  57815=>"111100011",
  57816=>"100001000",
  57817=>"010011100",
  57818=>"101110010",
  57819=>"100111101",
  57820=>"100000010",
  57821=>"000010010",
  57822=>"101010100",
  57823=>"010011010",
  57824=>"001001111",
  57825=>"000100001",
  57826=>"110100111",
  57827=>"000111110",
  57828=>"001000010",
  57829=>"101111111",
  57830=>"100110010",
  57831=>"100100111",
  57832=>"101010101",
  57833=>"100101010",
  57834=>"110100001",
  57835=>"010011100",
  57836=>"111101010",
  57837=>"000000111",
  57838=>"110000111",
  57839=>"000001010",
  57840=>"001011100",
  57841=>"000010010",
  57842=>"010010001",
  57843=>"001111111",
  57844=>"010110100",
  57845=>"100111000",
  57846=>"111101010",
  57847=>"100100110",
  57848=>"010011111",
  57849=>"010111011",
  57850=>"011111000",
  57851=>"010011001",
  57852=>"010000010",
  57853=>"101100000",
  57854=>"000000100",
  57855=>"111010001",
  57856=>"101111000",
  57857=>"011011101",
  57858=>"100010110",
  57859=>"001101001",
  57860=>"110010011",
  57861=>"110100010",
  57862=>"100100001",
  57863=>"011010010",
  57864=>"101001111",
  57865=>"000011111",
  57866=>"111101001",
  57867=>"100101101",
  57868=>"001010111",
  57869=>"100000110",
  57870=>"000000110",
  57871=>"111101010",
  57872=>"000000101",
  57873=>"100100011",
  57874=>"011001101",
  57875=>"111001011",
  57876=>"100010111",
  57877=>"101010111",
  57878=>"011000000",
  57879=>"010001110",
  57880=>"110101000",
  57881=>"001101010",
  57882=>"001011100",
  57883=>"100001010",
  57884=>"110110101",
  57885=>"000110100",
  57886=>"000101101",
  57887=>"010110110",
  57888=>"010000001",
  57889=>"110100011",
  57890=>"100000110",
  57891=>"101011101",
  57892=>"101111111",
  57893=>"111110100",
  57894=>"011010010",
  57895=>"100101011",
  57896=>"000100111",
  57897=>"101111011",
  57898=>"101111101",
  57899=>"010111011",
  57900=>"000111100",
  57901=>"010101001",
  57902=>"111101001",
  57903=>"100010000",
  57904=>"010100010",
  57905=>"110110111",
  57906=>"010111000",
  57907=>"111110100",
  57908=>"001001111",
  57909=>"010110001",
  57910=>"111101010",
  57911=>"110111000",
  57912=>"000001000",
  57913=>"000011000",
  57914=>"101011000",
  57915=>"001001100",
  57916=>"010000011",
  57917=>"010011011",
  57918=>"111000011",
  57919=>"010000000",
  57920=>"011101110",
  57921=>"011111111",
  57922=>"110011101",
  57923=>"100000101",
  57924=>"101110000",
  57925=>"100100010",
  57926=>"000100001",
  57927=>"100000111",
  57928=>"100001011",
  57929=>"011000100",
  57930=>"000100111",
  57931=>"011011011",
  57932=>"000010111",
  57933=>"101101000",
  57934=>"111001100",
  57935=>"001011111",
  57936=>"110100111",
  57937=>"011101111",
  57938=>"001010110",
  57939=>"100001110",
  57940=>"101000011",
  57941=>"100000001",
  57942=>"111011000",
  57943=>"111000011",
  57944=>"110000100",
  57945=>"110110111",
  57946=>"011111010",
  57947=>"011111111",
  57948=>"100101001",
  57949=>"000001001",
  57950=>"110110110",
  57951=>"111100111",
  57952=>"001110011",
  57953=>"011111001",
  57954=>"100111101",
  57955=>"010100000",
  57956=>"000100101",
  57957=>"010100001",
  57958=>"110001010",
  57959=>"100101001",
  57960=>"010100101",
  57961=>"101111001",
  57962=>"001000001",
  57963=>"111111111",
  57964=>"010010011",
  57965=>"110101101",
  57966=>"110011100",
  57967=>"000000000",
  57968=>"100101100",
  57969=>"000000001",
  57970=>"000010001",
  57971=>"100110011",
  57972=>"010001000",
  57973=>"000000000",
  57974=>"000111110",
  57975=>"011111101",
  57976=>"110001010",
  57977=>"101101101",
  57978=>"011101111",
  57979=>"011110111",
  57980=>"000001000",
  57981=>"100110110",
  57982=>"000000111",
  57983=>"011111000",
  57984=>"100001001",
  57985=>"110001001",
  57986=>"111010000",
  57987=>"100001000",
  57988=>"110100101",
  57989=>"011100000",
  57990=>"111110100",
  57991=>"100001010",
  57992=>"101110110",
  57993=>"110010001",
  57994=>"000110010",
  57995=>"000001110",
  57996=>"101011000",
  57997=>"000010000",
  57998=>"111010010",
  57999=>"100000111",
  58000=>"101010111",
  58001=>"110111110",
  58002=>"011110110",
  58003=>"010010111",
  58004=>"000010010",
  58005=>"111110010",
  58006=>"110001001",
  58007=>"100010010",
  58008=>"001010010",
  58009=>"100111111",
  58010=>"100011110",
  58011=>"010001011",
  58012=>"101011111",
  58013=>"000001011",
  58014=>"110010110",
  58015=>"100110000",
  58016=>"110000101",
  58017=>"001000110",
  58018=>"110111110",
  58019=>"110010000",
  58020=>"101110011",
  58021=>"000000010",
  58022=>"110001100",
  58023=>"000011000",
  58024=>"100101001",
  58025=>"011000000",
  58026=>"001101011",
  58027=>"010010101",
  58028=>"100100011",
  58029=>"111101100",
  58030=>"111010001",
  58031=>"100010000",
  58032=>"010000000",
  58033=>"111001111",
  58034=>"111101111",
  58035=>"001110111",
  58036=>"111110011",
  58037=>"100000101",
  58038=>"101010111",
  58039=>"011101101",
  58040=>"111100011",
  58041=>"011001110",
  58042=>"110100010",
  58043=>"001100000",
  58044=>"000101010",
  58045=>"110011101",
  58046=>"001100011",
  58047=>"001101101",
  58048=>"100010111",
  58049=>"000110100",
  58050=>"101101011",
  58051=>"011111101",
  58052=>"110110110",
  58053=>"000100110",
  58054=>"101101111",
  58055=>"011011001",
  58056=>"101000010",
  58057=>"111001001",
  58058=>"110000100",
  58059=>"111010100",
  58060=>"110011111",
  58061=>"110001100",
  58062=>"011001111",
  58063=>"111100001",
  58064=>"100111000",
  58065=>"101010101",
  58066=>"111000101",
  58067=>"100100100",
  58068=>"111001101",
  58069=>"001110111",
  58070=>"001101110",
  58071=>"010011011",
  58072=>"001000001",
  58073=>"111011010",
  58074=>"000001111",
  58075=>"110001001",
  58076=>"000000110",
  58077=>"110000000",
  58078=>"001001010",
  58079=>"001010001",
  58080=>"000000000",
  58081=>"111110101",
  58082=>"101101101",
  58083=>"101000100",
  58084=>"001101000",
  58085=>"010101011",
  58086=>"000111101",
  58087=>"111000110",
  58088=>"001011011",
  58089=>"110010100",
  58090=>"000010000",
  58091=>"101110001",
  58092=>"000001000",
  58093=>"001111111",
  58094=>"101110010",
  58095=>"111111111",
  58096=>"111001110",
  58097=>"110100000",
  58098=>"010101011",
  58099=>"110000110",
  58100=>"101000010",
  58101=>"101100011",
  58102=>"001001001",
  58103=>"110101110",
  58104=>"011000010",
  58105=>"000110110",
  58106=>"001010011",
  58107=>"011110101",
  58108=>"001011000",
  58109=>"101000100",
  58110=>"110101011",
  58111=>"000111100",
  58112=>"011101110",
  58113=>"000010010",
  58114=>"000101001",
  58115=>"111100111",
  58116=>"000100100",
  58117=>"000110011",
  58118=>"110000111",
  58119=>"001001111",
  58120=>"110001010",
  58121=>"110001110",
  58122=>"111100101",
  58123=>"000010010",
  58124=>"010111111",
  58125=>"010001011",
  58126=>"000111010",
  58127=>"110101111",
  58128=>"101100101",
  58129=>"110001110",
  58130=>"010000000",
  58131=>"001010110",
  58132=>"111001111",
  58133=>"100000001",
  58134=>"110110111",
  58135=>"111000011",
  58136=>"101001101",
  58137=>"000011011",
  58138=>"001001111",
  58139=>"000100001",
  58140=>"000000100",
  58141=>"110111110",
  58142=>"111000100",
  58143=>"010010001",
  58144=>"000001011",
  58145=>"101000111",
  58146=>"010111101",
  58147=>"101110010",
  58148=>"100101000",
  58149=>"010110000",
  58150=>"111111111",
  58151=>"001101001",
  58152=>"101001111",
  58153=>"110000111",
  58154=>"111101000",
  58155=>"100101100",
  58156=>"110001010",
  58157=>"000000011",
  58158=>"110111001",
  58159=>"110110011",
  58160=>"000010111",
  58161=>"000010110",
  58162=>"110111110",
  58163=>"000101000",
  58164=>"101000110",
  58165=>"111111101",
  58166=>"010010111",
  58167=>"000010001",
  58168=>"100100001",
  58169=>"100010000",
  58170=>"011111101",
  58171=>"001100111",
  58172=>"101100101",
  58173=>"001101011",
  58174=>"101011001",
  58175=>"101101011",
  58176=>"000100100",
  58177=>"110001011",
  58178=>"100100110",
  58179=>"011101100",
  58180=>"111010011",
  58181=>"001000110",
  58182=>"111011001",
  58183=>"010011001",
  58184=>"010111001",
  58185=>"101101111",
  58186=>"011011000",
  58187=>"001110000",
  58188=>"011001011",
  58189=>"000010100",
  58190=>"010011010",
  58191=>"100110010",
  58192=>"011101111",
  58193=>"000111001",
  58194=>"101110001",
  58195=>"001100000",
  58196=>"101110111",
  58197=>"001001101",
  58198=>"100101000",
  58199=>"100011110",
  58200=>"111111010",
  58201=>"000101111",
  58202=>"001000101",
  58203=>"101000111",
  58204=>"001000100",
  58205=>"010010101",
  58206=>"010010010",
  58207=>"000000011",
  58208=>"110011111",
  58209=>"100111110",
  58210=>"001100111",
  58211=>"001011000",
  58212=>"111010011",
  58213=>"111010001",
  58214=>"110101101",
  58215=>"001010000",
  58216=>"010101001",
  58217=>"010000101",
  58218=>"011000000",
  58219=>"101000001",
  58220=>"000000010",
  58221=>"101010000",
  58222=>"011110101",
  58223=>"101011110",
  58224=>"101011111",
  58225=>"011001001",
  58226=>"011100101",
  58227=>"110111110",
  58228=>"000010101",
  58229=>"101011010",
  58230=>"110100101",
  58231=>"011100000",
  58232=>"100011001",
  58233=>"100000010",
  58234=>"101111001",
  58235=>"100100100",
  58236=>"111111111",
  58237=>"000001100",
  58238=>"101010110",
  58239=>"111011110",
  58240=>"001111010",
  58241=>"001101010",
  58242=>"000011100",
  58243=>"110010100",
  58244=>"100000110",
  58245=>"101101011",
  58246=>"111000100",
  58247=>"100001000",
  58248=>"000000000",
  58249=>"100101010",
  58250=>"000100100",
  58251=>"110011101",
  58252=>"001100011",
  58253=>"000001111",
  58254=>"010110000",
  58255=>"101101000",
  58256=>"101001110",
  58257=>"111011110",
  58258=>"000101001",
  58259=>"000000011",
  58260=>"000010010",
  58261=>"101001101",
  58262=>"001011011",
  58263=>"101001000",
  58264=>"010100000",
  58265=>"000011010",
  58266=>"000000100",
  58267=>"101000001",
  58268=>"111100001",
  58269=>"101110000",
  58270=>"101110111",
  58271=>"100110110",
  58272=>"111111010",
  58273=>"011101101",
  58274=>"100000100",
  58275=>"010010101",
  58276=>"010000100",
  58277=>"110110001",
  58278=>"100001011",
  58279=>"000001000",
  58280=>"101011110",
  58281=>"000110101",
  58282=>"110111110",
  58283=>"111000111",
  58284=>"111101011",
  58285=>"111010101",
  58286=>"001000011",
  58287=>"011011101",
  58288=>"100000000",
  58289=>"101111001",
  58290=>"100110001",
  58291=>"001101111",
  58292=>"000000000",
  58293=>"101000110",
  58294=>"111111111",
  58295=>"000100111",
  58296=>"001010101",
  58297=>"001110011",
  58298=>"100101010",
  58299=>"011010111",
  58300=>"000100010",
  58301=>"001110111",
  58302=>"111010010",
  58303=>"011111011",
  58304=>"111111110",
  58305=>"101010100",
  58306=>"001001001",
  58307=>"000101001",
  58308=>"110001110",
  58309=>"111111111",
  58310=>"111001100",
  58311=>"111010111",
  58312=>"010101101",
  58313=>"011110111",
  58314=>"000110001",
  58315=>"111000101",
  58316=>"111001010",
  58317=>"100110110",
  58318=>"100100100",
  58319=>"001110100",
  58320=>"110111101",
  58321=>"000011010",
  58322=>"000110110",
  58323=>"100111110",
  58324=>"111011101",
  58325=>"111010111",
  58326=>"101110001",
  58327=>"101010100",
  58328=>"110001111",
  58329=>"011001101",
  58330=>"101111001",
  58331=>"101011101",
  58332=>"100001100",
  58333=>"010110000",
  58334=>"011111101",
  58335=>"010001010",
  58336=>"111110000",
  58337=>"011000110",
  58338=>"111001100",
  58339=>"111101001",
  58340=>"101111001",
  58341=>"111111111",
  58342=>"001001010",
  58343=>"110000001",
  58344=>"000101000",
  58345=>"000101011",
  58346=>"110100011",
  58347=>"100101011",
  58348=>"000100110",
  58349=>"100001101",
  58350=>"000111101",
  58351=>"110001000",
  58352=>"000110111",
  58353=>"111001101",
  58354=>"000010110",
  58355=>"000100101",
  58356=>"001100110",
  58357=>"110101100",
  58358=>"111001110",
  58359=>"100101100",
  58360=>"001011111",
  58361=>"111001110",
  58362=>"001000100",
  58363=>"110100101",
  58364=>"001111111",
  58365=>"101111001",
  58366=>"101011011",
  58367=>"011011111",
  58368=>"000011100",
  58369=>"001111101",
  58370=>"000100010",
  58371=>"000011001",
  58372=>"010100000",
  58373=>"010111111",
  58374=>"000001111",
  58375=>"111010100",
  58376=>"011001111",
  58377=>"010010001",
  58378=>"001010100",
  58379=>"001101101",
  58380=>"011100101",
  58381=>"010000100",
  58382=>"110010010",
  58383=>"001001101",
  58384=>"111100100",
  58385=>"000010111",
  58386=>"101001011",
  58387=>"110100110",
  58388=>"110000111",
  58389=>"100101000",
  58390=>"111110100",
  58391=>"001000101",
  58392=>"111011100",
  58393=>"011110001",
  58394=>"000001011",
  58395=>"001011010",
  58396=>"111000111",
  58397=>"010001011",
  58398=>"110101110",
  58399=>"010110110",
  58400=>"111111001",
  58401=>"100000111",
  58402=>"110011010",
  58403=>"000101011",
  58404=>"111110000",
  58405=>"000111011",
  58406=>"000101011",
  58407=>"001111000",
  58408=>"000110110",
  58409=>"101101000",
  58410=>"000000110",
  58411=>"101010101",
  58412=>"011101011",
  58413=>"001100001",
  58414=>"101111111",
  58415=>"111010100",
  58416=>"000010001",
  58417=>"100110111",
  58418=>"001110100",
  58419=>"100111110",
  58420=>"011001001",
  58421=>"010001010",
  58422=>"111010000",
  58423=>"001111010",
  58424=>"000110010",
  58425=>"100010101",
  58426=>"101110111",
  58427=>"001001100",
  58428=>"011110101",
  58429=>"000011101",
  58430=>"010100011",
  58431=>"110111101",
  58432=>"111111111",
  58433=>"011111011",
  58434=>"111100110",
  58435=>"101000000",
  58436=>"010100100",
  58437=>"000000010",
  58438=>"110101010",
  58439=>"100001000",
  58440=>"110101001",
  58441=>"000001100",
  58442=>"100100101",
  58443=>"011111110",
  58444=>"110010100",
  58445=>"100101111",
  58446=>"010100110",
  58447=>"010101100",
  58448=>"001011110",
  58449=>"010011011",
  58450=>"100010010",
  58451=>"101010111",
  58452=>"110111111",
  58453=>"111011111",
  58454=>"110001010",
  58455=>"000011010",
  58456=>"000110000",
  58457=>"010111100",
  58458=>"001100100",
  58459=>"111000010",
  58460=>"000100111",
  58461=>"111001010",
  58462=>"011111111",
  58463=>"001101001",
  58464=>"001100000",
  58465=>"100010001",
  58466=>"111101110",
  58467=>"010001111",
  58468=>"001100001",
  58469=>"101110011",
  58470=>"101111011",
  58471=>"110111100",
  58472=>"110000010",
  58473=>"111110011",
  58474=>"110011111",
  58475=>"101101111",
  58476=>"101111110",
  58477=>"111001001",
  58478=>"010100010",
  58479=>"000000000",
  58480=>"001010000",
  58481=>"010111110",
  58482=>"001110101",
  58483=>"101100011",
  58484=>"010011111",
  58485=>"111111010",
  58486=>"100001001",
  58487=>"010000010",
  58488=>"001011111",
  58489=>"010000011",
  58490=>"110001101",
  58491=>"111111101",
  58492=>"010101110",
  58493=>"001011001",
  58494=>"110101000",
  58495=>"001000010",
  58496=>"100000000",
  58497=>"110110011",
  58498=>"100011011",
  58499=>"011001110",
  58500=>"001001111",
  58501=>"010000111",
  58502=>"000001100",
  58503=>"011110001",
  58504=>"000101100",
  58505=>"110101101",
  58506=>"010000010",
  58507=>"001001011",
  58508=>"000100000",
  58509=>"100110100",
  58510=>"001011011",
  58511=>"111000111",
  58512=>"100110001",
  58513=>"001010001",
  58514=>"101101111",
  58515=>"111101101",
  58516=>"111100001",
  58517=>"100100001",
  58518=>"011110111",
  58519=>"000001110",
  58520=>"000110010",
  58521=>"101001100",
  58522=>"111100100",
  58523=>"100100101",
  58524=>"000110010",
  58525=>"111001001",
  58526=>"110010001",
  58527=>"110001000",
  58528=>"110011110",
  58529=>"000010111",
  58530=>"000010010",
  58531=>"001010110",
  58532=>"110000010",
  58533=>"100100101",
  58534=>"011110101",
  58535=>"001011011",
  58536=>"100100111",
  58537=>"010010011",
  58538=>"010010110",
  58539=>"000001101",
  58540=>"001000100",
  58541=>"100111110",
  58542=>"010101111",
  58543=>"101111001",
  58544=>"110101101",
  58545=>"010001111",
  58546=>"011011101",
  58547=>"001100111",
  58548=>"111001110",
  58549=>"000010111",
  58550=>"111001011",
  58551=>"110101011",
  58552=>"000111001",
  58553=>"001100110",
  58554=>"000111010",
  58555=>"000011111",
  58556=>"111010010",
  58557=>"110000000",
  58558=>"101000000",
  58559=>"111101001",
  58560=>"101010011",
  58561=>"001011000",
  58562=>"100100010",
  58563=>"001101011",
  58564=>"101001000",
  58565=>"111111000",
  58566=>"010010110",
  58567=>"011010010",
  58568=>"110110011",
  58569=>"001001000",
  58570=>"111001000",
  58571=>"100100010",
  58572=>"011101010",
  58573=>"101000010",
  58574=>"100011111",
  58575=>"111111001",
  58576=>"011101011",
  58577=>"110010110",
  58578=>"111000110",
  58579=>"100111000",
  58580=>"111111000",
  58581=>"110110101",
  58582=>"010011100",
  58583=>"001000110",
  58584=>"000111111",
  58585=>"001101000",
  58586=>"110111101",
  58587=>"101011001",
  58588=>"000011110",
  58589=>"111111001",
  58590=>"010000111",
  58591=>"110111011",
  58592=>"010000001",
  58593=>"000011011",
  58594=>"010011101",
  58595=>"011001001",
  58596=>"010011010",
  58597=>"100100111",
  58598=>"000001001",
  58599=>"001110000",
  58600=>"100000111",
  58601=>"110101111",
  58602=>"101000000",
  58603=>"100111100",
  58604=>"110001110",
  58605=>"101101110",
  58606=>"100110000",
  58607=>"100010000",
  58608=>"001010001",
  58609=>"011011110",
  58610=>"111001111",
  58611=>"100010010",
  58612=>"100100011",
  58613=>"000000001",
  58614=>"011001010",
  58615=>"010110011",
  58616=>"100101111",
  58617=>"010101101",
  58618=>"000110100",
  58619=>"010110000",
  58620=>"101101111",
  58621=>"010000010",
  58622=>"011110000",
  58623=>"111111111",
  58624=>"111001011",
  58625=>"111000100",
  58626=>"001010100",
  58627=>"101010111",
  58628=>"010111110",
  58629=>"000111111",
  58630=>"110100101",
  58631=>"010100011",
  58632=>"011011101",
  58633=>"111110100",
  58634=>"101011011",
  58635=>"011010000",
  58636=>"110010100",
  58637=>"000111000",
  58638=>"001010100",
  58639=>"010100100",
  58640=>"011011001",
  58641=>"111000101",
  58642=>"010001001",
  58643=>"111111110",
  58644=>"101000001",
  58645=>"101111101",
  58646=>"010101000",
  58647=>"010000100",
  58648=>"001110001",
  58649=>"011111010",
  58650=>"111010001",
  58651=>"101000101",
  58652=>"010101100",
  58653=>"000000111",
  58654=>"110110111",
  58655=>"000000100",
  58656=>"100011011",
  58657=>"011010001",
  58658=>"110011100",
  58659=>"101010010",
  58660=>"010101000",
  58661=>"111100111",
  58662=>"100000001",
  58663=>"001001001",
  58664=>"010001101",
  58665=>"000111101",
  58666=>"001010101",
  58667=>"110101001",
  58668=>"001101001",
  58669=>"001100100",
  58670=>"001111111",
  58671=>"100000001",
  58672=>"101011000",
  58673=>"101101111",
  58674=>"010011001",
  58675=>"001000111",
  58676=>"110000111",
  58677=>"100010110",
  58678=>"111000000",
  58679=>"001001000",
  58680=>"011001100",
  58681=>"001001011",
  58682=>"010000000",
  58683=>"100000101",
  58684=>"100000011",
  58685=>"101110111",
  58686=>"000101000",
  58687=>"111101101",
  58688=>"010111100",
  58689=>"100111101",
  58690=>"000000101",
  58691=>"100001100",
  58692=>"010011101",
  58693=>"010001010",
  58694=>"100101100",
  58695=>"111100010",
  58696=>"111110111",
  58697=>"010111001",
  58698=>"100110110",
  58699=>"110000101",
  58700=>"111000100",
  58701=>"000111011",
  58702=>"101001001",
  58703=>"111111100",
  58704=>"011011111",
  58705=>"100110010",
  58706=>"110100110",
  58707=>"100010101",
  58708=>"101011011",
  58709=>"000100010",
  58710=>"110111000",
  58711=>"000011100",
  58712=>"100110000",
  58713=>"010101111",
  58714=>"000100000",
  58715=>"100001110",
  58716=>"111000011",
  58717=>"011111111",
  58718=>"000010101",
  58719=>"110110110",
  58720=>"011000110",
  58721=>"011010000",
  58722=>"110000101",
  58723=>"000110110",
  58724=>"100101100",
  58725=>"010000001",
  58726=>"110011101",
  58727=>"111001000",
  58728=>"101000101",
  58729=>"001101100",
  58730=>"010011111",
  58731=>"000100000",
  58732=>"101000000",
  58733=>"111001100",
  58734=>"010001111",
  58735=>"110000001",
  58736=>"000100110",
  58737=>"100010110",
  58738=>"011111010",
  58739=>"111100101",
  58740=>"111111110",
  58741=>"111001111",
  58742=>"011000011",
  58743=>"001111000",
  58744=>"001000000",
  58745=>"010110001",
  58746=>"101010001",
  58747=>"110100000",
  58748=>"100000001",
  58749=>"101100110",
  58750=>"111101111",
  58751=>"000100010",
  58752=>"000111110",
  58753=>"101000111",
  58754=>"011001010",
  58755=>"110110100",
  58756=>"110100101",
  58757=>"001110110",
  58758=>"101001010",
  58759=>"000111110",
  58760=>"001111000",
  58761=>"101111111",
  58762=>"111111001",
  58763=>"000011100",
  58764=>"010001010",
  58765=>"000000110",
  58766=>"101001100",
  58767=>"111100010",
  58768=>"110011011",
  58769=>"000001101",
  58770=>"100010100",
  58771=>"101000110",
  58772=>"000111011",
  58773=>"000100001",
  58774=>"001001000",
  58775=>"111101110",
  58776=>"001111111",
  58777=>"010010111",
  58778=>"101101111",
  58779=>"001000001",
  58780=>"110111100",
  58781=>"000010010",
  58782=>"000101100",
  58783=>"110111101",
  58784=>"000100111",
  58785=>"101001100",
  58786=>"001011100",
  58787=>"100101111",
  58788=>"101101000",
  58789=>"111111001",
  58790=>"111111000",
  58791=>"001100000",
  58792=>"011010101",
  58793=>"011001000",
  58794=>"011011010",
  58795=>"000101111",
  58796=>"101100111",
  58797=>"011100100",
  58798=>"111101100",
  58799=>"011111101",
  58800=>"000100101",
  58801=>"010011000",
  58802=>"010001101",
  58803=>"000000101",
  58804=>"010100011",
  58805=>"111111010",
  58806=>"111111011",
  58807=>"001011110",
  58808=>"011111110",
  58809=>"100111000",
  58810=>"101110000",
  58811=>"000001011",
  58812=>"010101111",
  58813=>"011010000",
  58814=>"111001010",
  58815=>"111001100",
  58816=>"101001010",
  58817=>"100110110",
  58818=>"000010001",
  58819=>"001011000",
  58820=>"000110011",
  58821=>"101011111",
  58822=>"110011001",
  58823=>"001011100",
  58824=>"110101100",
  58825=>"011010110",
  58826=>"000101011",
  58827=>"110101110",
  58828=>"001111111",
  58829=>"001011100",
  58830=>"001000000",
  58831=>"000101010",
  58832=>"000000111",
  58833=>"111100110",
  58834=>"011101010",
  58835=>"110101100",
  58836=>"000100111",
  58837=>"110110000",
  58838=>"001011011",
  58839=>"001100010",
  58840=>"100001000",
  58841=>"111100110",
  58842=>"011010001",
  58843=>"010000101",
  58844=>"011100001",
  58845=>"111100010",
  58846=>"111011000",
  58847=>"110000010",
  58848=>"100010100",
  58849=>"010101101",
  58850=>"011000000",
  58851=>"001111110",
  58852=>"001011001",
  58853=>"010111101",
  58854=>"001101010",
  58855=>"010111100",
  58856=>"011000010",
  58857=>"011111111",
  58858=>"001110101",
  58859=>"101001011",
  58860=>"101010110",
  58861=>"101110000",
  58862=>"101011000",
  58863=>"110100011",
  58864=>"111111100",
  58865=>"110010010",
  58866=>"001100110",
  58867=>"001110001",
  58868=>"000011000",
  58869=>"100001010",
  58870=>"110010010",
  58871=>"101101101",
  58872=>"011110010",
  58873=>"001100101",
  58874=>"011001100",
  58875=>"111100001",
  58876=>"101011111",
  58877=>"101110011",
  58878=>"011011101",
  58879=>"110100101",
  58880=>"110011000",
  58881=>"010000101",
  58882=>"001010010",
  58883=>"110100110",
  58884=>"111000101",
  58885=>"111101011",
  58886=>"011010110",
  58887=>"010011111",
  58888=>"110000010",
  58889=>"001000111",
  58890=>"001101110",
  58891=>"000000000",
  58892=>"100100111",
  58893=>"000010000",
  58894=>"011001110",
  58895=>"001001110",
  58896=>"011110000",
  58897=>"100100111",
  58898=>"011010000",
  58899=>"000111111",
  58900=>"101011110",
  58901=>"011101010",
  58902=>"101101110",
  58903=>"000000100",
  58904=>"111111111",
  58905=>"000111110",
  58906=>"000110110",
  58907=>"011101000",
  58908=>"110111110",
  58909=>"000010000",
  58910=>"100111000",
  58911=>"110010101",
  58912=>"011111100",
  58913=>"110001011",
  58914=>"011101010",
  58915=>"000001111",
  58916=>"000001110",
  58917=>"111000011",
  58918=>"100110100",
  58919=>"110110101",
  58920=>"000010000",
  58921=>"000001010",
  58922=>"110111001",
  58923=>"000100010",
  58924=>"010101001",
  58925=>"111100101",
  58926=>"100100111",
  58927=>"010010110",
  58928=>"111001111",
  58929=>"010111000",
  58930=>"001101001",
  58931=>"010111100",
  58932=>"011011110",
  58933=>"011011010",
  58934=>"010100001",
  58935=>"111101111",
  58936=>"101100010",
  58937=>"001001101",
  58938=>"101101101",
  58939=>"100011100",
  58940=>"010100011",
  58941=>"001001010",
  58942=>"110100001",
  58943=>"100000010",
  58944=>"111001101",
  58945=>"101110101",
  58946=>"011110110",
  58947=>"000011111",
  58948=>"111010111",
  58949=>"010110101",
  58950=>"101001010",
  58951=>"000011001",
  58952=>"000101000",
  58953=>"011010110",
  58954=>"100100100",
  58955=>"111011110",
  58956=>"000100001",
  58957=>"001010010",
  58958=>"110001000",
  58959=>"110000111",
  58960=>"100111111",
  58961=>"101100101",
  58962=>"001100110",
  58963=>"000100000",
  58964=>"010010100",
  58965=>"010011010",
  58966=>"101010010",
  58967=>"010000001",
  58968=>"110011111",
  58969=>"100011111",
  58970=>"111001101",
  58971=>"011011010",
  58972=>"011100101",
  58973=>"001111101",
  58974=>"100111110",
  58975=>"000011001",
  58976=>"011111111",
  58977=>"100100110",
  58978=>"101000001",
  58979=>"101001000",
  58980=>"010011011",
  58981=>"011101101",
  58982=>"110001010",
  58983=>"000000111",
  58984=>"010000110",
  58985=>"111101111",
  58986=>"111111111",
  58987=>"100100011",
  58988=>"011111100",
  58989=>"001011100",
  58990=>"101000111",
  58991=>"010000011",
  58992=>"011011011",
  58993=>"111001111",
  58994=>"101101001",
  58995=>"001001000",
  58996=>"010110110",
  58997=>"000000011",
  58998=>"101101100",
  58999=>"010110001",
  59000=>"010111100",
  59001=>"000000101",
  59002=>"111000011",
  59003=>"100001011",
  59004=>"011010011",
  59005=>"011110111",
  59006=>"000010001",
  59007=>"011111110",
  59008=>"000111011",
  59009=>"100011110",
  59010=>"001010011",
  59011=>"111011010",
  59012=>"011100011",
  59013=>"100010001",
  59014=>"000011111",
  59015=>"100011110",
  59016=>"010101111",
  59017=>"011000101",
  59018=>"111110101",
  59019=>"101000011",
  59020=>"101011111",
  59021=>"110110110",
  59022=>"000100000",
  59023=>"100101011",
  59024=>"100100001",
  59025=>"000101010",
  59026=>"111000110",
  59027=>"101100100",
  59028=>"101011110",
  59029=>"100011110",
  59030=>"111000001",
  59031=>"011101011",
  59032=>"001011010",
  59033=>"110111111",
  59034=>"010101011",
  59035=>"110000100",
  59036=>"010001100",
  59037=>"100110100",
  59038=>"011011011",
  59039=>"100011000",
  59040=>"011100101",
  59041=>"110010011",
  59042=>"100101000",
  59043=>"111011100",
  59044=>"100101001",
  59045=>"001100101",
  59046=>"001101001",
  59047=>"000000010",
  59048=>"111100110",
  59049=>"111011101",
  59050=>"110110010",
  59051=>"100011110",
  59052=>"110000101",
  59053=>"001011000",
  59054=>"100101001",
  59055=>"010011000",
  59056=>"011011010",
  59057=>"101000010",
  59058=>"110010000",
  59059=>"000010111",
  59060=>"000111101",
  59061=>"001101011",
  59062=>"001111100",
  59063=>"110110110",
  59064=>"100001001",
  59065=>"101010001",
  59066=>"101001010",
  59067=>"111000011",
  59068=>"111010000",
  59069=>"000111111",
  59070=>"000100000",
  59071=>"110000001",
  59072=>"111111011",
  59073=>"101110100",
  59074=>"110010010",
  59075=>"101010001",
  59076=>"011101110",
  59077=>"111110001",
  59078=>"011001001",
  59079=>"110011100",
  59080=>"101111000",
  59081=>"011100111",
  59082=>"010101010",
  59083=>"101110101",
  59084=>"111111011",
  59085=>"000000000",
  59086=>"001000001",
  59087=>"000011101",
  59088=>"110000100",
  59089=>"010011000",
  59090=>"111101101",
  59091=>"100011101",
  59092=>"000000110",
  59093=>"001110010",
  59094=>"001100001",
  59095=>"110100000",
  59096=>"111010100",
  59097=>"000111011",
  59098=>"110010000",
  59099=>"111000111",
  59100=>"000011101",
  59101=>"110100011",
  59102=>"001110011",
  59103=>"110101000",
  59104=>"101010110",
  59105=>"000010110",
  59106=>"101111011",
  59107=>"110010100",
  59108=>"011101110",
  59109=>"110100100",
  59110=>"101101111",
  59111=>"011111110",
  59112=>"001000101",
  59113=>"101110111",
  59114=>"100010000",
  59115=>"011010000",
  59116=>"001010011",
  59117=>"000100101",
  59118=>"110110110",
  59119=>"010100001",
  59120=>"011000000",
  59121=>"001010010",
  59122=>"111011110",
  59123=>"101111101",
  59124=>"100000111",
  59125=>"001000001",
  59126=>"001101010",
  59127=>"111101110",
  59128=>"010110000",
  59129=>"111101011",
  59130=>"111010001",
  59131=>"000101001",
  59132=>"010000100",
  59133=>"100001001",
  59134=>"001010010",
  59135=>"010000111",
  59136=>"001110101",
  59137=>"100010001",
  59138=>"001100011",
  59139=>"000101101",
  59140=>"001110101",
  59141=>"100110111",
  59142=>"100110000",
  59143=>"111111111",
  59144=>"101100000",
  59145=>"001000101",
  59146=>"100111111",
  59147=>"000011011",
  59148=>"111100001",
  59149=>"001001111",
  59150=>"000000010",
  59151=>"011101101",
  59152=>"000110001",
  59153=>"010100001",
  59154=>"101010010",
  59155=>"100001101",
  59156=>"011110011",
  59157=>"010010111",
  59158=>"010111000",
  59159=>"110011001",
  59160=>"100110101",
  59161=>"001101110",
  59162=>"010110001",
  59163=>"110101110",
  59164=>"001100110",
  59165=>"010001111",
  59166=>"110011100",
  59167=>"111010111",
  59168=>"100000011",
  59169=>"011111000",
  59170=>"001010001",
  59171=>"100011100",
  59172=>"100001100",
  59173=>"011000001",
  59174=>"110110000",
  59175=>"110100011",
  59176=>"110111001",
  59177=>"000000001",
  59178=>"011011010",
  59179=>"011010010",
  59180=>"100101001",
  59181=>"000010001",
  59182=>"100111110",
  59183=>"010010011",
  59184=>"111100001",
  59185=>"011101000",
  59186=>"101001000",
  59187=>"110011001",
  59188=>"000000000",
  59189=>"101100000",
  59190=>"010100111",
  59191=>"111101101",
  59192=>"000000011",
  59193=>"001111010",
  59194=>"101011011",
  59195=>"001000010",
  59196=>"100011010",
  59197=>"111100111",
  59198=>"110110011",
  59199=>"001111101",
  59200=>"111101101",
  59201=>"111110100",
  59202=>"111010111",
  59203=>"100100001",
  59204=>"011011000",
  59205=>"100111010",
  59206=>"100011101",
  59207=>"011111101",
  59208=>"001010001",
  59209=>"110000010",
  59210=>"100101111",
  59211=>"010010010",
  59212=>"001100111",
  59213=>"010010001",
  59214=>"011110010",
  59215=>"110110111",
  59216=>"000110000",
  59217=>"111011110",
  59218=>"001010000",
  59219=>"100000100",
  59220=>"000011110",
  59221=>"011110100",
  59222=>"001111000",
  59223=>"110111100",
  59224=>"100010001",
  59225=>"010110000",
  59226=>"011000110",
  59227=>"011101011",
  59228=>"011000000",
  59229=>"110101011",
  59230=>"101010100",
  59231=>"100011111",
  59232=>"000011011",
  59233=>"000011100",
  59234=>"101011010",
  59235=>"000010010",
  59236=>"101101011",
  59237=>"111001011",
  59238=>"100001000",
  59239=>"111111100",
  59240=>"001101100",
  59241=>"110000101",
  59242=>"111000101",
  59243=>"011000000",
  59244=>"110101110",
  59245=>"000011000",
  59246=>"111010110",
  59247=>"111110001",
  59248=>"011001001",
  59249=>"011100001",
  59250=>"001101000",
  59251=>"101000011",
  59252=>"011100110",
  59253=>"101101101",
  59254=>"011110001",
  59255=>"100000001",
  59256=>"010111001",
  59257=>"010101100",
  59258=>"110101111",
  59259=>"111011110",
  59260=>"010000000",
  59261=>"011111000",
  59262=>"101110100",
  59263=>"001111010",
  59264=>"110110101",
  59265=>"110110000",
  59266=>"110001110",
  59267=>"110000000",
  59268=>"001011000",
  59269=>"110100000",
  59270=>"001001000",
  59271=>"100011010",
  59272=>"101110111",
  59273=>"100000011",
  59274=>"100101001",
  59275=>"001101111",
  59276=>"011110010",
  59277=>"110010110",
  59278=>"000101100",
  59279=>"111011011",
  59280=>"010010100",
  59281=>"011100010",
  59282=>"010000000",
  59283=>"111011010",
  59284=>"100110110",
  59285=>"100101001",
  59286=>"100100110",
  59287=>"011100111",
  59288=>"011011001",
  59289=>"100000000",
  59290=>"010111001",
  59291=>"101001110",
  59292=>"110011000",
  59293=>"110000011",
  59294=>"000111100",
  59295=>"001011100",
  59296=>"011001101",
  59297=>"111111011",
  59298=>"111110101",
  59299=>"000101111",
  59300=>"010111010",
  59301=>"110011000",
  59302=>"011011010",
  59303=>"100000001",
  59304=>"011100001",
  59305=>"001001001",
  59306=>"110000011",
  59307=>"111100010",
  59308=>"101001010",
  59309=>"110001110",
  59310=>"001111100",
  59311=>"010110000",
  59312=>"100101010",
  59313=>"000010110",
  59314=>"011111101",
  59315=>"000011111",
  59316=>"011110000",
  59317=>"111101000",
  59318=>"110010100",
  59319=>"111001000",
  59320=>"101100101",
  59321=>"011001100",
  59322=>"001011010",
  59323=>"110010001",
  59324=>"100111001",
  59325=>"011010001",
  59326=>"011000010",
  59327=>"111111101",
  59328=>"111010100",
  59329=>"010111100",
  59330=>"111011100",
  59331=>"110101010",
  59332=>"000000110",
  59333=>"000000001",
  59334=>"011001100",
  59335=>"100010001",
  59336=>"100110000",
  59337=>"010010100",
  59338=>"100111111",
  59339=>"110001000",
  59340=>"111001101",
  59341=>"101011111",
  59342=>"010101111",
  59343=>"100111111",
  59344=>"001110111",
  59345=>"100010111",
  59346=>"000010011",
  59347=>"101010010",
  59348=>"110000101",
  59349=>"000110110",
  59350=>"001110111",
  59351=>"101111101",
  59352=>"001001010",
  59353=>"110110010",
  59354=>"001001000",
  59355=>"111001000",
  59356=>"111001010",
  59357=>"111100010",
  59358=>"110000011",
  59359=>"000001001",
  59360=>"111101111",
  59361=>"100010101",
  59362=>"001101101",
  59363=>"111101011",
  59364=>"100001000",
  59365=>"000101000",
  59366=>"011110101",
  59367=>"001010110",
  59368=>"100111111",
  59369=>"101001110",
  59370=>"000011000",
  59371=>"111111010",
  59372=>"111011111",
  59373=>"111010000",
  59374=>"010110100",
  59375=>"000010111",
  59376=>"111010010",
  59377=>"011000110",
  59378=>"100000100",
  59379=>"101011000",
  59380=>"001111001",
  59381=>"100111100",
  59382=>"001111100",
  59383=>"001110011",
  59384=>"110110011",
  59385=>"011011101",
  59386=>"111001111",
  59387=>"100000111",
  59388=>"111110000",
  59389=>"110000000",
  59390=>"100010100",
  59391=>"010000100",
  59392=>"110110101",
  59393=>"001101111",
  59394=>"011011110",
  59395=>"110101111",
  59396=>"111011111",
  59397=>"101000110",
  59398=>"000011000",
  59399=>"001010101",
  59400=>"110100111",
  59401=>"001010101",
  59402=>"010000010",
  59403=>"110110101",
  59404=>"010000000",
  59405=>"001010011",
  59406=>"100001010",
  59407=>"000010001",
  59408=>"100000101",
  59409=>"111011110",
  59410=>"101111111",
  59411=>"001100101",
  59412=>"011111010",
  59413=>"010000110",
  59414=>"000110000",
  59415=>"100101100",
  59416=>"100011000",
  59417=>"101110101",
  59418=>"010100100",
  59419=>"101110011",
  59420=>"000011010",
  59421=>"111011101",
  59422=>"111101101",
  59423=>"000101000",
  59424=>"100111111",
  59425=>"110110110",
  59426=>"111001110",
  59427=>"001110000",
  59428=>"100000001",
  59429=>"001011011",
  59430=>"111001111",
  59431=>"000010111",
  59432=>"110110100",
  59433=>"000001001",
  59434=>"111111111",
  59435=>"010111001",
  59436=>"011000000",
  59437=>"010001100",
  59438=>"110001110",
  59439=>"110100010",
  59440=>"001100101",
  59441=>"101111001",
  59442=>"100000000",
  59443=>"110000000",
  59444=>"101010110",
  59445=>"000001010",
  59446=>"111001010",
  59447=>"000010000",
  59448=>"011101000",
  59449=>"011000000",
  59450=>"111110000",
  59451=>"010101000",
  59452=>"000001110",
  59453=>"111000100",
  59454=>"111111111",
  59455=>"100101001",
  59456=>"001010001",
  59457=>"010100000",
  59458=>"001001010",
  59459=>"100100010",
  59460=>"111010111",
  59461=>"100010110",
  59462=>"100110000",
  59463=>"100000101",
  59464=>"011111100",
  59465=>"000110110",
  59466=>"001100000",
  59467=>"000000100",
  59468=>"101011101",
  59469=>"111010110",
  59470=>"111100001",
  59471=>"101010101",
  59472=>"011011111",
  59473=>"110001101",
  59474=>"010100110",
  59475=>"100111011",
  59476=>"010010110",
  59477=>"011000001",
  59478=>"100101110",
  59479=>"000001111",
  59480=>"110110100",
  59481=>"110010111",
  59482=>"011000010",
  59483=>"100011101",
  59484=>"011111100",
  59485=>"110111010",
  59486=>"101001010",
  59487=>"111011000",
  59488=>"100000001",
  59489=>"111011111",
  59490=>"000110101",
  59491=>"011000111",
  59492=>"111110010",
  59493=>"000011111",
  59494=>"101111001",
  59495=>"110111101",
  59496=>"110011111",
  59497=>"000001111",
  59498=>"101001011",
  59499=>"001100110",
  59500=>"011110011",
  59501=>"111001001",
  59502=>"011110010",
  59503=>"100111110",
  59504=>"111110101",
  59505=>"001100000",
  59506=>"110011000",
  59507=>"111100110",
  59508=>"010111100",
  59509=>"000111110",
  59510=>"000011010",
  59511=>"101111100",
  59512=>"011101010",
  59513=>"100000010",
  59514=>"111111100",
  59515=>"001111011",
  59516=>"110011110",
  59517=>"111111111",
  59518=>"001101011",
  59519=>"110010100",
  59520=>"111001100",
  59521=>"111001111",
  59522=>"101110010",
  59523=>"100001000",
  59524=>"101010100",
  59525=>"000000111",
  59526=>"011010100",
  59527=>"101101001",
  59528=>"100110010",
  59529=>"011011100",
  59530=>"100011101",
  59531=>"110100101",
  59532=>"100100101",
  59533=>"100010001",
  59534=>"000111001",
  59535=>"001011010",
  59536=>"010001100",
  59537=>"111111111",
  59538=>"011001101",
  59539=>"010101011",
  59540=>"100101011",
  59541=>"100010110",
  59542=>"001001011",
  59543=>"111101101",
  59544=>"101000101",
  59545=>"000111011",
  59546=>"110110011",
  59547=>"111110111",
  59548=>"111011100",
  59549=>"000100111",
  59550=>"011011110",
  59551=>"000101101",
  59552=>"001100001",
  59553=>"001011111",
  59554=>"010001010",
  59555=>"000110111",
  59556=>"010010100",
  59557=>"010000010",
  59558=>"001010101",
  59559=>"100010010",
  59560=>"110001000",
  59561=>"010000011",
  59562=>"000010100",
  59563=>"100001000",
  59564=>"000010000",
  59565=>"111101110",
  59566=>"000101100",
  59567=>"011001111",
  59568=>"000001010",
  59569=>"111000101",
  59570=>"110100010",
  59571=>"010110101",
  59572=>"100100111",
  59573=>"101111011",
  59574=>"111010011",
  59575=>"111000101",
  59576=>"010010100",
  59577=>"101001001",
  59578=>"110111100",
  59579=>"010100001",
  59580=>"001111101",
  59581=>"010001011",
  59582=>"001101000",
  59583=>"000010001",
  59584=>"100001100",
  59585=>"011000011",
  59586=>"011001001",
  59587=>"100010100",
  59588=>"111101111",
  59589=>"010110000",
  59590=>"000100010",
  59591=>"000101000",
  59592=>"101001111",
  59593=>"111010010",
  59594=>"110110011",
  59595=>"001011001",
  59596=>"101000001",
  59597=>"011110100",
  59598=>"010010110",
  59599=>"001010100",
  59600=>"001111100",
  59601=>"001111110",
  59602=>"100110110",
  59603=>"000111110",
  59604=>"100000011",
  59605=>"110100001",
  59606=>"100111011",
  59607=>"000100101",
  59608=>"101110011",
  59609=>"011110110",
  59610=>"111100110",
  59611=>"000101110",
  59612=>"100000001",
  59613=>"110100110",
  59614=>"011111011",
  59615=>"101011100",
  59616=>"111110011",
  59617=>"000110100",
  59618=>"110010000",
  59619=>"111110011",
  59620=>"111000111",
  59621=>"000001001",
  59622=>"100101101",
  59623=>"110000010",
  59624=>"001000110",
  59625=>"101010011",
  59626=>"100010100",
  59627=>"100000010",
  59628=>"011100000",
  59629=>"001100010",
  59630=>"010111010",
  59631=>"111100010",
  59632=>"101101100",
  59633=>"010011110",
  59634=>"110100100",
  59635=>"010000001",
  59636=>"000001001",
  59637=>"111011010",
  59638=>"010110111",
  59639=>"001011010",
  59640=>"001101001",
  59641=>"100010000",
  59642=>"001100011",
  59643=>"101111011",
  59644=>"110011100",
  59645=>"101111011",
  59646=>"100111000",
  59647=>"101111101",
  59648=>"111110001",
  59649=>"110111100",
  59650=>"100101111",
  59651=>"111110011",
  59652=>"111001110",
  59653=>"010100000",
  59654=>"000011111",
  59655=>"011100101",
  59656=>"001010001",
  59657=>"110010010",
  59658=>"010100100",
  59659=>"111110110",
  59660=>"010011000",
  59661=>"111111001",
  59662=>"010111011",
  59663=>"110010011",
  59664=>"000011100",
  59665=>"111011110",
  59666=>"111010111",
  59667=>"101001101",
  59668=>"000111101",
  59669=>"010001011",
  59670=>"000001111",
  59671=>"110010100",
  59672=>"000100101",
  59673=>"100110001",
  59674=>"111110100",
  59675=>"111001001",
  59676=>"100001110",
  59677=>"110010010",
  59678=>"101100001",
  59679=>"111100100",
  59680=>"010010101",
  59681=>"000010101",
  59682=>"011000110",
  59683=>"000001010",
  59684=>"010011100",
  59685=>"001110111",
  59686=>"100011001",
  59687=>"010100000",
  59688=>"000001000",
  59689=>"111010110",
  59690=>"100101001",
  59691=>"000000111",
  59692=>"000111100",
  59693=>"110000000",
  59694=>"000111000",
  59695=>"000010100",
  59696=>"001110101",
  59697=>"100001101",
  59698=>"010100011",
  59699=>"100010111",
  59700=>"100001100",
  59701=>"000000011",
  59702=>"011001101",
  59703=>"011101011",
  59704=>"111010011",
  59705=>"111010110",
  59706=>"111000111",
  59707=>"100011101",
  59708=>"000110101",
  59709=>"111000011",
  59710=>"100010110",
  59711=>"001101101",
  59712=>"001111000",
  59713=>"101010110",
  59714=>"001011000",
  59715=>"101101011",
  59716=>"000010000",
  59717=>"010010100",
  59718=>"110001001",
  59719=>"001011011",
  59720=>"111110100",
  59721=>"000011100",
  59722=>"000111110",
  59723=>"010100000",
  59724=>"100100000",
  59725=>"000001110",
  59726=>"101101001",
  59727=>"000010010",
  59728=>"111111001",
  59729=>"011010001",
  59730=>"101110111",
  59731=>"000010010",
  59732=>"101100101",
  59733=>"010101000",
  59734=>"101100110",
  59735=>"011011110",
  59736=>"010110001",
  59737=>"110110101",
  59738=>"000000010",
  59739=>"010011010",
  59740=>"111001000",
  59741=>"100111111",
  59742=>"010101101",
  59743=>"010101110",
  59744=>"101000011",
  59745=>"111111001",
  59746=>"001110111",
  59747=>"000101100",
  59748=>"111110100",
  59749=>"011011110",
  59750=>"001100000",
  59751=>"010100011",
  59752=>"110101001",
  59753=>"001100000",
  59754=>"110110011",
  59755=>"001111011",
  59756=>"010000010",
  59757=>"111110011",
  59758=>"001111001",
  59759=>"100110100",
  59760=>"000111000",
  59761=>"110011011",
  59762=>"001111110",
  59763=>"000111011",
  59764=>"110011101",
  59765=>"111111110",
  59766=>"101010000",
  59767=>"010110110",
  59768=>"011010111",
  59769=>"000101010",
  59770=>"101101111",
  59771=>"101010110",
  59772=>"010011101",
  59773=>"010101001",
  59774=>"100101001",
  59775=>"001010010",
  59776=>"110011100",
  59777=>"010101001",
  59778=>"001010011",
  59779=>"111100011",
  59780=>"001010101",
  59781=>"001010000",
  59782=>"000001111",
  59783=>"010111000",
  59784=>"101000100",
  59785=>"110000010",
  59786=>"101101001",
  59787=>"111011010",
  59788=>"011111110",
  59789=>"001000011",
  59790=>"100110001",
  59791=>"101000111",
  59792=>"011011001",
  59793=>"001011111",
  59794=>"101101000",
  59795=>"010000110",
  59796=>"110011100",
  59797=>"011010100",
  59798=>"111100100",
  59799=>"000010101",
  59800=>"001011010",
  59801=>"100010110",
  59802=>"010111110",
  59803=>"001111111",
  59804=>"000110010",
  59805=>"000101000",
  59806=>"110001010",
  59807=>"010101110",
  59808=>"000110101",
  59809=>"010101111",
  59810=>"001000011",
  59811=>"000001100",
  59812=>"011010011",
  59813=>"011001001",
  59814=>"100000000",
  59815=>"010011101",
  59816=>"000111011",
  59817=>"110001111",
  59818=>"110010001",
  59819=>"110100011",
  59820=>"010000000",
  59821=>"110010110",
  59822=>"100100110",
  59823=>"000101100",
  59824=>"101100100",
  59825=>"000000110",
  59826=>"100010010",
  59827=>"001010011",
  59828=>"101100000",
  59829=>"101000100",
  59830=>"001111011",
  59831=>"010100001",
  59832=>"010000010",
  59833=>"101101010",
  59834=>"101001011",
  59835=>"100011101",
  59836=>"100100100",
  59837=>"111100110",
  59838=>"010011100",
  59839=>"010100001",
  59840=>"010000001",
  59841=>"010110110",
  59842=>"100101101",
  59843=>"111010111",
  59844=>"110000010",
  59845=>"110100111",
  59846=>"001000100",
  59847=>"011011111",
  59848=>"100100100",
  59849=>"010100110",
  59850=>"011001000",
  59851=>"110111001",
  59852=>"001001100",
  59853=>"011111111",
  59854=>"110011110",
  59855=>"001001111",
  59856=>"110001111",
  59857=>"010010010",
  59858=>"001011110",
  59859=>"010000100",
  59860=>"001111100",
  59861=>"001000001",
  59862=>"000010000",
  59863=>"111100111",
  59864=>"010110000",
  59865=>"100100001",
  59866=>"000111001",
  59867=>"001010010",
  59868=>"100011001",
  59869=>"010010000",
  59870=>"001111100",
  59871=>"110010010",
  59872=>"011000010",
  59873=>"110111110",
  59874=>"111110110",
  59875=>"011111100",
  59876=>"001001101",
  59877=>"001100001",
  59878=>"100000100",
  59879=>"100111110",
  59880=>"011011100",
  59881=>"101101100",
  59882=>"000010011",
  59883=>"011010001",
  59884=>"010110000",
  59885=>"001101001",
  59886=>"110010100",
  59887=>"100100001",
  59888=>"110010000",
  59889=>"110101001",
  59890=>"011011111",
  59891=>"010011010",
  59892=>"101001011",
  59893=>"011101111",
  59894=>"010101010",
  59895=>"100010000",
  59896=>"110010110",
  59897=>"001010001",
  59898=>"000110000",
  59899=>"101000000",
  59900=>"001100111",
  59901=>"101001101",
  59902=>"010100100",
  59903=>"011011000",
  59904=>"100110111",
  59905=>"010001110",
  59906=>"100000010",
  59907=>"001011001",
  59908=>"100010100",
  59909=>"110001110",
  59910=>"111110001",
  59911=>"010100010",
  59912=>"100101000",
  59913=>"001001001",
  59914=>"011000101",
  59915=>"011001101",
  59916=>"000110000",
  59917=>"110010010",
  59918=>"100011100",
  59919=>"100110000",
  59920=>"001000111",
  59921=>"001011000",
  59922=>"011000111",
  59923=>"100010101",
  59924=>"001000001",
  59925=>"111000010",
  59926=>"001000000",
  59927=>"100101101",
  59928=>"100110000",
  59929=>"000010110",
  59930=>"011011101",
  59931=>"010000010",
  59932=>"110010001",
  59933=>"011010000",
  59934=>"111111101",
  59935=>"001011011",
  59936=>"101101000",
  59937=>"110000100",
  59938=>"010111110",
  59939=>"100011111",
  59940=>"111110111",
  59941=>"100110111",
  59942=>"101110010",
  59943=>"001010000",
  59944=>"001000011",
  59945=>"010001010",
  59946=>"000011111",
  59947=>"010100110",
  59948=>"110000100",
  59949=>"000100111",
  59950=>"111001000",
  59951=>"010110000",
  59952=>"010101010",
  59953=>"110001011",
  59954=>"110000001",
  59955=>"110101010",
  59956=>"111001111",
  59957=>"011010111",
  59958=>"100111101",
  59959=>"010110011",
  59960=>"000110011",
  59961=>"001111111",
  59962=>"101010111",
  59963=>"101101001",
  59964=>"101101000",
  59965=>"100001110",
  59966=>"000100101",
  59967=>"100001100",
  59968=>"110100010",
  59969=>"101010111",
  59970=>"101010000",
  59971=>"101010111",
  59972=>"010010101",
  59973=>"011111101",
  59974=>"101100100",
  59975=>"011011011",
  59976=>"111101110",
  59977=>"100011111",
  59978=>"001001011",
  59979=>"101111111",
  59980=>"000011101",
  59981=>"000101100",
  59982=>"001100000",
  59983=>"110001111",
  59984=>"000000110",
  59985=>"011111010",
  59986=>"100101100",
  59987=>"011000010",
  59988=>"000011101",
  59989=>"110010000",
  59990=>"011011010",
  59991=>"001100111",
  59992=>"110010011",
  59993=>"100001010",
  59994=>"010000111",
  59995=>"011011011",
  59996=>"100100101",
  59997=>"110110101",
  59998=>"000001101",
  59999=>"001101011",
  60000=>"010011001",
  60001=>"001011010",
  60002=>"010011111",
  60003=>"111100010",
  60004=>"111110111",
  60005=>"101100101",
  60006=>"101100011",
  60007=>"000110111",
  60008=>"101101001",
  60009=>"001011001",
  60010=>"111000100",
  60011=>"111110100",
  60012=>"011001110",
  60013=>"110101010",
  60014=>"110100101",
  60015=>"110111010",
  60016=>"101000111",
  60017=>"110111111",
  60018=>"000110010",
  60019=>"001010110",
  60020=>"000111111",
  60021=>"000100100",
  60022=>"000100000",
  60023=>"001110000",
  60024=>"101000101",
  60025=>"000100111",
  60026=>"000011010",
  60027=>"111101110",
  60028=>"001100101",
  60029=>"011101000",
  60030=>"101011111",
  60031=>"101101000",
  60032=>"011100010",
  60033=>"011111010",
  60034=>"000000101",
  60035=>"111111001",
  60036=>"111011100",
  60037=>"010110111",
  60038=>"001010011",
  60039=>"010011110",
  60040=>"001100100",
  60041=>"011010100",
  60042=>"101101110",
  60043=>"010001100",
  60044=>"000000011",
  60045=>"100101010",
  60046=>"010001001",
  60047=>"000010101",
  60048=>"111101100",
  60049=>"111010001",
  60050=>"110110101",
  60051=>"010010101",
  60052=>"001100001",
  60053=>"000101111",
  60054=>"011011000",
  60055=>"111010100",
  60056=>"011011011",
  60057=>"001010010",
  60058=>"101010001",
  60059=>"101001101",
  60060=>"110010001",
  60061=>"101010100",
  60062=>"100100101",
  60063=>"010001101",
  60064=>"100110011",
  60065=>"100101001",
  60066=>"010000011",
  60067=>"001011011",
  60068=>"001010101",
  60069=>"001011001",
  60070=>"110011000",
  60071=>"000100101",
  60072=>"101111011",
  60073=>"100101101",
  60074=>"101000001",
  60075=>"010110110",
  60076=>"111101111",
  60077=>"011110101",
  60078=>"000111001",
  60079=>"010111101",
  60080=>"001010000",
  60081=>"110010001",
  60082=>"010111011",
  60083=>"100101001",
  60084=>"001010011",
  60085=>"110111111",
  60086=>"100011001",
  60087=>"010000001",
  60088=>"111111101",
  60089=>"110000110",
  60090=>"001011001",
  60091=>"010000001",
  60092=>"111101111",
  60093=>"001001001",
  60094=>"001100011",
  60095=>"011011111",
  60096=>"011011001",
  60097=>"110011011",
  60098=>"010100000",
  60099=>"001010101",
  60100=>"000000110",
  60101=>"111001100",
  60102=>"110011110",
  60103=>"100110001",
  60104=>"010001001",
  60105=>"100111000",
  60106=>"110011111",
  60107=>"011101011",
  60108=>"010010010",
  60109=>"100000100",
  60110=>"101001000",
  60111=>"101101101",
  60112=>"011001001",
  60113=>"101111100",
  60114=>"010101000",
  60115=>"001100011",
  60116=>"000001001",
  60117=>"011000101",
  60118=>"101011110",
  60119=>"001110010",
  60120=>"010100001",
  60121=>"001110110",
  60122=>"110000100",
  60123=>"001111001",
  60124=>"000000010",
  60125=>"100000110",
  60126=>"100111100",
  60127=>"101111001",
  60128=>"011100011",
  60129=>"000001101",
  60130=>"101100010",
  60131=>"110000101",
  60132=>"000001100",
  60133=>"010101101",
  60134=>"111000111",
  60135=>"111100100",
  60136=>"111101001",
  60137=>"010111010",
  60138=>"100111110",
  60139=>"110010010",
  60140=>"100000111",
  60141=>"001000011",
  60142=>"111101110",
  60143=>"101111000",
  60144=>"100010000",
  60145=>"110100011",
  60146=>"111101101",
  60147=>"101100001",
  60148=>"110010100",
  60149=>"100001101",
  60150=>"011011111",
  60151=>"110100001",
  60152=>"010011110",
  60153=>"100010101",
  60154=>"010010111",
  60155=>"010011101",
  60156=>"100111111",
  60157=>"111101010",
  60158=>"101011011",
  60159=>"010000011",
  60160=>"001100001",
  60161=>"111000011",
  60162=>"101110110",
  60163=>"101101000",
  60164=>"110011010",
  60165=>"111011001",
  60166=>"000010010",
  60167=>"110101010",
  60168=>"111111101",
  60169=>"000010010",
  60170=>"001001000",
  60171=>"101001000",
  60172=>"100111110",
  60173=>"010000011",
  60174=>"110011111",
  60175=>"010111100",
  60176=>"011001101",
  60177=>"010110111",
  60178=>"011000011",
  60179=>"101101111",
  60180=>"001010100",
  60181=>"000111011",
  60182=>"100100100",
  60183=>"111000101",
  60184=>"000000001",
  60185=>"001000110",
  60186=>"101111101",
  60187=>"110100111",
  60188=>"100100100",
  60189=>"100000010",
  60190=>"110110100",
  60191=>"011110011",
  60192=>"111111011",
  60193=>"101110011",
  60194=>"001011011",
  60195=>"000111010",
  60196=>"110010110",
  60197=>"011010100",
  60198=>"101011111",
  60199=>"001101100",
  60200=>"001010010",
  60201=>"000101110",
  60202=>"111000110",
  60203=>"011100011",
  60204=>"111100011",
  60205=>"101101011",
  60206=>"111100111",
  60207=>"100101010",
  60208=>"000110010",
  60209=>"010001010",
  60210=>"101000010",
  60211=>"010000100",
  60212=>"010001001",
  60213=>"001100100",
  60214=>"110100010",
  60215=>"001100111",
  60216=>"001010100",
  60217=>"011000100",
  60218=>"110100011",
  60219=>"111101001",
  60220=>"001100011",
  60221=>"000001100",
  60222=>"111101111",
  60223=>"000111011",
  60224=>"111110101",
  60225=>"100100101",
  60226=>"010001010",
  60227=>"101111101",
  60228=>"101100101",
  60229=>"010001111",
  60230=>"000101111",
  60231=>"100001101",
  60232=>"000100101",
  60233=>"100110111",
  60234=>"000011101",
  60235=>"000000001",
  60236=>"100010011",
  60237=>"100011110",
  60238=>"010011101",
  60239=>"111001001",
  60240=>"111111100",
  60241=>"110001101",
  60242=>"010001001",
  60243=>"100110001",
  60244=>"101000110",
  60245=>"101011010",
  60246=>"011111001",
  60247=>"110001000",
  60248=>"011110111",
  60249=>"100100001",
  60250=>"100011011",
  60251=>"010100000",
  60252=>"000010111",
  60253=>"100110100",
  60254=>"010001010",
  60255=>"100111010",
  60256=>"010100100",
  60257=>"010100110",
  60258=>"110101100",
  60259=>"000011010",
  60260=>"100100011",
  60261=>"010100001",
  60262=>"111111000",
  60263=>"111000110",
  60264=>"000000000",
  60265=>"101010011",
  60266=>"111100100",
  60267=>"000100001",
  60268=>"011100001",
  60269=>"000101101",
  60270=>"000101000",
  60271=>"011001011",
  60272=>"000000000",
  60273=>"100100011",
  60274=>"100001110",
  60275=>"011010100",
  60276=>"101100001",
  60277=>"010011010",
  60278=>"010000000",
  60279=>"010100110",
  60280=>"000010111",
  60281=>"001011011",
  60282=>"001010011",
  60283=>"111011100",
  60284=>"000100011",
  60285=>"011100110",
  60286=>"010110000",
  60287=>"110010011",
  60288=>"101100100",
  60289=>"011011000",
  60290=>"111000000",
  60291=>"001100010",
  60292=>"001110010",
  60293=>"100000010",
  60294=>"010111011",
  60295=>"100001100",
  60296=>"100100010",
  60297=>"101101011",
  60298=>"101000001",
  60299=>"011100101",
  60300=>"111011001",
  60301=>"101100110",
  60302=>"110000011",
  60303=>"101100001",
  60304=>"100101111",
  60305=>"101001101",
  60306=>"100101111",
  60307=>"000001001",
  60308=>"011010010",
  60309=>"001110111",
  60310=>"001011101",
  60311=>"011011010",
  60312=>"000001001",
  60313=>"010100111",
  60314=>"011010000",
  60315=>"001101010",
  60316=>"110001101",
  60317=>"111101000",
  60318=>"101101110",
  60319=>"110110110",
  60320=>"101011001",
  60321=>"101001011",
  60322=>"100010000",
  60323=>"000111100",
  60324=>"001000110",
  60325=>"011010010",
  60326=>"001111111",
  60327=>"001100000",
  60328=>"101110000",
  60329=>"100110000",
  60330=>"001111100",
  60331=>"010111101",
  60332=>"001010111",
  60333=>"000011001",
  60334=>"110010111",
  60335=>"100010000",
  60336=>"111100101",
  60337=>"001101010",
  60338=>"100111100",
  60339=>"100110100",
  60340=>"111001101",
  60341=>"100011000",
  60342=>"011110000",
  60343=>"000110110",
  60344=>"010111000",
  60345=>"110100011",
  60346=>"110100100",
  60347=>"010101010",
  60348=>"101010010",
  60349=>"100111101",
  60350=>"100010000",
  60351=>"000110011",
  60352=>"111001110",
  60353=>"011001010",
  60354=>"011011101",
  60355=>"001100011",
  60356=>"111000100",
  60357=>"110000010",
  60358=>"000111110",
  60359=>"010110100",
  60360=>"001011100",
  60361=>"011011110",
  60362=>"000100000",
  60363=>"010100100",
  60364=>"010000001",
  60365=>"100111110",
  60366=>"110110101",
  60367=>"011000101",
  60368=>"110000110",
  60369=>"101110000",
  60370=>"000100000",
  60371=>"101010111",
  60372=>"000100010",
  60373=>"111000101",
  60374=>"010110100",
  60375=>"001100010",
  60376=>"101111110",
  60377=>"011110110",
  60378=>"011111001",
  60379=>"111111101",
  60380=>"101100110",
  60381=>"111100010",
  60382=>"101110001",
  60383=>"000100101",
  60384=>"001010001",
  60385=>"110101111",
  60386=>"111110001",
  60387=>"011001000",
  60388=>"101000000",
  60389=>"001100101",
  60390=>"100010100",
  60391=>"010111110",
  60392=>"000111100",
  60393=>"110011010",
  60394=>"101011110",
  60395=>"101100100",
  60396=>"111111010",
  60397=>"101000001",
  60398=>"110101001",
  60399=>"100011100",
  60400=>"000001010",
  60401=>"010010110",
  60402=>"000000010",
  60403=>"000101010",
  60404=>"111011001",
  60405=>"111110001",
  60406=>"110110011",
  60407=>"010011011",
  60408=>"001010100",
  60409=>"000101011",
  60410=>"101000010",
  60411=>"111101010",
  60412=>"111111111",
  60413=>"111101010",
  60414=>"111110101",
  60415=>"000011111",
  60416=>"100100101",
  60417=>"000010000",
  60418=>"111000110",
  60419=>"011110000",
  60420=>"111011001",
  60421=>"100110111",
  60422=>"100111011",
  60423=>"101010110",
  60424=>"110000110",
  60425=>"000100000",
  60426=>"110000010",
  60427=>"001110110",
  60428=>"000010101",
  60429=>"110111111",
  60430=>"000000010",
  60431=>"001011011",
  60432=>"000011010",
  60433=>"011111111",
  60434=>"110101100",
  60435=>"101001001",
  60436=>"011110011",
  60437=>"100100001",
  60438=>"110100110",
  60439=>"000001000",
  60440=>"011111101",
  60441=>"100101100",
  60442=>"111001111",
  60443=>"101011110",
  60444=>"001000011",
  60445=>"001010000",
  60446=>"011100000",
  60447=>"001101111",
  60448=>"100000100",
  60449=>"001010001",
  60450=>"110100100",
  60451=>"010010000",
  60452=>"100000001",
  60453=>"111001101",
  60454=>"011111100",
  60455=>"101001001",
  60456=>"010010001",
  60457=>"000010010",
  60458=>"100011110",
  60459=>"010100000",
  60460=>"111001110",
  60461=>"000110010",
  60462=>"101000000",
  60463=>"110101110",
  60464=>"001011001",
  60465=>"100101100",
  60466=>"101000001",
  60467=>"011010010",
  60468=>"101101011",
  60469=>"101001111",
  60470=>"000100101",
  60471=>"111010000",
  60472=>"100111001",
  60473=>"101001110",
  60474=>"001000011",
  60475=>"011010001",
  60476=>"100100111",
  60477=>"001010010",
  60478=>"110011101",
  60479=>"011001000",
  60480=>"111101110",
  60481=>"001101111",
  60482=>"011000001",
  60483=>"100111101",
  60484=>"001000010",
  60485=>"101011010",
  60486=>"111111011",
  60487=>"001001110",
  60488=>"111011000",
  60489=>"110010011",
  60490=>"110110111",
  60491=>"001101000",
  60492=>"011010110",
  60493=>"111011100",
  60494=>"100111001",
  60495=>"010111000",
  60496=>"110011111",
  60497=>"000110011",
  60498=>"110101110",
  60499=>"001100101",
  60500=>"101111111",
  60501=>"100010000",
  60502=>"100001111",
  60503=>"000000100",
  60504=>"110110110",
  60505=>"001010010",
  60506=>"110101100",
  60507=>"000111100",
  60508=>"001001111",
  60509=>"110011010",
  60510=>"110011110",
  60511=>"001011110",
  60512=>"111011111",
  60513=>"000111001",
  60514=>"110100101",
  60515=>"001010001",
  60516=>"010100100",
  60517=>"111101001",
  60518=>"111001011",
  60519=>"101001011",
  60520=>"010111100",
  60521=>"000010110",
  60522=>"000000000",
  60523=>"010110001",
  60524=>"001011101",
  60525=>"111001111",
  60526=>"110101101",
  60527=>"000110000",
  60528=>"010110000",
  60529=>"010110100",
  60530=>"100101100",
  60531=>"000110010",
  60532=>"000100101",
  60533=>"000011110",
  60534=>"110110010",
  60535=>"011110110",
  60536=>"101101011",
  60537=>"100010110",
  60538=>"110101111",
  60539=>"100100101",
  60540=>"011110110",
  60541=>"001111101",
  60542=>"101010111",
  60543=>"000101100",
  60544=>"111101111",
  60545=>"010000100",
  60546=>"010110011",
  60547=>"111101101",
  60548=>"000011110",
  60549=>"011011011",
  60550=>"111110100",
  60551=>"001110011",
  60552=>"011011000",
  60553=>"100001110",
  60554=>"101101000",
  60555=>"010001111",
  60556=>"111100001",
  60557=>"100011110",
  60558=>"001111011",
  60559=>"111000000",
  60560=>"000000000",
  60561=>"100000001",
  60562=>"101100111",
  60563=>"011000000",
  60564=>"001101100",
  60565=>"111100001",
  60566=>"110000010",
  60567=>"111010101",
  60568=>"111010101",
  60569=>"011110001",
  60570=>"111100101",
  60571=>"100011010",
  60572=>"010000101",
  60573=>"000011110",
  60574=>"001001001",
  60575=>"001111101",
  60576=>"000101000",
  60577=>"111110110",
  60578=>"101100111",
  60579=>"010010010",
  60580=>"111010110",
  60581=>"100010101",
  60582=>"011010000",
  60583=>"100110111",
  60584=>"011110100",
  60585=>"001100000",
  60586=>"110000100",
  60587=>"111110000",
  60588=>"100100001",
  60589=>"001110001",
  60590=>"010110001",
  60591=>"010100111",
  60592=>"010100100",
  60593=>"101111101",
  60594=>"110101100",
  60595=>"011001100",
  60596=>"110110101",
  60597=>"010001000",
  60598=>"100110111",
  60599=>"000100111",
  60600=>"000101100",
  60601=>"100011010",
  60602=>"111000111",
  60603=>"110111101",
  60604=>"110000101",
  60605=>"010000011",
  60606=>"011010010",
  60607=>"011100000",
  60608=>"111101110",
  60609=>"011101000",
  60610=>"000001100",
  60611=>"101010010",
  60612=>"001001011",
  60613=>"101011011",
  60614=>"110010101",
  60615=>"101010001",
  60616=>"111101100",
  60617=>"001101101",
  60618=>"111111101",
  60619=>"011110001",
  60620=>"011000010",
  60621=>"011101000",
  60622=>"001100101",
  60623=>"001111001",
  60624=>"001100001",
  60625=>"010110010",
  60626=>"100011100",
  60627=>"111101000",
  60628=>"110110100",
  60629=>"011000101",
  60630=>"100001110",
  60631=>"101010110",
  60632=>"100111100",
  60633=>"111001000",
  60634=>"111110010",
  60635=>"001001010",
  60636=>"010000000",
  60637=>"001011000",
  60638=>"011010000",
  60639=>"000111011",
  60640=>"000111100",
  60641=>"000110110",
  60642=>"111001000",
  60643=>"100110011",
  60644=>"110011001",
  60645=>"101010111",
  60646=>"101100010",
  60647=>"000001000",
  60648=>"111111011",
  60649=>"010100000",
  60650=>"100101101",
  60651=>"010100000",
  60652=>"110011110",
  60653=>"000111010",
  60654=>"100111001",
  60655=>"000001101",
  60656=>"100100011",
  60657=>"011010001",
  60658=>"000001011",
  60659=>"110011111",
  60660=>"101101000",
  60661=>"010011000",
  60662=>"110100101",
  60663=>"000000000",
  60664=>"101011111",
  60665=>"111100010",
  60666=>"010100011",
  60667=>"100011000",
  60668=>"111000111",
  60669=>"110101000",
  60670=>"011110010",
  60671=>"000011011",
  60672=>"001111011",
  60673=>"000111010",
  60674=>"011010101",
  60675=>"001011111",
  60676=>"111101001",
  60677=>"010001011",
  60678=>"001010111",
  60679=>"101110001",
  60680=>"010110100",
  60681=>"100101100",
  60682=>"101110000",
  60683=>"110100110",
  60684=>"111011100",
  60685=>"010111100",
  60686=>"111010100",
  60687=>"000110000",
  60688=>"010100001",
  60689=>"110000100",
  60690=>"000101101",
  60691=>"111111100",
  60692=>"110111010",
  60693=>"010001111",
  60694=>"001010101",
  60695=>"101101110",
  60696=>"100101011",
  60697=>"111000001",
  60698=>"010110000",
  60699=>"000000111",
  60700=>"000001010",
  60701=>"000000001",
  60702=>"111111101",
  60703=>"000111001",
  60704=>"000001010",
  60705=>"110100101",
  60706=>"101100000",
  60707=>"000000111",
  60708=>"101011111",
  60709=>"111111110",
  60710=>"000010001",
  60711=>"100110000",
  60712=>"011110100",
  60713=>"110110000",
  60714=>"010011010",
  60715=>"101000101",
  60716=>"000010110",
  60717=>"010000101",
  60718=>"010110111",
  60719=>"010010011",
  60720=>"011010101",
  60721=>"100001110",
  60722=>"010011010",
  60723=>"010000111",
  60724=>"100000010",
  60725=>"100011010",
  60726=>"110110100",
  60727=>"110100011",
  60728=>"010110110",
  60729=>"101001011",
  60730=>"101101001",
  60731=>"101000100",
  60732=>"000010110",
  60733=>"000110111",
  60734=>"011001100",
  60735=>"011011000",
  60736=>"010100100",
  60737=>"010000101",
  60738=>"101001000",
  60739=>"101010001",
  60740=>"100100110",
  60741=>"111101111",
  60742=>"011100011",
  60743=>"100101000",
  60744=>"011111010",
  60745=>"110101100",
  60746=>"101101100",
  60747=>"000001110",
  60748=>"000000010",
  60749=>"000111000",
  60750=>"001011111",
  60751=>"011101100",
  60752=>"011111010",
  60753=>"000111010",
  60754=>"101011001",
  60755=>"000011001",
  60756=>"101111001",
  60757=>"000001000",
  60758=>"011000001",
  60759=>"011100100",
  60760=>"010111001",
  60761=>"011110111",
  60762=>"110001010",
  60763=>"100011010",
  60764=>"101100011",
  60765=>"001000011",
  60766=>"111101001",
  60767=>"100010101",
  60768=>"010100000",
  60769=>"110001100",
  60770=>"001000011",
  60771=>"101111100",
  60772=>"111010101",
  60773=>"110111111",
  60774=>"101110001",
  60775=>"000000111",
  60776=>"001101110",
  60777=>"011011111",
  60778=>"110100001",
  60779=>"000001101",
  60780=>"111101100",
  60781=>"101101111",
  60782=>"010100001",
  60783=>"101011010",
  60784=>"000111101",
  60785=>"110110110",
  60786=>"011111101",
  60787=>"100010110",
  60788=>"010101101",
  60789=>"110011111",
  60790=>"101011001",
  60791=>"111100101",
  60792=>"101001000",
  60793=>"100000101",
  60794=>"111111100",
  60795=>"000011000",
  60796=>"111001001",
  60797=>"000011000",
  60798=>"001001001",
  60799=>"000001100",
  60800=>"000010000",
  60801=>"000000011",
  60802=>"001100100",
  60803=>"101111011",
  60804=>"101111001",
  60805=>"111011001",
  60806=>"111001100",
  60807=>"100011010",
  60808=>"101010101",
  60809=>"001010100",
  60810=>"010011100",
  60811=>"000000001",
  60812=>"011100100",
  60813=>"110001111",
  60814=>"101000111",
  60815=>"111011001",
  60816=>"000000000",
  60817=>"011011100",
  60818=>"101010000",
  60819=>"001011011",
  60820=>"110100101",
  60821=>"110010000",
  60822=>"000111010",
  60823=>"000011111",
  60824=>"101111100",
  60825=>"010010101",
  60826=>"011001100",
  60827=>"101011001",
  60828=>"111010001",
  60829=>"010011100",
  60830=>"111001111",
  60831=>"111001111",
  60832=>"111010001",
  60833=>"001011011",
  60834=>"110011110",
  60835=>"111110010",
  60836=>"011000000",
  60837=>"000000000",
  60838=>"010000110",
  60839=>"001101011",
  60840=>"100101001",
  60841=>"110111111",
  60842=>"101011101",
  60843=>"000001101",
  60844=>"000010000",
  60845=>"000011110",
  60846=>"111100000",
  60847=>"100000100",
  60848=>"011111101",
  60849=>"011010000",
  60850=>"000010001",
  60851=>"101001011",
  60852=>"001111000",
  60853=>"101101101",
  60854=>"010110101",
  60855=>"000101100",
  60856=>"110110010",
  60857=>"011111001",
  60858=>"001111010",
  60859=>"100111011",
  60860=>"100101100",
  60861=>"110011011",
  60862=>"001111111",
  60863=>"110000111",
  60864=>"001101000",
  60865=>"100100010",
  60866=>"011101110",
  60867=>"011100110",
  60868=>"110010010",
  60869=>"110110000",
  60870=>"001000001",
  60871=>"111110010",
  60872=>"001011010",
  60873=>"101010011",
  60874=>"110000111",
  60875=>"011010010",
  60876=>"111000101",
  60877=>"010000110",
  60878=>"110100001",
  60879=>"000001001",
  60880=>"101011010",
  60881=>"000100010",
  60882=>"001110000",
  60883=>"011011110",
  60884=>"100101001",
  60885=>"111011011",
  60886=>"111001101",
  60887=>"110110011",
  60888=>"110011110",
  60889=>"111101011",
  60890=>"110000001",
  60891=>"100001110",
  60892=>"011101110",
  60893=>"001010000",
  60894=>"100000011",
  60895=>"001010000",
  60896=>"110101100",
  60897=>"111101100",
  60898=>"011111000",
  60899=>"001101111",
  60900=>"001101011",
  60901=>"011010011",
  60902=>"001100100",
  60903=>"010101111",
  60904=>"010010111",
  60905=>"100110110",
  60906=>"110110010",
  60907=>"100011101",
  60908=>"110001101",
  60909=>"001001101",
  60910=>"010001111",
  60911=>"001101010",
  60912=>"010001111",
  60913=>"100101111",
  60914=>"100101110",
  60915=>"001001011",
  60916=>"100111110",
  60917=>"111001011",
  60918=>"001000000",
  60919=>"010111001",
  60920=>"000001010",
  60921=>"111100110",
  60922=>"101000011",
  60923=>"101001101",
  60924=>"000100000",
  60925=>"011101100",
  60926=>"001101100",
  60927=>"100001111",
  60928=>"110000001",
  60929=>"011000000",
  60930=>"011010110",
  60931=>"011011010",
  60932=>"000010010",
  60933=>"111110111",
  60934=>"101010010",
  60935=>"110000001",
  60936=>"000000010",
  60937=>"110110010",
  60938=>"101001001",
  60939=>"011101000",
  60940=>"111111110",
  60941=>"000000101",
  60942=>"001010101",
  60943=>"111101111",
  60944=>"110110010",
  60945=>"100110001",
  60946=>"110011000",
  60947=>"010101100",
  60948=>"101101111",
  60949=>"001101100",
  60950=>"111110100",
  60951=>"001000111",
  60952=>"111111101",
  60953=>"000101111",
  60954=>"010111101",
  60955=>"001100000",
  60956=>"011000010",
  60957=>"001001111",
  60958=>"010011111",
  60959=>"011011011",
  60960=>"000101111",
  60961=>"101100110",
  60962=>"001000010",
  60963=>"110000101",
  60964=>"010110111",
  60965=>"110101001",
  60966=>"111111001",
  60967=>"001001001",
  60968=>"100001110",
  60969=>"001000100",
  60970=>"101011010",
  60971=>"100011101",
  60972=>"111100000",
  60973=>"100011100",
  60974=>"100100110",
  60975=>"011001011",
  60976=>"000110110",
  60977=>"110101111",
  60978=>"010101011",
  60979=>"111110111",
  60980=>"101010001",
  60981=>"101011101",
  60982=>"100101010",
  60983=>"000011000",
  60984=>"111110010",
  60985=>"110101111",
  60986=>"000000110",
  60987=>"110011000",
  60988=>"010011100",
  60989=>"010010001",
  60990=>"001111000",
  60991=>"100000010",
  60992=>"001010010",
  60993=>"101010010",
  60994=>"110000111",
  60995=>"111011001",
  60996=>"111001110",
  60997=>"001000101",
  60998=>"101110001",
  60999=>"000111011",
  61000=>"111111101",
  61001=>"110110001",
  61002=>"010010001",
  61003=>"100100011",
  61004=>"010101000",
  61005=>"000010010",
  61006=>"101011111",
  61007=>"111100100",
  61008=>"101010011",
  61009=>"001011101",
  61010=>"000010010",
  61011=>"000100011",
  61012=>"101000101",
  61013=>"100010000",
  61014=>"111010000",
  61015=>"110101110",
  61016=>"101101100",
  61017=>"101010101",
  61018=>"111110100",
  61019=>"101110000",
  61020=>"001101101",
  61021=>"110010100",
  61022=>"111011010",
  61023=>"000101101",
  61024=>"011001000",
  61025=>"111011001",
  61026=>"001011000",
  61027=>"110101110",
  61028=>"010110011",
  61029=>"001000011",
  61030=>"100110011",
  61031=>"100111000",
  61032=>"011101100",
  61033=>"010110000",
  61034=>"001000001",
  61035=>"100001100",
  61036=>"000000001",
  61037=>"110111011",
  61038=>"111010010",
  61039=>"011000000",
  61040=>"001000111",
  61041=>"001011001",
  61042=>"011100011",
  61043=>"010001111",
  61044=>"101111111",
  61045=>"011010101",
  61046=>"010100100",
  61047=>"000001110",
  61048=>"111010100",
  61049=>"011000011",
  61050=>"111001011",
  61051=>"101100000",
  61052=>"100010000",
  61053=>"000000111",
  61054=>"000000100",
  61055=>"111111011",
  61056=>"111111110",
  61057=>"001000110",
  61058=>"111001100",
  61059=>"110111011",
  61060=>"100000110",
  61061=>"011100001",
  61062=>"100111001",
  61063=>"110011111",
  61064=>"111111100",
  61065=>"001011010",
  61066=>"111111110",
  61067=>"001000001",
  61068=>"101111111",
  61069=>"110011100",
  61070=>"001011000",
  61071=>"000100100",
  61072=>"100001001",
  61073=>"000110001",
  61074=>"001001000",
  61075=>"001111001",
  61076=>"000110100",
  61077=>"010111000",
  61078=>"101110011",
  61079=>"011010010",
  61080=>"110110010",
  61081=>"000011000",
  61082=>"011010000",
  61083=>"001011110",
  61084=>"000100010",
  61085=>"011101101",
  61086=>"101111101",
  61087=>"100100100",
  61088=>"001001001",
  61089=>"111000011",
  61090=>"111001000",
  61091=>"000111100",
  61092=>"000101101",
  61093=>"111001001",
  61094=>"010000111",
  61095=>"000010110",
  61096=>"111011101",
  61097=>"000010110",
  61098=>"100111101",
  61099=>"000100111",
  61100=>"110001100",
  61101=>"101010110",
  61102=>"001110111",
  61103=>"010001000",
  61104=>"100101111",
  61105=>"100110100",
  61106=>"000101000",
  61107=>"011000100",
  61108=>"101111010",
  61109=>"010110101",
  61110=>"110111011",
  61111=>"010001000",
  61112=>"101110000",
  61113=>"100110111",
  61114=>"001001111",
  61115=>"011100001",
  61116=>"000010001",
  61117=>"001011100",
  61118=>"001011101",
  61119=>"011011011",
  61120=>"110111101",
  61121=>"000110111",
  61122=>"110110100",
  61123=>"001100010",
  61124=>"111001111",
  61125=>"111100000",
  61126=>"010001001",
  61127=>"001100110",
  61128=>"000011110",
  61129=>"110100100",
  61130=>"110001001",
  61131=>"010100000",
  61132=>"010011101",
  61133=>"000100010",
  61134=>"110100111",
  61135=>"000101100",
  61136=>"001011110",
  61137=>"101000111",
  61138=>"111111101",
  61139=>"000000111",
  61140=>"010000010",
  61141=>"110011110",
  61142=>"110100001",
  61143=>"010000101",
  61144=>"000101110",
  61145=>"100101011",
  61146=>"010001101",
  61147=>"000100000",
  61148=>"001110100",
  61149=>"110001100",
  61150=>"001000101",
  61151=>"001110101",
  61152=>"000100011",
  61153=>"100000001",
  61154=>"001110111",
  61155=>"100111010",
  61156=>"011111110",
  61157=>"011101000",
  61158=>"110110100",
  61159=>"001011010",
  61160=>"000010100",
  61161=>"111110100",
  61162=>"010001010",
  61163=>"101000111",
  61164=>"100010101",
  61165=>"111111111",
  61166=>"001111001",
  61167=>"000000001",
  61168=>"000111000",
  61169=>"111101010",
  61170=>"100111110",
  61171=>"000001010",
  61172=>"000010100",
  61173=>"010110110",
  61174=>"111111010",
  61175=>"001000110",
  61176=>"100001000",
  61177=>"010001000",
  61178=>"100100111",
  61179=>"000001111",
  61180=>"011111101",
  61181=>"001100000",
  61182=>"100101000",
  61183=>"011100000",
  61184=>"100110011",
  61185=>"010111001",
  61186=>"101000011",
  61187=>"000011100",
  61188=>"111001110",
  61189=>"011011110",
  61190=>"010000010",
  61191=>"101000000",
  61192=>"000010011",
  61193=>"001011011",
  61194=>"101001101",
  61195=>"000100101",
  61196=>"100111010",
  61197=>"000010100",
  61198=>"111001110",
  61199=>"110110001",
  61200=>"110000000",
  61201=>"100000000",
  61202=>"110111101",
  61203=>"000100100",
  61204=>"010000010",
  61205=>"010101101",
  61206=>"111010000",
  61207=>"000110011",
  61208=>"000010001",
  61209=>"101011001",
  61210=>"111111000",
  61211=>"111010010",
  61212=>"100001101",
  61213=>"011001001",
  61214=>"111100110",
  61215=>"101110010",
  61216=>"011110101",
  61217=>"110001010",
  61218=>"110100100",
  61219=>"100001100",
  61220=>"011001010",
  61221=>"001100100",
  61222=>"000010000",
  61223=>"111001101",
  61224=>"110101111",
  61225=>"111100111",
  61226=>"111011100",
  61227=>"111010110",
  61228=>"010111010",
  61229=>"001010101",
  61230=>"000010100",
  61231=>"111010010",
  61232=>"100111111",
  61233=>"110011100",
  61234=>"010111111",
  61235=>"100111110",
  61236=>"011000110",
  61237=>"000000110",
  61238=>"110110110",
  61239=>"011111000",
  61240=>"101101110",
  61241=>"011011000",
  61242=>"100111001",
  61243=>"011010101",
  61244=>"100111111",
  61245=>"101110001",
  61246=>"000100101",
  61247=>"100010111",
  61248=>"011111110",
  61249=>"110110011",
  61250=>"111000010",
  61251=>"111000010",
  61252=>"011110110",
  61253=>"011100100",
  61254=>"111111001",
  61255=>"001111000",
  61256=>"010011001",
  61257=>"001110100",
  61258=>"110011001",
  61259=>"110000001",
  61260=>"011100101",
  61261=>"010101111",
  61262=>"110110000",
  61263=>"010110110",
  61264=>"110110111",
  61265=>"100010100",
  61266=>"001000000",
  61267=>"101111011",
  61268=>"110001100",
  61269=>"010000111",
  61270=>"101101101",
  61271=>"011100111",
  61272=>"010011010",
  61273=>"110100001",
  61274=>"100001100",
  61275=>"000101011",
  61276=>"111000011",
  61277=>"001010000",
  61278=>"101001000",
  61279=>"000111011",
  61280=>"011101101",
  61281=>"111001110",
  61282=>"011110101",
  61283=>"001011101",
  61284=>"110111010",
  61285=>"101000110",
  61286=>"101010010",
  61287=>"110100111",
  61288=>"110100011",
  61289=>"011110110",
  61290=>"011011001",
  61291=>"110000000",
  61292=>"100100000",
  61293=>"110111101",
  61294=>"000001010",
  61295=>"100001010",
  61296=>"101011000",
  61297=>"101010010",
  61298=>"110111011",
  61299=>"000111010",
  61300=>"011110000",
  61301=>"000111111",
  61302=>"000000010",
  61303=>"101000000",
  61304=>"111100010",
  61305=>"111101001",
  61306=>"010000011",
  61307=>"010100110",
  61308=>"000011010",
  61309=>"000000111",
  61310=>"000110001",
  61311=>"011000011",
  61312=>"001010111",
  61313=>"000011010",
  61314=>"111110101",
  61315=>"110111100",
  61316=>"001100000",
  61317=>"011011101",
  61318=>"101000110",
  61319=>"000111110",
  61320=>"101001011",
  61321=>"000110111",
  61322=>"011001111",
  61323=>"100000001",
  61324=>"100011000",
  61325=>"100000100",
  61326=>"101010100",
  61327=>"000100011",
  61328=>"000010101",
  61329=>"101101101",
  61330=>"001100000",
  61331=>"101001010",
  61332=>"001011011",
  61333=>"100100101",
  61334=>"101110001",
  61335=>"100110000",
  61336=>"000111001",
  61337=>"101010000",
  61338=>"010111100",
  61339=>"001001101",
  61340=>"100100101",
  61341=>"000000111",
  61342=>"111000010",
  61343=>"001100000",
  61344=>"011011100",
  61345=>"101001000",
  61346=>"010111100",
  61347=>"110010100",
  61348=>"010100011",
  61349=>"100111110",
  61350=>"101000100",
  61351=>"100110111",
  61352=>"011010001",
  61353=>"000111100",
  61354=>"111001101",
  61355=>"010001000",
  61356=>"011101011",
  61357=>"011010011",
  61358=>"001011011",
  61359=>"110011110",
  61360=>"100001000",
  61361=>"011000100",
  61362=>"101001011",
  61363=>"010000011",
  61364=>"010001000",
  61365=>"100111100",
  61366=>"011101011",
  61367=>"001000111",
  61368=>"000010000",
  61369=>"000101111",
  61370=>"011111100",
  61371=>"110100111",
  61372=>"000011001",
  61373=>"111010100",
  61374=>"100100110",
  61375=>"111100000",
  61376=>"110000111",
  61377=>"000000110",
  61378=>"011110101",
  61379=>"110011111",
  61380=>"000011110",
  61381=>"110001000",
  61382=>"010000001",
  61383=>"110100011",
  61384=>"100110110",
  61385=>"111000001",
  61386=>"101001010",
  61387=>"111011011",
  61388=>"111101111",
  61389=>"000110101",
  61390=>"111100001",
  61391=>"010101101",
  61392=>"100100000",
  61393=>"000111010",
  61394=>"011001110",
  61395=>"100100001",
  61396=>"001101101",
  61397=>"100010110",
  61398=>"010000100",
  61399=>"101100001",
  61400=>"001000000",
  61401=>"111100011",
  61402=>"001001110",
  61403=>"101001001",
  61404=>"010001000",
  61405=>"101001000",
  61406=>"011000010",
  61407=>"100111110",
  61408=>"100111011",
  61409=>"011111000",
  61410=>"000100101",
  61411=>"110010000",
  61412=>"111101111",
  61413=>"011101100",
  61414=>"110000111",
  61415=>"000110111",
  61416=>"000100010",
  61417=>"000000011",
  61418=>"111011111",
  61419=>"100110100",
  61420=>"110010111",
  61421=>"100101010",
  61422=>"011100011",
  61423=>"010111111",
  61424=>"001000001",
  61425=>"011110111",
  61426=>"111110110",
  61427=>"101110011",
  61428=>"001000111",
  61429=>"001010010",
  61430=>"011100111",
  61431=>"100001111",
  61432=>"100100100",
  61433=>"100001000",
  61434=>"010110011",
  61435=>"101111110",
  61436=>"010111100",
  61437=>"100101110",
  61438=>"111100011",
  61439=>"010101101",
  61440=>"101111000",
  61441=>"100001110",
  61442=>"100000110",
  61443=>"111011011",
  61444=>"010110110",
  61445=>"000100011",
  61446=>"000110001",
  61447=>"000000001",
  61448=>"110001000",
  61449=>"100010100",
  61450=>"111100000",
  61451=>"010100001",
  61452=>"010001111",
  61453=>"000001110",
  61454=>"010010011",
  61455=>"111101110",
  61456=>"101011011",
  61457=>"011010100",
  61458=>"110001001",
  61459=>"101111001",
  61460=>"001010110",
  61461=>"011100111",
  61462=>"110110010",
  61463=>"010101101",
  61464=>"110000010",
  61465=>"100001011",
  61466=>"111111111",
  61467=>"101011011",
  61468=>"101100010",
  61469=>"100111011",
  61470=>"011101101",
  61471=>"111000001",
  61472=>"000100110",
  61473=>"101101001",
  61474=>"100010000",
  61475=>"101111010",
  61476=>"001101110",
  61477=>"010010100",
  61478=>"110001001",
  61479=>"000011001",
  61480=>"110000011",
  61481=>"101110001",
  61482=>"001111111",
  61483=>"111011100",
  61484=>"101101101",
  61485=>"010100000",
  61486=>"001011001",
  61487=>"111110100",
  61488=>"001000011",
  61489=>"101111100",
  61490=>"001001100",
  61491=>"011101001",
  61492=>"001100110",
  61493=>"000110000",
  61494=>"100000110",
  61495=>"100111111",
  61496=>"000101001",
  61497=>"110110011",
  61498=>"010101101",
  61499=>"011101000",
  61500=>"101110110",
  61501=>"001101110",
  61502=>"001010101",
  61503=>"000101000",
  61504=>"100000011",
  61505=>"000010000",
  61506=>"111000110",
  61507=>"001111101",
  61508=>"001100101",
  61509=>"111001101",
  61510=>"010110011",
  61511=>"001011111",
  61512=>"111101100",
  61513=>"000001110",
  61514=>"100001101",
  61515=>"101110110",
  61516=>"000010001",
  61517=>"001111010",
  61518=>"011011101",
  61519=>"100001010",
  61520=>"101001100",
  61521=>"100111011",
  61522=>"001100001",
  61523=>"100001111",
  61524=>"000010001",
  61525=>"011111111",
  61526=>"110011111",
  61527=>"000011001",
  61528=>"110001111",
  61529=>"111110101",
  61530=>"011000001",
  61531=>"010001111",
  61532=>"111101000",
  61533=>"011100001",
  61534=>"110111110",
  61535=>"000000000",
  61536=>"111000010",
  61537=>"101010000",
  61538=>"011101101",
  61539=>"110001100",
  61540=>"011110001",
  61541=>"001010011",
  61542=>"101100111",
  61543=>"110010010",
  61544=>"010101111",
  61545=>"111010001",
  61546=>"100100001",
  61547=>"100100100",
  61548=>"000100101",
  61549=>"000100010",
  61550=>"001011100",
  61551=>"101100101",
  61552=>"100101011",
  61553=>"101011111",
  61554=>"111101100",
  61555=>"110110101",
  61556=>"001011010",
  61557=>"011100001",
  61558=>"011010100",
  61559=>"000011101",
  61560=>"111111101",
  61561=>"000110001",
  61562=>"110101000",
  61563=>"001010001",
  61564=>"100101010",
  61565=>"000010111",
  61566=>"001100011",
  61567=>"010000000",
  61568=>"000001110",
  61569=>"100100111",
  61570=>"000011000",
  61571=>"010111011",
  61572=>"110001011",
  61573=>"101011111",
  61574=>"001010000",
  61575=>"111110011",
  61576=>"100101011",
  61577=>"010101110",
  61578=>"100101111",
  61579=>"000011111",
  61580=>"111101011",
  61581=>"100000001",
  61582=>"000101011",
  61583=>"000000000",
  61584=>"100000111",
  61585=>"000110001",
  61586=>"100000001",
  61587=>"010011110",
  61588=>"000110101",
  61589=>"011100011",
  61590=>"000000101",
  61591=>"110111111",
  61592=>"001111110",
  61593=>"011101000",
  61594=>"001010110",
  61595=>"101110101",
  61596=>"000110011",
  61597=>"010010111",
  61598=>"000011110",
  61599=>"011110001",
  61600=>"111010010",
  61601=>"010011101",
  61602=>"001100000",
  61603=>"101110011",
  61604=>"000100101",
  61605=>"101111100",
  61606=>"000101000",
  61607=>"000110001",
  61608=>"101111000",
  61609=>"000011110",
  61610=>"000010000",
  61611=>"001011001",
  61612=>"110110101",
  61613=>"101011110",
  61614=>"001001101",
  61615=>"101100100",
  61616=>"000101100",
  61617=>"000110101",
  61618=>"100010011",
  61619=>"001001111",
  61620=>"100111011",
  61621=>"011011001",
  61622=>"001010101",
  61623=>"100111111",
  61624=>"110010011",
  61625=>"101000111",
  61626=>"101101000",
  61627=>"100101101",
  61628=>"000100111",
  61629=>"101000010",
  61630=>"001111001",
  61631=>"100001101",
  61632=>"001011110",
  61633=>"100000100",
  61634=>"001000101",
  61635=>"011011111",
  61636=>"100000001",
  61637=>"000111111",
  61638=>"110000011",
  61639=>"101100101",
  61640=>"011101011",
  61641=>"111100000",
  61642=>"000001110",
  61643=>"000111111",
  61644=>"011111000",
  61645=>"010010111",
  61646=>"110111101",
  61647=>"110000101",
  61648=>"100101010",
  61649=>"110001111",
  61650=>"011001011",
  61651=>"011010011",
  61652=>"000111110",
  61653=>"100011111",
  61654=>"100100110",
  61655=>"111001110",
  61656=>"110001010",
  61657=>"011100100",
  61658=>"011001100",
  61659=>"111011010",
  61660=>"011011001",
  61661=>"001101100",
  61662=>"110100001",
  61663=>"100100110",
  61664=>"000011010",
  61665=>"111100001",
  61666=>"010100001",
  61667=>"011101101",
  61668=>"100001001",
  61669=>"000000000",
  61670=>"110000000",
  61671=>"000101111",
  61672=>"111100101",
  61673=>"111001111",
  61674=>"100001111",
  61675=>"011000000",
  61676=>"010101100",
  61677=>"100000101",
  61678=>"011000101",
  61679=>"011111010",
  61680=>"011011101",
  61681=>"100000110",
  61682=>"001110100",
  61683=>"001100011",
  61684=>"011000011",
  61685=>"101100000",
  61686=>"101110001",
  61687=>"000010110",
  61688=>"001110010",
  61689=>"001011110",
  61690=>"000101010",
  61691=>"000100100",
  61692=>"111011101",
  61693=>"111100010",
  61694=>"111100010",
  61695=>"111100110",
  61696=>"000010110",
  61697=>"110101101",
  61698=>"111110011",
  61699=>"111111011",
  61700=>"000101000",
  61701=>"101100000",
  61702=>"111001101",
  61703=>"100001100",
  61704=>"100001111",
  61705=>"000000110",
  61706=>"100001100",
  61707=>"111101001",
  61708=>"101000100",
  61709=>"001000100",
  61710=>"001110000",
  61711=>"101101110",
  61712=>"111010100",
  61713=>"111110101",
  61714=>"110010100",
  61715=>"110101010",
  61716=>"100000001",
  61717=>"011010011",
  61718=>"001101110",
  61719=>"101100000",
  61720=>"001000000",
  61721=>"011000101",
  61722=>"101111011",
  61723=>"011011100",
  61724=>"001000111",
  61725=>"101011111",
  61726=>"111110100",
  61727=>"111101010",
  61728=>"101100000",
  61729=>"001100111",
  61730=>"011101100",
  61731=>"011010000",
  61732=>"001000100",
  61733=>"110110010",
  61734=>"000000011",
  61735=>"011100101",
  61736=>"101000000",
  61737=>"011110000",
  61738=>"101011001",
  61739=>"010011100",
  61740=>"000011010",
  61741=>"010000110",
  61742=>"011000000",
  61743=>"001000010",
  61744=>"111010001",
  61745=>"110000100",
  61746=>"011111110",
  61747=>"010010110",
  61748=>"010110010",
  61749=>"011100011",
  61750=>"010010110",
  61751=>"010010011",
  61752=>"101000001",
  61753=>"011101011",
  61754=>"011110110",
  61755=>"000000011",
  61756=>"111001111",
  61757=>"111110011",
  61758=>"000111100",
  61759=>"110110000",
  61760=>"100001001",
  61761=>"001111001",
  61762=>"100100011",
  61763=>"010000010",
  61764=>"011000100",
  61765=>"111001100",
  61766=>"100001110",
  61767=>"001011001",
  61768=>"111100000",
  61769=>"010001000",
  61770=>"011010001",
  61771=>"100110001",
  61772=>"111000111",
  61773=>"101111101",
  61774=>"001001001",
  61775=>"011101101",
  61776=>"110010010",
  61777=>"100111011",
  61778=>"000101100",
  61779=>"011000011",
  61780=>"100111001",
  61781=>"000010101",
  61782=>"101100111",
  61783=>"000011110",
  61784=>"001000101",
  61785=>"101101000",
  61786=>"101010101",
  61787=>"011001100",
  61788=>"001111110",
  61789=>"010111111",
  61790=>"111111010",
  61791=>"011111001",
  61792=>"000001000",
  61793=>"100010111",
  61794=>"001011000",
  61795=>"110000011",
  61796=>"010110010",
  61797=>"001001111",
  61798=>"111000000",
  61799=>"010011000",
  61800=>"001000001",
  61801=>"000111010",
  61802=>"001101100",
  61803=>"111010100",
  61804=>"101011001",
  61805=>"011101001",
  61806=>"010111110",
  61807=>"111000111",
  61808=>"010000100",
  61809=>"000010100",
  61810=>"011110111",
  61811=>"100110000",
  61812=>"011101000",
  61813=>"001101000",
  61814=>"111010101",
  61815=>"110011111",
  61816=>"100011111",
  61817=>"010001011",
  61818=>"111000000",
  61819=>"001010000",
  61820=>"101111111",
  61821=>"101010011",
  61822=>"001100011",
  61823=>"000010110",
  61824=>"100101100",
  61825=>"100010001",
  61826=>"011011011",
  61827=>"000100001",
  61828=>"010011100",
  61829=>"111100110",
  61830=>"001110011",
  61831=>"100000100",
  61832=>"010010011",
  61833=>"000111000",
  61834=>"101101110",
  61835=>"001000111",
  61836=>"000111000",
  61837=>"111000101",
  61838=>"110101100",
  61839=>"110010111",
  61840=>"111000101",
  61841=>"001001101",
  61842=>"111101111",
  61843=>"110101000",
  61844=>"100101011",
  61845=>"001100101",
  61846=>"011000000",
  61847=>"110101000",
  61848=>"001111110",
  61849=>"000110101",
  61850=>"101010111",
  61851=>"001000110",
  61852=>"111110010",
  61853=>"000100100",
  61854=>"011111110",
  61855=>"011001100",
  61856=>"100100011",
  61857=>"011001000",
  61858=>"000010111",
  61859=>"111000011",
  61860=>"111011000",
  61861=>"101000101",
  61862=>"001110010",
  61863=>"101111000",
  61864=>"000101110",
  61865=>"111011001",
  61866=>"011101101",
  61867=>"010111000",
  61868=>"110111001",
  61869=>"010000101",
  61870=>"100111101",
  61871=>"101101101",
  61872=>"111011110",
  61873=>"110111100",
  61874=>"000100111",
  61875=>"010101111",
  61876=>"010010100",
  61877=>"101110110",
  61878=>"101011011",
  61879=>"011111100",
  61880=>"001011000",
  61881=>"010000000",
  61882=>"111010010",
  61883=>"100011100",
  61884=>"001100100",
  61885=>"011001011",
  61886=>"000010100",
  61887=>"010111011",
  61888=>"110111011",
  61889=>"001101111",
  61890=>"001110101",
  61891=>"100001110",
  61892=>"110010111",
  61893=>"110011101",
  61894=>"111110001",
  61895=>"000010001",
  61896=>"101011111",
  61897=>"001100110",
  61898=>"010111110",
  61899=>"111011100",
  61900=>"111110110",
  61901=>"101101010",
  61902=>"001010101",
  61903=>"000011010",
  61904=>"101001101",
  61905=>"000001111",
  61906=>"001011001",
  61907=>"110001001",
  61908=>"101000101",
  61909=>"100101001",
  61910=>"101000000",
  61911=>"001010000",
  61912=>"000101011",
  61913=>"110000000",
  61914=>"001101011",
  61915=>"100100000",
  61916=>"111100110",
  61917=>"010100101",
  61918=>"010011000",
  61919=>"110110110",
  61920=>"100010011",
  61921=>"101000011",
  61922=>"010000001",
  61923=>"111011111",
  61924=>"100010011",
  61925=>"000010011",
  61926=>"101101100",
  61927=>"110011100",
  61928=>"110111001",
  61929=>"110101011",
  61930=>"101010000",
  61931=>"110011111",
  61932=>"001110010",
  61933=>"101011011",
  61934=>"100110000",
  61935=>"111001011",
  61936=>"101111111",
  61937=>"110011101",
  61938=>"101100111",
  61939=>"100000000",
  61940=>"110000111",
  61941=>"001000101",
  61942=>"001111001",
  61943=>"101111000",
  61944=>"011000011",
  61945=>"001011100",
  61946=>"101110110",
  61947=>"000010010",
  61948=>"010101001",
  61949=>"011111101",
  61950=>"101110001",
  61951=>"100100000",
  61952=>"111111000",
  61953=>"010011011",
  61954=>"010100101",
  61955=>"100011100",
  61956=>"011011110",
  61957=>"010010001",
  61958=>"001001011",
  61959=>"110011010",
  61960=>"100000000",
  61961=>"101010011",
  61962=>"010111100",
  61963=>"001111100",
  61964=>"000001010",
  61965=>"011011010",
  61966=>"010011010",
  61967=>"001000110",
  61968=>"110101100",
  61969=>"111111001",
  61970=>"000011000",
  61971=>"110100001",
  61972=>"111100100",
  61973=>"110011110",
  61974=>"100110000",
  61975=>"111101100",
  61976=>"100111010",
  61977=>"110101011",
  61978=>"001110111",
  61979=>"001011010",
  61980=>"010001111",
  61981=>"011001101",
  61982=>"010110001",
  61983=>"111001010",
  61984=>"111010011",
  61985=>"001110110",
  61986=>"101100100",
  61987=>"010011100",
  61988=>"110011110",
  61989=>"000100000",
  61990=>"111000001",
  61991=>"000011011",
  61992=>"110011001",
  61993=>"110000100",
  61994=>"000001000",
  61995=>"110101111",
  61996=>"000011100",
  61997=>"111100000",
  61998=>"001000010",
  61999=>"110100101",
  62000=>"111101100",
  62001=>"110011100",
  62002=>"101001001",
  62003=>"010001000",
  62004=>"001011011",
  62005=>"111100101",
  62006=>"101001010",
  62007=>"011101111",
  62008=>"011011100",
  62009=>"010010101",
  62010=>"000111001",
  62011=>"010100001",
  62012=>"001011011",
  62013=>"100111110",
  62014=>"110010101",
  62015=>"101100101",
  62016=>"010001111",
  62017=>"010110001",
  62018=>"000001010",
  62019=>"001011100",
  62020=>"011001111",
  62021=>"011101001",
  62022=>"101010100",
  62023=>"011010001",
  62024=>"000000000",
  62025=>"000001001",
  62026=>"001000010",
  62027=>"000000000",
  62028=>"010101001",
  62029=>"010100111",
  62030=>"011110111",
  62031=>"111101110",
  62032=>"000100110",
  62033=>"100101110",
  62034=>"101000011",
  62035=>"011001110",
  62036=>"100000011",
  62037=>"011000111",
  62038=>"001000101",
  62039=>"010110010",
  62040=>"111010101",
  62041=>"000110010",
  62042=>"010000011",
  62043=>"010000010",
  62044=>"100010001",
  62045=>"011100000",
  62046=>"000101100",
  62047=>"011010010",
  62048=>"101111001",
  62049=>"000101100",
  62050=>"101001010",
  62051=>"100100110",
  62052=>"001010011",
  62053=>"011100011",
  62054=>"110001101",
  62055=>"001001100",
  62056=>"111000010",
  62057=>"100001110",
  62058=>"000100001",
  62059=>"100101110",
  62060=>"100001111",
  62061=>"010000000",
  62062=>"101111100",
  62063=>"111010001",
  62064=>"101100011",
  62065=>"001010110",
  62066=>"101101101",
  62067=>"011100001",
  62068=>"001110010",
  62069=>"111000100",
  62070=>"101000001",
  62071=>"010010000",
  62072=>"111100111",
  62073=>"110001111",
  62074=>"001010010",
  62075=>"101111010",
  62076=>"101010100",
  62077=>"001110010",
  62078=>"010100011",
  62079=>"110111100",
  62080=>"001101010",
  62081=>"100001010",
  62082=>"001001000",
  62083=>"011101010",
  62084=>"011100111",
  62085=>"110100001",
  62086=>"101000010",
  62087=>"100101100",
  62088=>"010100011",
  62089=>"110010000",
  62090=>"001111110",
  62091=>"110010010",
  62092=>"110101011",
  62093=>"011101011",
  62094=>"101110000",
  62095=>"000011011",
  62096=>"010000110",
  62097=>"101110010",
  62098=>"110011100",
  62099=>"010101000",
  62100=>"101101101",
  62101=>"110010110",
  62102=>"010010010",
  62103=>"011100000",
  62104=>"011111000",
  62105=>"010011101",
  62106=>"110000010",
  62107=>"101110100",
  62108=>"000110100",
  62109=>"010110000",
  62110=>"010101000",
  62111=>"000001001",
  62112=>"011000100",
  62113=>"000101100",
  62114=>"101111100",
  62115=>"110010001",
  62116=>"001100011",
  62117=>"011001111",
  62118=>"011000100",
  62119=>"100010000",
  62120=>"010010100",
  62121=>"110000011",
  62122=>"100000011",
  62123=>"111110101",
  62124=>"001010100",
  62125=>"001000000",
  62126=>"010010100",
  62127=>"001101111",
  62128=>"010010001",
  62129=>"001010100",
  62130=>"100000101",
  62131=>"111100110",
  62132=>"001101001",
  62133=>"111100010",
  62134=>"110000100",
  62135=>"010110011",
  62136=>"000111110",
  62137=>"111000011",
  62138=>"011101010",
  62139=>"100000101",
  62140=>"111111110",
  62141=>"001111100",
  62142=>"000110101",
  62143=>"111101101",
  62144=>"011011010",
  62145=>"011010010",
  62146=>"101111010",
  62147=>"110010101",
  62148=>"111110000",
  62149=>"111101110",
  62150=>"001110111",
  62151=>"100101001",
  62152=>"110101000",
  62153=>"000100000",
  62154=>"111110100",
  62155=>"111001101",
  62156=>"110100011",
  62157=>"101111010",
  62158=>"010100010",
  62159=>"000100000",
  62160=>"100110000",
  62161=>"001010010",
  62162=>"100101101",
  62163=>"001011010",
  62164=>"011001001",
  62165=>"010000010",
  62166=>"011011111",
  62167=>"110000100",
  62168=>"100110111",
  62169=>"000110011",
  62170=>"100000000",
  62171=>"001000011",
  62172=>"101001100",
  62173=>"010010001",
  62174=>"100011101",
  62175=>"111110010",
  62176=>"001011010",
  62177=>"001100001",
  62178=>"110111001",
  62179=>"100100101",
  62180=>"001011001",
  62181=>"001101010",
  62182=>"101010001",
  62183=>"001100011",
  62184=>"010001001",
  62185=>"101011000",
  62186=>"001011110",
  62187=>"011001000",
  62188=>"110100010",
  62189=>"110011101",
  62190=>"110110110",
  62191=>"101101110",
  62192=>"011110110",
  62193=>"010000000",
  62194=>"100110010",
  62195=>"000011001",
  62196=>"011100001",
  62197=>"010000101",
  62198=>"100011000",
  62199=>"001000101",
  62200=>"001011000",
  62201=>"110011101",
  62202=>"010100001",
  62203=>"100111010",
  62204=>"101111010",
  62205=>"011000010",
  62206=>"101111110",
  62207=>"011010111",
  62208=>"011110010",
  62209=>"000100010",
  62210=>"001001000",
  62211=>"000000110",
  62212=>"110010010",
  62213=>"111101101",
  62214=>"100011011",
  62215=>"010001011",
  62216=>"001001111",
  62217=>"101000100",
  62218=>"010001010",
  62219=>"010010000",
  62220=>"010100011",
  62221=>"110101000",
  62222=>"100010010",
  62223=>"100111000",
  62224=>"011001000",
  62225=>"001010111",
  62226=>"001010011",
  62227=>"011100010",
  62228=>"111011101",
  62229=>"000101100",
  62230=>"110001110",
  62231=>"101000100",
  62232=>"010011001",
  62233=>"101011001",
  62234=>"011111101",
  62235=>"100000100",
  62236=>"000101110",
  62237=>"100000100",
  62238=>"100010110",
  62239=>"010010111",
  62240=>"110100011",
  62241=>"001001101",
  62242=>"100010011",
  62243=>"101010011",
  62244=>"011000011",
  62245=>"000001110",
  62246=>"010001001",
  62247=>"011110101",
  62248=>"001100001",
  62249=>"010000010",
  62250=>"001111011",
  62251=>"111111100",
  62252=>"100100101",
  62253=>"111011000",
  62254=>"011010010",
  62255=>"000011000",
  62256=>"100000101",
  62257=>"100100101",
  62258=>"000010100",
  62259=>"100100010",
  62260=>"111000001",
  62261=>"111000101",
  62262=>"101011011",
  62263=>"101010110",
  62264=>"001111111",
  62265=>"000000101",
  62266=>"011001111",
  62267=>"000111001",
  62268=>"000101100",
  62269=>"100100111",
  62270=>"010111000",
  62271=>"001100001",
  62272=>"110010011",
  62273=>"101011010",
  62274=>"000000001",
  62275=>"001101001",
  62276=>"111011011",
  62277=>"100001011",
  62278=>"110110011",
  62279=>"011101010",
  62280=>"000101100",
  62281=>"011011011",
  62282=>"110010101",
  62283=>"000011011",
  62284=>"100101101",
  62285=>"001110010",
  62286=>"010110011",
  62287=>"111011111",
  62288=>"110000010",
  62289=>"000101010",
  62290=>"000010010",
  62291=>"100111111",
  62292=>"011011001",
  62293=>"011101001",
  62294=>"010011000",
  62295=>"010100000",
  62296=>"011001101",
  62297=>"111110011",
  62298=>"101111001",
  62299=>"011100101",
  62300=>"001000111",
  62301=>"101010011",
  62302=>"111001111",
  62303=>"000101111",
  62304=>"101101000",
  62305=>"000101010",
  62306=>"011001110",
  62307=>"111110000",
  62308=>"101010111",
  62309=>"111011001",
  62310=>"000010001",
  62311=>"011111111",
  62312=>"000111000",
  62313=>"001100010",
  62314=>"010001110",
  62315=>"000100010",
  62316=>"101001010",
  62317=>"001001101",
  62318=>"100111011",
  62319=>"110110111",
  62320=>"111011110",
  62321=>"011000100",
  62322=>"101011110",
  62323=>"010110110",
  62324=>"000100001",
  62325=>"111000110",
  62326=>"000001001",
  62327=>"010100001",
  62328=>"111011011",
  62329=>"110111001",
  62330=>"111101101",
  62331=>"111001010",
  62332=>"010011001",
  62333=>"011101101",
  62334=>"110101111",
  62335=>"101001000",
  62336=>"011110110",
  62337=>"000000011",
  62338=>"100100001",
  62339=>"110001111",
  62340=>"010011100",
  62341=>"110001111",
  62342=>"000000000",
  62343=>"010101001",
  62344=>"001110101",
  62345=>"110001101",
  62346=>"110011010",
  62347=>"001011010",
  62348=>"000100000",
  62349=>"011010010",
  62350=>"100011111",
  62351=>"111100000",
  62352=>"101111110",
  62353=>"011010111",
  62354=>"000000000",
  62355=>"000101101",
  62356=>"010010100",
  62357=>"110001001",
  62358=>"100101011",
  62359=>"001101000",
  62360=>"111111110",
  62361=>"000011111",
  62362=>"001101101",
  62363=>"011101100",
  62364=>"111101011",
  62365=>"011011011",
  62366=>"100011010",
  62367=>"110110101",
  62368=>"111100000",
  62369=>"101100100",
  62370=>"100101001",
  62371=>"010000100",
  62372=>"001000010",
  62373=>"111010011",
  62374=>"010100011",
  62375=>"011111000",
  62376=>"011101010",
  62377=>"101001100",
  62378=>"000100111",
  62379=>"010001110",
  62380=>"000100101",
  62381=>"001001010",
  62382=>"000010000",
  62383=>"010000101",
  62384=>"111001010",
  62385=>"011110111",
  62386=>"010100011",
  62387=>"111010000",
  62388=>"101001100",
  62389=>"110110010",
  62390=>"111001101",
  62391=>"000001001",
  62392=>"000000101",
  62393=>"000010100",
  62394=>"111010100",
  62395=>"011111101",
  62396=>"101100111",
  62397=>"000111001",
  62398=>"110111000",
  62399=>"011100000",
  62400=>"110011011",
  62401=>"001010000",
  62402=>"011110100",
  62403=>"110101011",
  62404=>"000110010",
  62405=>"101000000",
  62406=>"111111101",
  62407=>"101100001",
  62408=>"100101010",
  62409=>"100110000",
  62410=>"001011100",
  62411=>"100101101",
  62412=>"010010110",
  62413=>"100000100",
  62414=>"100101010",
  62415=>"000110001",
  62416=>"101111000",
  62417=>"000001001",
  62418=>"000011100",
  62419=>"000111011",
  62420=>"011101111",
  62421=>"011010001",
  62422=>"011010010",
  62423=>"101010000",
  62424=>"100000011",
  62425=>"101001011",
  62426=>"010000010",
  62427=>"111011000",
  62428=>"001010101",
  62429=>"111001110",
  62430=>"001111110",
  62431=>"010001001",
  62432=>"000011100",
  62433=>"110000011",
  62434=>"101000111",
  62435=>"101000100",
  62436=>"000100010",
  62437=>"000001111",
  62438=>"001100100",
  62439=>"000011111",
  62440=>"011010100",
  62441=>"011000110",
  62442=>"111110001",
  62443=>"101000010",
  62444=>"010100100",
  62445=>"001001010",
  62446=>"001001100",
  62447=>"110111010",
  62448=>"000001011",
  62449=>"100010100",
  62450=>"010110111",
  62451=>"011010110",
  62452=>"001111001",
  62453=>"101010100",
  62454=>"111100011",
  62455=>"111010010",
  62456=>"111100010",
  62457=>"000001110",
  62458=>"001000000",
  62459=>"000001100",
  62460=>"001000010",
  62461=>"010111001",
  62462=>"100001111",
  62463=>"001100001",
  62464=>"111000100",
  62465=>"010010011",
  62466=>"100011001",
  62467=>"110101010",
  62468=>"001111110",
  62469=>"001110001",
  62470=>"001000010",
  62471=>"101000000",
  62472=>"101101101",
  62473=>"101111101",
  62474=>"011001110",
  62475=>"010011001",
  62476=>"001101111",
  62477=>"001001111",
  62478=>"110110001",
  62479=>"100000011",
  62480=>"010101100",
  62481=>"001111000",
  62482=>"111111101",
  62483=>"101101001",
  62484=>"111011111",
  62485=>"100010100",
  62486=>"001011011",
  62487=>"110011011",
  62488=>"011101100",
  62489=>"101101011",
  62490=>"010011101",
  62491=>"000001100",
  62492=>"111111010",
  62493=>"000111001",
  62494=>"101011100",
  62495=>"010000000",
  62496=>"111001000",
  62497=>"000101111",
  62498=>"000110001",
  62499=>"010010010",
  62500=>"101111001",
  62501=>"100011101",
  62502=>"000011001",
  62503=>"111101100",
  62504=>"001111000",
  62505=>"000111101",
  62506=>"111000100",
  62507=>"100010111",
  62508=>"101001110",
  62509=>"110001110",
  62510=>"100001101",
  62511=>"000100001",
  62512=>"001011111",
  62513=>"110111110",
  62514=>"001011000",
  62515=>"101101011",
  62516=>"100100011",
  62517=>"011001100",
  62518=>"110010101",
  62519=>"001010111",
  62520=>"100000010",
  62521=>"011110110",
  62522=>"000000010",
  62523=>"110011100",
  62524=>"100001101",
  62525=>"100101011",
  62526=>"100000011",
  62527=>"001100001",
  62528=>"000110111",
  62529=>"000000100",
  62530=>"101010010",
  62531=>"010010010",
  62532=>"001010110",
  62533=>"100001111",
  62534=>"000010111",
  62535=>"011101011",
  62536=>"100101001",
  62537=>"001001110",
  62538=>"101101010",
  62539=>"101010110",
  62540=>"000001110",
  62541=>"111100110",
  62542=>"110111110",
  62543=>"111001100",
  62544=>"101110100",
  62545=>"111001100",
  62546=>"110010100",
  62547=>"101111010",
  62548=>"101101100",
  62549=>"000100000",
  62550=>"000010110",
  62551=>"001101100",
  62552=>"110101000",
  62553=>"001110010",
  62554=>"001011010",
  62555=>"011001110",
  62556=>"000010001",
  62557=>"100011001",
  62558=>"000000010",
  62559=>"110100011",
  62560=>"111100111",
  62561=>"111010000",
  62562=>"000100100",
  62563=>"001000011",
  62564=>"000001000",
  62565=>"001010001",
  62566=>"011110010",
  62567=>"111000101",
  62568=>"001110111",
  62569=>"101111000",
  62570=>"111011001",
  62571=>"110001110",
  62572=>"010100111",
  62573=>"001111010",
  62574=>"110101011",
  62575=>"110010011",
  62576=>"110000000",
  62577=>"110010011",
  62578=>"111100011",
  62579=>"110010000",
  62580=>"101001111",
  62581=>"100001110",
  62582=>"001111111",
  62583=>"101010001",
  62584=>"110010100",
  62585=>"100101110",
  62586=>"011011001",
  62587=>"101111000",
  62588=>"011001101",
  62589=>"001000010",
  62590=>"010100100",
  62591=>"101001010",
  62592=>"001111100",
  62593=>"011011110",
  62594=>"010100000",
  62595=>"011000010",
  62596=>"010010011",
  62597=>"001111111",
  62598=>"000000000",
  62599=>"110101010",
  62600=>"110001110",
  62601=>"000000100",
  62602=>"001001111",
  62603=>"010000000",
  62604=>"110011000",
  62605=>"100001111",
  62606=>"001011111",
  62607=>"010011010",
  62608=>"001110010",
  62609=>"011100011",
  62610=>"011100010",
  62611=>"111010011",
  62612=>"011010011",
  62613=>"001000101",
  62614=>"100100011",
  62615=>"111100110",
  62616=>"001010111",
  62617=>"101111011",
  62618=>"001001111",
  62619=>"000011010",
  62620=>"111011001",
  62621=>"010010000",
  62622=>"110101000",
  62623=>"110001100",
  62624=>"101000110",
  62625=>"010100110",
  62626=>"101111111",
  62627=>"110001001",
  62628=>"100101010",
  62629=>"010100100",
  62630=>"001001101",
  62631=>"000010011",
  62632=>"010110101",
  62633=>"011001000",
  62634=>"010011101",
  62635=>"010111100",
  62636=>"111011101",
  62637=>"110101011",
  62638=>"100001010",
  62639=>"011111110",
  62640=>"010010011",
  62641=>"000010100",
  62642=>"011001010",
  62643=>"100010110",
  62644=>"001101011",
  62645=>"101101111",
  62646=>"101111000",
  62647=>"010000001",
  62648=>"111101100",
  62649=>"011101101",
  62650=>"001111000",
  62651=>"001000111",
  62652=>"110110111",
  62653=>"001010010",
  62654=>"100000110",
  62655=>"110001111",
  62656=>"101011011",
  62657=>"111111011",
  62658=>"111111100",
  62659=>"011110010",
  62660=>"011000000",
  62661=>"000110111",
  62662=>"100110111",
  62663=>"000010101",
  62664=>"101110001",
  62665=>"100001110",
  62666=>"101010111",
  62667=>"011000001",
  62668=>"001000110",
  62669=>"000011000",
  62670=>"000011100",
  62671=>"000101111",
  62672=>"110010000",
  62673=>"010010110",
  62674=>"110101010",
  62675=>"010011010",
  62676=>"101101011",
  62677=>"101111011",
  62678=>"101100011",
  62679=>"111011111",
  62680=>"100111011",
  62681=>"110001001",
  62682=>"000100110",
  62683=>"011001101",
  62684=>"110110111",
  62685=>"110101010",
  62686=>"110111000",
  62687=>"011101010",
  62688=>"000001001",
  62689=>"101010111",
  62690=>"011000110",
  62691=>"110001001",
  62692=>"001001101",
  62693=>"101010111",
  62694=>"010100110",
  62695=>"010110000",
  62696=>"011010011",
  62697=>"101000110",
  62698=>"111101101",
  62699=>"011101010",
  62700=>"101000001",
  62701=>"110100000",
  62702=>"000111001",
  62703=>"110000100",
  62704=>"101010101",
  62705=>"110100011",
  62706=>"000001000",
  62707=>"110111110",
  62708=>"101001001",
  62709=>"100101101",
  62710=>"101011111",
  62711=>"101000100",
  62712=>"101110011",
  62713=>"100100100",
  62714=>"001010110",
  62715=>"011111011",
  62716=>"011010000",
  62717=>"101110101",
  62718=>"011101011",
  62719=>"011001100",
  62720=>"110001100",
  62721=>"100101111",
  62722=>"110001000",
  62723=>"000100001",
  62724=>"010110010",
  62725=>"100010000",
  62726=>"001110000",
  62727=>"110000000",
  62728=>"001000010",
  62729=>"110000111",
  62730=>"000000010",
  62731=>"111000100",
  62732=>"110101001",
  62733=>"001000110",
  62734=>"100100000",
  62735=>"001110011",
  62736=>"111100101",
  62737=>"110011111",
  62738=>"000110010",
  62739=>"100001001",
  62740=>"010111111",
  62741=>"001010010",
  62742=>"101110111",
  62743=>"111111110",
  62744=>"110001000",
  62745=>"110110110",
  62746=>"101010010",
  62747=>"101101011",
  62748=>"110110001",
  62749=>"011101011",
  62750=>"110101100",
  62751=>"011000110",
  62752=>"000110010",
  62753=>"001011110",
  62754=>"111100101",
  62755=>"000011010",
  62756=>"000111101",
  62757=>"110110010",
  62758=>"100001011",
  62759=>"001110010",
  62760=>"010000101",
  62761=>"011001110",
  62762=>"101110000",
  62763=>"010000001",
  62764=>"110101010",
  62765=>"110001101",
  62766=>"001000110",
  62767=>"100000111",
  62768=>"000110111",
  62769=>"111101111",
  62770=>"000000110",
  62771=>"000100110",
  62772=>"010101000",
  62773=>"011010000",
  62774=>"001001110",
  62775=>"110011000",
  62776=>"000010100",
  62777=>"000010001",
  62778=>"010010011",
  62779=>"000001000",
  62780=>"001100111",
  62781=>"011111011",
  62782=>"001101111",
  62783=>"011100010",
  62784=>"111011000",
  62785=>"000101000",
  62786=>"001110111",
  62787=>"110011011",
  62788=>"100001100",
  62789=>"111111010",
  62790=>"011101010",
  62791=>"010010011",
  62792=>"110010101",
  62793=>"001100101",
  62794=>"010000110",
  62795=>"010101010",
  62796=>"000011110",
  62797=>"000010101",
  62798=>"110111111",
  62799=>"100001011",
  62800=>"100011110",
  62801=>"001000000",
  62802=>"101111010",
  62803=>"000100001",
  62804=>"100001001",
  62805=>"010010110",
  62806=>"010011111",
  62807=>"110110100",
  62808=>"101110110",
  62809=>"101111111",
  62810=>"010000010",
  62811=>"010101001",
  62812=>"110110101",
  62813=>"001010110",
  62814=>"000011010",
  62815=>"000110011",
  62816=>"010001011",
  62817=>"001101111",
  62818=>"100000100",
  62819=>"111001111",
  62820=>"000110000",
  62821=>"110000101",
  62822=>"111100111",
  62823=>"000111011",
  62824=>"110011001",
  62825=>"111000111",
  62826=>"011111011",
  62827=>"110100110",
  62828=>"010000000",
  62829=>"101101110",
  62830=>"110111000",
  62831=>"001101010",
  62832=>"110000111",
  62833=>"011011000",
  62834=>"001001101",
  62835=>"010000111",
  62836=>"001101001",
  62837=>"011010000",
  62838=>"011001111",
  62839=>"000110001",
  62840=>"110110011",
  62841=>"010110101",
  62842=>"010111010",
  62843=>"111101111",
  62844=>"100100001",
  62845=>"110011111",
  62846=>"010110101",
  62847=>"101111111",
  62848=>"100111111",
  62849=>"110000111",
  62850=>"111001111",
  62851=>"111111000",
  62852=>"000000000",
  62853=>"110001010",
  62854=>"010000011",
  62855=>"110011111",
  62856=>"000000101",
  62857=>"111101110",
  62858=>"010111001",
  62859=>"101100000",
  62860=>"011001010",
  62861=>"111011011",
  62862=>"001111100",
  62863=>"110110100",
  62864=>"000011010",
  62865=>"000001001",
  62866=>"000001100",
  62867=>"110011000",
  62868=>"100001001",
  62869=>"001010001",
  62870=>"111111101",
  62871=>"101001110",
  62872=>"001000000",
  62873=>"110101111",
  62874=>"011101100",
  62875=>"000101111",
  62876=>"111110001",
  62877=>"110010101",
  62878=>"100101100",
  62879=>"001111111",
  62880=>"001011101",
  62881=>"000000101",
  62882=>"011100000",
  62883=>"011101001",
  62884=>"011001000",
  62885=>"100111100",
  62886=>"011011001",
  62887=>"011001101",
  62888=>"110111110",
  62889=>"100011011",
  62890=>"100001000",
  62891=>"001010001",
  62892=>"000001000",
  62893=>"010110100",
  62894=>"111111000",
  62895=>"111110111",
  62896=>"001000000",
  62897=>"100110110",
  62898=>"000110001",
  62899=>"111011101",
  62900=>"011111001",
  62901=>"011110010",
  62902=>"000000100",
  62903=>"100001011",
  62904=>"011100101",
  62905=>"101011111",
  62906=>"110110010",
  62907=>"011010111",
  62908=>"110101000",
  62909=>"010011011",
  62910=>"110000100",
  62911=>"000011010",
  62912=>"011001100",
  62913=>"111011111",
  62914=>"110000010",
  62915=>"011001001",
  62916=>"100010000",
  62917=>"110111111",
  62918=>"001000101",
  62919=>"111000110",
  62920=>"000101010",
  62921=>"010000100",
  62922=>"001000110",
  62923=>"110100101",
  62924=>"111101100",
  62925=>"011011000",
  62926=>"100010000",
  62927=>"101010110",
  62928=>"111111101",
  62929=>"000100101",
  62930=>"100100111",
  62931=>"101000111",
  62932=>"001110110",
  62933=>"011101100",
  62934=>"011011111",
  62935=>"110000001",
  62936=>"000001111",
  62937=>"111100100",
  62938=>"010111000",
  62939=>"000000101",
  62940=>"011011011",
  62941=>"100110111",
  62942=>"100110011",
  62943=>"010001000",
  62944=>"100101100",
  62945=>"100110111",
  62946=>"001011011",
  62947=>"111010000",
  62948=>"101001011",
  62949=>"101111111",
  62950=>"010010101",
  62951=>"010100000",
  62952=>"001010101",
  62953=>"000010011",
  62954=>"000110111",
  62955=>"100000110",
  62956=>"000001000",
  62957=>"100101100",
  62958=>"010010010",
  62959=>"011011010",
  62960=>"101000101",
  62961=>"010100101",
  62962=>"011010000",
  62963=>"100001100",
  62964=>"010000010",
  62965=>"010111111",
  62966=>"001011111",
  62967=>"110000000",
  62968=>"000001100",
  62969=>"110010110",
  62970=>"100001100",
  62971=>"100010001",
  62972=>"111011011",
  62973=>"110110100",
  62974=>"110111111",
  62975=>"011000010",
  62976=>"111001000",
  62977=>"100110001",
  62978=>"100010110",
  62979=>"010011000",
  62980=>"011001000",
  62981=>"001100010",
  62982=>"000110101",
  62983=>"110011100",
  62984=>"101010011",
  62985=>"110100100",
  62986=>"010011000",
  62987=>"001010111",
  62988=>"101110011",
  62989=>"000000110",
  62990=>"110010110",
  62991=>"011001101",
  62992=>"101010101",
  62993=>"010101101",
  62994=>"000001110",
  62995=>"100001000",
  62996=>"110010001",
  62997=>"011010101",
  62998=>"010110001",
  62999=>"111011101",
  63000=>"101001001",
  63001=>"011011001",
  63002=>"000010011",
  63003=>"001000111",
  63004=>"010001000",
  63005=>"111101101",
  63006=>"100001001",
  63007=>"000010011",
  63008=>"000000000",
  63009=>"110011101",
  63010=>"001011111",
  63011=>"010111110",
  63012=>"110000010",
  63013=>"100100000",
  63014=>"001011001",
  63015=>"100001100",
  63016=>"001000111",
  63017=>"001000111",
  63018=>"010011000",
  63019=>"110101000",
  63020=>"011100101",
  63021=>"100110011",
  63022=>"111101001",
  63023=>"010010100",
  63024=>"000111010",
  63025=>"000011010",
  63026=>"100101101",
  63027=>"001001101",
  63028=>"101011011",
  63029=>"100101111",
  63030=>"110010001",
  63031=>"001000101",
  63032=>"101011111",
  63033=>"111100100",
  63034=>"111010000",
  63035=>"010010010",
  63036=>"011110101",
  63037=>"010011011",
  63038=>"011101110",
  63039=>"000000001",
  63040=>"100010101",
  63041=>"100011000",
  63042=>"110000000",
  63043=>"100110001",
  63044=>"010001010",
  63045=>"010110110",
  63046=>"110000001",
  63047=>"010010010",
  63048=>"100010011",
  63049=>"101100101",
  63050=>"010101011",
  63051=>"001100001",
  63052=>"101011010",
  63053=>"110110110",
  63054=>"111000100",
  63055=>"100111001",
  63056=>"100110000",
  63057=>"011001010",
  63058=>"111111001",
  63059=>"111001111",
  63060=>"111001011",
  63061=>"000001111",
  63062=>"111000010",
  63063=>"000100110",
  63064=>"010110101",
  63065=>"110000111",
  63066=>"011110000",
  63067=>"000001000",
  63068=>"001110000",
  63069=>"101100001",
  63070=>"000101110",
  63071=>"000000101",
  63072=>"001111000",
  63073=>"110110001",
  63074=>"101110011",
  63075=>"110011110",
  63076=>"101110101",
  63077=>"000110111",
  63078=>"111010010",
  63079=>"111010001",
  63080=>"101001000",
  63081=>"000000111",
  63082=>"010110101",
  63083=>"000010100",
  63084=>"000110000",
  63085=>"001101010",
  63086=>"101110100",
  63087=>"010101010",
  63088=>"011001110",
  63089=>"100111111",
  63090=>"101000000",
  63091=>"000100010",
  63092=>"010000101",
  63093=>"011011110",
  63094=>"000000111",
  63095=>"001000111",
  63096=>"101111011",
  63097=>"100101100",
  63098=>"010011000",
  63099=>"001010110",
  63100=>"110001000",
  63101=>"100010000",
  63102=>"000011010",
  63103=>"010101011",
  63104=>"011110101",
  63105=>"011010101",
  63106=>"000111100",
  63107=>"100101101",
  63108=>"110111101",
  63109=>"101010000",
  63110=>"001000010",
  63111=>"001010010",
  63112=>"001101100",
  63113=>"111110100",
  63114=>"110010100",
  63115=>"001000100",
  63116=>"111110110",
  63117=>"110011011",
  63118=>"011110001",
  63119=>"011001101",
  63120=>"011000000",
  63121=>"101010000",
  63122=>"100010010",
  63123=>"010110011",
  63124=>"100101110",
  63125=>"110101010",
  63126=>"010110000",
  63127=>"010110010",
  63128=>"011101010",
  63129=>"001101100",
  63130=>"001011010",
  63131=>"000101111",
  63132=>"111000000",
  63133=>"100101010",
  63134=>"001010001",
  63135=>"001011011",
  63136=>"011111100",
  63137=>"011111100",
  63138=>"011001101",
  63139=>"101001100",
  63140=>"111111010",
  63141=>"000010010",
  63142=>"011000101",
  63143=>"001101110",
  63144=>"101000010",
  63145=>"100001101",
  63146=>"000111101",
  63147=>"110011001",
  63148=>"001111011",
  63149=>"010110101",
  63150=>"010110011",
  63151=>"101100011",
  63152=>"001010010",
  63153=>"110010110",
  63154=>"100100100",
  63155=>"110111010",
  63156=>"101111101",
  63157=>"100101110",
  63158=>"100001011",
  63159=>"000111011",
  63160=>"100010110",
  63161=>"110111101",
  63162=>"110001110",
  63163=>"100010000",
  63164=>"011001110",
  63165=>"010001100",
  63166=>"001101101",
  63167=>"111101110",
  63168=>"100101101",
  63169=>"110101001",
  63170=>"100101100",
  63171=>"011001011",
  63172=>"010001100",
  63173=>"101110100",
  63174=>"110100100",
  63175=>"000001010",
  63176=>"011001010",
  63177=>"001100110",
  63178=>"001010111",
  63179=>"000101010",
  63180=>"011100010",
  63181=>"110010101",
  63182=>"011101110",
  63183=>"100100010",
  63184=>"100111111",
  63185=>"011010000",
  63186=>"100000110",
  63187=>"100011010",
  63188=>"010100000",
  63189=>"111101111",
  63190=>"101001101",
  63191=>"111111011",
  63192=>"000001110",
  63193=>"101000010",
  63194=>"111101000",
  63195=>"001111101",
  63196=>"001011000",
  63197=>"111100001",
  63198=>"011101111",
  63199=>"010100010",
  63200=>"001110001",
  63201=>"110100010",
  63202=>"000111110",
  63203=>"001101011",
  63204=>"100100010",
  63205=>"110111111",
  63206=>"110100011",
  63207=>"101000010",
  63208=>"010000010",
  63209=>"001011111",
  63210=>"000110010",
  63211=>"110100010",
  63212=>"000001001",
  63213=>"100101100",
  63214=>"011101000",
  63215=>"101011010",
  63216=>"001111100",
  63217=>"110101110",
  63218=>"110101100",
  63219=>"110111001",
  63220=>"001011001",
  63221=>"000110101",
  63222=>"000011010",
  63223=>"001110001",
  63224=>"010000111",
  63225=>"010110110",
  63226=>"111010100",
  63227=>"111100101",
  63228=>"110100011",
  63229=>"110100110",
  63230=>"100010001",
  63231=>"001001111",
  63232=>"101111110",
  63233=>"011001111",
  63234=>"100010011",
  63235=>"000000010",
  63236=>"010110000",
  63237=>"000111010",
  63238=>"000101011",
  63239=>"111101001",
  63240=>"011111010",
  63241=>"111001000",
  63242=>"101100111",
  63243=>"001100110",
  63244=>"110111010",
  63245=>"010111010",
  63246=>"101011010",
  63247=>"100010011",
  63248=>"011000111",
  63249=>"111101110",
  63250=>"001101101",
  63251=>"100010110",
  63252=>"011111000",
  63253=>"001010000",
  63254=>"011110101",
  63255=>"111111110",
  63256=>"000000111",
  63257=>"000000111",
  63258=>"100100011",
  63259=>"101110001",
  63260=>"111101101",
  63261=>"011110110",
  63262=>"110111111",
  63263=>"001110011",
  63264=>"101101000",
  63265=>"100100100",
  63266=>"001100010",
  63267=>"001100111",
  63268=>"010100111",
  63269=>"111010011",
  63270=>"000001011",
  63271=>"001010001",
  63272=>"100100001",
  63273=>"000011101",
  63274=>"001000100",
  63275=>"111010110",
  63276=>"111100000",
  63277=>"101100010",
  63278=>"110000011",
  63279=>"000000000",
  63280=>"111100001",
  63281=>"010000111",
  63282=>"110111000",
  63283=>"111010011",
  63284=>"011111000",
  63285=>"111100000",
  63286=>"000010000",
  63287=>"001000010",
  63288=>"100101010",
  63289=>"001001111",
  63290=>"111100100",
  63291=>"110100101",
  63292=>"111111101",
  63293=>"100110010",
  63294=>"001100101",
  63295=>"111011111",
  63296=>"001011011",
  63297=>"001110000",
  63298=>"000100101",
  63299=>"110001101",
  63300=>"111110011",
  63301=>"010110101",
  63302=>"101111110",
  63303=>"010001011",
  63304=>"001000011",
  63305=>"011101110",
  63306=>"110001100",
  63307=>"100000011",
  63308=>"000101100",
  63309=>"000101101",
  63310=>"110011000",
  63311=>"111011110",
  63312=>"101010100",
  63313=>"110100001",
  63314=>"010011011",
  63315=>"000001011",
  63316=>"110101010",
  63317=>"001001010",
  63318=>"110011100",
  63319=>"011101000",
  63320=>"101010111",
  63321=>"000101101",
  63322=>"100110010",
  63323=>"111111010",
  63324=>"110000010",
  63325=>"000100000",
  63326=>"110011101",
  63327=>"101100000",
  63328=>"101000001",
  63329=>"101100100",
  63330=>"110001111",
  63331=>"011000000",
  63332=>"101110110",
  63333=>"000000000",
  63334=>"110010110",
  63335=>"000011000",
  63336=>"111000001",
  63337=>"000011110",
  63338=>"100011100",
  63339=>"011111111",
  63340=>"100000011",
  63341=>"010110011",
  63342=>"101000100",
  63343=>"111111100",
  63344=>"010101000",
  63345=>"000011010",
  63346=>"110100101",
  63347=>"011101000",
  63348=>"000111100",
  63349=>"100111011",
  63350=>"010100100",
  63351=>"100100100",
  63352=>"000110101",
  63353=>"110010010",
  63354=>"100001110",
  63355=>"110101110",
  63356=>"011110000",
  63357=>"011010110",
  63358=>"111101001",
  63359=>"110111010",
  63360=>"010110001",
  63361=>"101010010",
  63362=>"110000100",
  63363=>"001110010",
  63364=>"101111010",
  63365=>"000111110",
  63366=>"100111111",
  63367=>"010010100",
  63368=>"000010001",
  63369=>"010000101",
  63370=>"000100111",
  63371=>"001010011",
  63372=>"000101010",
  63373=>"101111001",
  63374=>"000011010",
  63375=>"010001001",
  63376=>"111101111",
  63377=>"000001110",
  63378=>"010100110",
  63379=>"000001111",
  63380=>"011101011",
  63381=>"100011000",
  63382=>"001111110",
  63383=>"000011001",
  63384=>"010111110",
  63385=>"011110101",
  63386=>"011100111",
  63387=>"010011000",
  63388=>"011100000",
  63389=>"011011101",
  63390=>"000110001",
  63391=>"010011010",
  63392=>"000111010",
  63393=>"111100011",
  63394=>"000011011",
  63395=>"000101101",
  63396=>"100000100",
  63397=>"100101100",
  63398=>"101011000",
  63399=>"011101100",
  63400=>"000110011",
  63401=>"101110111",
  63402=>"001100011",
  63403=>"011101011",
  63404=>"010110100",
  63405=>"110101111",
  63406=>"001110001",
  63407=>"000010111",
  63408=>"001001011",
  63409=>"110111000",
  63410=>"110001110",
  63411=>"001101110",
  63412=>"011110001",
  63413=>"011000101",
  63414=>"000001000",
  63415=>"011001110",
  63416=>"011110101",
  63417=>"000001111",
  63418=>"111101000",
  63419=>"101001101",
  63420=>"001101111",
  63421=>"011001111",
  63422=>"101101110",
  63423=>"100111111",
  63424=>"001110011",
  63425=>"010011110",
  63426=>"101000010",
  63427=>"111100110",
  63428=>"101101000",
  63429=>"000011001",
  63430=>"011010000",
  63431=>"010010000",
  63432=>"010110011",
  63433=>"001000101",
  63434=>"001001011",
  63435=>"010111001",
  63436=>"101101010",
  63437=>"110011011",
  63438=>"000110010",
  63439=>"011111000",
  63440=>"001110111",
  63441=>"010111110",
  63442=>"001001000",
  63443=>"010110100",
  63444=>"101101111",
  63445=>"010110111",
  63446=>"011001010",
  63447=>"101110101",
  63448=>"111001101",
  63449=>"010110110",
  63450=>"000110010",
  63451=>"111000011",
  63452=>"001011000",
  63453=>"000100010",
  63454=>"000011100",
  63455=>"001000000",
  63456=>"010000001",
  63457=>"111011101",
  63458=>"101110101",
  63459=>"000011110",
  63460=>"100000111",
  63461=>"000010011",
  63462=>"111010001",
  63463=>"011001110",
  63464=>"101101011",
  63465=>"110001001",
  63466=>"001011000",
  63467=>"010010011",
  63468=>"001111000",
  63469=>"000101100",
  63470=>"110110001",
  63471=>"000001000",
  63472=>"100111011",
  63473=>"000100011",
  63474=>"110000111",
  63475=>"010111111",
  63476=>"110111000",
  63477=>"010001011",
  63478=>"111110111",
  63479=>"000101111",
  63480=>"010101101",
  63481=>"100111001",
  63482=>"010000011",
  63483=>"011011001",
  63484=>"101010111",
  63485=>"010001000",
  63486=>"011000100",
  63487=>"000001111",
  63488=>"100100101",
  63489=>"101111111",
  63490=>"011011111",
  63491=>"110011111",
  63492=>"000000001",
  63493=>"011000100",
  63494=>"000000111",
  63495=>"100111110",
  63496=>"100111110",
  63497=>"101011110",
  63498=>"111100001",
  63499=>"011011000",
  63500=>"000010101",
  63501=>"111110000",
  63502=>"000000101",
  63503=>"110000000",
  63504=>"100010011",
  63505=>"111110010",
  63506=>"011111011",
  63507=>"000100010",
  63508=>"011011010",
  63509=>"110101110",
  63510=>"000110111",
  63511=>"010001000",
  63512=>"110000000",
  63513=>"110101010",
  63514=>"111011000",
  63515=>"001100001",
  63516=>"101111011",
  63517=>"111110110",
  63518=>"110111001",
  63519=>"010010010",
  63520=>"111101000",
  63521=>"110000001",
  63522=>"100110100",
  63523=>"000000001",
  63524=>"011101110",
  63525=>"110110010",
  63526=>"011111011",
  63527=>"101000011",
  63528=>"111000000",
  63529=>"101000000",
  63530=>"101111100",
  63531=>"001100000",
  63532=>"111101111",
  63533=>"110111101",
  63534=>"100100001",
  63535=>"110011100",
  63536=>"101101000",
  63537=>"010010010",
  63538=>"101111000",
  63539=>"111101000",
  63540=>"110010011",
  63541=>"100101000",
  63542=>"001010001",
  63543=>"101100010",
  63544=>"011010110",
  63545=>"000101010",
  63546=>"010011010",
  63547=>"001011010",
  63548=>"100000010",
  63549=>"110001110",
  63550=>"111100111",
  63551=>"111001111",
  63552=>"001111100",
  63553=>"001000001",
  63554=>"100000001",
  63555=>"101100011",
  63556=>"010001110",
  63557=>"000011101",
  63558=>"010000110",
  63559=>"100100110",
  63560=>"110101100",
  63561=>"101101101",
  63562=>"001100110",
  63563=>"110000001",
  63564=>"010111110",
  63565=>"011010000",
  63566=>"000101111",
  63567=>"000000100",
  63568=>"001111001",
  63569=>"100100101",
  63570=>"100110000",
  63571=>"010001001",
  63572=>"011101100",
  63573=>"000110110",
  63574=>"010101011",
  63575=>"110110111",
  63576=>"111110010",
  63577=>"111111111",
  63578=>"100000110",
  63579=>"000111000",
  63580=>"100000010",
  63581=>"110010010",
  63582=>"101010001",
  63583=>"010111001",
  63584=>"001011000",
  63585=>"011000011",
  63586=>"001101011",
  63587=>"101001000",
  63588=>"110111100",
  63589=>"100110110",
  63590=>"111000010",
  63591=>"011100100",
  63592=>"110111100",
  63593=>"001110100",
  63594=>"111101110",
  63595=>"110000010",
  63596=>"010011000",
  63597=>"010000001",
  63598=>"111110010",
  63599=>"010011111",
  63600=>"000000111",
  63601=>"011010100",
  63602=>"101111101",
  63603=>"111101010",
  63604=>"011001000",
  63605=>"110100100",
  63606=>"000010011",
  63607=>"111011011",
  63608=>"011111110",
  63609=>"001011011",
  63610=>"010010101",
  63611=>"001000010",
  63612=>"111010101",
  63613=>"111011110",
  63614=>"101101100",
  63615=>"100101001",
  63616=>"001000000",
  63617=>"000111011",
  63618=>"000010110",
  63619=>"101010000",
  63620=>"011010010",
  63621=>"111110100",
  63622=>"011000100",
  63623=>"000110000",
  63624=>"101111001",
  63625=>"011110001",
  63626=>"100101010",
  63627=>"101111100",
  63628=>"111100111",
  63629=>"101010100",
  63630=>"011100010",
  63631=>"111110111",
  63632=>"000010001",
  63633=>"000100100",
  63634=>"100111010",
  63635=>"001111101",
  63636=>"110100001",
  63637=>"011010010",
  63638=>"111001111",
  63639=>"101101100",
  63640=>"000011101",
  63641=>"110100110",
  63642=>"000001010",
  63643=>"010001000",
  63644=>"010111110",
  63645=>"111000000",
  63646=>"010111010",
  63647=>"110000111",
  63648=>"111000100",
  63649=>"101010011",
  63650=>"011111111",
  63651=>"110111010",
  63652=>"111110010",
  63653=>"110110000",
  63654=>"110010101",
  63655=>"011100110",
  63656=>"001010100",
  63657=>"101011101",
  63658=>"110101101",
  63659=>"111010111",
  63660=>"001100001",
  63661=>"111101111",
  63662=>"101101000",
  63663=>"100001011",
  63664=>"000011011",
  63665=>"001000111",
  63666=>"001110010",
  63667=>"100101100",
  63668=>"000001010",
  63669=>"001010010",
  63670=>"010110110",
  63671=>"111101111",
  63672=>"010110110",
  63673=>"101001010",
  63674=>"010101101",
  63675=>"101111100",
  63676=>"111110110",
  63677=>"111101101",
  63678=>"111101000",
  63679=>"111111100",
  63680=>"110000010",
  63681=>"111100001",
  63682=>"001111010",
  63683=>"010111101",
  63684=>"111010101",
  63685=>"011111101",
  63686=>"111110000",
  63687=>"000100000",
  63688=>"000000101",
  63689=>"000010010",
  63690=>"001101011",
  63691=>"100111010",
  63692=>"000111000",
  63693=>"001010110",
  63694=>"100010111",
  63695=>"110111011",
  63696=>"111001000",
  63697=>"000001001",
  63698=>"000011111",
  63699=>"110000011",
  63700=>"010111011",
  63701=>"100010100",
  63702=>"000001011",
  63703=>"110011011",
  63704=>"111010001",
  63705=>"110101101",
  63706=>"110000010",
  63707=>"011011101",
  63708=>"111111011",
  63709=>"110101000",
  63710=>"111111100",
  63711=>"101100001",
  63712=>"001100100",
  63713=>"100001111",
  63714=>"001111110",
  63715=>"000000101",
  63716=>"101100000",
  63717=>"010101101",
  63718=>"110100101",
  63719=>"000100110",
  63720=>"100100000",
  63721=>"101010010",
  63722=>"011111011",
  63723=>"001010010",
  63724=>"011111011",
  63725=>"000100100",
  63726=>"101010010",
  63727=>"110111111",
  63728=>"010111011",
  63729=>"001011010",
  63730=>"011000010",
  63731=>"001101000",
  63732=>"101001100",
  63733=>"110110100",
  63734=>"010010011",
  63735=>"011100000",
  63736=>"010011111",
  63737=>"101011100",
  63738=>"010011100",
  63739=>"000000011",
  63740=>"000101111",
  63741=>"101100100",
  63742=>"101000111",
  63743=>"000000100",
  63744=>"111100010",
  63745=>"011010110",
  63746=>"110011111",
  63747=>"010001000",
  63748=>"010111001",
  63749=>"000110000",
  63750=>"111000010",
  63751=>"101100100",
  63752=>"000001000",
  63753=>"000001010",
  63754=>"111110001",
  63755=>"101100010",
  63756=>"011110000",
  63757=>"110101110",
  63758=>"100001001",
  63759=>"111010110",
  63760=>"011001010",
  63761=>"111000011",
  63762=>"001110101",
  63763=>"000101010",
  63764=>"011010111",
  63765=>"001100110",
  63766=>"100010111",
  63767=>"010110110",
  63768=>"111100101",
  63769=>"110100011",
  63770=>"101110011",
  63771=>"011011011",
  63772=>"101001111",
  63773=>"111111001",
  63774=>"000010100",
  63775=>"011000000",
  63776=>"100100011",
  63777=>"111000101",
  63778=>"101110111",
  63779=>"101000010",
  63780=>"011111100",
  63781=>"110111110",
  63782=>"000101001",
  63783=>"111111110",
  63784=>"100100010",
  63785=>"010111100",
  63786=>"011000100",
  63787=>"101110000",
  63788=>"010111101",
  63789=>"000000001",
  63790=>"100110100",
  63791=>"101001011",
  63792=>"000100010",
  63793=>"110110011",
  63794=>"100100110",
  63795=>"111001010",
  63796=>"100111010",
  63797=>"011110010",
  63798=>"000010000",
  63799=>"011111111",
  63800=>"000100001",
  63801=>"100111110",
  63802=>"011010101",
  63803=>"101100001",
  63804=>"110100011",
  63805=>"111010100",
  63806=>"001101111",
  63807=>"111111101",
  63808=>"101101001",
  63809=>"101011011",
  63810=>"011111000",
  63811=>"011110100",
  63812=>"111010011",
  63813=>"011000111",
  63814=>"011010010",
  63815=>"111011110",
  63816=>"000110010",
  63817=>"101011101",
  63818=>"111100001",
  63819=>"001111100",
  63820=>"111101110",
  63821=>"011101001",
  63822=>"110001011",
  63823=>"110001000",
  63824=>"000111000",
  63825=>"110101011",
  63826=>"111010011",
  63827=>"111111100",
  63828=>"111011001",
  63829=>"000001101",
  63830=>"010001111",
  63831=>"010111011",
  63832=>"001100000",
  63833=>"000110010",
  63834=>"100010011",
  63835=>"010111111",
  63836=>"000110011",
  63837=>"111010001",
  63838=>"101001100",
  63839=>"010000000",
  63840=>"101101000",
  63841=>"010001000",
  63842=>"000100011",
  63843=>"100100100",
  63844=>"101110000",
  63845=>"000111010",
  63846=>"110101100",
  63847=>"000100000",
  63848=>"101101010",
  63849=>"100001100",
  63850=>"001001101",
  63851=>"111011101",
  63852=>"101000000",
  63853=>"001011101",
  63854=>"111001000",
  63855=>"101110010",
  63856=>"001100001",
  63857=>"001001010",
  63858=>"001101011",
  63859=>"010101111",
  63860=>"110110000",
  63861=>"010100110",
  63862=>"101001101",
  63863=>"010000000",
  63864=>"100000000",
  63865=>"100110100",
  63866=>"001010111",
  63867=>"101010011",
  63868=>"101111101",
  63869=>"111110101",
  63870=>"011001001",
  63871=>"001011111",
  63872=>"101000111",
  63873=>"010010100",
  63874=>"010000000",
  63875=>"100010100",
  63876=>"000110011",
  63877=>"010100010",
  63878=>"110110010",
  63879=>"011100010",
  63880=>"000000001",
  63881=>"000010101",
  63882=>"001001001",
  63883=>"001001010",
  63884=>"000110000",
  63885=>"011001100",
  63886=>"011011111",
  63887=>"100101000",
  63888=>"100110010",
  63889=>"011110000",
  63890=>"101011010",
  63891=>"010000100",
  63892=>"000011011",
  63893=>"101011101",
  63894=>"110110101",
  63895=>"111011001",
  63896=>"011001101",
  63897=>"001000110",
  63898=>"010110111",
  63899=>"110101000",
  63900=>"001111101",
  63901=>"011001000",
  63902=>"011111110",
  63903=>"100010110",
  63904=>"100110010",
  63905=>"000100101",
  63906=>"100100000",
  63907=>"001010010",
  63908=>"000010110",
  63909=>"100100011",
  63910=>"010001001",
  63911=>"110111100",
  63912=>"010110101",
  63913=>"010000010",
  63914=>"000101001",
  63915=>"101010000",
  63916=>"100110110",
  63917=>"110110110",
  63918=>"100010101",
  63919=>"000100011",
  63920=>"000010000",
  63921=>"111001011",
  63922=>"110111001",
  63923=>"100111001",
  63924=>"010110010",
  63925=>"011110000",
  63926=>"001000111",
  63927=>"000100111",
  63928=>"100100101",
  63929=>"101110001",
  63930=>"111011110",
  63931=>"100101101",
  63932=>"110000000",
  63933=>"010011101",
  63934=>"110000010",
  63935=>"001100010",
  63936=>"001111000",
  63937=>"101101100",
  63938=>"011000000",
  63939=>"001000010",
  63940=>"001000111",
  63941=>"101111100",
  63942=>"100100111",
  63943=>"100111001",
  63944=>"111010001",
  63945=>"101100000",
  63946=>"001100000",
  63947=>"110100101",
  63948=>"011100101",
  63949=>"100011001",
  63950=>"010101100",
  63951=>"010101000",
  63952=>"100101101",
  63953=>"001011001",
  63954=>"000000100",
  63955=>"111100010",
  63956=>"111001001",
  63957=>"111111100",
  63958=>"110001000",
  63959=>"101000101",
  63960=>"111001100",
  63961=>"010110011",
  63962=>"101100000",
  63963=>"001100111",
  63964=>"010110011",
  63965=>"011101101",
  63966=>"100001001",
  63967=>"100111001",
  63968=>"001100001",
  63969=>"110110101",
  63970=>"011111010",
  63971=>"010011000",
  63972=>"110011001",
  63973=>"100011110",
  63974=>"101000100",
  63975=>"110000010",
  63976=>"101011011",
  63977=>"010000111",
  63978=>"001011111",
  63979=>"000010101",
  63980=>"111011010",
  63981=>"111100010",
  63982=>"000011010",
  63983=>"110001100",
  63984=>"110010000",
  63985=>"011010000",
  63986=>"111100011",
  63987=>"001000100",
  63988=>"100011001",
  63989=>"110111001",
  63990=>"111110111",
  63991=>"111110010",
  63992=>"001010001",
  63993=>"101100011",
  63994=>"011111110",
  63995=>"000100101",
  63996=>"010101101",
  63997=>"011100000",
  63998=>"111100000",
  63999=>"111101110",
  64000=>"100100000",
  64001=>"011011010",
  64002=>"010100110",
  64003=>"101101101",
  64004=>"100110100",
  64005=>"001011110",
  64006=>"001110110",
  64007=>"000010000",
  64008=>"001000011",
  64009=>"111000110",
  64010=>"001011011",
  64011=>"000000011",
  64012=>"111111111",
  64013=>"011010001",
  64014=>"111111000",
  64015=>"111111001",
  64016=>"110011001",
  64017=>"000001000",
  64018=>"001101110",
  64019=>"000110000",
  64020=>"000111000",
  64021=>"001110000",
  64022=>"000110011",
  64023=>"000111101",
  64024=>"111001111",
  64025=>"100011010",
  64026=>"011000101",
  64027=>"101010000",
  64028=>"010111011",
  64029=>"000110111",
  64030=>"001001101",
  64031=>"001001100",
  64032=>"010001000",
  64033=>"001000110",
  64034=>"100111011",
  64035=>"110000101",
  64036=>"010000000",
  64037=>"100101110",
  64038=>"010011101",
  64039=>"110101100",
  64040=>"110011101",
  64041=>"010010010",
  64042=>"100101011",
  64043=>"011110110",
  64044=>"000000101",
  64045=>"001000000",
  64046=>"000011010",
  64047=>"101101010",
  64048=>"010011100",
  64049=>"000011010",
  64050=>"011110111",
  64051=>"110101001",
  64052=>"001000111",
  64053=>"111100001",
  64054=>"000100000",
  64055=>"000111111",
  64056=>"100110110",
  64057=>"011111011",
  64058=>"011110111",
  64059=>"101001101",
  64060=>"110010010",
  64061=>"000001111",
  64062=>"000010110",
  64063=>"101010000",
  64064=>"101001000",
  64065=>"001000101",
  64066=>"001011011",
  64067=>"111111101",
  64068=>"000010001",
  64069=>"100100011",
  64070=>"000011000",
  64071=>"110110111",
  64072=>"110111000",
  64073=>"010000001",
  64074=>"111011110",
  64075=>"111110011",
  64076=>"000001010",
  64077=>"010011100",
  64078=>"111111000",
  64079=>"000111111",
  64080=>"111111010",
  64081=>"011010000",
  64082=>"011100110",
  64083=>"010100001",
  64084=>"001110010",
  64085=>"101100000",
  64086=>"000111100",
  64087=>"010011110",
  64088=>"110100011",
  64089=>"100010111",
  64090=>"000110011",
  64091=>"000100100",
  64092=>"000110000",
  64093=>"000010001",
  64094=>"111100110",
  64095=>"010111111",
  64096=>"011010101",
  64097=>"100010001",
  64098=>"011110101",
  64099=>"111000100",
  64100=>"100111001",
  64101=>"110010100",
  64102=>"001111010",
  64103=>"111101011",
  64104=>"010111001",
  64105=>"101000001",
  64106=>"101000111",
  64107=>"000001000",
  64108=>"101001000",
  64109=>"010000111",
  64110=>"101011110",
  64111=>"010011111",
  64112=>"101111001",
  64113=>"000111010",
  64114=>"000011011",
  64115=>"110001000",
  64116=>"111101111",
  64117=>"000100101",
  64118=>"001000101",
  64119=>"011101011",
  64120=>"010110101",
  64121=>"101110110",
  64122=>"001110101",
  64123=>"011011111",
  64124=>"011110011",
  64125=>"000001001",
  64126=>"110100000",
  64127=>"111010001",
  64128=>"010000010",
  64129=>"010100010",
  64130=>"010010000",
  64131=>"000000011",
  64132=>"100100000",
  64133=>"001101010",
  64134=>"110001101",
  64135=>"010000101",
  64136=>"100110111",
  64137=>"010100011",
  64138=>"011111000",
  64139=>"110101101",
  64140=>"000110000",
  64141=>"110001111",
  64142=>"001100001",
  64143=>"110000111",
  64144=>"100010110",
  64145=>"110001001",
  64146=>"101001110",
  64147=>"101100011",
  64148=>"100000111",
  64149=>"010000011",
  64150=>"100101101",
  64151=>"011110111",
  64152=>"101100101",
  64153=>"001100110",
  64154=>"101100001",
  64155=>"010100101",
  64156=>"011010001",
  64157=>"101010110",
  64158=>"010100101",
  64159=>"111010001",
  64160=>"100010000",
  64161=>"001100001",
  64162=>"111110000",
  64163=>"010001010",
  64164=>"111101101",
  64165=>"011100110",
  64166=>"111010001",
  64167=>"010000001",
  64168=>"001100101",
  64169=>"110011111",
  64170=>"010001110",
  64171=>"000000000",
  64172=>"100001110",
  64173=>"100111101",
  64174=>"101111111",
  64175=>"000010011",
  64176=>"010111100",
  64177=>"010110000",
  64178=>"011101111",
  64179=>"111000011",
  64180=>"101011110",
  64181=>"001000001",
  64182=>"000100000",
  64183=>"111010010",
  64184=>"101011110",
  64185=>"010110010",
  64186=>"111111110",
  64187=>"110111110",
  64188=>"101011110",
  64189=>"110100100",
  64190=>"000110110",
  64191=>"010100000",
  64192=>"111000000",
  64193=>"000000100",
  64194=>"101111101",
  64195=>"010101111",
  64196=>"101111000",
  64197=>"001111000",
  64198=>"101111100",
  64199=>"101000101",
  64200=>"100000100",
  64201=>"111110010",
  64202=>"101000101",
  64203=>"101110101",
  64204=>"000001000",
  64205=>"110011111",
  64206=>"011101001",
  64207=>"100000000",
  64208=>"111101101",
  64209=>"011110100",
  64210=>"100010001",
  64211=>"101010011",
  64212=>"000011110",
  64213=>"001000111",
  64214=>"000001001",
  64215=>"000010011",
  64216=>"110011000",
  64217=>"011001001",
  64218=>"000111111",
  64219=>"111010100",
  64220=>"011110111",
  64221=>"001001111",
  64222=>"010100110",
  64223=>"100000101",
  64224=>"001111010",
  64225=>"000101000",
  64226=>"001011010",
  64227=>"011011111",
  64228=>"001000001",
  64229=>"011101011",
  64230=>"101000100",
  64231=>"100000001",
  64232=>"011100110",
  64233=>"111011000",
  64234=>"010100101",
  64235=>"011011001",
  64236=>"100110000",
  64237=>"001010110",
  64238=>"110011011",
  64239=>"010010101",
  64240=>"010010110",
  64241=>"001011100",
  64242=>"000000000",
  64243=>"111111100",
  64244=>"100001110",
  64245=>"001101010",
  64246=>"110100111",
  64247=>"010000000",
  64248=>"101010111",
  64249=>"100110010",
  64250=>"000010000",
  64251=>"000101110",
  64252=>"110001101",
  64253=>"101010011",
  64254=>"011100011",
  64255=>"101011110",
  64256=>"000100001",
  64257=>"110011111",
  64258=>"011001111",
  64259=>"001101100",
  64260=>"011100100",
  64261=>"101101010",
  64262=>"011111010",
  64263=>"001000010",
  64264=>"011111000",
  64265=>"100101011",
  64266=>"110010110",
  64267=>"110000011",
  64268=>"011111001",
  64269=>"111100101",
  64270=>"101111000",
  64271=>"010011101",
  64272=>"101011100",
  64273=>"110101000",
  64274=>"001000101",
  64275=>"000000010",
  64276=>"000000010",
  64277=>"111011000",
  64278=>"101001010",
  64279=>"000100010",
  64280=>"010111011",
  64281=>"000010101",
  64282=>"100011010",
  64283=>"110110011",
  64284=>"001111111",
  64285=>"000100100",
  64286=>"001000000",
  64287=>"111011011",
  64288=>"010011111",
  64289=>"110110101",
  64290=>"110110100",
  64291=>"001000011",
  64292=>"100111110",
  64293=>"111001100",
  64294=>"110111010",
  64295=>"011011011",
  64296=>"111111011",
  64297=>"100011100",
  64298=>"010010110",
  64299=>"101001101",
  64300=>"111101111",
  64301=>"000000110",
  64302=>"110100110",
  64303=>"001110110",
  64304=>"000100101",
  64305=>"010010110",
  64306=>"000011011",
  64307=>"011101110",
  64308=>"010010101",
  64309=>"101000001",
  64310=>"100000010",
  64311=>"101111011",
  64312=>"001000110",
  64313=>"001100110",
  64314=>"000011010",
  64315=>"110001010",
  64316=>"011000100",
  64317=>"001111111",
  64318=>"010101101",
  64319=>"101110111",
  64320=>"010100101",
  64321=>"110001011",
  64322=>"010001110",
  64323=>"111100101",
  64324=>"011101011",
  64325=>"100101100",
  64326=>"100011001",
  64327=>"000100000",
  64328=>"101111110",
  64329=>"111111011",
  64330=>"110100111",
  64331=>"001100110",
  64332=>"111100000",
  64333=>"001100101",
  64334=>"000011011",
  64335=>"000011100",
  64336=>"101000011",
  64337=>"111001001",
  64338=>"101010011",
  64339=>"100000101",
  64340=>"011110101",
  64341=>"110000011",
  64342=>"110011111",
  64343=>"011010100",
  64344=>"001111000",
  64345=>"111011101",
  64346=>"001101000",
  64347=>"000000101",
  64348=>"111110100",
  64349=>"110101111",
  64350=>"000101011",
  64351=>"100011010",
  64352=>"010010010",
  64353=>"000000101",
  64354=>"000011111",
  64355=>"100000100",
  64356=>"000010101",
  64357=>"101000111",
  64358=>"010111010",
  64359=>"111111110",
  64360=>"001111111",
  64361=>"011011100",
  64362=>"000010011",
  64363=>"011010011",
  64364=>"111011010",
  64365=>"100000000",
  64366=>"110111000",
  64367=>"100101100",
  64368=>"111100101",
  64369=>"001110101",
  64370=>"111000110",
  64371=>"000111001",
  64372=>"110000000",
  64373=>"010011001",
  64374=>"011000011",
  64375=>"001000000",
  64376=>"011101110",
  64377=>"010010000",
  64378=>"011111111",
  64379=>"010111111",
  64380=>"000010100",
  64381=>"110111111",
  64382=>"101011101",
  64383=>"001110001",
  64384=>"010110110",
  64385=>"001101010",
  64386=>"100010010",
  64387=>"010000010",
  64388=>"101011110",
  64389=>"111100101",
  64390=>"010110000",
  64391=>"101100100",
  64392=>"001110100",
  64393=>"101011000",
  64394=>"111100111",
  64395=>"101111100",
  64396=>"001001000",
  64397=>"101010100",
  64398=>"000110111",
  64399=>"001110010",
  64400=>"111011111",
  64401=>"011011001",
  64402=>"101010001",
  64403=>"011111011",
  64404=>"101100100",
  64405=>"111011110",
  64406=>"111111000",
  64407=>"101100000",
  64408=>"010100011",
  64409=>"100101011",
  64410=>"101100111",
  64411=>"101011001",
  64412=>"000111111",
  64413=>"111010110",
  64414=>"000100101",
  64415=>"110000010",
  64416=>"110000000",
  64417=>"100100100",
  64418=>"111110000",
  64419=>"000100010",
  64420=>"001110011",
  64421=>"010110111",
  64422=>"010111101",
  64423=>"011111111",
  64424=>"011100001",
  64425=>"010110000",
  64426=>"110111000",
  64427=>"000101000",
  64428=>"000000100",
  64429=>"100000101",
  64430=>"001101101",
  64431=>"010000111",
  64432=>"110001100",
  64433=>"110111110",
  64434=>"000001010",
  64435=>"101100010",
  64436=>"101010000",
  64437=>"000010010",
  64438=>"100101101",
  64439=>"101000101",
  64440=>"011011000",
  64441=>"110001010",
  64442=>"100110110",
  64443=>"111101010",
  64444=>"111010111",
  64445=>"110010000",
  64446=>"110010100",
  64447=>"001001110",
  64448=>"100010111",
  64449=>"100011000",
  64450=>"111111100",
  64451=>"000111001",
  64452=>"110110010",
  64453=>"100011111",
  64454=>"101011011",
  64455=>"100001101",
  64456=>"100001110",
  64457=>"001111101",
  64458=>"100000110",
  64459=>"010001011",
  64460=>"110110110",
  64461=>"001100011",
  64462=>"000111000",
  64463=>"101101001",
  64464=>"110001001",
  64465=>"011111001",
  64466=>"011010010",
  64467=>"011000110",
  64468=>"111000011",
  64469=>"100100111",
  64470=>"100010000",
  64471=>"001001100",
  64472=>"101101110",
  64473=>"010111000",
  64474=>"100110101",
  64475=>"100110110",
  64476=>"100111000",
  64477=>"110011011",
  64478=>"111101101",
  64479=>"010011100",
  64480=>"011110110",
  64481=>"011000000",
  64482=>"001000111",
  64483=>"000011110",
  64484=>"101101100",
  64485=>"000000001",
  64486=>"010011101",
  64487=>"100001111",
  64488=>"011110000",
  64489=>"111001011",
  64490=>"110000101",
  64491=>"111000010",
  64492=>"101010011",
  64493=>"110000101",
  64494=>"110101001",
  64495=>"111101001",
  64496=>"000001010",
  64497=>"101000101",
  64498=>"100111010",
  64499=>"000111011",
  64500=>"010101011",
  64501=>"110000110",
  64502=>"111100011",
  64503=>"110001010",
  64504=>"010011001",
  64505=>"111101101",
  64506=>"100010110",
  64507=>"101000010",
  64508=>"010001100",
  64509=>"011011101",
  64510=>"001000111",
  64511=>"010010000",
  64512=>"011000011",
  64513=>"110101001",
  64514=>"110000100",
  64515=>"000111010",
  64516=>"011010100",
  64517=>"011001111",
  64518=>"001110111",
  64519=>"111001000",
  64520=>"011001101",
  64521=>"010101100",
  64522=>"001110011",
  64523=>"110000100",
  64524=>"101101100",
  64525=>"100000000",
  64526=>"110011010",
  64527=>"110101010",
  64528=>"011001100",
  64529=>"010001011",
  64530=>"111100011",
  64531=>"111010000",
  64532=>"001000011",
  64533=>"011100010",
  64534=>"010011011",
  64535=>"100100010",
  64536=>"100011100",
  64537=>"001010000",
  64538=>"000111000",
  64539=>"000100101",
  64540=>"101100100",
  64541=>"010110111",
  64542=>"010101111",
  64543=>"010100101",
  64544=>"000011001",
  64545=>"101000101",
  64546=>"101101101",
  64547=>"011100110",
  64548=>"110110001",
  64549=>"100110000",
  64550=>"110010000",
  64551=>"011000111",
  64552=>"001011011",
  64553=>"111111110",
  64554=>"000010101",
  64555=>"010001000",
  64556=>"110111000",
  64557=>"010111100",
  64558=>"110100000",
  64559=>"100011011",
  64560=>"000101010",
  64561=>"111111001",
  64562=>"000010101",
  64563=>"111010010",
  64564=>"010011110",
  64565=>"010010000",
  64566=>"010001101",
  64567=>"110010111",
  64568=>"010100101",
  64569=>"001000111",
  64570=>"100001000",
  64571=>"010010100",
  64572=>"100101110",
  64573=>"001110110",
  64574=>"101100110",
  64575=>"000011000",
  64576=>"011000011",
  64577=>"111010101",
  64578=>"000001001",
  64579=>"100010100",
  64580=>"110100101",
  64581=>"111001000",
  64582=>"110011011",
  64583=>"001111010",
  64584=>"100010010",
  64585=>"010010000",
  64586=>"110010100",
  64587=>"101100011",
  64588=>"010010111",
  64589=>"101101111",
  64590=>"011110101",
  64591=>"111010010",
  64592=>"010011001",
  64593=>"110100110",
  64594=>"101110001",
  64595=>"001111010",
  64596=>"100110110",
  64597=>"001001101",
  64598=>"000111111",
  64599=>"000000101",
  64600=>"110101010",
  64601=>"100011010",
  64602=>"000010101",
  64603=>"000010110",
  64604=>"100011011",
  64605=>"100101111",
  64606=>"110110101",
  64607=>"010101100",
  64608=>"110000111",
  64609=>"111000010",
  64610=>"010010100",
  64611=>"001011111",
  64612=>"001010110",
  64613=>"000100011",
  64614=>"000010000",
  64615=>"110101000",
  64616=>"100110001",
  64617=>"000001110",
  64618=>"111011011",
  64619=>"111010111",
  64620=>"011110100",
  64621=>"111101110",
  64622=>"011111110",
  64623=>"101001000",
  64624=>"001010011",
  64625=>"100000011",
  64626=>"001100101",
  64627=>"001100011",
  64628=>"010010111",
  64629=>"111111001",
  64630=>"000001001",
  64631=>"011000101",
  64632=>"011100111",
  64633=>"000010101",
  64634=>"010011111",
  64635=>"110111110",
  64636=>"000100010",
  64637=>"000010111",
  64638=>"111000000",
  64639=>"011101110",
  64640=>"101010101",
  64641=>"111101010",
  64642=>"100101001",
  64643=>"011010011",
  64644=>"010001100",
  64645=>"101101111",
  64646=>"101100110",
  64647=>"110101100",
  64648=>"100110010",
  64649=>"010100001",
  64650=>"011010010",
  64651=>"010110000",
  64652=>"011010010",
  64653=>"001101011",
  64654=>"000100100",
  64655=>"001000010",
  64656=>"101000001",
  64657=>"110000101",
  64658=>"101001010",
  64659=>"000110100",
  64660=>"000110100",
  64661=>"000011100",
  64662=>"110000000",
  64663=>"111111011",
  64664=>"010010011",
  64665=>"010000010",
  64666=>"110110010",
  64667=>"001100100",
  64668=>"100101010",
  64669=>"011101001",
  64670=>"110100111",
  64671=>"111110111",
  64672=>"100010101",
  64673=>"100110010",
  64674=>"000110101",
  64675=>"111101101",
  64676=>"100110000",
  64677=>"111110111",
  64678=>"110111001",
  64679=>"111111110",
  64680=>"000001000",
  64681=>"001011001",
  64682=>"011001011",
  64683=>"111111000",
  64684=>"110000010",
  64685=>"001111111",
  64686=>"001000101",
  64687=>"101110101",
  64688=>"000000001",
  64689=>"100001100",
  64690=>"100001011",
  64691=>"111010001",
  64692=>"101110000",
  64693=>"111110100",
  64694=>"100110100",
  64695=>"110001001",
  64696=>"111000010",
  64697=>"100000010",
  64698=>"001000101",
  64699=>"110001100",
  64700=>"010000000",
  64701=>"110001100",
  64702=>"000011011",
  64703=>"100101010",
  64704=>"010110000",
  64705=>"110001100",
  64706=>"001000000",
  64707=>"000000001",
  64708=>"001101011",
  64709=>"001000100",
  64710=>"010111100",
  64711=>"100111111",
  64712=>"011001000",
  64713=>"011111001",
  64714=>"111010110",
  64715=>"001000110",
  64716=>"011110011",
  64717=>"011111111",
  64718=>"000100001",
  64719=>"000100101",
  64720=>"111110110",
  64721=>"000000011",
  64722=>"100111110",
  64723=>"100110001",
  64724=>"101001001",
  64725=>"111100011",
  64726=>"100000110",
  64727=>"101101000",
  64728=>"000010001",
  64729=>"010011011",
  64730=>"011111010",
  64731=>"000010010",
  64732=>"101010011",
  64733=>"001011100",
  64734=>"101101100",
  64735=>"000011000",
  64736=>"000010011",
  64737=>"111100101",
  64738=>"000110010",
  64739=>"100010000",
  64740=>"010101000",
  64741=>"100011010",
  64742=>"100100001",
  64743=>"010111111",
  64744=>"000110011",
  64745=>"100011010",
  64746=>"011001010",
  64747=>"100110010",
  64748=>"110010001",
  64749=>"100000111",
  64750=>"000100000",
  64751=>"011101101",
  64752=>"111101010",
  64753=>"101010110",
  64754=>"111101110",
  64755=>"001000110",
  64756=>"100111000",
  64757=>"100010011",
  64758=>"100110000",
  64759=>"100010010",
  64760=>"100000000",
  64761=>"010100101",
  64762=>"010001101",
  64763=>"000101000",
  64764=>"101000000",
  64765=>"100100000",
  64766=>"110010110",
  64767=>"111111001",
  64768=>"011110001",
  64769=>"001001001",
  64770=>"000010101",
  64771=>"100011101",
  64772=>"011111101",
  64773=>"110110011",
  64774=>"000100000",
  64775=>"101100100",
  64776=>"001110111",
  64777=>"001110100",
  64778=>"011100011",
  64779=>"000100000",
  64780=>"010111010",
  64781=>"111000111",
  64782=>"001110001",
  64783=>"101111111",
  64784=>"101010011",
  64785=>"111010111",
  64786=>"001000001",
  64787=>"000100010",
  64788=>"101010011",
  64789=>"111110100",
  64790=>"111100110",
  64791=>"000010001",
  64792=>"001000100",
  64793=>"111001101",
  64794=>"101001011",
  64795=>"111000101",
  64796=>"001101100",
  64797=>"110100011",
  64798=>"010100110",
  64799=>"100010110",
  64800=>"000110101",
  64801=>"001111001",
  64802=>"001111111",
  64803=>"001010110",
  64804=>"000111100",
  64805=>"111100011",
  64806=>"010001101",
  64807=>"110111010",
  64808=>"001000000",
  64809=>"000101001",
  64810=>"101111010",
  64811=>"100001011",
  64812=>"111100001",
  64813=>"101001001",
  64814=>"101001000",
  64815=>"101111110",
  64816=>"110101010",
  64817=>"110101011",
  64818=>"111110110",
  64819=>"001101110",
  64820=>"111110000",
  64821=>"110000000",
  64822=>"000110001",
  64823=>"001001100",
  64824=>"001000001",
  64825=>"010100110",
  64826=>"100100100",
  64827=>"001110010",
  64828=>"011000100",
  64829=>"100100000",
  64830=>"110100111",
  64831=>"011001000",
  64832=>"111101100",
  64833=>"010000100",
  64834=>"001011101",
  64835=>"100111010",
  64836=>"010010101",
  64837=>"110011010",
  64838=>"111100101",
  64839=>"111110100",
  64840=>"110000110",
  64841=>"101101000",
  64842=>"100110011",
  64843=>"101100010",
  64844=>"101110111",
  64845=>"001010101",
  64846=>"001110110",
  64847=>"001000010",
  64848=>"001111101",
  64849=>"101100100",
  64850=>"100111011",
  64851=>"110101000",
  64852=>"011011010",
  64853=>"000010111",
  64854=>"001111000",
  64855=>"110000001",
  64856=>"100001011",
  64857=>"100110110",
  64858=>"010111100",
  64859=>"100100001",
  64860=>"111111111",
  64861=>"000010000",
  64862=>"101011100",
  64863=>"001101100",
  64864=>"011101100",
  64865=>"011011001",
  64866=>"010101100",
  64867=>"011100000",
  64868=>"011011000",
  64869=>"111111111",
  64870=>"100010101",
  64871=>"011111101",
  64872=>"011110000",
  64873=>"001110100",
  64874=>"100000111",
  64875=>"100001110",
  64876=>"111001001",
  64877=>"001101110",
  64878=>"111101100",
  64879=>"110010101",
  64880=>"001010001",
  64881=>"000001111",
  64882=>"110010011",
  64883=>"110100000",
  64884=>"100100011",
  64885=>"010010011",
  64886=>"000000011",
  64887=>"110111110",
  64888=>"011011110",
  64889=>"100001011",
  64890=>"010100110",
  64891=>"011111111",
  64892=>"001011100",
  64893=>"001010111",
  64894=>"010101011",
  64895=>"101101111",
  64896=>"000110000",
  64897=>"111110100",
  64898=>"110111011",
  64899=>"001110000",
  64900=>"110111001",
  64901=>"100001000",
  64902=>"110011011",
  64903=>"111101010",
  64904=>"000110111",
  64905=>"100010101",
  64906=>"000000001",
  64907=>"111111111",
  64908=>"000101000",
  64909=>"001011101",
  64910=>"100011010",
  64911=>"100001101",
  64912=>"010111101",
  64913=>"000000000",
  64914=>"100110001",
  64915=>"000001101",
  64916=>"001110010",
  64917=>"000100110",
  64918=>"011111110",
  64919=>"110011010",
  64920=>"100100110",
  64921=>"000100110",
  64922=>"100001111",
  64923=>"011101101",
  64924=>"111000011",
  64925=>"100001101",
  64926=>"111000101",
  64927=>"110101000",
  64928=>"111110110",
  64929=>"100110100",
  64930=>"101110100",
  64931=>"110111110",
  64932=>"101001001",
  64933=>"101101000",
  64934=>"001001101",
  64935=>"000001001",
  64936=>"001100111",
  64937=>"001010001",
  64938=>"101011101",
  64939=>"000111011",
  64940=>"101011011",
  64941=>"000110100",
  64942=>"110110101",
  64943=>"010101100",
  64944=>"000010010",
  64945=>"100110101",
  64946=>"010011111",
  64947=>"000000000",
  64948=>"010100100",
  64949=>"001100111",
  64950=>"101001111",
  64951=>"010110100",
  64952=>"001001100",
  64953=>"001010001",
  64954=>"011000011",
  64955=>"101011100",
  64956=>"111111100",
  64957=>"110000000",
  64958=>"011100110",
  64959=>"110101011",
  64960=>"001001110",
  64961=>"110000111",
  64962=>"100111111",
  64963=>"001110001",
  64964=>"111111110",
  64965=>"011101011",
  64966=>"011111100",
  64967=>"101010000",
  64968=>"000001100",
  64969=>"111110010",
  64970=>"101011111",
  64971=>"000000000",
  64972=>"101010000",
  64973=>"101100110",
  64974=>"000001011",
  64975=>"101111110",
  64976=>"101010000",
  64977=>"011000100",
  64978=>"100101000",
  64979=>"110010111",
  64980=>"100011100",
  64981=>"011010111",
  64982=>"110110011",
  64983=>"001001000",
  64984=>"000000000",
  64985=>"111111100",
  64986=>"000101110",
  64987=>"110101010",
  64988=>"011110101",
  64989=>"000100101",
  64990=>"110100001",
  64991=>"000010101",
  64992=>"011010000",
  64993=>"100110111",
  64994=>"110010100",
  64995=>"101111011",
  64996=>"010110011",
  64997=>"110101010",
  64998=>"111111100",
  64999=>"000110100",
  65000=>"111111111",
  65001=>"110100101",
  65002=>"101100100",
  65003=>"101101101",
  65004=>"011000001",
  65005=>"111110101",
  65006=>"110111100",
  65007=>"000100001",
  65008=>"110100010",
  65009=>"110110000",
  65010=>"110000011",
  65011=>"011100100",
  65012=>"111011110",
  65013=>"111010111",
  65014=>"011001100",
  65015=>"001101111",
  65016=>"100100001",
  65017=>"111011001",
  65018=>"110100101",
  65019=>"001110000",
  65020=>"010011001",
  65021=>"011011001",
  65022=>"110100100",
  65023=>"101011010",
  65024=>"001101011",
  65025=>"101111011",
  65026=>"010110111",
  65027=>"000001110",
  65028=>"100100000",
  65029=>"000011000",
  65030=>"110110001",
  65031=>"101001110",
  65032=>"100100100",
  65033=>"100000011",
  65034=>"011011110",
  65035=>"001001000",
  65036=>"100011010",
  65037=>"011001110",
  65038=>"100100001",
  65039=>"010010011",
  65040=>"100010111",
  65041=>"010111110",
  65042=>"000011001",
  65043=>"000101001",
  65044=>"101000110",
  65045=>"101110011",
  65046=>"110110110",
  65047=>"001010100",
  65048=>"100111000",
  65049=>"000010000",
  65050=>"011000001",
  65051=>"001100111",
  65052=>"100001000",
  65053=>"111100100",
  65054=>"100111101",
  65055=>"101111010",
  65056=>"001011011",
  65057=>"010000001",
  65058=>"001000001",
  65059=>"001000010",
  65060=>"111101001",
  65061=>"111001011",
  65062=>"011111110",
  65063=>"100100010",
  65064=>"000110110",
  65065=>"010001000",
  65066=>"010000101",
  65067=>"111011111",
  65068=>"010110101",
  65069=>"101101010",
  65070=>"100100011",
  65071=>"001100000",
  65072=>"100001000",
  65073=>"111110100",
  65074=>"001000101",
  65075=>"011100011",
  65076=>"010100101",
  65077=>"100101001",
  65078=>"100001010",
  65079=>"000001111",
  65080=>"101111111",
  65081=>"110100110",
  65082=>"010101101",
  65083=>"111011101",
  65084=>"001000010",
  65085=>"110111000",
  65086=>"000000101",
  65087=>"111101010",
  65088=>"101110010",
  65089=>"111100000",
  65090=>"100001111",
  65091=>"110001100",
  65092=>"000100001",
  65093=>"110100000",
  65094=>"101111010",
  65095=>"011110110",
  65096=>"011110110",
  65097=>"011010001",
  65098=>"011111000",
  65099=>"101101110",
  65100=>"011111101",
  65101=>"111100110",
  65102=>"100011111",
  65103=>"001101110",
  65104=>"100000010",
  65105=>"101111011",
  65106=>"110100111",
  65107=>"110001001",
  65108=>"011101101",
  65109=>"000000000",
  65110=>"000101100",
  65111=>"111100001",
  65112=>"111000100",
  65113=>"000000101",
  65114=>"001111000",
  65115=>"000011100",
  65116=>"000101110",
  65117=>"000110100",
  65118=>"101011010",
  65119=>"011001110",
  65120=>"011000000",
  65121=>"000001011",
  65122=>"101010101",
  65123=>"010100101",
  65124=>"000000111",
  65125=>"011001111",
  65126=>"000011110",
  65127=>"011011011",
  65128=>"000000001",
  65129=>"000110101",
  65130=>"111111010",
  65131=>"000100100",
  65132=>"100111001",
  65133=>"101000010",
  65134=>"100000101",
  65135=>"010110001",
  65136=>"100001011",
  65137=>"001010000",
  65138=>"111111111",
  65139=>"011111000",
  65140=>"100100000",
  65141=>"011111001",
  65142=>"001100100",
  65143=>"100000110",
  65144=>"001100001",
  65145=>"000110000",
  65146=>"100101001",
  65147=>"011001010",
  65148=>"000001001",
  65149=>"100000010",
  65150=>"111010101",
  65151=>"101111110",
  65152=>"101000000",
  65153=>"111111010",
  65154=>"110101100",
  65155=>"000101011",
  65156=>"111100000",
  65157=>"111001100",
  65158=>"110001100",
  65159=>"011001010",
  65160=>"000100001",
  65161=>"011000111",
  65162=>"001010000",
  65163=>"000010000",
  65164=>"111010111",
  65165=>"010111001",
  65166=>"111000000",
  65167=>"100111100",
  65168=>"010101011",
  65169=>"001100101",
  65170=>"001011111",
  65171=>"001111011",
  65172=>"001100110",
  65173=>"010011110",
  65174=>"001110100",
  65175=>"010000010",
  65176=>"011010111",
  65177=>"001010010",
  65178=>"001111101",
  65179=>"000000011",
  65180=>"010000110",
  65181=>"011110001",
  65182=>"101001110",
  65183=>"010111110",
  65184=>"111101101",
  65185=>"100000110",
  65186=>"100001101",
  65187=>"001011001",
  65188=>"110100101",
  65189=>"100001001",
  65190=>"111001001",
  65191=>"001101001",
  65192=>"100000001",
  65193=>"110000000",
  65194=>"011100111",
  65195=>"111000100",
  65196=>"011000000",
  65197=>"011100010",
  65198=>"111000011",
  65199=>"010011111",
  65200=>"000000000",
  65201=>"110101110",
  65202=>"000101111",
  65203=>"100100111",
  65204=>"100011010",
  65205=>"001101110",
  65206=>"011000001",
  65207=>"111111100",
  65208=>"100110100",
  65209=>"100110111",
  65210=>"101100010",
  65211=>"010101110",
  65212=>"111001001",
  65213=>"110011100",
  65214=>"111101011",
  65215=>"111010011",
  65216=>"101110101",
  65217=>"010000110",
  65218=>"100011100",
  65219=>"000101011",
  65220=>"001101101",
  65221=>"001011011",
  65222=>"011110110",
  65223=>"110000100",
  65224=>"111000000",
  65225=>"110111101",
  65226=>"100111110",
  65227=>"000000000",
  65228=>"101101111",
  65229=>"001000010",
  65230=>"111010000",
  65231=>"111100010",
  65232=>"110010000",
  65233=>"000100000",
  65234=>"011100000",
  65235=>"000111101",
  65236=>"001111001",
  65237=>"010011111",
  65238=>"000011111",
  65239=>"000111001",
  65240=>"010001011",
  65241=>"110111100",
  65242=>"111110001",
  65243=>"000101101",
  65244=>"101100001",
  65245=>"101001110",
  65246=>"111111111",
  65247=>"010011100",
  65248=>"111101001",
  65249=>"100100011",
  65250=>"000011100",
  65251=>"011110001",
  65252=>"101100000",
  65253=>"011010000",
  65254=>"010100101",
  65255=>"100001001",
  65256=>"101111110",
  65257=>"101111101",
  65258=>"011010001",
  65259=>"101000110",
  65260=>"001000001",
  65261=>"100101101",
  65262=>"001100110",
  65263=>"000011000",
  65264=>"110010000",
  65265=>"111111000",
  65266=>"001110000",
  65267=>"101110111",
  65268=>"011110010",
  65269=>"011000000",
  65270=>"100111010",
  65271=>"011111101",
  65272=>"010011000",
  65273=>"110100100",
  65274=>"001010010",
  65275=>"001000010",
  65276=>"000011110",
  65277=>"110001111",
  65278=>"000001101",
  65279=>"011011001",
  65280=>"011010100",
  65281=>"110110101",
  65282=>"010010100",
  65283=>"100111101",
  65284=>"100001110",
  65285=>"000110000",
  65286=>"000101110",
  65287=>"101001011",
  65288=>"100001000",
  65289=>"101111101",
  65290=>"011001111",
  65291=>"010100011",
  65292=>"101010100",
  65293=>"010010001",
  65294=>"000101001",
  65295=>"100100100",
  65296=>"000000110",
  65297=>"100100001",
  65298=>"010101011",
  65299=>"110110010",
  65300=>"000100110",
  65301=>"000100101",
  65302=>"001010010",
  65303=>"100111101",
  65304=>"100001101",
  65305=>"001110010",
  65306=>"010100000",
  65307=>"101111001",
  65308=>"001000001",
  65309=>"011001000",
  65310=>"110100110",
  65311=>"010001101",
  65312=>"001011100",
  65313=>"010001100",
  65314=>"011001100",
  65315=>"100001000",
  65316=>"101010101",
  65317=>"111101111",
  65318=>"001110001",
  65319=>"000100000",
  65320=>"100010010",
  65321=>"101001101",
  65322=>"111010110",
  65323=>"111101101",
  65324=>"000000001",
  65325=>"010011001",
  65326=>"001101011",
  65327=>"010110100",
  65328=>"001001011",
  65329=>"011000010",
  65330=>"000001101",
  65331=>"011000000",
  65332=>"010111100",
  65333=>"000110101",
  65334=>"101111111",
  65335=>"011100101",
  65336=>"110001010",
  65337=>"100001100",
  65338=>"011101100",
  65339=>"100010000",
  65340=>"101010100",
  65341=>"010010010",
  65342=>"001101101",
  65343=>"111110111",
  65344=>"101111001",
  65345=>"111111111",
  65346=>"000000100",
  65347=>"110100100",
  65348=>"100010110",
  65349=>"011011010",
  65350=>"110001000",
  65351=>"110100000",
  65352=>"010001110",
  65353=>"100111100",
  65354=>"100110011",
  65355=>"110000000",
  65356=>"101100010",
  65357=>"110110001",
  65358=>"110000100",
  65359=>"101011010",
  65360=>"111101100",
  65361=>"111000010",
  65362=>"110101001",
  65363=>"001011000",
  65364=>"001100000",
  65365=>"010101001",
  65366=>"001110000",
  65367=>"111001110",
  65368=>"011100101",
  65369=>"001101100",
  65370=>"110000110",
  65371=>"101111001",
  65372=>"101100000",
  65373=>"110111010",
  65374=>"001000011",
  65375=>"100100001",
  65376=>"110010111",
  65377=>"111110000",
  65378=>"011011001",
  65379=>"101100101",
  65380=>"111100110",
  65381=>"101010110",
  65382=>"101101011",
  65383=>"000110111",
  65384=>"110001100",
  65385=>"010010100",
  65386=>"101110101",
  65387=>"100000101",
  65388=>"011101100",
  65389=>"000111000",
  65390=>"101100110",
  65391=>"100000010",
  65392=>"111000110",
  65393=>"010000011",
  65394=>"010000110",
  65395=>"100111000",
  65396=>"100011000",
  65397=>"100111010",
  65398=>"000010010",
  65399=>"001001110",
  65400=>"100101110",
  65401=>"101001011",
  65402=>"001101010",
  65403=>"101010000",
  65404=>"000000100",
  65405=>"100010011",
  65406=>"110101000",
  65407=>"010011011",
  65408=>"010001011",
  65409=>"011001111",
  65410=>"000101011",
  65411=>"100111100",
  65412=>"011101100",
  65413=>"111011011",
  65414=>"010111101",
  65415=>"111000100",
  65416=>"101110010",
  65417=>"000101010",
  65418=>"010010011",
  65419=>"110110111",
  65420=>"110100101",
  65421=>"111001101",
  65422=>"001010010",
  65423=>"101011110",
  65424=>"110010110",
  65425=>"110101001",
  65426=>"111101000",
  65427=>"010010111",
  65428=>"111110000",
  65429=>"111110111",
  65430=>"111100100",
  65431=>"010100101",
  65432=>"110000010",
  65433=>"110100010",
  65434=>"110010110",
  65435=>"101101011",
  65436=>"100011000",
  65437=>"001001110",
  65438=>"100000001",
  65439=>"101001100",
  65440=>"111100110",
  65441=>"010110101",
  65442=>"000101011",
  65443=>"100010100",
  65444=>"100000010",
  65445=>"111010110",
  65446=>"001010101",
  65447=>"010110011",
  65448=>"011110101",
  65449=>"110000011",
  65450=>"011111011",
  65451=>"010110101",
  65452=>"101101001",
  65453=>"101001001",
  65454=>"100011110",
  65455=>"101011001",
  65456=>"100110001",
  65457=>"001100011",
  65458=>"110110110",
  65459=>"000001011",
  65460=>"101010110",
  65461=>"001110110",
  65462=>"000110111",
  65463=>"010101001",
  65464=>"000101001",
  65465=>"101101100",
  65466=>"011101011",
  65467=>"100111100",
  65468=>"111001100",
  65469=>"100100100",
  65470=>"110001110",
  65471=>"110000110",
  65472=>"011100010",
  65473=>"011100101",
  65474=>"000001100",
  65475=>"100011001",
  65476=>"000110100",
  65477=>"001100100",
  65478=>"111011000",
  65479=>"110111010",
  65480=>"001101110",
  65481=>"110011111",
  65482=>"101110010",
  65483=>"110101100",
  65484=>"011111010",
  65485=>"101111011",
  65486=>"000000111",
  65487=>"101111110",
  65488=>"110110110",
  65489=>"010000011",
  65490=>"111000001",
  65491=>"000110101",
  65492=>"111101100",
  65493=>"011100000",
  65494=>"101011101",
  65495=>"101111111",
  65496=>"001011011",
  65497=>"101110111",
  65498=>"000001000",
  65499=>"101100110",
  65500=>"011111110",
  65501=>"100011100",
  65502=>"000101110",
  65503=>"000011010",
  65504=>"001100110",
  65505=>"100010101",
  65506=>"010111110",
  65507=>"100101111",
  65508=>"110100100",
  65509=>"110000111",
  65510=>"011111101",
  65511=>"110001110",
  65512=>"101000111",
  65513=>"101110001",
  65514=>"011000110",
  65515=>"101100100",
  65516=>"000111010",
  65517=>"100100110",
  65518=>"100011000",
  65519=>"000001001",
  65520=>"110110001",
  65521=>"111110101",
  65522=>"000011000",
  65523=>"100000000",
  65524=>"010110110",
  65525=>"100111001",
  65526=>"111100111",
  65527=>"110111010",
  65528=>"000101110",
  65529=>"100111010",
  65530=>"101110110",
  65531=>"111000010",
  65532=>"110111001",
  65533=>"010001110",
  65534=>"100101100",
  65535=>"110000111");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;