LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L7_6_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(7) - 1 DOWNTO 0));
END L7_6_WROM;

ARCHITECTURE RTL OF L7_6_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"111010000",
  1=>"111111101",
  2=>"011011011",
  3=>"110110111",
  4=>"100111111",
  5=>"110000000",
  6=>"000000000",
  7=>"000001011",
  8=>"101000000",
  9=>"100000000",
  10=>"000001001",
  11=>"111111111",
  12=>"111011101",
  13=>"000000000",
  14=>"010000100",
  15=>"000000000",
  16=>"110000011",
  17=>"111001000",
  18=>"011011011",
  19=>"111111111",
  20=>"000100110",
  21=>"000100111",
  22=>"000110110",
  23=>"101000001",
  24=>"111111111",
  25=>"101101101",
  26=>"011111000",
  27=>"111111000",
  28=>"000000000",
  29=>"111111000",
  30=>"000000000",
  31=>"001000000",
  32=>"101000000",
  33=>"000000011",
  34=>"111111111",
  35=>"000000000",
  36=>"001000000",
  37=>"000010111",
  38=>"111111010",
  39=>"000000001",
  40=>"000000110",
  41=>"000000000",
  42=>"101000101",
  43=>"110100000",
  44=>"000000110",
  45=>"000010000",
  46=>"001010000",
  47=>"000010110",
  48=>"110111111",
  49=>"111111111",
  50=>"011101111",
  51=>"011010010",
  52=>"010010011",
  53=>"001001000",
  54=>"000100100",
  55=>"111101000",
  56=>"100111000",
  57=>"100100000",
  58=>"000000000",
  59=>"000011000",
  60=>"000000000",
  61=>"000000000",
  62=>"000001011",
  63=>"000000111",
  64=>"011111011",
  65=>"111110111",
  66=>"100000000",
  67=>"000100100",
  68=>"110110000",
  69=>"001001011",
  70=>"000000000",
  71=>"000000000",
  72=>"000000000",
  73=>"000000100",
  74=>"111001000",
  75=>"111111111",
  76=>"000000000",
  77=>"111111000",
  78=>"011100100",
  79=>"111111111",
  80=>"000000000",
  81=>"000000000",
  82=>"110110100",
  83=>"000000000",
  84=>"001001011",
  85=>"000000000",
  86=>"111111100",
  87=>"110100001",
  88=>"111111110",
  89=>"110000000",
  90=>"011111111",
  91=>"000000001",
  92=>"111111110",
  93=>"000000000",
  94=>"000000001",
  95=>"011011011",
  96=>"000001111",
  97=>"000000000",
  98=>"000000000",
  99=>"111011111",
  100=>"100000000",
  101=>"111111101",
  102=>"010000111",
  103=>"001001101",
  104=>"110111111",
  105=>"000001001",
  106=>"111111111",
  107=>"011011111",
  108=>"100110010",
  109=>"000000000",
  110=>"001100000",
  111=>"111111111",
  112=>"111111111",
  113=>"111111110",
  114=>"000000000",
  115=>"111111111",
  116=>"000000001",
  117=>"111111111",
  118=>"111111111",
  119=>"000000001",
  120=>"110110110",
  121=>"000000000",
  122=>"111011001",
  123=>"111111100",
  124=>"000000000",
  125=>"111111111",
  126=>"111101000",
  127=>"000000000",
  128=>"000000000",
  129=>"011011000",
  130=>"111111000",
  131=>"000010000",
  132=>"000000111",
  133=>"111101111",
  134=>"111111111",
  135=>"000000000",
  136=>"000000111",
  137=>"000000000",
  138=>"111111111",
  139=>"000000000",
  140=>"000000111",
  141=>"110111000",
  142=>"111111111",
  143=>"001000000",
  144=>"111110111",
  145=>"010011111",
  146=>"000000000",
  147=>"111101001",
  148=>"000000000",
  149=>"001111111",
  150=>"000000111",
  151=>"000000000",
  152=>"111111111",
  153=>"110110000",
  154=>"110111111",
  155=>"111000001",
  156=>"001111100",
  157=>"111111111",
  158=>"000000000",
  159=>"000111111",
  160=>"000100000",
  161=>"111111000",
  162=>"111011000",
  163=>"111111111",
  164=>"000101111",
  165=>"111111111",
  166=>"000000000",
  167=>"000000000",
  168=>"000001111",
  169=>"110110111",
  170=>"001000000",
  171=>"110000111",
  172=>"000101111",
  173=>"111111111",
  174=>"111111111",
  175=>"111111100",
  176=>"111111000",
  177=>"000100000",
  178=>"000000111",
  179=>"000000100",
  180=>"000101111",
  181=>"000000000",
  182=>"111111111",
  183=>"001101111",
  184=>"111111101",
  185=>"000000000",
  186=>"000100100",
  187=>"100110100",
  188=>"111101000",
  189=>"101100111",
  190=>"010011011",
  191=>"111111111",
  192=>"111111111",
  193=>"000000001",
  194=>"000000000",
  195=>"000111100",
  196=>"000000101",
  197=>"000000000",
  198=>"111001101",
  199=>"000000000",
  200=>"111111010",
  201=>"100000000",
  202=>"111001101",
  203=>"001011000",
  204=>"110111000",
  205=>"000000000",
  206=>"111110111",
  207=>"111110111",
  208=>"011011111",
  209=>"001000001",
  210=>"111111110",
  211=>"001001001",
  212=>"111111001",
  213=>"000000000",
  214=>"001001111",
  215=>"111111111",
  216=>"111111111",
  217=>"000000000",
  218=>"000000000",
  219=>"001111010",
  220=>"110100111",
  221=>"000001101",
  222=>"111010110",
  223=>"111110010",
  224=>"111111001",
  225=>"010010010",
  226=>"111111111",
  227=>"000000000",
  228=>"111111111",
  229=>"000000100",
  230=>"001111111",
  231=>"000000000",
  232=>"111110111",
  233=>"101111001",
  234=>"000000000",
  235=>"000000000",
  236=>"110111000",
  237=>"011011010",
  238=>"111111111",
  239=>"111000000",
  240=>"111111000",
  241=>"000000000",
  242=>"001000110",
  243=>"000000000",
  244=>"001000111",
  245=>"010010100",
  246=>"111001000",
  247=>"000000000",
  248=>"010011111",
  249=>"000110010",
  250=>"000100000",
  251=>"000000000",
  252=>"001011111",
  253=>"101111111",
  254=>"000000000",
  255=>"011011010",
  256=>"000000001",
  257=>"011001011",
  258=>"001001001",
  259=>"111111110",
  260=>"000001111",
  261=>"000000111",
  262=>"000101000",
  263=>"111111111",
  264=>"001111000",
  265=>"000001011",
  266=>"001101000",
  267=>"000000000",
  268=>"100100110",
  269=>"111111111",
  270=>"000000000",
  271=>"000011111",
  272=>"111111100",
  273=>"100100100",
  274=>"111100100",
  275=>"000111111",
  276=>"111011101",
  277=>"100000000",
  278=>"001001001",
  279=>"000000000",
  280=>"111111011",
  281=>"111001000",
  282=>"101111111",
  283=>"000000000",
  284=>"000000110",
  285=>"111111111",
  286=>"111101111",
  287=>"111111100",
  288=>"000000000",
  289=>"111111111",
  290=>"001001000",
  291=>"111111111",
  292=>"000000001",
  293=>"111111110",
  294=>"011011000",
  295=>"101000000",
  296=>"111111111",
  297=>"111111111",
  298=>"110001000",
  299=>"111111111",
  300=>"111111000",
  301=>"111010011",
  302=>"101010111",
  303=>"111111111",
  304=>"111111111",
  305=>"000000000",
  306=>"111111111",
  307=>"000001101",
  308=>"000011111",
  309=>"000000000",
  310=>"000011111",
  311=>"100000000",
  312=>"000000000",
  313=>"001010000",
  314=>"111111111",
  315=>"100111110",
  316=>"000010011",
  317=>"010000000",
  318=>"101101111",
  319=>"111111110",
  320=>"000000101",
  321=>"000010010",
  322=>"100100000",
  323=>"010010111",
  324=>"000000000",
  325=>"111000000",
  326=>"011010111",
  327=>"000000000",
  328=>"000000000",
  329=>"010000000",
  330=>"000111110",
  331=>"111111001",
  332=>"000000001",
  333=>"110111101",
  334=>"111111111",
  335=>"111111111",
  336=>"001001001",
  337=>"110110110",
  338=>"110000000",
  339=>"001111110",
  340=>"000000000",
  341=>"001011001",
  342=>"000000000",
  343=>"111111100",
  344=>"100111101",
  345=>"000000111",
  346=>"000000100",
  347=>"000000000",
  348=>"010000000",
  349=>"100000000",
  350=>"111110110",
  351=>"000111010",
  352=>"111111111",
  353=>"000000000",
  354=>"000011111",
  355=>"111111010",
  356=>"101111101",
  357=>"000000000",
  358=>"001000000",
  359=>"001011011",
  360=>"011011101",
  361=>"000001000",
  362=>"000000000",
  363=>"110111111",
  364=>"100000000",
  365=>"000000001",
  366=>"011111111",
  367=>"010000000",
  368=>"000000000",
  369=>"010000000",
  370=>"000000001",
  371=>"010001000",
  372=>"100111111",
  373=>"001000001",
  374=>"000001000",
  375=>"000010010",
  376=>"000010111",
  377=>"000000000",
  378=>"000000100",
  379=>"111001111",
  380=>"010000000",
  381=>"111111111",
  382=>"100000000",
  383=>"101000001",
  384=>"000000000",
  385=>"110111100",
  386=>"100100111",
  387=>"111111111",
  388=>"111100110",
  389=>"011000000",
  390=>"110000100",
  391=>"011011111",
  392=>"000000111",
  393=>"000000000",
  394=>"001000001",
  395=>"000011000",
  396=>"111111111",
  397=>"010110110",
  398=>"011000001",
  399=>"000000000",
  400=>"000111111",
  401=>"111101000",
  402=>"000000000",
  403=>"100110110",
  404=>"001000000",
  405=>"001101111",
  406=>"000000000",
  407=>"011110000",
  408=>"000000000",
  409=>"110110000",
  410=>"000000000",
  411=>"111111111",
  412=>"111111011",
  413=>"100000100",
  414=>"000000010",
  415=>"110000000",
  416=>"111111111",
  417=>"111111011",
  418=>"000100000",
  419=>"000000010",
  420=>"000000010",
  421=>"111111011",
  422=>"111111111",
  423=>"010011001",
  424=>"000110011",
  425=>"000000000",
  426=>"000000000",
  427=>"000000010",
  428=>"000000111",
  429=>"011101101",
  430=>"000000010",
  431=>"000000000",
  432=>"111011000",
  433=>"000000000",
  434=>"000000000",
  435=>"111111111",
  436=>"011110111",
  437=>"000000100",
  438=>"111101111",
  439=>"110100000",
  440=>"000000110",
  441=>"000001001",
  442=>"100000000",
  443=>"110110111",
  444=>"100111111",
  445=>"111000000",
  446=>"000000000",
  447=>"010000000",
  448=>"111111111",
  449=>"111001101",
  450=>"000000000",
  451=>"111000111",
  452=>"001001010",
  453=>"100101101",
  454=>"000111000",
  455=>"010110111",
  456=>"000000000",
  457=>"111111111",
  458=>"000100100",
  459=>"110111111",
  460=>"111111111",
  461=>"000000000",
  462=>"000011011",
  463=>"000110111",
  464=>"000000000",
  465=>"000111100",
  466=>"011111111",
  467=>"011001001",
  468=>"001001000",
  469=>"111111111",
  470=>"100100000",
  471=>"010010000",
  472=>"111111111",
  473=>"100000000",
  474=>"000000100",
  475=>"111111111",
  476=>"000000001",
  477=>"111100000",
  478=>"111111100",
  479=>"110110100",
  480=>"000000000",
  481=>"000000111",
  482=>"000000000",
  483=>"000000100",
  484=>"110111111",
  485=>"111111001",
  486=>"111111111",
  487=>"000000000",
  488=>"000000101",
  489=>"011111111",
  490=>"111011001",
  491=>"111111111",
  492=>"100100110",
  493=>"011011011",
  494=>"000110100",
  495=>"100100000",
  496=>"111010111",
  497=>"101000110",
  498=>"111100100",
  499=>"111111000",
  500=>"101001000",
  501=>"100111111",
  502=>"111111111",
  503=>"110111110",
  504=>"000000010",
  505=>"000000111",
  506=>"001000110",
  507=>"000000000",
  508=>"111111111",
  509=>"000000000",
  510=>"000000000",
  511=>"111111111",
  512=>"000000000",
  513=>"000000000",
  514=>"000000000",
  515=>"011011000",
  516=>"100111110",
  517=>"000000000",
  518=>"000110110",
  519=>"111111111",
  520=>"111111111",
  521=>"100100110",
  522=>"111101101",
  523=>"101111111",
  524=>"000100111",
  525=>"000100100",
  526=>"001001001",
  527=>"000000000",
  528=>"011000000",
  529=>"010110011",
  530=>"000000000",
  531=>"111111000",
  532=>"111111011",
  533=>"000000000",
  534=>"000000000",
  535=>"111110111",
  536=>"000000000",
  537=>"100100100",
  538=>"000000000",
  539=>"110111111",
  540=>"110000000",
  541=>"100011000",
  542=>"101111111",
  543=>"000110110",
  544=>"110110110",
  545=>"111111111",
  546=>"011011001",
  547=>"100001001",
  548=>"111111111",
  549=>"011111111",
  550=>"000000110",
  551=>"110000000",
  552=>"111000000",
  553=>"111111111",
  554=>"011111011",
  555=>"111111111",
  556=>"000101101",
  557=>"000000000",
  558=>"111111110",
  559=>"000000000",
  560=>"100000000",
  561=>"000000000",
  562=>"010110110",
  563=>"001001000",
  564=>"000000000",
  565=>"100000000",
  566=>"111000001",
  567=>"111101000",
  568=>"000000000",
  569=>"000000000",
  570=>"000111111",
  571=>"000000000",
  572=>"111100100",
  573=>"000100100",
  574=>"000001011",
  575=>"000000000",
  576=>"001001100",
  577=>"000000000",
  578=>"111111111",
  579=>"000000000",
  580=>"000000000",
  581=>"111110000",
  582=>"111111011",
  583=>"111111000",
  584=>"111110110",
  585=>"000000110",
  586=>"111111100",
  587=>"111111000",
  588=>"000001101",
  589=>"000110000",
  590=>"111110000",
  591=>"111111111",
  592=>"000001000",
  593=>"101001001",
  594=>"100000000",
  595=>"000000000",
  596=>"111111111",
  597=>"000000000",
  598=>"011000000",
  599=>"000000111",
  600=>"000000111",
  601=>"111011000",
  602=>"000111111",
  603=>"011111110",
  604=>"000000011",
  605=>"000000000",
  606=>"111111111",
  607=>"100100110",
  608=>"000000000",
  609=>"111111011",
  610=>"111111111",
  611=>"000000000",
  612=>"000000001",
  613=>"000000000",
  614=>"111111111",
  615=>"000000000",
  616=>"001111111",
  617=>"111111111",
  618=>"011011110",
  619=>"111111111",
  620=>"000100110",
  621=>"000000111",
  622=>"111111000",
  623=>"101001111",
  624=>"101111110",
  625=>"000001000",
  626=>"000000000",
  627=>"100001111",
  628=>"111011111",
  629=>"001000000",
  630=>"111001001",
  631=>"001000000",
  632=>"000000111",
  633=>"000000100",
  634=>"111111111",
  635=>"001001001",
  636=>"000010000",
  637=>"000000110",
  638=>"010000000",
  639=>"011000000",
  640=>"111111111",
  641=>"000001111",
  642=>"111111000",
  643=>"011011001",
  644=>"011111011",
  645=>"101000111",
  646=>"000001000",
  647=>"111111111",
  648=>"111111000",
  649=>"000000001",
  650=>"000000000",
  651=>"000110111",
  652=>"010000000",
  653=>"110010000",
  654=>"111110001",
  655=>"000000110",
  656=>"000111110",
  657=>"000110110",
  658=>"110111111",
  659=>"000000000",
  660=>"000000110",
  661=>"111110111",
  662=>"111111111",
  663=>"111000000",
  664=>"000000000",
  665=>"000000110",
  666=>"111111111",
  667=>"100100111",
  668=>"000111000",
  669=>"000100001",
  670=>"000100111",
  671=>"011111111",
  672=>"010111101",
  673=>"000000000",
  674=>"111111111",
  675=>"000110110",
  676=>"000000101",
  677=>"111110100",
  678=>"000010000",
  679=>"100110110",
  680=>"000000011",
  681=>"110111011",
  682=>"011000000",
  683=>"110111111",
  684=>"000000000",
  685=>"100000000",
  686=>"111111111",
  687=>"000001101",
  688=>"000000000",
  689=>"111111101",
  690=>"110110110",
  691=>"000000111",
  692=>"111111111",
  693=>"111111000",
  694=>"000001111",
  695=>"111111100",
  696=>"100100101",
  697=>"000111110",
  698=>"000000101",
  699=>"111111100",
  700=>"111111111",
  701=>"000000000",
  702=>"000000000",
  703=>"000000000",
  704=>"111111000",
  705=>"000000000",
  706=>"000101111",
  707=>"110110000",
  708=>"111111000",
  709=>"001000001",
  710=>"100100000",
  711=>"111111111",
  712=>"111111111",
  713=>"101100000",
  714=>"000000011",
  715=>"001111111",
  716=>"000000000",
  717=>"000111001",
  718=>"111111111",
  719=>"000000001",
  720=>"111111111",
  721=>"001001011",
  722=>"000000000",
  723=>"010000011",
  724=>"000000001",
  725=>"111111111",
  726=>"000000000",
  727=>"111101111",
  728=>"011000010",
  729=>"100100111",
  730=>"111111111",
  731=>"000000000",
  732=>"000000001",
  733=>"111000000",
  734=>"000010111",
  735=>"111111111",
  736=>"000000110",
  737=>"000000000",
  738=>"111111111",
  739=>"111101101",
  740=>"000000000",
  741=>"100100000",
  742=>"000000011",
  743=>"111000000",
  744=>"000000000",
  745=>"000001000",
  746=>"111111001",
  747=>"110000000",
  748=>"000001011",
  749=>"000000000",
  750=>"000111111",
  751=>"000000000",
  752=>"010000100",
  753=>"111111111",
  754=>"111111001",
  755=>"000001111",
  756=>"010111111",
  757=>"001001111",
  758=>"011001101",
  759=>"111111000",
  760=>"000001111",
  761=>"000000000",
  762=>"110111000",
  763=>"000000000",
  764=>"011011011",
  765=>"000000000",
  766=>"010000000",
  767=>"000000111",
  768=>"000001111",
  769=>"000101111",
  770=>"000000000",
  771=>"000000000",
  772=>"111101000",
  773=>"000000100",
  774=>"000000000",
  775=>"000000000",
  776=>"111111111",
  777=>"101001000",
  778=>"111111111",
  779=>"000000000",
  780=>"000110110",
  781=>"100100100",
  782=>"111111111",
  783=>"001011111",
  784=>"011000000",
  785=>"001000011",
  786=>"111000111",
  787=>"000000001",
  788=>"110100100",
  789=>"110011011",
  790=>"111111111",
  791=>"000000000",
  792=>"100100110",
  793=>"000000100",
  794=>"111111111",
  795=>"000000000",
  796=>"001001011",
  797=>"000111111",
  798=>"000000011",
  799=>"000000111",
  800=>"000000000",
  801=>"111111110",
  802=>"011011001",
  803=>"110111111",
  804=>"000001001",
  805=>"100000111",
  806=>"100111111",
  807=>"000000001",
  808=>"000000000",
  809=>"000000000",
  810=>"000000000",
  811=>"000000000",
  812=>"000110111",
  813=>"100111111",
  814=>"000000000",
  815=>"001000111",
  816=>"010111111",
  817=>"111111110",
  818=>"111111111",
  819=>"111111010",
  820=>"111111000",
  821=>"111111111",
  822=>"011011111",
  823=>"111000000",
  824=>"000111000",
  825=>"001001111",
  826=>"011111111",
  827=>"111111111",
  828=>"000000111",
  829=>"000000000",
  830=>"000001111",
  831=>"010111111",
  832=>"000000000",
  833=>"011011111",
  834=>"000000000",
  835=>"000000000",
  836=>"000000000",
  837=>"000000001",
  838=>"000000000",
  839=>"001011111",
  840=>"000000000",
  841=>"111000000",
  842=>"000000000",
  843=>"000011000",
  844=>"111110111",
  845=>"111011111",
  846=>"000000011",
  847=>"000000000",
  848=>"110110110",
  849=>"000000000",
  850=>"100110111",
  851=>"111111000",
  852=>"100000101",
  853=>"001011011",
  854=>"100100000",
  855=>"100000000",
  856=>"000000000",
  857=>"000000000",
  858=>"111010000",
  859=>"001001000",
  860=>"000110110",
  861=>"000101111",
  862=>"000000000",
  863=>"111111111",
  864=>"100000110",
  865=>"111111111",
  866=>"011001001",
  867=>"000000001",
  868=>"100000101",
  869=>"111000001",
  870=>"111111011",
  871=>"000000000",
  872=>"111110100",
  873=>"000000000",
  874=>"000000000",
  875=>"000000011",
  876=>"000000010",
  877=>"001111101",
  878=>"000000000",
  879=>"100000000",
  880=>"100101111",
  881=>"000000000",
  882=>"000000000",
  883=>"001001000",
  884=>"000000000",
  885=>"111110110",
  886=>"000000000",
  887=>"111111111",
  888=>"111111001",
  889=>"111000000",
  890=>"111111111",
  891=>"000010000",
  892=>"111111000",
  893=>"111010111",
  894=>"000000100",
  895=>"000111111",
  896=>"110100100",
  897=>"010100111",
  898=>"111111001",
  899=>"001000000",
  900=>"000000000",
  901=>"000000000",
  902=>"100000000",
  903=>"100001111",
  904=>"000000111",
  905=>"111111111",
  906=>"000000000",
  907=>"110111111",
  908=>"110111111",
  909=>"000000000",
  910=>"001000000",
  911=>"011011011",
  912=>"111100000",
  913=>"111000000",
  914=>"100100111",
  915=>"000000111",
  916=>"111111000",
  917=>"000000001",
  918=>"110110111",
  919=>"000000100",
  920=>"000000000",
  921=>"110000000",
  922=>"000111111",
  923=>"111000100",
  924=>"001111111",
  925=>"000000000",
  926=>"000001001",
  927=>"000000000",
  928=>"001001000",
  929=>"111111111",
  930=>"000000101",
  931=>"111111011",
  932=>"110000000",
  933=>"000001011",
  934=>"000000000",
  935=>"111111111",
  936=>"000001011",
  937=>"000000000",
  938=>"000000111",
  939=>"000000000",
  940=>"001001000",
  941=>"000100110",
  942=>"111111000",
  943=>"011010000",
  944=>"111101000",
  945=>"111101100",
  946=>"000111111",
  947=>"111111111",
  948=>"000000000",
  949=>"111111111",
  950=>"110000110",
  951=>"111111000",
  952=>"110000000",
  953=>"111111111",
  954=>"100000111",
  955=>"111111111",
  956=>"111111111",
  957=>"101101111",
  958=>"000000100",
  959=>"001001001",
  960=>"111111000",
  961=>"111111111",
  962=>"111111111",
  963=>"000000101",
  964=>"011001001",
  965=>"000000100",
  966=>"111111100",
  967=>"001000000",
  968=>"000000000",
  969=>"000000000",
  970=>"000000000",
  971=>"110110000",
  972=>"001101100",
  973=>"000000000",
  974=>"000000001",
  975=>"000111001",
  976=>"000000000",
  977=>"000000111",
  978=>"001001011",
  979=>"111011000",
  980=>"001000000",
  981=>"000000000",
  982=>"110111110",
  983=>"000011001",
  984=>"000000101",
  985=>"000000000",
  986=>"111111111",
  987=>"111111111",
  988=>"001001001",
  989=>"110111000",
  990=>"111111011",
  991=>"000000000",
  992=>"100100100",
  993=>"111111111",
  994=>"111111111",
  995=>"000000000",
  996=>"111101100",
  997=>"001000100",
  998=>"000000111",
  999=>"001000000",
  1000=>"000000000",
  1001=>"111111110",
  1002=>"110000111",
  1003=>"010000000",
  1004=>"111111111",
  1005=>"011011001",
  1006=>"000000000",
  1007=>"000000101",
  1008=>"000000000",
  1009=>"011111100",
  1010=>"111000000",
  1011=>"100000100",
  1012=>"111111111",
  1013=>"100000000",
  1014=>"000000000",
  1015=>"111111111",
  1016=>"000000101",
  1017=>"000000000",
  1018=>"111111111",
  1019=>"111111111",
  1020=>"011000111",
  1021=>"110000110",
  1022=>"111111111",
  1023=>"101110000",
  1024=>"110010000",
  1025=>"011001100",
  1026=>"010010010",
  1027=>"000111000",
  1028=>"111101001",
  1029=>"010000110",
  1030=>"001000000",
  1031=>"000000100",
  1032=>"111111010",
  1033=>"111110110",
  1034=>"100000111",
  1035=>"001001111",
  1036=>"000000000",
  1037=>"011001000",
  1038=>"110110000",
  1039=>"111111110",
  1040=>"111111011",
  1041=>"000110111",
  1042=>"100000010",
  1043=>"111100000",
  1044=>"011001111",
  1045=>"100111000",
  1046=>"001011011",
  1047=>"100000111",
  1048=>"011111110",
  1049=>"100001000",
  1050=>"110100101",
  1051=>"111111111",
  1052=>"111111111",
  1053=>"111010010",
  1054=>"000000001",
  1055=>"111000000",
  1056=>"000000000",
  1057=>"000000001",
  1058=>"100000111",
  1059=>"111111111",
  1060=>"011111111",
  1061=>"111100100",
  1062=>"110010110",
  1063=>"001000000",
  1064=>"111111111",
  1065=>"000100111",
  1066=>"111111111",
  1067=>"001001000",
  1068=>"011001111",
  1069=>"000100100",
  1070=>"011111111",
  1071=>"000010000",
  1072=>"000000111",
  1073=>"000000000",
  1074=>"000000101",
  1075=>"100110100",
  1076=>"000000000",
  1077=>"000100011",
  1078=>"100110111",
  1079=>"011010010",
  1080=>"101000111",
  1081=>"000011111",
  1082=>"111101001",
  1083=>"011011011",
  1084=>"000000111",
  1085=>"111111111",
  1086=>"110110111",
  1087=>"011111111",
  1088=>"001011111",
  1089=>"000010000",
  1090=>"011101111",
  1091=>"111111110",
  1092=>"000111110",
  1093=>"001101100",
  1094=>"000000111",
  1095=>"010010000",
  1096=>"001001011",
  1097=>"100100100",
  1098=>"000000000",
  1099=>"110110111",
  1100=>"000000110",
  1101=>"101101111",
  1102=>"111000000",
  1103=>"111111111",
  1104=>"111001000",
  1105=>"111111011",
  1106=>"000000000",
  1107=>"110110100",
  1108=>"000000000",
  1109=>"111111000",
  1110=>"111111001",
  1111=>"100000000",
  1112=>"111111000",
  1113=>"000000100",
  1114=>"001011000",
  1115=>"100000000",
  1116=>"111111111",
  1117=>"000000000",
  1118=>"000000011",
  1119=>"001011111",
  1120=>"000000000",
  1121=>"111010000",
  1122=>"111101101",
  1123=>"111001000",
  1124=>"000000100",
  1125=>"000001011",
  1126=>"111000000",
  1127=>"111110111",
  1128=>"111111001",
  1129=>"110110110",
  1130=>"000000000",
  1131=>"001111110",
  1132=>"100010001",
  1133=>"000000111",
  1134=>"001101111",
  1135=>"101000000",
  1136=>"011000000",
  1137=>"000001011",
  1138=>"011011011",
  1139=>"111111111",
  1140=>"111110000",
  1141=>"000000000",
  1142=>"111111111",
  1143=>"000111011",
  1144=>"001000000",
  1145=>"111111111",
  1146=>"100110000",
  1147=>"011111011",
  1148=>"101001101",
  1149=>"000000000",
  1150=>"100110110",
  1151=>"000101100",
  1152=>"111000111",
  1153=>"111110110",
  1154=>"110110010",
  1155=>"011011001",
  1156=>"100000000",
  1157=>"000000000",
  1158=>"000000000",
  1159=>"001001000",
  1160=>"111111000",
  1161=>"000110010",
  1162=>"111111101",
  1163=>"000000000",
  1164=>"111111111",
  1165=>"001111111",
  1166=>"111111101",
  1167=>"111101111",
  1168=>"011011111",
  1169=>"000100100",
  1170=>"011001000",
  1171=>"011000000",
  1172=>"000000000",
  1173=>"000000011",
  1174=>"001001001",
  1175=>"010010000",
  1176=>"000010110",
  1177=>"010000110",
  1178=>"101000000",
  1179=>"000000000",
  1180=>"001011111",
  1181=>"111100110",
  1182=>"111110110",
  1183=>"111110110",
  1184=>"100000110",
  1185=>"110010000",
  1186=>"000000000",
  1187=>"000000001",
  1188=>"000000001",
  1189=>"011000000",
  1190=>"000001111",
  1191=>"101001000",
  1192=>"000000000",
  1193=>"111111111",
  1194=>"001011001",
  1195=>"111000111",
  1196=>"111101101",
  1197=>"000000000",
  1198=>"100100111",
  1199=>"110111000",
  1200=>"000111111",
  1201=>"000001001",
  1202=>"000101101",
  1203=>"111111000",
  1204=>"000000100",
  1205=>"000111000",
  1206=>"101101000",
  1207=>"111010000",
  1208=>"110000000",
  1209=>"000010010",
  1210=>"000000110",
  1211=>"000011011",
  1212=>"101101101",
  1213=>"001001000",
  1214=>"000110100",
  1215=>"001000000",
  1216=>"110100100",
  1217=>"000000001",
  1218=>"000000000",
  1219=>"111101000",
  1220=>"111111000",
  1221=>"000010110",
  1222=>"100010010",
  1223=>"110111111",
  1224=>"101111111",
  1225=>"111111111",
  1226=>"111111111",
  1227=>"011111111",
  1228=>"011111001",
  1229=>"000111011",
  1230=>"000101000",
  1231=>"001001000",
  1232=>"000000000",
  1233=>"101101111",
  1234=>"000010000",
  1235=>"101001101",
  1236=>"000011011",
  1237=>"111111111",
  1238=>"000010010",
  1239=>"000100100",
  1240=>"001000111",
  1241=>"111111001",
  1242=>"000000000",
  1243=>"001111111",
  1244=>"000000000",
  1245=>"100001111",
  1246=>"000000000",
  1247=>"010011000",
  1248=>"111111110",
  1249=>"011111111",
  1250=>"111111011",
  1251=>"011011000",
  1252=>"111111000",
  1253=>"001001001",
  1254=>"011010001",
  1255=>"111111011",
  1256=>"000000101",
  1257=>"101001000",
  1258=>"111101111",
  1259=>"111111101",
  1260=>"110000000",
  1261=>"001001001",
  1262=>"111111111",
  1263=>"111010000",
  1264=>"110110001",
  1265=>"000000100",
  1266=>"111010000",
  1267=>"111111001",
  1268=>"111111111",
  1269=>"100110111",
  1270=>"100100001",
  1271=>"111011011",
  1272=>"111101111",
  1273=>"100100100",
  1274=>"001001000",
  1275=>"111110000",
  1276=>"101000001",
  1277=>"000011010",
  1278=>"000000000",
  1279=>"010000000",
  1280=>"000000000",
  1281=>"000000100",
  1282=>"000000000",
  1283=>"000111111",
  1284=>"000000000",
  1285=>"001000010",
  1286=>"100111111",
  1287=>"111111001",
  1288=>"001001100",
  1289=>"111111100",
  1290=>"111011111",
  1291=>"100000110",
  1292=>"110100000",
  1293=>"000000000",
  1294=>"111011111",
  1295=>"000000000",
  1296=>"000101001",
  1297=>"111111000",
  1298=>"000000000",
  1299=>"111000110",
  1300=>"111111001",
  1301=>"100100111",
  1302=>"000100100",
  1303=>"000000110",
  1304=>"001101100",
  1305=>"011101000",
  1306=>"111110000",
  1307=>"001111111",
  1308=>"000000001",
  1309=>"111001001",
  1310=>"000000000",
  1311=>"110000111",
  1312=>"010010001",
  1313=>"111111001",
  1314=>"001000000",
  1315=>"100111111",
  1316=>"000000101",
  1317=>"111111111",
  1318=>"101001001",
  1319=>"011110110",
  1320=>"001000100",
  1321=>"110111110",
  1322=>"010011001",
  1323=>"011010111",
  1324=>"101101000",
  1325=>"110000000",
  1326=>"011000000",
  1327=>"000000000",
  1328=>"111111000",
  1329=>"111111000",
  1330=>"111011111",
  1331=>"111000011",
  1332=>"000010000",
  1333=>"000110111",
  1334=>"000000000",
  1335=>"111111111",
  1336=>"000000000",
  1337=>"001100111",
  1338=>"001001111",
  1339=>"111110010",
  1340=>"111111011",
  1341=>"011110000",
  1342=>"101101101",
  1343=>"001000001",
  1344=>"000000000",
  1345=>"100000000",
  1346=>"111111111",
  1347=>"000000000",
  1348=>"001000000",
  1349=>"101101110",
  1350=>"000000000",
  1351=>"000010011",
  1352=>"100111111",
  1353=>"000010011",
  1354=>"011111111",
  1355=>"101001001",
  1356=>"100011000",
  1357=>"111000111",
  1358=>"110000000",
  1359=>"111101101",
  1360=>"001001001",
  1361=>"001000000",
  1362=>"000010111",
  1363=>"111000100",
  1364=>"101000100",
  1365=>"011011011",
  1366=>"101111111",
  1367=>"111111000",
  1368=>"111000100",
  1369=>"111111011",
  1370=>"000000000",
  1371=>"000000000",
  1372=>"111000000",
  1373=>"110110110",
  1374=>"000110100",
  1375=>"000000111",
  1376=>"010011111",
  1377=>"000001101",
  1378=>"000000000",
  1379=>"111000000",
  1380=>"000000000",
  1381=>"111011111",
  1382=>"010010110",
  1383=>"001000000",
  1384=>"001000100",
  1385=>"000000000",
  1386=>"001011111",
  1387=>"111111111",
  1388=>"010011001",
  1389=>"000000000",
  1390=>"111101111",
  1391=>"111111011",
  1392=>"000000111",
  1393=>"000000000",
  1394=>"111111010",
  1395=>"110001001",
  1396=>"111111111",
  1397=>"000000001",
  1398=>"101011111",
  1399=>"111111100",
  1400=>"000000011",
  1401=>"111011101",
  1402=>"001000100",
  1403=>"000011001",
  1404=>"100101111",
  1405=>"111011101",
  1406=>"111111111",
  1407=>"111101101",
  1408=>"001001001",
  1409=>"011000111",
  1410=>"100001001",
  1411=>"111111111",
  1412=>"111000000",
  1413=>"000000000",
  1414=>"000000010",
  1415=>"000011111",
  1416=>"000000000",
  1417=>"000000101",
  1418=>"101000000",
  1419=>"010111111",
  1420=>"111111111",
  1421=>"100010100",
  1422=>"100100101",
  1423=>"100000110",
  1424=>"000100101",
  1425=>"111111111",
  1426=>"111111001",
  1427=>"101111110",
  1428=>"101101111",
  1429=>"000000001",
  1430=>"101101000",
  1431=>"000010010",
  1432=>"111010100",
  1433=>"000000000",
  1434=>"111001110",
  1435=>"000000000",
  1436=>"000001101",
  1437=>"111110110",
  1438=>"000010010",
  1439=>"111111111",
  1440=>"100100111",
  1441=>"111111111",
  1442=>"110010001",
  1443=>"111000000",
  1444=>"011011111",
  1445=>"111111000",
  1446=>"000000000",
  1447=>"111111111",
  1448=>"000000000",
  1449=>"000111111",
  1450=>"000011000",
  1451=>"000000000",
  1452=>"101111111",
  1453=>"000001000",
  1454=>"111011111",
  1455=>"000000000",
  1456=>"000111111",
  1457=>"101101111",
  1458=>"111110110",
  1459=>"111111100",
  1460=>"110000010",
  1461=>"110110111",
  1462=>"000000100",
  1463=>"111111111",
  1464=>"011011010",
  1465=>"111000001",
  1466=>"001111101",
  1467=>"000000000",
  1468=>"101100110",
  1469=>"111111111",
  1470=>"110010000",
  1471=>"000000000",
  1472=>"010111000",
  1473=>"111111111",
  1474=>"111001000",
  1475=>"111111111",
  1476=>"111011010",
  1477=>"000000000",
  1478=>"011000000",
  1479=>"111110000",
  1480=>"000011000",
  1481=>"000000000",
  1482=>"010110010",
  1483=>"000000111",
  1484=>"000000000",
  1485=>"111111010",
  1486=>"010010010",
  1487=>"000010111",
  1488=>"010011001",
  1489=>"000000000",
  1490=>"001001011",
  1491=>"111101111",
  1492=>"110110110",
  1493=>"000000000",
  1494=>"000011010",
  1495=>"111111100",
  1496=>"000000011",
  1497=>"011111001",
  1498=>"111111111",
  1499=>"000000100",
  1500=>"100100111",
  1501=>"111001111",
  1502=>"111100000",
  1503=>"110100000",
  1504=>"000000111",
  1505=>"100000101",
  1506=>"111000001",
  1507=>"011000100",
  1508=>"110111111",
  1509=>"010000000",
  1510=>"111110010",
  1511=>"001001111",
  1512=>"111111111",
  1513=>"111111111",
  1514=>"111011111",
  1515=>"100100100",
  1516=>"011001111",
  1517=>"010000000",
  1518=>"101111111",
  1519=>"100100000",
  1520=>"111111000",
  1521=>"110110110",
  1522=>"111111111",
  1523=>"010000000",
  1524=>"111111000",
  1525=>"000000000",
  1526=>"010110111",
  1527=>"011011011",
  1528=>"011000000",
  1529=>"000100000",
  1530=>"000100110",
  1531=>"000000000",
  1532=>"111111110",
  1533=>"000010111",
  1534=>"011010000",
  1535=>"000000000",
  1536=>"110110110",
  1537=>"101001001",
  1538=>"111111111",
  1539=>"111011011",
  1540=>"101000000",
  1541=>"010111010",
  1542=>"100100111",
  1543=>"011111111",
  1544=>"101101111",
  1545=>"000000010",
  1546=>"000000000",
  1547=>"000000101",
  1548=>"001001111",
  1549=>"111111111",
  1550=>"010010111",
  1551=>"000111110",
  1552=>"100000000",
  1553=>"000000000",
  1554=>"111110110",
  1555=>"000000100",
  1556=>"000100101",
  1557=>"101101111",
  1558=>"101111011",
  1559=>"100001001",
  1560=>"100000000",
  1561=>"110011011",
  1562=>"001101111",
  1563=>"110010000",
  1564=>"001001101",
  1565=>"111000000",
  1566=>"001001001",
  1567=>"111101110",
  1568=>"000111111",
  1569=>"110000000",
  1570=>"011111111",
  1571=>"001011111",
  1572=>"101001000",
  1573=>"101001000",
  1574=>"010000000",
  1575=>"000000000",
  1576=>"100000000",
  1577=>"101101101",
  1578=>"011001011",
  1579=>"010011001",
  1580=>"001101111",
  1581=>"010001010",
  1582=>"010010010",
  1583=>"101101000",
  1584=>"011001111",
  1585=>"001000000",
  1586=>"001001100",
  1587=>"111111111",
  1588=>"001100100",
  1589=>"010010000",
  1590=>"000010011",
  1591=>"000001111",
  1592=>"110110101",
  1593=>"000000100",
  1594=>"101001001",
  1595=>"000000000",
  1596=>"100000000",
  1597=>"011001100",
  1598=>"010001000",
  1599=>"001000100",
  1600=>"000000001",
  1601=>"101101101",
  1602=>"101000000",
  1603=>"101001001",
  1604=>"000000010",
  1605=>"000000000",
  1606=>"100101111",
  1607=>"011010000",
  1608=>"000001001",
  1609=>"000000100",
  1610=>"111111111",
  1611=>"110110110",
  1612=>"000100100",
  1613=>"000101111",
  1614=>"011011011",
  1615=>"000111000",
  1616=>"111010000",
  1617=>"000101001",
  1618=>"111111111",
  1619=>"010110110",
  1620=>"010010000",
  1621=>"011111111",
  1622=>"001001111",
  1623=>"001001000",
  1624=>"101001000",
  1625=>"101101101",
  1626=>"111111100",
  1627=>"100110111",
  1628=>"101111000",
  1629=>"111111111",
  1630=>"111001111",
  1631=>"011011011",
  1632=>"100100111",
  1633=>"001001111",
  1634=>"111111111",
  1635=>"101101111",
  1636=>"100000001",
  1637=>"110110010",
  1638=>"111111110",
  1639=>"100000000",
  1640=>"111111111",
  1641=>"000000111",
  1642=>"000100101",
  1643=>"111111111",
  1644=>"110110100",
  1645=>"111111000",
  1646=>"100000000",
  1647=>"101001001",
  1648=>"001011111",
  1649=>"111000101",
  1650=>"010011010",
  1651=>"111111100",
  1652=>"000000000",
  1653=>"010000010",
  1654=>"000000101",
  1655=>"010000000",
  1656=>"000101110",
  1657=>"001001000",
  1658=>"101000000",
  1659=>"001011000",
  1660=>"000100100",
  1661=>"100100000",
  1662=>"111101100",
  1663=>"000010000",
  1664=>"101000000",
  1665=>"001111111",
  1666=>"000101100",
  1667=>"011111110",
  1668=>"111011011",
  1669=>"100001001",
  1670=>"100000110",
  1671=>"100100100",
  1672=>"100100000",
  1673=>"111111111",
  1674=>"100100100",
  1675=>"111001101",
  1676=>"111111000",
  1677=>"000000000",
  1678=>"000001101",
  1679=>"000000000",
  1680=>"000001101",
  1681=>"010110000",
  1682=>"000111111",
  1683=>"111100000",
  1684=>"101001100",
  1685=>"100111110",
  1686=>"101111111",
  1687=>"000000000",
  1688=>"001000100",
  1689=>"111011011",
  1690=>"001101111",
  1691=>"011011111",
  1692=>"101111111",
  1693=>"110110110",
  1694=>"001111100",
  1695=>"111111111",
  1696=>"001001101",
  1697=>"000000101",
  1698=>"101101111",
  1699=>"000000000",
  1700=>"001001001",
  1701=>"100100000",
  1702=>"111111110",
  1703=>"011011000",
  1704=>"101101101",
  1705=>"001111111",
  1706=>"111000000",
  1707=>"101111000",
  1708=>"100000000",
  1709=>"001000000",
  1710=>"111111111",
  1711=>"000010010",
  1712=>"000111111",
  1713=>"100100000",
  1714=>"111111010",
  1715=>"111111100",
  1716=>"001100000",
  1717=>"100100111",
  1718=>"001001000",
  1719=>"111101111",
  1720=>"100000001",
  1721=>"101101000",
  1722=>"101001101",
  1723=>"101101111",
  1724=>"000000001",
  1725=>"111001111",
  1726=>"010110011",
  1727=>"110110110",
  1728=>"111111011",
  1729=>"011101001",
  1730=>"111110100",
  1731=>"000001000",
  1732=>"111010111",
  1733=>"011011010",
  1734=>"110000000",
  1735=>"000010011",
  1736=>"101101001",
  1737=>"101111011",
  1738=>"000000000",
  1739=>"101101101",
  1740=>"001001111",
  1741=>"100101000",
  1742=>"100101111",
  1743=>"101001001",
  1744=>"100111111",
  1745=>"111111111",
  1746=>"101101000",
  1747=>"101100101",
  1748=>"111001000",
  1749=>"001000111",
  1750=>"010010110",
  1751=>"100101001",
  1752=>"000000000",
  1753=>"111101001",
  1754=>"000000111",
  1755=>"100000101",
  1756=>"000000000",
  1757=>"010110110",
  1758=>"101101101",
  1759=>"000001001",
  1760=>"111101101",
  1761=>"111000111",
  1762=>"101101110",
  1763=>"000000111",
  1764=>"110110110",
  1765=>"000001111",
  1766=>"111011010",
  1767=>"101110100",
  1768=>"100000000",
  1769=>"110110110",
  1770=>"111111100",
  1771=>"101001101",
  1772=>"101100111",
  1773=>"101111111",
  1774=>"101001111",
  1775=>"000111011",
  1776=>"011011011",
  1777=>"000010111",
  1778=>"111111111",
  1779=>"111001101",
  1780=>"000001111",
  1781=>"110110110",
  1782=>"110010010",
  1783=>"000110110",
  1784=>"111001101",
  1785=>"000000000",
  1786=>"111111111",
  1787=>"000100110",
  1788=>"101001001",
  1789=>"100110011",
  1790=>"100100100",
  1791=>"001100101",
  1792=>"000000100",
  1793=>"100100000",
  1794=>"111111111",
  1795=>"001111111",
  1796=>"111111111",
  1797=>"111111111",
  1798=>"001000000",
  1799=>"001000101",
  1800=>"001001101",
  1801=>"101100100",
  1802=>"101000010",
  1803=>"111111111",
  1804=>"110100110",
  1805=>"110110010",
  1806=>"100000111",
  1807=>"000010000",
  1808=>"101000000",
  1809=>"000001001",
  1810=>"000000000",
  1811=>"000100101",
  1812=>"101111001",
  1813=>"100000000",
  1814=>"001001001",
  1815=>"110110110",
  1816=>"110110000",
  1817=>"111111111",
  1818=>"001001000",
  1819=>"001101111",
  1820=>"100101001",
  1821=>"001000100",
  1822=>"111111111",
  1823=>"111111000",
  1824=>"011010110",
  1825=>"010110010",
  1826=>"011111111",
  1827=>"000000000",
  1828=>"000010010",
  1829=>"000101101",
  1830=>"100111100",
  1831=>"110110010",
  1832=>"111100010",
  1833=>"110111111",
  1834=>"011111101",
  1835=>"001011000",
  1836=>"000000000",
  1837=>"110110010",
  1838=>"111010011",
  1839=>"111000011",
  1840=>"010110010",
  1841=>"000000000",
  1842=>"111111111",
  1843=>"100000000",
  1844=>"111111111",
  1845=>"001111010",
  1846=>"000000000",
  1847=>"110110111",
  1848=>"111001000",
  1849=>"101000101",
  1850=>"101101101",
  1851=>"101101001",
  1852=>"111111111",
  1853=>"110000010",
  1854=>"000000000",
  1855=>"111111111",
  1856=>"011111111",
  1857=>"011111111",
  1858=>"000101101",
  1859=>"011110010",
  1860=>"001111111",
  1861=>"111101111",
  1862=>"101101000",
  1863=>"000000010",
  1864=>"101101101",
  1865=>"001100111",
  1866=>"000000001",
  1867=>"101100000",
  1868=>"000111111",
  1869=>"101101111",
  1870=>"101101001",
  1871=>"111110110",
  1872=>"001111110",
  1873=>"000100001",
  1874=>"000000000",
  1875=>"100101111",
  1876=>"000111111",
  1877=>"101011011",
  1878=>"101111111",
  1879=>"001001000",
  1880=>"000000101",
  1881=>"111111111",
  1882=>"000000000",
  1883=>"001000101",
  1884=>"011000010",
  1885=>"111111111",
  1886=>"000110110",
  1887=>"110110110",
  1888=>"000000000",
  1889=>"010010011",
  1890=>"100100100",
  1891=>"101000001",
  1892=>"000000000",
  1893=>"111111010",
  1894=>"010011111",
  1895=>"111011011",
  1896=>"101001000",
  1897=>"001001101",
  1898=>"000110111",
  1899=>"101110110",
  1900=>"111110011",
  1901=>"111111000",
  1902=>"101101101",
  1903=>"000000000",
  1904=>"000101111",
  1905=>"000000100",
  1906=>"101100100",
  1907=>"111011111",
  1908=>"001100000",
  1909=>"101110111",
  1910=>"111101101",
  1911=>"001001000",
  1912=>"111001000",
  1913=>"111100100",
  1914=>"000100100",
  1915=>"001000000",
  1916=>"000000000",
  1917=>"110100000",
  1918=>"000011111",
  1919=>"111101101",
  1920=>"001000110",
  1921=>"101101111",
  1922=>"000000000",
  1923=>"000101101",
  1924=>"111111111",
  1925=>"000100110",
  1926=>"010010010",
  1927=>"101101100",
  1928=>"101001101",
  1929=>"000010000",
  1930=>"010111000",
  1931=>"001000000",
  1932=>"000000000",
  1933=>"000000000",
  1934=>"111001111",
  1935=>"011011010",
  1936=>"101111110",
  1937=>"000100111",
  1938=>"000000000",
  1939=>"000101111",
  1940=>"010010011",
  1941=>"000000001",
  1942=>"110111000",
  1943=>"110111011",
  1944=>"001111111",
  1945=>"001000000",
  1946=>"001001001",
  1947=>"111110110",
  1948=>"000000000",
  1949=>"000000001",
  1950=>"001011001",
  1951=>"000101111",
  1952=>"101101111",
  1953=>"011011011",
  1954=>"111111001",
  1955=>"111101100",
  1956=>"011011011",
  1957=>"111101000",
  1958=>"111110010",
  1959=>"101111111",
  1960=>"101000000",
  1961=>"001001001",
  1962=>"110110111",
  1963=>"000100000",
  1964=>"001000000",
  1965=>"101101100",
  1966=>"000000000",
  1967=>"010000000",
  1968=>"111001000",
  1969=>"011111111",
  1970=>"111111111",
  1971=>"000100000",
  1972=>"001111101",
  1973=>"101101001",
  1974=>"111111111",
  1975=>"001000001",
  1976=>"101001101",
  1977=>"000000001",
  1978=>"101100110",
  1979=>"000110110",
  1980=>"111111101",
  1981=>"111111111",
  1982=>"000010111",
  1983=>"011001001",
  1984=>"000000101",
  1985=>"111111111",
  1986=>"111111111",
  1987=>"000101110",
  1988=>"000000000",
  1989=>"001001011",
  1990=>"001001001",
  1991=>"001001100",
  1992=>"001101100",
  1993=>"100000000",
  1994=>"101001001",
  1995=>"111111100",
  1996=>"001001100",
  1997=>"010110010",
  1998=>"001001001",
  1999=>"000101111",
  2000=>"001001111",
  2001=>"111111011",
  2002=>"000000000",
  2003=>"001001000",
  2004=>"001001100",
  2005=>"010010010",
  2006=>"100010010",
  2007=>"100111111",
  2008=>"011011010",
  2009=>"010010000",
  2010=>"111000001",
  2011=>"101111110",
  2012=>"111111111",
  2013=>"101100101",
  2014=>"010011111",
  2015=>"100110100",
  2016=>"101001111",
  2017=>"111110100",
  2018=>"111111111",
  2019=>"100000000",
  2020=>"001001000",
  2021=>"100000000",
  2022=>"000000000",
  2023=>"000001001",
  2024=>"000000000",
  2025=>"001001000",
  2026=>"111000000",
  2027=>"000010010",
  2028=>"101111111",
  2029=>"100111001",
  2030=>"000001111",
  2031=>"101001001",
  2032=>"101101101",
  2033=>"000011011",
  2034=>"111001001",
  2035=>"000101101",
  2036=>"111111000",
  2037=>"000000000",
  2038=>"101101111",
  2039=>"000110110",
  2040=>"100100100",
  2041=>"110110100",
  2042=>"111001010",
  2043=>"000110100",
  2044=>"011001111",
  2045=>"000000000",
  2046=>"001011011",
  2047=>"111111111",
  2048=>"001000000",
  2049=>"111110000",
  2050=>"100000111",
  2051=>"110110010",
  2052=>"011011001",
  2053=>"001011111",
  2054=>"000110000",
  2055=>"001000000",
  2056=>"111111001",
  2057=>"000000010",
  2058=>"100000101",
  2059=>"111111111",
  2060=>"000001000",
  2061=>"001000010",
  2062=>"001001010",
  2063=>"000000000",
  2064=>"110111111",
  2065=>"111100101",
  2066=>"111111111",
  2067=>"010011111",
  2068=>"111101111",
  2069=>"000000000",
  2070=>"001001111",
  2071=>"100000000",
  2072=>"100110111",
  2073=>"000110110",
  2074=>"000000101",
  2075=>"110011000",
  2076=>"111000001",
  2077=>"001001111",
  2078=>"100101111",
  2079=>"000100000",
  2080=>"111110110",
  2081=>"000011011",
  2082=>"101111111",
  2083=>"000110011",
  2084=>"001001101",
  2085=>"111001001",
  2086=>"100000100",
  2087=>"000000111",
  2088=>"110000001",
  2089=>"101000000",
  2090=>"000001111",
  2091=>"000000001",
  2092=>"000000101",
  2093=>"110110110",
  2094=>"111000001",
  2095=>"000000000",
  2096=>"001011000",
  2097=>"011111000",
  2098=>"011011011",
  2099=>"110100010",
  2100=>"000000000",
  2101=>"001001111",
  2102=>"100001111",
  2103=>"001001001",
  2104=>"000001111",
  2105=>"001001101",
  2106=>"000000000",
  2107=>"000000000",
  2108=>"001101111",
  2109=>"111111111",
  2110=>"000000001",
  2111=>"010000010",
  2112=>"111111111",
  2113=>"011011010",
  2114=>"000000110",
  2115=>"111111010",
  2116=>"001011111",
  2117=>"001101100",
  2118=>"111111111",
  2119=>"100000100",
  2120=>"010000011",
  2121=>"001000111",
  2122=>"110110000",
  2123=>"000001101",
  2124=>"001001001",
  2125=>"001111001",
  2126=>"000000000",
  2127=>"100100000",
  2128=>"101111111",
  2129=>"000000010",
  2130=>"111111111",
  2131=>"100100100",
  2132=>"010110000",
  2133=>"010111110",
  2134=>"100000000",
  2135=>"111000000",
  2136=>"000000000",
  2137=>"001001111",
  2138=>"001001001",
  2139=>"100000000",
  2140=>"101001011",
  2141=>"100111111",
  2142=>"001000000",
  2143=>"001001000",
  2144=>"111111111",
  2145=>"100001001",
  2146=>"101111111",
  2147=>"111101110",
  2148=>"000000000",
  2149=>"000000010",
  2150=>"111111011",
  2151=>"000000001",
  2152=>"111110101",
  2153=>"111000010",
  2154=>"111011011",
  2155=>"111111110",
  2156=>"111101111",
  2157=>"110000000",
  2158=>"000000000",
  2159=>"010111111",
  2160=>"001000010",
  2161=>"011010000",
  2162=>"000011111",
  2163=>"111000000",
  2164=>"111110000",
  2165=>"000000110",
  2166=>"001000000",
  2167=>"001000101",
  2168=>"101000111",
  2169=>"000001111",
  2170=>"011011011",
  2171=>"101111101",
  2172=>"001111111",
  2173=>"000000011",
  2174=>"000000000",
  2175=>"000000111",
  2176=>"001000000",
  2177=>"100100100",
  2178=>"101111011",
  2179=>"000000011",
  2180=>"111111101",
  2181=>"111111000",
  2182=>"110110000",
  2183=>"111011111",
  2184=>"000000000",
  2185=>"000000000",
  2186=>"111111110",
  2187=>"110111010",
  2188=>"110111111",
  2189=>"111111111",
  2190=>"000010101",
  2191=>"000000000",
  2192=>"101000101",
  2193=>"110000100",
  2194=>"111000000",
  2195=>"000000110",
  2196=>"001000000",
  2197=>"111100000",
  2198=>"111110111",
  2199=>"000000000",
  2200=>"001000000",
  2201=>"111111010",
  2202=>"100000000",
  2203=>"011011011",
  2204=>"001101111",
  2205=>"011001101",
  2206=>"101111011",
  2207=>"000000000",
  2208=>"001000000",
  2209=>"000000111",
  2210=>"100100000",
  2211=>"000000100",
  2212=>"111001001",
  2213=>"111111111",
  2214=>"001000000",
  2215=>"110100111",
  2216=>"000001000",
  2217=>"001011000",
  2218=>"011000000",
  2219=>"001001001",
  2220=>"111111110",
  2221=>"111111011",
  2222=>"110111111",
  2223=>"111111111",
  2224=>"111001001",
  2225=>"111111001",
  2226=>"101000001",
  2227=>"011100111",
  2228=>"000000110",
  2229=>"000111110",
  2230=>"001001000",
  2231=>"000000100",
  2232=>"101001100",
  2233=>"011011011",
  2234=>"111101001",
  2235=>"111111111",
  2236=>"001000011",
  2237=>"000100000",
  2238=>"000000010",
  2239=>"001001000",
  2240=>"000000000",
  2241=>"100100100",
  2242=>"111111111",
  2243=>"001000000",
  2244=>"011111111",
  2245=>"000000000",
  2246=>"000000001",
  2247=>"001000001",
  2248=>"010110110",
  2249=>"000000000",
  2250=>"000000101",
  2251=>"111111110",
  2252=>"110111101",
  2253=>"010100000",
  2254=>"000110111",
  2255=>"111111100",
  2256=>"111110100",
  2257=>"111001000",
  2258=>"000100000",
  2259=>"001001001",
  2260=>"111111000",
  2261=>"011011011",
  2262=>"111000000",
  2263=>"111010000",
  2264=>"001111000",
  2265=>"000010010",
  2266=>"011000111",
  2267=>"101111111",
  2268=>"000000000",
  2269=>"111111111",
  2270=>"001000001",
  2271=>"000010100",
  2272=>"111011011",
  2273=>"010010000",
  2274=>"001000101",
  2275=>"110110001",
  2276=>"001011011",
  2277=>"100100100",
  2278=>"110111111",
  2279=>"101001111",
  2280=>"001000111",
  2281=>"000010111",
  2282=>"001101111",
  2283=>"111100111",
  2284=>"000000000",
  2285=>"001001111",
  2286=>"111101111",
  2287=>"001010111",
  2288=>"000000000",
  2289=>"001111001",
  2290=>"101001001",
  2291=>"101000000",
  2292=>"000000011",
  2293=>"000101011",
  2294=>"100000100",
  2295=>"011000001",
  2296=>"111111110",
  2297=>"000111010",
  2298=>"000000001",
  2299=>"110110000",
  2300=>"001001101",
  2301=>"100101001",
  2302=>"100111111",
  2303=>"111000000",
  2304=>"000000000",
  2305=>"101001000",
  2306=>"110110111",
  2307=>"000000000",
  2308=>"001000000",
  2309=>"000011111",
  2310=>"001000100",
  2311=>"000010010",
  2312=>"000000000",
  2313=>"011111111",
  2314=>"110111111",
  2315=>"111001000",
  2316=>"001000001",
  2317=>"011000111",
  2318=>"000010011",
  2319=>"111111111",
  2320=>"001001011",
  2321=>"111111111",
  2322=>"111101111",
  2323=>"110000000",
  2324=>"000000000",
  2325=>"000001011",
  2326=>"001100110",
  2327=>"000000001",
  2328=>"000001100",
  2329=>"001001011",
  2330=>"101001000",
  2331=>"000101111",
  2332=>"100000100",
  2333=>"111110100",
  2334=>"111111000",
  2335=>"000000000",
  2336=>"011001000",
  2337=>"100001111",
  2338=>"111111111",
  2339=>"001011011",
  2340=>"011111101",
  2341=>"000000010",
  2342=>"000000000",
  2343=>"000000000",
  2344=>"000000000",
  2345=>"110111010",
  2346=>"111011111",
  2347=>"110110011",
  2348=>"001011111",
  2349=>"101111111",
  2350=>"000001000",
  2351=>"100101111",
  2352=>"001000001",
  2353=>"101001000",
  2354=>"111111101",
  2355=>"000011010",
  2356=>"000100011",
  2357=>"111111111",
  2358=>"001000100",
  2359=>"111111000",
  2360=>"001001101",
  2361=>"111000000",
  2362=>"001001001",
  2363=>"000000000",
  2364=>"001001001",
  2365=>"001001000",
  2366=>"111101001",
  2367=>"000000100",
  2368=>"001011111",
  2369=>"000000000",
  2370=>"111111111",
  2371=>"000000000",
  2372=>"000000100",
  2373=>"011011111",
  2374=>"000000010",
  2375=>"100111110",
  2376=>"000000100",
  2377=>"111110110",
  2378=>"011001111",
  2379=>"000000000",
  2380=>"001001000",
  2381=>"001000000",
  2382=>"001001011",
  2383=>"011001001",
  2384=>"101101001",
  2385=>"001001001",
  2386=>"000000100",
  2387=>"111111111",
  2388=>"101001001",
  2389=>"001011011",
  2390=>"101100100",
  2391=>"000000000",
  2392=>"000000001",
  2393=>"010000011",
  2394=>"001001100",
  2395=>"000001111",
  2396=>"011010010",
  2397=>"111010000",
  2398=>"001001000",
  2399=>"000000000",
  2400=>"000000000",
  2401=>"000000000",
  2402=>"001000100",
  2403=>"111000000",
  2404=>"111000000",
  2405=>"001000101",
  2406=>"011000111",
  2407=>"110110111",
  2408=>"000100111",
  2409=>"000000000",
  2410=>"001000001",
  2411=>"010110110",
  2412=>"001000000",
  2413=>"111011100",
  2414=>"000000000",
  2415=>"111111000",
  2416=>"111111111",
  2417=>"111111001",
  2418=>"001111000",
  2419=>"111111011",
  2420=>"111111111",
  2421=>"100000000",
  2422=>"111111111",
  2423=>"000001011",
  2424=>"111111111",
  2425=>"011111111",
  2426=>"000001111",
  2427=>"110111011",
  2428=>"111001000",
  2429=>"001001111",
  2430=>"011000000",
  2431=>"111101101",
  2432=>"000010100",
  2433=>"101011101",
  2434=>"000000000",
  2435=>"111000001",
  2436=>"100000000",
  2437=>"110000110",
  2438=>"111111111",
  2439=>"111111001",
  2440=>"101001101",
  2441=>"111111000",
  2442=>"000000000",
  2443=>"010000111",
  2444=>"110111101",
  2445=>"011110001",
  2446=>"000000000",
  2447=>"000000000",
  2448=>"001000100",
  2449=>"000000000",
  2450=>"000010111",
  2451=>"000000000",
  2452=>"101001111",
  2453=>"010010000",
  2454=>"110111111",
  2455=>"001001111",
  2456=>"111111111",
  2457=>"011101001",
  2458=>"110110000",
  2459=>"001000101",
  2460=>"011010010",
  2461=>"000000000",
  2462=>"000111111",
  2463=>"110010111",
  2464=>"001000000",
  2465=>"011001001",
  2466=>"101001000",
  2467=>"001001000",
  2468=>"000000000",
  2469=>"000000000",
  2470=>"111111111",
  2471=>"000110111",
  2472=>"110110010",
  2473=>"001001000",
  2474=>"000000111",
  2475=>"001001111",
  2476=>"000110000",
  2477=>"001001100",
  2478=>"111111111",
  2479=>"101000001",
  2480=>"001011111",
  2481=>"111111111",
  2482=>"000101110",
  2483=>"111111111",
  2484=>"001000000",
  2485=>"001011011",
  2486=>"000010000",
  2487=>"000000011",
  2488=>"001000000",
  2489=>"111010010",
  2490=>"100000000",
  2491=>"010110111",
  2492=>"100000000",
  2493=>"001001001",
  2494=>"000000000",
  2495=>"111011001",
  2496=>"001001011",
  2497=>"100111111",
  2498=>"000000000",
  2499=>"000000010",
  2500=>"100000000",
  2501=>"001000000",
  2502=>"001011111",
  2503=>"000110110",
  2504=>"011111111",
  2505=>"101110011",
  2506=>"101001000",
  2507=>"010010000",
  2508=>"001000110",
  2509=>"000000000",
  2510=>"110110100",
  2511=>"000001111",
  2512=>"001001111",
  2513=>"001001100",
  2514=>"001011111",
  2515=>"000110010",
  2516=>"000000000",
  2517=>"100000000",
  2518=>"101000111",
  2519=>"000000000",
  2520=>"001000101",
  2521=>"000000011",
  2522=>"110011111",
  2523=>"100000000",
  2524=>"011010000",
  2525=>"011110010",
  2526=>"000000111",
  2527=>"110110111",
  2528=>"110110111",
  2529=>"100000001",
  2530=>"000000001",
  2531=>"111111111",
  2532=>"111100111",
  2533=>"000000000",
  2534=>"110110011",
  2535=>"000000000",
  2536=>"110110111",
  2537=>"001101000",
  2538=>"000110011",
  2539=>"111111111",
  2540=>"011111111",
  2541=>"111001000",
  2542=>"111111111",
  2543=>"000000111",
  2544=>"001001001",
  2545=>"100110111",
  2546=>"111111000",
  2547=>"101011111",
  2548=>"000111111",
  2549=>"000000000",
  2550=>"111111001",
  2551=>"111101100",
  2552=>"110110110",
  2553=>"100001001",
  2554=>"101101000",
  2555=>"111111101",
  2556=>"110000010",
  2557=>"001000111",
  2558=>"110100111",
  2559=>"000111111",
  2560=>"111000100",
  2561=>"000001000",
  2562=>"111111111",
  2563=>"111000000",
  2564=>"100100100",
  2565=>"000010000",
  2566=>"111000100",
  2567=>"000000000",
  2568=>"111000001",
  2569=>"111111011",
  2570=>"000000000",
  2571=>"000000000",
  2572=>"110010000",
  2573=>"000110000",
  2574=>"000000011",
  2575=>"000001011",
  2576=>"111111111",
  2577=>"111111110",
  2578=>"001000000",
  2579=>"100110100",
  2580=>"111111111",
  2581=>"111111000",
  2582=>"000000000",
  2583=>"000100000",
  2584=>"100100000",
  2585=>"000111111",
  2586=>"000000000",
  2587=>"101011011",
  2588=>"000000000",
  2589=>"001000000",
  2590=>"001011111",
  2591=>"110111111",
  2592=>"000000000",
  2593=>"000010111",
  2594=>"111110000",
  2595=>"001001101",
  2596=>"101111111",
  2597=>"111111100",
  2598=>"000000000",
  2599=>"111111111",
  2600=>"000000000",
  2601=>"111001000",
  2602=>"000100111",
  2603=>"110100101",
  2604=>"101111111",
  2605=>"000000000",
  2606=>"110100000",
  2607=>"111001111",
  2608=>"000000100",
  2609=>"000000000",
  2610=>"100110110",
  2611=>"001000000",
  2612=>"110110110",
  2613=>"111111111",
  2614=>"111100110",
  2615=>"111000000",
  2616=>"100100000",
  2617=>"001000000",
  2618=>"100111111",
  2619=>"000000111",
  2620=>"000010111",
  2621=>"001000101",
  2622=>"001011011",
  2623=>"111111111",
  2624=>"111111111",
  2625=>"000110110",
  2626=>"111111111",
  2627=>"000000111",
  2628=>"000000100",
  2629=>"000001111",
  2630=>"100001000",
  2631=>"111111111",
  2632=>"101111111",
  2633=>"001000111",
  2634=>"111111111",
  2635=>"000111111",
  2636=>"111111000",
  2637=>"111111111",
  2638=>"111111100",
  2639=>"010000000",
  2640=>"011011111",
  2641=>"101111111",
  2642=>"100110110",
  2643=>"101111100",
  2644=>"111111111",
  2645=>"010110000",
  2646=>"000111111",
  2647=>"101000000",
  2648=>"000111100",
  2649=>"111111111",
  2650=>"001000000",
  2651=>"111111110",
  2652=>"000010110",
  2653=>"111111111",
  2654=>"100111000",
  2655=>"000000110",
  2656=>"111000000",
  2657=>"000011001",
  2658=>"000000000",
  2659=>"000000000",
  2660=>"110111000",
  2661=>"100110111",
  2662=>"011001111",
  2663=>"111111100",
  2664=>"111111111",
  2665=>"111110010",
  2666=>"000111111",
  2667=>"000001001",
  2668=>"001000100",
  2669=>"111111111",
  2670=>"000000111",
  2671=>"000011111",
  2672=>"111110000",
  2673=>"000000001",
  2674=>"011111010",
  2675=>"000000000",
  2676=>"111111111",
  2677=>"110111111",
  2678=>"010010000",
  2679=>"000010000",
  2680=>"000000000",
  2681=>"110111111",
  2682=>"000000100",
  2683=>"101101111",
  2684=>"100101111",
  2685=>"111111111",
  2686=>"000000000",
  2687=>"111111111",
  2688=>"100111111",
  2689=>"110111111",
  2690=>"000001111",
  2691=>"000111111",
  2692=>"110110111",
  2693=>"111111011",
  2694=>"000000000",
  2695=>"000000000",
  2696=>"001101111",
  2697=>"000001011",
  2698=>"000000000",
  2699=>"100000000",
  2700=>"000111111",
  2701=>"000000000",
  2702=>"111111011",
  2703=>"000100111",
  2704=>"111111111",
  2705=>"111010000",
  2706=>"000000000",
  2707=>"001000000",
  2708=>"000110000",
  2709=>"011001100",
  2710=>"101111111",
  2711=>"001000000",
  2712=>"000000001",
  2713=>"000000000",
  2714=>"101111111",
  2715=>"000111111",
  2716=>"001000101",
  2717=>"110110110",
  2718=>"111111111",
  2719=>"100111111",
  2720=>"100000000",
  2721=>"111001101",
  2722=>"111111111",
  2723=>"111111111",
  2724=>"000000000",
  2725=>"000000001",
  2726=>"111111010",
  2727=>"011001001",
  2728=>"110000111",
  2729=>"111111111",
  2730=>"100000001",
  2731=>"000000000",
  2732=>"000000000",
  2733=>"000000110",
  2734=>"111101101",
  2735=>"110110111",
  2736=>"111100111",
  2737=>"011000000",
  2738=>"010000010",
  2739=>"000000000",
  2740=>"000011010",
  2741=>"011001000",
  2742=>"000000000",
  2743=>"111111111",
  2744=>"000000110",
  2745=>"111111111",
  2746=>"010010000",
  2747=>"111010000",
  2748=>"101111111",
  2749=>"111111000",
  2750=>"111000000",
  2751=>"111000000",
  2752=>"111110110",
  2753=>"001101101",
  2754=>"111000000",
  2755=>"000000000",
  2756=>"000000111",
  2757=>"000000111",
  2758=>"000010000",
  2759=>"111011000",
  2760=>"100000100",
  2761=>"101101111",
  2762=>"111110011",
  2763=>"111111111",
  2764=>"001011101",
  2765=>"111100000",
  2766=>"000000000",
  2767=>"110111111",
  2768=>"111111111",
  2769=>"111111110",
  2770=>"000000100",
  2771=>"000000101",
  2772=>"000000001",
  2773=>"000000000",
  2774=>"111111111",
  2775=>"110111000",
  2776=>"000000000",
  2777=>"111100000",
  2778=>"110110100",
  2779=>"010110000",
  2780=>"000000000",
  2781=>"000000000",
  2782=>"000000010",
  2783=>"001011011",
  2784=>"011010001",
  2785=>"111001001",
  2786=>"001000000",
  2787=>"101001000",
  2788=>"111011000",
  2789=>"111111011",
  2790=>"111111001",
  2791=>"111111111",
  2792=>"000000000",
  2793=>"011111000",
  2794=>"111111100",
  2795=>"000000000",
  2796=>"000000000",
  2797=>"000000000",
  2798=>"111001111",
  2799=>"011111111",
  2800=>"111111111",
  2801=>"111100000",
  2802=>"111011001",
  2803=>"111100000",
  2804=>"000000000",
  2805=>"100000000",
  2806=>"111111100",
  2807=>"001001111",
  2808=>"111111111",
  2809=>"111111111",
  2810=>"100101111",
  2811=>"000110111",
  2812=>"001001100",
  2813=>"110110110",
  2814=>"101100111",
  2815=>"111111111",
  2816=>"000000011",
  2817=>"000011010",
  2818=>"111111111",
  2819=>"000000000",
  2820=>"111111111",
  2821=>"111110100",
  2822=>"100100000",
  2823=>"000000000",
  2824=>"000100000",
  2825=>"111111111",
  2826=>"101000000",
  2827=>"000110111",
  2828=>"000000000",
  2829=>"100111011",
  2830=>"000000001",
  2831=>"000111111",
  2832=>"111111101",
  2833=>"011111111",
  2834=>"111111000",
  2835=>"111110000",
  2836=>"001111101",
  2837=>"000000111",
  2838=>"001000100",
  2839=>"100000111",
  2840=>"000000000",
  2841=>"110000000",
  2842=>"000011111",
  2843=>"000000001",
  2844=>"111111111",
  2845=>"111000000",
  2846=>"000001011",
  2847=>"000000000",
  2848=>"000000000",
  2849=>"010010010",
  2850=>"100000000",
  2851=>"111110100",
  2852=>"111111111",
  2853=>"000001111",
  2854=>"111111101",
  2855=>"111110000",
  2856=>"111111000",
  2857=>"111111111",
  2858=>"000000000",
  2859=>"010000000",
  2860=>"111111001",
  2861=>"001000000",
  2862=>"000000000",
  2863=>"100110110",
  2864=>"101011011",
  2865=>"000000111",
  2866=>"001000000",
  2867=>"000101001",
  2868=>"000000000",
  2869=>"011011110",
  2870=>"001001001",
  2871=>"000111111",
  2872=>"000000111",
  2873=>"000000000",
  2874=>"111111111",
  2875=>"000000000",
  2876=>"001001111",
  2877=>"110111001",
  2878=>"000000000",
  2879=>"101100001",
  2880=>"000111111",
  2881=>"111100101",
  2882=>"000000000",
  2883=>"111010010",
  2884=>"000101001",
  2885=>"111111111",
  2886=>"111111111",
  2887=>"001000000",
  2888=>"111010011",
  2889=>"000000000",
  2890=>"000111111",
  2891=>"000000000",
  2892=>"001001111",
  2893=>"000000000",
  2894=>"110111111",
  2895=>"110110100",
  2896=>"101000100",
  2897=>"111111111",
  2898=>"000000000",
  2899=>"111111111",
  2900=>"000000100",
  2901=>"101111111",
  2902=>"001111111",
  2903=>"100111111",
  2904=>"000000001",
  2905=>"000000000",
  2906=>"111010111",
  2907=>"000000000",
  2908=>"111111111",
  2909=>"111111111",
  2910=>"000000101",
  2911=>"111111011",
  2912=>"111000011",
  2913=>"000000000",
  2914=>"111111000",
  2915=>"000000000",
  2916=>"110110000",
  2917=>"011111000",
  2918=>"000000000",
  2919=>"111111111",
  2920=>"000001011",
  2921=>"111111111",
  2922=>"111111000",
  2923=>"110110110",
  2924=>"111111111",
  2925=>"100000011",
  2926=>"110111111",
  2927=>"111000000",
  2928=>"001001001",
  2929=>"000000000",
  2930=>"110010000",
  2931=>"011001001",
  2932=>"000000000",
  2933=>"101000111",
  2934=>"000000101",
  2935=>"100000111",
  2936=>"001000101",
  2937=>"101111111",
  2938=>"111111111",
  2939=>"000000000",
  2940=>"110010110",
  2941=>"000000001",
  2942=>"000111101",
  2943=>"101000111",
  2944=>"000000000",
  2945=>"111001111",
  2946=>"111111111",
  2947=>"101000000",
  2948=>"111111111",
  2949=>"000000000",
  2950=>"000100000",
  2951=>"000001000",
  2952=>"000000000",
  2953=>"000000011",
  2954=>"111111111",
  2955=>"000001111",
  2956=>"101111111",
  2957=>"011011011",
  2958=>"000001111",
  2959=>"000000000",
  2960=>"101101001",
  2961=>"000000111",
  2962=>"110110100",
  2963=>"111110111",
  2964=>"000000000",
  2965=>"000000011",
  2966=>"111000110",
  2967=>"111111111",
  2968=>"110111001",
  2969=>"111111100",
  2970=>"111111111",
  2971=>"010111111",
  2972=>"101100100",
  2973=>"000000000",
  2974=>"111111111",
  2975=>"000000000",
  2976=>"111001001",
  2977=>"110110011",
  2978=>"111111011",
  2979=>"000000001",
  2980=>"111111000",
  2981=>"000000000",
  2982=>"000110000",
  2983=>"111111000",
  2984=>"000000111",
  2985=>"111111111",
  2986=>"011000000",
  2987=>"000100110",
  2988=>"000000000",
  2989=>"000100100",
  2990=>"000000010",
  2991=>"011001001",
  2992=>"000000000",
  2993=>"000000000",
  2994=>"111111111",
  2995=>"000000001",
  2996=>"111111111",
  2997=>"101111111",
  2998=>"000110110",
  2999=>"100110100",
  3000=>"110110100",
  3001=>"101111111",
  3002=>"000001001",
  3003=>"111111111",
  3004=>"111111000",
  3005=>"100000000",
  3006=>"111111111",
  3007=>"111011011",
  3008=>"100111111",
  3009=>"111111101",
  3010=>"000000000",
  3011=>"000000000",
  3012=>"010010000",
  3013=>"000000101",
  3014=>"111111111",
  3015=>"111111111",
  3016=>"001000000",
  3017=>"111111110",
  3018=>"110000111",
  3019=>"000000000",
  3020=>"110111101",
  3021=>"111111111",
  3022=>"110010110",
  3023=>"111000000",
  3024=>"111111111",
  3025=>"111011001",
  3026=>"111101000",
  3027=>"111000000",
  3028=>"000000101",
  3029=>"000100110",
  3030=>"110111001",
  3031=>"000000000",
  3032=>"100000000",
  3033=>"111001111",
  3034=>"111000000",
  3035=>"001001000",
  3036=>"111111111",
  3037=>"000000111",
  3038=>"000000000",
  3039=>"110111000",
  3040=>"111111111",
  3041=>"111111101",
  3042=>"000000000",
  3043=>"111111111",
  3044=>"001001000",
  3045=>"010011011",
  3046=>"010110110",
  3047=>"111111111",
  3048=>"111111111",
  3049=>"111011111",
  3050=>"000000000",
  3051=>"111111111",
  3052=>"111111111",
  3053=>"011011111",
  3054=>"010100100",
  3055=>"010010000",
  3056=>"111111100",
  3057=>"111111111",
  3058=>"111111000",
  3059=>"111111110",
  3060=>"000000110",
  3061=>"111001000",
  3062=>"011000000",
  3063=>"001001000",
  3064=>"000000111",
  3065=>"111100100",
  3066=>"111000000",
  3067=>"111000000",
  3068=>"111111001",
  3069=>"110000000",
  3070=>"111111111",
  3071=>"000000000",
  3072=>"111000000",
  3073=>"110000000",
  3074=>"111010000",
  3075=>"000000000",
  3076=>"000000000",
  3077=>"111011001",
  3078=>"000000000",
  3079=>"111111101",
  3080=>"000000001",
  3081=>"111111111",
  3082=>"000000000",
  3083=>"000000001",
  3084=>"101111111",
  3085=>"111110110",
  3086=>"000000000",
  3087=>"000000000",
  3088=>"000000000",
  3089=>"000111111",
  3090=>"000000000",
  3091=>"000000000",
  3092=>"000000000",
  3093=>"001000001",
  3094=>"000001011",
  3095=>"000000111",
  3096=>"111111111",
  3097=>"111110000",
  3098=>"111111111",
  3099=>"111111000",
  3100=>"101101111",
  3101=>"000000000",
  3102=>"000000011",
  3103=>"000000000",
  3104=>"111101111",
  3105=>"111001101",
  3106=>"111111111",
  3107=>"000000000",
  3108=>"001001100",
  3109=>"100000000",
  3110=>"111111111",
  3111=>"011000000",
  3112=>"000000000",
  3113=>"110100000",
  3114=>"000000000",
  3115=>"000000100",
  3116=>"001000000",
  3117=>"001000000",
  3118=>"000000000",
  3119=>"011011011",
  3120=>"000000000",
  3121=>"111001001",
  3122=>"000000000",
  3123=>"111111000",
  3124=>"001111111",
  3125=>"101111111",
  3126=>"000000000",
  3127=>"111111111",
  3128=>"000000000",
  3129=>"111111111",
  3130=>"111000000",
  3131=>"110110000",
  3132=>"111101111",
  3133=>"000000000",
  3134=>"011001001",
  3135=>"000000000",
  3136=>"011011000",
  3137=>"111111111",
  3138=>"111001000",
  3139=>"111111111",
  3140=>"110000000",
  3141=>"111111111",
  3142=>"111111111",
  3143=>"000111111",
  3144=>"011111111",
  3145=>"000000110",
  3146=>"111111111",
  3147=>"000000000",
  3148=>"111111111",
  3149=>"010111101",
  3150=>"111111000",
  3151=>"000000000",
  3152=>"111111110",
  3153=>"111011111",
  3154=>"000000000",
  3155=>"000000100",
  3156=>"110000000",
  3157=>"111111111",
  3158=>"111001100",
  3159=>"111101001",
  3160=>"110111011",
  3161=>"111111111",
  3162=>"000000000",
  3163=>"000000011",
  3164=>"000000001",
  3165=>"100000001",
  3166=>"011001111",
  3167=>"000000000",
  3168=>"000000000",
  3169=>"110111111",
  3170=>"000000000",
  3171=>"111111010",
  3172=>"000000000",
  3173=>"001011001",
  3174=>"001000000",
  3175=>"110111011",
  3176=>"111111111",
  3177=>"111100111",
  3178=>"110101000",
  3179=>"000000000",
  3180=>"000010100",
  3181=>"111111001",
  3182=>"000000000",
  3183=>"100111000",
  3184=>"011111111",
  3185=>"000000001",
  3186=>"000111111",
  3187=>"111111111",
  3188=>"111000000",
  3189=>"000100000",
  3190=>"111111111",
  3191=>"000000000",
  3192=>"101011000",
  3193=>"011110100",
  3194=>"000011111",
  3195=>"000000000",
  3196=>"100100100",
  3197=>"000010000",
  3198=>"001001000",
  3199=>"000000100",
  3200=>"010000000",
  3201=>"000000011",
  3202=>"001111111",
  3203=>"111101111",
  3204=>"111000000",
  3205=>"111000000",
  3206=>"110000000",
  3207=>"011000000",
  3208=>"000000000",
  3209=>"111111111",
  3210=>"111111111",
  3211=>"111111011",
  3212=>"111111100",
  3213=>"110100001",
  3214=>"000000000",
  3215=>"000110110",
  3216=>"111100100",
  3217=>"000011111",
  3218=>"000000101",
  3219=>"100000010",
  3220=>"110000000",
  3221=>"000111111",
  3222=>"101100000",
  3223=>"000000000",
  3224=>"011111111",
  3225=>"100000000",
  3226=>"110111100",
  3227=>"001000000",
  3228=>"111111111",
  3229=>"000010001",
  3230=>"101001000",
  3231=>"110000111",
  3232=>"000000000",
  3233=>"111011111",
  3234=>"000000000",
  3235=>"010111110",
  3236=>"000100100",
  3237=>"111100111",
  3238=>"100000000",
  3239=>"001011011",
  3240=>"111111101",
  3241=>"111111111",
  3242=>"000100111",
  3243=>"111111111",
  3244=>"100000111",
  3245=>"111011010",
  3246=>"000001100",
  3247=>"110000011",
  3248=>"111110111",
  3249=>"000000111",
  3250=>"100000000",
  3251=>"000000000",
  3252=>"000000100",
  3253=>"111111111",
  3254=>"000110111",
  3255=>"000110111",
  3256=>"111111111",
  3257=>"111111110",
  3258=>"000010010",
  3259=>"000001101",
  3260=>"111111111",
  3261=>"111111001",
  3262=>"001000000",
  3263=>"000000000",
  3264=>"000000000",
  3265=>"111001000",
  3266=>"111111111",
  3267=>"111000000",
  3268=>"101100000",
  3269=>"111111111",
  3270=>"100111111",
  3271=>"101111111",
  3272=>"011111110",
  3273=>"111111111",
  3274=>"110110000",
  3275=>"111111111",
  3276=>"111111111",
  3277=>"111111000",
  3278=>"101100110",
  3279=>"000000000",
  3280=>"000010010",
  3281=>"111111111",
  3282=>"110100000",
  3283=>"111111111",
  3284=>"000111010",
  3285=>"001010011",
  3286=>"111111010",
  3287=>"010000000",
  3288=>"000000000",
  3289=>"000000000",
  3290=>"000000000",
  3291=>"001001111",
  3292=>"111111111",
  3293=>"000000111",
  3294=>"001000000",
  3295=>"100000100",
  3296=>"000000000",
  3297=>"011011111",
  3298=>"000000000",
  3299=>"111111101",
  3300=>"010000000",
  3301=>"001001001",
  3302=>"111111111",
  3303=>"000000000",
  3304=>"111110100",
  3305=>"000000000",
  3306=>"000000000",
  3307=>"111111111",
  3308=>"111000000",
  3309=>"010110011",
  3310=>"101111100",
  3311=>"000000000",
  3312=>"111101110",
  3313=>"000000010",
  3314=>"111111111",
  3315=>"110111011",
  3316=>"001111111",
  3317=>"001000000",
  3318=>"001001111",
  3319=>"111111111",
  3320=>"101111001",
  3321=>"000000000",
  3322=>"000000000",
  3323=>"000000100",
  3324=>"110011011",
  3325=>"100000100",
  3326=>"111111110",
  3327=>"100100101",
  3328=>"111111000",
  3329=>"001111111",
  3330=>"111111111",
  3331=>"100100111",
  3332=>"011111111",
  3333=>"000000000",
  3334=>"111111111",
  3335=>"100100111",
  3336=>"111111110",
  3337=>"111111111",
  3338=>"000000000",
  3339=>"011111110",
  3340=>"111111111",
  3341=>"111111111",
  3342=>"111011011",
  3343=>"101001000",
  3344=>"000000001",
  3345=>"000000011",
  3346=>"000000100",
  3347=>"111111011",
  3348=>"000011000",
  3349=>"111111111",
  3350=>"001101111",
  3351=>"111111111",
  3352=>"000000100",
  3353=>"000100000",
  3354=>"111110000",
  3355=>"111111011",
  3356=>"000000010",
  3357=>"111000000",
  3358=>"111111101",
  3359=>"000000000",
  3360=>"100001001",
  3361=>"011011000",
  3362=>"111111111",
  3363=>"101001111",
  3364=>"000000000",
  3365=>"111111111",
  3366=>"000000111",
  3367=>"111111011",
  3368=>"110111001",
  3369=>"111111111",
  3370=>"111000100",
  3371=>"100000000",
  3372=>"000000000",
  3373=>"100100000",
  3374=>"111000000",
  3375=>"000000000",
  3376=>"111111100",
  3377=>"000000101",
  3378=>"111111011",
  3379=>"000000000",
  3380=>"111111011",
  3381=>"111011000",
  3382=>"000000000",
  3383=>"110000010",
  3384=>"000000001",
  3385=>"001001000",
  3386=>"000000000",
  3387=>"111111000",
  3388=>"000001000",
  3389=>"000110111",
  3390=>"111101000",
  3391=>"000100100",
  3392=>"111011111",
  3393=>"100100110",
  3394=>"111111110",
  3395=>"000000000",
  3396=>"001000000",
  3397=>"100111111",
  3398=>"000000000",
  3399=>"000000100",
  3400=>"000000000",
  3401=>"110000000",
  3402=>"001001001",
  3403=>"000000000",
  3404=>"111111011",
  3405=>"111110000",
  3406=>"110110101",
  3407=>"100100000",
  3408=>"000001101",
  3409=>"111001000",
  3410=>"111111111",
  3411=>"000000000",
  3412=>"000000000",
  3413=>"011001011",
  3414=>"111111100",
  3415=>"111111111",
  3416=>"100000000",
  3417=>"111111111",
  3418=>"110000111",
  3419=>"001000000",
  3420=>"111111011",
  3421=>"111111111",
  3422=>"111111111",
  3423=>"001011001",
  3424=>"111000110",
  3425=>"000000000",
  3426=>"010010110",
  3427=>"110111111",
  3428=>"000000000",
  3429=>"000000000",
  3430=>"000000000",
  3431=>"000000000",
  3432=>"100000101",
  3433=>"000011111",
  3434=>"000000000",
  3435=>"000000011",
  3436=>"111110000",
  3437=>"000110110",
  3438=>"111111111",
  3439=>"110110110",
  3440=>"110010000",
  3441=>"000000001",
  3442=>"111111100",
  3443=>"111111111",
  3444=>"000001000",
  3445=>"011111111",
  3446=>"000000000",
  3447=>"000000000",
  3448=>"111111111",
  3449=>"100000000",
  3450=>"000000100",
  3451=>"000000110",
  3452=>"111111111",
  3453=>"111000110",
  3454=>"001000000",
  3455=>"111111111",
  3456=>"101111100",
  3457=>"110000110",
  3458=>"111111111",
  3459=>"000000000",
  3460=>"010111111",
  3461=>"001000000",
  3462=>"000000111",
  3463=>"111111111",
  3464=>"111111111",
  3465=>"000000110",
  3466=>"111111001",
  3467=>"111111011",
  3468=>"111111111",
  3469=>"000110011",
  3470=>"001001000",
  3471=>"000000000",
  3472=>"000000000",
  3473=>"111010000",
  3474=>"000000000",
  3475=>"000010000",
  3476=>"111101100",
  3477=>"000000000",
  3478=>"111110000",
  3479=>"101000100",
  3480=>"001111111",
  3481=>"000000000",
  3482=>"111111110",
  3483=>"000000000",
  3484=>"000000000",
  3485=>"000000000",
  3486=>"001001000",
  3487=>"111111111",
  3488=>"000000000",
  3489=>"111101101",
  3490=>"000000100",
  3491=>"111111011",
  3492=>"101111111",
  3493=>"000010000",
  3494=>"111001010",
  3495=>"100000000",
  3496=>"101000000",
  3497=>"111010000",
  3498=>"010111111",
  3499=>"000001000",
  3500=>"000000000",
  3501=>"110110110",
  3502=>"000001111",
  3503=>"111111111",
  3504=>"010110111",
  3505=>"000000000",
  3506=>"111111110",
  3507=>"000000000",
  3508=>"111111111",
  3509=>"001000000",
  3510=>"001001100",
  3511=>"111000000",
  3512=>"111111111",
  3513=>"000000000",
  3514=>"000000000",
  3515=>"100111111",
  3516=>"111111111",
  3517=>"111110111",
  3518=>"001000000",
  3519=>"000000000",
  3520=>"111111111",
  3521=>"111000000",
  3522=>"000000000",
  3523=>"101101000",
  3524=>"111111111",
  3525=>"100110100",
  3526=>"111111001",
  3527=>"000000000",
  3528=>"111111110",
  3529=>"100000000",
  3530=>"110110110",
  3531=>"000000001",
  3532=>"010111011",
  3533=>"000000000",
  3534=>"110111010",
  3535=>"000000000",
  3536=>"000000000",
  3537=>"110111111",
  3538=>"111111000",
  3539=>"011111011",
  3540=>"100000000",
  3541=>"000001000",
  3542=>"000000001",
  3543=>"001001001",
  3544=>"101000111",
  3545=>"101001111",
  3546=>"111111000",
  3547=>"000001101",
  3548=>"000000000",
  3549=>"111001001",
  3550=>"011000000",
  3551=>"000000100",
  3552=>"111111111",
  3553=>"000000000",
  3554=>"000000011",
  3555=>"000001001",
  3556=>"000000010",
  3557=>"100000001",
  3558=>"111111111",
  3559=>"111111110",
  3560=>"000000001",
  3561=>"001111010",
  3562=>"000010110",
  3563=>"000000000",
  3564=>"000000000",
  3565=>"000000000",
  3566=>"000000000",
  3567=>"110111111",
  3568=>"000011001",
  3569=>"000000100",
  3570=>"111111111",
  3571=>"000000000",
  3572=>"111000000",
  3573=>"111011000",
  3574=>"111101111",
  3575=>"100000000",
  3576=>"000110110",
  3577=>"000010010",
  3578=>"000001001",
  3579=>"000000000",
  3580=>"100000000",
  3581=>"110111111",
  3582=>"111111111",
  3583=>"111001011",
  3584=>"001101111",
  3585=>"001000001",
  3586=>"101101101",
  3587=>"101101111",
  3588=>"111111111",
  3589=>"101001001",
  3590=>"000000000",
  3591=>"111111111",
  3592=>"001011101",
  3593=>"111000000",
  3594=>"111001101",
  3595=>"101101101",
  3596=>"010010010",
  3597=>"111100100",
  3598=>"000011010",
  3599=>"110101101",
  3600=>"101101101",
  3601=>"111111000",
  3602=>"000000000",
  3603=>"101001000",
  3604=>"001101101",
  3605=>"101000000",
  3606=>"000000001",
  3607=>"111001000",
  3608=>"111111111",
  3609=>"110010010",
  3610=>"111000000",
  3611=>"101101000",
  3612=>"001001111",
  3613=>"000000000",
  3614=>"111111010",
  3615=>"000000101",
  3616=>"011001000",
  3617=>"111111110",
  3618=>"100110111",
  3619=>"000101101",
  3620=>"001011111",
  3621=>"111101000",
  3622=>"000101000",
  3623=>"000011001",
  3624=>"001000100",
  3625=>"101001001",
  3626=>"101001101",
  3627=>"000000100",
  3628=>"100110011",
  3629=>"000000100",
  3630=>"101100111",
  3631=>"101101101",
  3632=>"111111100",
  3633=>"110010010",
  3634=>"111111111",
  3635=>"010100100",
  3636=>"010010110",
  3637=>"110110111",
  3638=>"110100100",
  3639=>"001001101",
  3640=>"001001101",
  3641=>"000000110",
  3642=>"000000000",
  3643=>"110000000",
  3644=>"111000001",
  3645=>"000000100",
  3646=>"111111100",
  3647=>"000000111",
  3648=>"001111111",
  3649=>"100001101",
  3650=>"010010010",
  3651=>"111011001",
  3652=>"000111111",
  3653=>"000000000",
  3654=>"000001000",
  3655=>"001000000",
  3656=>"110110000",
  3657=>"001001001",
  3658=>"110110010",
  3659=>"101001100",
  3660=>"110110111",
  3661=>"111111010",
  3662=>"111011110",
  3663=>"000110110",
  3664=>"001001111",
  3665=>"110011111",
  3666=>"100100100",
  3667=>"000110000",
  3668=>"000000000",
  3669=>"000110010",
  3670=>"100100000",
  3671=>"011001011",
  3672=>"000001111",
  3673=>"101100100",
  3674=>"101101101",
  3675=>"000000000",
  3676=>"000000000",
  3677=>"100000000",
  3678=>"000001001",
  3679=>"001001101",
  3680=>"110110110",
  3681=>"111111111",
  3682=>"101101101",
  3683=>"110010111",
  3684=>"010011111",
  3685=>"001000100",
  3686=>"001111101",
  3687=>"001101111",
  3688=>"001011111",
  3689=>"000000001",
  3690=>"010010011",
  3691=>"101101101",
  3692=>"000000001",
  3693=>"000001000",
  3694=>"101101101",
  3695=>"010111111",
  3696=>"011010010",
  3697=>"011001001",
  3698=>"010010011",
  3699=>"101101001",
  3700=>"101111111",
  3701=>"000110110",
  3702=>"101101101",
  3703=>"010010010",
  3704=>"001001011",
  3705=>"011010010",
  3706=>"010010000",
  3707=>"101101101",
  3708=>"000000100",
  3709=>"111111011",
  3710=>"010010010",
  3711=>"011011000",
  3712=>"011111111",
  3713=>"100001001",
  3714=>"001001000",
  3715=>"111011011",
  3716=>"001000100",
  3717=>"101001100",
  3718=>"011001000",
  3719=>"100100100",
  3720=>"111000010",
  3721=>"111011111",
  3722=>"000010010",
  3723=>"101001000",
  3724=>"101101101",
  3725=>"010010010",
  3726=>"111111001",
  3727=>"101111011",
  3728=>"000000010",
  3729=>"000000010",
  3730=>"101001011",
  3731=>"000000010",
  3732=>"000000000",
  3733=>"010000000",
  3734=>"101000000",
  3735=>"101001001",
  3736=>"001101111",
  3737=>"001001001",
  3738=>"101100000",
  3739=>"100101101",
  3740=>"001001001",
  3741=>"101111111",
  3742=>"101111001",
  3743=>"100100000",
  3744=>"111000000",
  3745=>"100100111",
  3746=>"001101111",
  3747=>"100111111",
  3748=>"100100100",
  3749=>"001111001",
  3750=>"000010010",
  3751=>"011010011",
  3752=>"000000101",
  3753=>"011000010",
  3754=>"000000000",
  3755=>"010010110",
  3756=>"101101000",
  3757=>"001111110",
  3758=>"111111101",
  3759=>"001111110",
  3760=>"000000111",
  3761=>"010111010",
  3762=>"110110110",
  3763=>"010010010",
  3764=>"111010000",
  3765=>"111111101",
  3766=>"010000011",
  3767=>"011111010",
  3768=>"011101111",
  3769=>"010010011",
  3770=>"000000000",
  3771=>"101111000",
  3772=>"011001001",
  3773=>"000010111",
  3774=>"111001101",
  3775=>"001011011",
  3776=>"111011111",
  3777=>"100111101",
  3778=>"001001001",
  3779=>"000000000",
  3780=>"001110110",
  3781=>"101101101",
  3782=>"101001101",
  3783=>"001001000",
  3784=>"110110100",
  3785=>"000101101",
  3786=>"001101101",
  3787=>"010010000",
  3788=>"101101000",
  3789=>"000000100",
  3790=>"110111110",
  3791=>"000010010",
  3792=>"101000000",
  3793=>"011111111",
  3794=>"000001111",
  3795=>"000000000",
  3796=>"000000011",
  3797=>"100100000",
  3798=>"101101101",
  3799=>"101101001",
  3800=>"001101110",
  3801=>"111111111",
  3802=>"101101101",
  3803=>"010011001",
  3804=>"000010010",
  3805=>"111111010",
  3806=>"110110111",
  3807=>"101011000",
  3808=>"001001000",
  3809=>"000011001",
  3810=>"101101101",
  3811=>"101101001",
  3812=>"001101101",
  3813=>"010010110",
  3814=>"000110111",
  3815=>"111111101",
  3816=>"000000000",
  3817=>"100101111",
  3818=>"101101101",
  3819=>"000000100",
  3820=>"010010010",
  3821=>"001101101",
  3822=>"111011011",
  3823=>"110000000",
  3824=>"111110110",
  3825=>"100111100",
  3826=>"111101101",
  3827=>"000000000",
  3828=>"000100010",
  3829=>"100100001",
  3830=>"111110110",
  3831=>"000000000",
  3832=>"110111111",
  3833=>"000010000",
  3834=>"000101000",
  3835=>"111111101",
  3836=>"010011011",
  3837=>"001101101",
  3838=>"011000000",
  3839=>"001111111",
  3840=>"000000000",
  3841=>"111011001",
  3842=>"000000100",
  3843=>"111111100",
  3844=>"101101101",
  3845=>"000000111",
  3846=>"001101101",
  3847=>"100101000",
  3848=>"111111111",
  3849=>"000111111",
  3850=>"101101101",
  3851=>"001101000",
  3852=>"110110110",
  3853=>"000100111",
  3854=>"111111111",
  3855=>"100100100",
  3856=>"011111101",
  3857=>"111111101",
  3858=>"111000101",
  3859=>"110000101",
  3860=>"010000000",
  3861=>"000001001",
  3862=>"010010011",
  3863=>"010000000",
  3864=>"000000110",
  3865=>"001000000",
  3866=>"001000000",
  3867=>"110110110",
  3868=>"010000000",
  3869=>"000000111",
  3870=>"101111111",
  3871=>"000000000",
  3872=>"101101011",
  3873=>"111111111",
  3874=>"001001011",
  3875=>"111101000",
  3876=>"001101100",
  3877=>"100010000",
  3878=>"000010000",
  3879=>"001001110",
  3880=>"111001000",
  3881=>"010100010",
  3882=>"101101110",
  3883=>"111000000",
  3884=>"001001001",
  3885=>"110000100",
  3886=>"000000000",
  3887=>"000000010",
  3888=>"001000000",
  3889=>"000010000",
  3890=>"000000111",
  3891=>"111101000",
  3892=>"111001001",
  3893=>"111111101",
  3894=>"101001001",
  3895=>"001101111",
  3896=>"000010110",
  3897=>"001101101",
  3898=>"010010001",
  3899=>"101101111",
  3900=>"000000111",
  3901=>"100110000",
  3902=>"000100000",
  3903=>"100000001",
  3904=>"111101000",
  3905=>"110111110",
  3906=>"111001101",
  3907=>"111101101",
  3908=>"000000000",
  3909=>"000001011",
  3910=>"000000101",
  3911=>"111101101",
  3912=>"000000100",
  3913=>"000000001",
  3914=>"001100100",
  3915=>"110110010",
  3916=>"000000100",
  3917=>"010011011",
  3918=>"010110111",
  3919=>"000110110",
  3920=>"100110100",
  3921=>"101101101",
  3922=>"110110111",
  3923=>"010010010",
  3924=>"000000000",
  3925=>"001001001",
  3926=>"101101111",
  3927=>"110000000",
  3928=>"101111101",
  3929=>"000000000",
  3930=>"111110110",
  3931=>"000000111",
  3932=>"101000100",
  3933=>"000100110",
  3934=>"001001100",
  3935=>"100111111",
  3936=>"101101101",
  3937=>"001000100",
  3938=>"110110110",
  3939=>"000000000",
  3940=>"110110110",
  3941=>"001001000",
  3942=>"000000000",
  3943=>"100110111",
  3944=>"011111111",
  3945=>"111110111",
  3946=>"010110111",
  3947=>"110100111",
  3948=>"010001111",
  3949=>"001011001",
  3950=>"000010010",
  3951=>"000000001",
  3952=>"001100101",
  3953=>"111111111",
  3954=>"111111000",
  3955=>"111110110",
  3956=>"110111010",
  3957=>"100111111",
  3958=>"001100100",
  3959=>"000000000",
  3960=>"000000101",
  3961=>"000011111",
  3962=>"000000000",
  3963=>"000010000",
  3964=>"000101100",
  3965=>"100111111",
  3966=>"001001000",
  3967=>"000010010",
  3968=>"111111100",
  3969=>"001001111",
  3970=>"000000000",
  3971=>"101101101",
  3972=>"000000100",
  3973=>"001000000",
  3974=>"101000100",
  3975=>"010000000",
  3976=>"000000000",
  3977=>"010010011",
  3978=>"001000101",
  3979=>"001001101",
  3980=>"000000000",
  3981=>"111111010",
  3982=>"000000000",
  3983=>"110110110",
  3984=>"110010110",
  3985=>"110100100",
  3986=>"000000110",
  3987=>"100000011",
  3988=>"000100100",
  3989=>"010010000",
  3990=>"111101101",
  3991=>"110111000",
  3992=>"111111001",
  3993=>"101101100",
  3994=>"101111111",
  3995=>"010001001",
  3996=>"000000000",
  3997=>"010011010",
  3998=>"010011010",
  3999=>"000000000",
  4000=>"101101000",
  4001=>"101001001",
  4002=>"000111111",
  4003=>"001101100",
  4004=>"001101101",
  4005=>"010010000",
  4006=>"000000111",
  4007=>"000000110",
  4008=>"111111111",
  4009=>"100101001",
  4010=>"101101001",
  4011=>"010110110",
  4012=>"001000001",
  4013=>"001100101",
  4014=>"101111010",
  4015=>"011011011",
  4016=>"000001000",
  4017=>"010010110",
  4018=>"001101101",
  4019=>"000001001",
  4020=>"000000110",
  4021=>"111111110",
  4022=>"000001001",
  4023=>"111001000",
  4024=>"111111100",
  4025=>"111011111",
  4026=>"101001001",
  4027=>"101101101",
  4028=>"110000000",
  4029=>"001101100",
  4030=>"101000000",
  4031=>"011010011",
  4032=>"111111111",
  4033=>"010010010",
  4034=>"010010010",
  4035=>"110010000",
  4036=>"111111111",
  4037=>"101101111",
  4038=>"101100000",
  4039=>"101101101",
  4040=>"000000111",
  4041=>"010010100",
  4042=>"000000000",
  4043=>"000000110",
  4044=>"010000000",
  4045=>"000110000",
  4046=>"001001001",
  4047=>"111101101",
  4048=>"011110110",
  4049=>"000100000",
  4050=>"000000111",
  4051=>"010010110",
  4052=>"010111111",
  4053=>"101001001",
  4054=>"111011000",
  4055=>"001111001",
  4056=>"000101001",
  4057=>"010111111",
  4058=>"101111101",
  4059=>"000001001",
  4060=>"001101111",
  4061=>"110010110",
  4062=>"111111111",
  4063=>"001011011",
  4064=>"000010110",
  4065=>"000010010",
  4066=>"110100001",
  4067=>"100111110",
  4068=>"111100100",
  4069=>"101101101",
  4070=>"011000011",
  4071=>"101101000",
  4072=>"111010000",
  4073=>"000000000",
  4074=>"011001101",
  4075=>"100110010",
  4076=>"001101101",
  4077=>"100000000",
  4078=>"110000010",
  4079=>"101100000",
  4080=>"010111010",
  4081=>"110011000",
  4082=>"111000000",
  4083=>"000000010",
  4084=>"000100111",
  4085=>"100101000",
  4086=>"100100010",
  4087=>"111011000",
  4088=>"111111001",
  4089=>"000000100",
  4090=>"000001101",
  4091=>"000000000",
  4092=>"000100110",
  4093=>"111111001",
  4094=>"110000000",
  4095=>"000000000",
  4096=>"001001001",
  4097=>"000000100",
  4098=>"100111111",
  4099=>"000000000",
  4100=>"000011011",
  4101=>"100100111",
  4102=>"000110111",
  4103=>"111111111",
  4104=>"100011111",
  4105=>"000000000",
  4106=>"110100111",
  4107=>"000000010",
  4108=>"000100100",
  4109=>"100100111",
  4110=>"011000000",
  4111=>"001011000",
  4112=>"111000000",
  4113=>"111111111",
  4114=>"011000000",
  4115=>"111010000",
  4116=>"011000000",
  4117=>"000001000",
  4118=>"110110111",
  4119=>"001001000",
  4120=>"100000100",
  4121=>"100000000",
  4122=>"000010111",
  4123=>"111111010",
  4124=>"000000100",
  4125=>"111111111",
  4126=>"000000000",
  4127=>"000000111",
  4128=>"000000000",
  4129=>"010010111",
  4130=>"111111111",
  4131=>"000000000",
  4132=>"000000000",
  4133=>"111101111",
  4134=>"011011100",
  4135=>"000000100",
  4136=>"111000101",
  4137=>"001000111",
  4138=>"111110110",
  4139=>"111100100",
  4140=>"111111111",
  4141=>"001000000",
  4142=>"100001001",
  4143=>"000000111",
  4144=>"000010111",
  4145=>"000000001",
  4146=>"110010010",
  4147=>"000000111",
  4148=>"000011111",
  4149=>"000001001",
  4150=>"000000101",
  4151=>"111111111",
  4152=>"011001011",
  4153=>"101000011",
  4154=>"101000111",
  4155=>"111000000",
  4156=>"001001111",
  4157=>"000000100",
  4158=>"000000000",
  4159=>"111111111",
  4160=>"111110111",
  4161=>"000000000",
  4162=>"111111111",
  4163=>"110000001",
  4164=>"000000000",
  4165=>"000000110",
  4166=>"000000000",
  4167=>"000000000",
  4168=>"111111111",
  4169=>"000001001",
  4170=>"000000000",
  4171=>"111010111",
  4172=>"000000001",
  4173=>"111100000",
  4174=>"111100100",
  4175=>"000000000",
  4176=>"111000111",
  4177=>"111111000",
  4178=>"010110100",
  4179=>"000000000",
  4180=>"111111111",
  4181=>"000000100",
  4182=>"001001111",
  4183=>"000000000",
  4184=>"000000000",
  4185=>"101001001",
  4186=>"011000110",
  4187=>"100010011",
  4188=>"111111111",
  4189=>"000000101",
  4190=>"001000100",
  4191=>"000000100",
  4192=>"011011000",
  4193=>"111111000",
  4194=>"000000000",
  4195=>"000000000",
  4196=>"111011111",
  4197=>"111100001",
  4198=>"000000000",
  4199=>"000111011",
  4200=>"110000011",
  4201=>"111111100",
  4202=>"000000000",
  4203=>"011010011",
  4204=>"000000000",
  4205=>"111111111",
  4206=>"000000000",
  4207=>"000000000",
  4208=>"000000000",
  4209=>"111001000",
  4210=>"000000001",
  4211=>"000000000",
  4212=>"000011011",
  4213=>"000000110",
  4214=>"100100000",
  4215=>"000000000",
  4216=>"111010001",
  4217=>"111111011",
  4218=>"101000000",
  4219=>"110000100",
  4220=>"100110111",
  4221=>"000000000",
  4222=>"000000000",
  4223=>"000000000",
  4224=>"000000000",
  4225=>"000000000",
  4226=>"111110110",
  4227=>"111111111",
  4228=>"001000000",
  4229=>"001000001",
  4230=>"100000000",
  4231=>"110110110",
  4232=>"111111100",
  4233=>"111111000",
  4234=>"000100101",
  4235=>"111111111",
  4236=>"000000101",
  4237=>"111111111",
  4238=>"111001011",
  4239=>"000111111",
  4240=>"000000001",
  4241=>"000000001",
  4242=>"101000000",
  4243=>"111100111",
  4244=>"000000111",
  4245=>"000010111",
  4246=>"111111111",
  4247=>"000000000",
  4248=>"000000000",
  4249=>"000000000",
  4250=>"000000000",
  4251=>"000100110",
  4252=>"000000111",
  4253=>"111110100",
  4254=>"011110111",
  4255=>"000000000",
  4256=>"100110111",
  4257=>"100111100",
  4258=>"111111011",
  4259=>"111111111",
  4260=>"000000000",
  4261=>"000001111",
  4262=>"111111111",
  4263=>"001000000",
  4264=>"111100000",
  4265=>"011011001",
  4266=>"000110111",
  4267=>"000000001",
  4268=>"001011111",
  4269=>"100100110",
  4270=>"111111111",
  4271=>"111111111",
  4272=>"000011000",
  4273=>"111111111",
  4274=>"111111011",
  4275=>"111111111",
  4276=>"111011000",
  4277=>"111110000",
  4278=>"000110111",
  4279=>"011111111",
  4280=>"011011111",
  4281=>"011111111",
  4282=>"000000000",
  4283=>"111111001",
  4284=>"111000000",
  4285=>"111111111",
  4286=>"111111111",
  4287=>"000000000",
  4288=>"000000000",
  4289=>"001000000",
  4290=>"000000000",
  4291=>"111111111",
  4292=>"001111111",
  4293=>"000000000",
  4294=>"001000001",
  4295=>"011110111",
  4296=>"110000010",
  4297=>"000001001",
  4298=>"111111101",
  4299=>"000000111",
  4300=>"110010000",
  4301=>"111111111",
  4302=>"111111111",
  4303=>"000000101",
  4304=>"000000000",
  4305=>"000000000",
  4306=>"110000000",
  4307=>"000000000",
  4308=>"000000001",
  4309=>"110000000",
  4310=>"001001001",
  4311=>"000000011",
  4312=>"110000011",
  4313=>"110111111",
  4314=>"111111111",
  4315=>"001010010",
  4316=>"111110110",
  4317=>"110110111",
  4318=>"001000000",
  4319=>"000100000",
  4320=>"011001100",
  4321=>"000100111",
  4322=>"111111111",
  4323=>"111111111",
  4324=>"100000000",
  4325=>"001000000",
  4326=>"001000000",
  4327=>"111111111",
  4328=>"110110111",
  4329=>"100100000",
  4330=>"001000000",
  4331=>"011111111",
  4332=>"111111000",
  4333=>"000000010",
  4334=>"000111111",
  4335=>"000000000",
  4336=>"111111111",
  4337=>"000000000",
  4338=>"000000001",
  4339=>"001000000",
  4340=>"001111101",
  4341=>"111000000",
  4342=>"111111000",
  4343=>"000000000",
  4344=>"000000000",
  4345=>"000000000",
  4346=>"000000000",
  4347=>"001011111",
  4348=>"000001101",
  4349=>"101110111",
  4350=>"001111111",
  4351=>"110100100",
  4352=>"111111111",
  4353=>"100100101",
  4354=>"010100001",
  4355=>"111110101",
  4356=>"111111111",
  4357=>"011001000",
  4358=>"100000110",
  4359=>"111111111",
  4360=>"111001111",
  4361=>"111111011",
  4362=>"000000000",
  4363=>"001000000",
  4364=>"000000011",
  4365=>"000000000",
  4366=>"111111111",
  4367=>"111111110",
  4368=>"000100110",
  4369=>"111111111",
  4370=>"111111111",
  4371=>"000000000",
  4372=>"000000000",
  4373=>"000000000",
  4374=>"110111101",
  4375=>"000110111",
  4376=>"111111101",
  4377=>"000000000",
  4378=>"000000001",
  4379=>"111011100",
  4380=>"011111111",
  4381=>"111111111",
  4382=>"000000000",
  4383=>"111111111",
  4384=>"111100000",
  4385=>"000000001",
  4386=>"111000000",
  4387=>"111111111",
  4388=>"000100100",
  4389=>"011110111",
  4390=>"011000000",
  4391=>"000001111",
  4392=>"000100000",
  4393=>"000001000",
  4394=>"111111111",
  4395=>"111101110",
  4396=>"000000100",
  4397=>"111111001",
  4398=>"000000101",
  4399=>"000000000",
  4400=>"111111110",
  4401=>"111100111",
  4402=>"110000100",
  4403=>"000000111",
  4404=>"111101001",
  4405=>"011100000",
  4406=>"111111111",
  4407=>"000000000",
  4408=>"110111111",
  4409=>"111000111",
  4410=>"000111110",
  4411=>"001000110",
  4412=>"000000111",
  4413=>"110111111",
  4414=>"110100001",
  4415=>"000000011",
  4416=>"000000000",
  4417=>"100100111",
  4418=>"111110111",
  4419=>"111111111",
  4420=>"000000000",
  4421=>"111000000",
  4422=>"000000000",
  4423=>"110110110",
  4424=>"011111111",
  4425=>"110000000",
  4426=>"111111111",
  4427=>"110110110",
  4428=>"001000110",
  4429=>"111011111",
  4430=>"001000000",
  4431=>"000001001",
  4432=>"010110110",
  4433=>"111010111",
  4434=>"111000000",
  4435=>"111111011",
  4436=>"111111110",
  4437=>"011011011",
  4438=>"111111000",
  4439=>"111111111",
  4440=>"110000000",
  4441=>"001001111",
  4442=>"100000000",
  4443=>"111111111",
  4444=>"111111011",
  4445=>"000000000",
  4446=>"000000111",
  4447=>"111111111",
  4448=>"000001001",
  4449=>"111111111",
  4450=>"110010000",
  4451=>"101101111",
  4452=>"111111111",
  4453=>"011000000",
  4454=>"000000000",
  4455=>"111000110",
  4456=>"001000000",
  4457=>"100111001",
  4458=>"111111111",
  4459=>"111111110",
  4460=>"111111101",
  4461=>"000000000",
  4462=>"011111111",
  4463=>"110001000",
  4464=>"001000000",
  4465=>"001111111",
  4466=>"000111111",
  4467=>"100100000",
  4468=>"111111111",
  4469=>"001000000",
  4470=>"101111101",
  4471=>"111111110",
  4472=>"000110111",
  4473=>"111111111",
  4474=>"111111111",
  4475=>"000110000",
  4476=>"000000110",
  4477=>"100000000",
  4478=>"100000000",
  4479=>"111111111",
  4480=>"111001001",
  4481=>"011010111",
  4482=>"110100011",
  4483=>"011001000",
  4484=>"000100101",
  4485=>"000111111",
  4486=>"001000000",
  4487=>"111011000",
  4488=>"010000111",
  4489=>"001111111",
  4490=>"111101000",
  4491=>"111110000",
  4492=>"101001111",
  4493=>"000100111",
  4494=>"011111111",
  4495=>"000011000",
  4496=>"000010000",
  4497=>"000000000",
  4498=>"000011000",
  4499=>"100100001",
  4500=>"000011000",
  4501=>"000000001",
  4502=>"011011000",
  4503=>"000000000",
  4504=>"111011111",
  4505=>"001000110",
  4506=>"111111111",
  4507=>"111011111",
  4508=>"100110000",
  4509=>"000000000",
  4510=>"000000000",
  4511=>"000000000",
  4512=>"011011000",
  4513=>"000000111",
  4514=>"111111111",
  4515=>"111111111",
  4516=>"111100111",
  4517=>"001001000",
  4518=>"111111101",
  4519=>"111100111",
  4520=>"000000000",
  4521=>"001111111",
  4522=>"011111111",
  4523=>"000000000",
  4524=>"000000000",
  4525=>"111111111",
  4526=>"000010000",
  4527=>"110111111",
  4528=>"011001111",
  4529=>"010000000",
  4530=>"001111111",
  4531=>"011011110",
  4532=>"111111111",
  4533=>"010001110",
  4534=>"111111111",
  4535=>"011111100",
  4536=>"111110111",
  4537=>"111111111",
  4538=>"100100000",
  4539=>"110000101",
  4540=>"111111111",
  4541=>"110110000",
  4542=>"111111111",
  4543=>"100100101",
  4544=>"000000000",
  4545=>"111011111",
  4546=>"111111111",
  4547=>"000000001",
  4548=>"001000111",
  4549=>"100111111",
  4550=>"100000000",
  4551=>"000001011",
  4552=>"000000000",
  4553=>"000001001",
  4554=>"000000000",
  4555=>"111111000",
  4556=>"110000000",
  4557=>"100000000",
  4558=>"000000000",
  4559=>"101100000",
  4560=>"000000000",
  4561=>"111111111",
  4562=>"111101000",
  4563=>"000111011",
  4564=>"000000001",
  4565=>"111111111",
  4566=>"000000000",
  4567=>"001111111",
  4568=>"001000000",
  4569=>"000000000",
  4570=>"000000000",
  4571=>"000000001",
  4572=>"011011000",
  4573=>"001001000",
  4574=>"010000000",
  4575=>"000000000",
  4576=>"111111111",
  4577=>"000000000",
  4578=>"111110000",
  4579=>"000000000",
  4580=>"011011011",
  4581=>"011111111",
  4582=>"001000000",
  4583=>"000010000",
  4584=>"111111001",
  4585=>"100010010",
  4586=>"010000000",
  4587=>"000100111",
  4588=>"110000000",
  4589=>"011011111",
  4590=>"000000000",
  4591=>"000000000",
  4592=>"000000000",
  4593=>"100000000",
  4594=>"111111111",
  4595=>"000000000",
  4596=>"000000100",
  4597=>"111000000",
  4598=>"000000100",
  4599=>"111110001",
  4600=>"000000000",
  4601=>"001001011",
  4602=>"111111111",
  4603=>"111111111",
  4604=>"111110111",
  4605=>"110101101",
  4606=>"111111000",
  4607=>"000000000",
  4608=>"110110110",
  4609=>"111111110",
  4610=>"111001000",
  4611=>"111100000",
  4612=>"111111111",
  4613=>"111111111",
  4614=>"111111111",
  4615=>"000001011",
  4616=>"001001101",
  4617=>"110011111",
  4618=>"001001101",
  4619=>"000010011",
  4620=>"110111101",
  4621=>"101001101",
  4622=>"110111111",
  4623=>"101101101",
  4624=>"000001000",
  4625=>"110110010",
  4626=>"000000101",
  4627=>"111111001",
  4628=>"001000000",
  4629=>"111111000",
  4630=>"000010010",
  4631=>"010000001",
  4632=>"110110000",
  4633=>"101001101",
  4634=>"111011010",
  4635=>"111111011",
  4636=>"101001111",
  4637=>"000010110",
  4638=>"100101100",
  4639=>"111000101",
  4640=>"000100000",
  4641=>"111111111",
  4642=>"100110111",
  4643=>"001000000",
  4644=>"000000011",
  4645=>"111000111",
  4646=>"000110111",
  4647=>"000000000",
  4648=>"000000000",
  4649=>"001001001",
  4650=>"111111111",
  4651=>"111111010",
  4652=>"100100110",
  4653=>"110010010",
  4654=>"001001000",
  4655=>"000010111",
  4656=>"111111111",
  4657=>"000000001",
  4658=>"011110111",
  4659=>"000000101",
  4660=>"100000000",
  4661=>"001001011",
  4662=>"111000000",
  4663=>"111011000",
  4664=>"000000111",
  4665=>"111111010",
  4666=>"111111111",
  4667=>"101001001",
  4668=>"000000001",
  4669=>"110110010",
  4670=>"100111111",
  4671=>"111111110",
  4672=>"011011111",
  4673=>"100101001",
  4674=>"000000101",
  4675=>"010110000",
  4676=>"001001100",
  4677=>"000000000",
  4678=>"111111110",
  4679=>"000000110",
  4680=>"011011000",
  4681=>"111111110",
  4682=>"000011111",
  4683=>"001001011",
  4684=>"100111001",
  4685=>"110000100",
  4686=>"100000100",
  4687=>"000110110",
  4688=>"001001001",
  4689=>"000110000",
  4690=>"000000001",
  4691=>"000000000",
  4692=>"001000001",
  4693=>"110100010",
  4694=>"000111111",
  4695=>"111001000",
  4696=>"001001111",
  4697=>"101101111",
  4698=>"010010000",
  4699=>"011111111",
  4700=>"000000000",
  4701=>"000000000",
  4702=>"111111011",
  4703=>"001101011",
  4704=>"100000100",
  4705=>"110111000",
  4706=>"111101011",
  4707=>"111111111",
  4708=>"010010011",
  4709=>"111111111",
  4710=>"000000000",
  4711=>"010111111",
  4712=>"000000000",
  4713=>"000001111",
  4714=>"111101111",
  4715=>"000011001",
  4716=>"111110110",
  4717=>"111111010",
  4718=>"001001000",
  4719=>"000010010",
  4720=>"000001001",
  4721=>"001001100",
  4722=>"110100000",
  4723=>"011000101",
  4724=>"111111010",
  4725=>"110000000",
  4726=>"111111011",
  4727=>"111111111",
  4728=>"000000001",
  4729=>"010001001",
  4730=>"000000110",
  4731=>"000000000",
  4732=>"100000010",
  4733=>"000000001",
  4734=>"000000101",
  4735=>"001111111",
  4736=>"111101111",
  4737=>"110111000",
  4738=>"110111111",
  4739=>"010011001",
  4740=>"011111111",
  4741=>"101001001",
  4742=>"111111001",
  4743=>"111011000",
  4744=>"000000111",
  4745=>"000000001",
  4746=>"111111111",
  4747=>"111111111",
  4748=>"001001110",
  4749=>"001000001",
  4750=>"111111111",
  4751=>"111111111",
  4752=>"001001001",
  4753=>"000000000",
  4754=>"110110000",
  4755=>"000000100",
  4756=>"111111111",
  4757=>"111111001",
  4758=>"000000000",
  4759=>"110000000",
  4760=>"001001001",
  4761=>"001001111",
  4762=>"000000001",
  4763=>"111100000",
  4764=>"111001000",
  4765=>"011001001",
  4766=>"111000000",
  4767=>"111101001",
  4768=>"111011000",
  4769=>"111101101",
  4770=>"001111111",
  4771=>"000000000",
  4772=>"000001001",
  4773=>"111100100",
  4774=>"001001111",
  4775=>"000000110",
  4776=>"000000011",
  4777=>"111100111",
  4778=>"001001001",
  4779=>"111111100",
  4780=>"011111111",
  4781=>"000000000",
  4782=>"101111111",
  4783=>"000000110",
  4784=>"111111111",
  4785=>"101100110",
  4786=>"011011010",
  4787=>"111101000",
  4788=>"110000000",
  4789=>"000110111",
  4790=>"001111111",
  4791=>"000000000",
  4792=>"101001111",
  4793=>"000111011",
  4794=>"000000000",
  4795=>"000101100",
  4796=>"000111111",
  4797=>"000000111",
  4798=>"000000111",
  4799=>"111101101",
  4800=>"100000100",
  4801=>"111111110",
  4802=>"111001111",
  4803=>"110000000",
  4804=>"000000110",
  4805=>"001001111",
  4806=>"111110010",
  4807=>"000000001",
  4808=>"110011010",
  4809=>"000101111",
  4810=>"110011111",
  4811=>"001000000",
  4812=>"111011101",
  4813=>"000110000",
  4814=>"111111000",
  4815=>"110100000",
  4816=>"110110010",
  4817=>"011111111",
  4818=>"000000001",
  4819=>"001001111",
  4820=>"100000111",
  4821=>"000101001",
  4822=>"111010010",
  4823=>"111101011",
  4824=>"111111000",
  4825=>"101101111",
  4826=>"000000000",
  4827=>"000000000",
  4828=>"100111111",
  4829=>"000100111",
  4830=>"000000000",
  4831=>"001001101",
  4832=>"000000000",
  4833=>"000001001",
  4834=>"000011111",
  4835=>"111111000",
  4836=>"101001101",
  4837=>"100111011",
  4838=>"000000111",
  4839=>"110110110",
  4840=>"000110000",
  4841=>"000000101",
  4842=>"000000001",
  4843=>"111111000",
  4844=>"111111111",
  4845=>"111010000",
  4846=>"000100100",
  4847=>"101001000",
  4848=>"000000000",
  4849=>"000000011",
  4850=>"000000000",
  4851=>"000101101",
  4852=>"101001001",
  4853=>"110110110",
  4854=>"011111001",
  4855=>"000000000",
  4856=>"011001011",
  4857=>"111010000",
  4858=>"000000001",
  4859=>"101001111",
  4860=>"111111000",
  4861=>"110111110",
  4862=>"001100100",
  4863=>"111101111",
  4864=>"111110000",
  4865=>"000110110",
  4866=>"110100110",
  4867=>"100010000",
  4868=>"000000101",
  4869=>"111111100",
  4870=>"000111111",
  4871=>"000011011",
  4872=>"111111111",
  4873=>"101101111",
  4874=>"000001101",
  4875=>"110111010",
  4876=>"001000000",
  4877=>"000000000",
  4878=>"001001111",
  4879=>"000110101",
  4880=>"100110000",
  4881=>"001101101",
  4882=>"011011010",
  4883=>"000000111",
  4884=>"111111111",
  4885=>"110100011",
  4886=>"111111110",
  4887=>"110100111",
  4888=>"001000000",
  4889=>"010000000",
  4890=>"100100100",
  4891=>"000000100",
  4892=>"001001111",
  4893=>"110000111",
  4894=>"000110111",
  4895=>"000000000",
  4896=>"000100000",
  4897=>"001100100",
  4898=>"111111000",
  4899=>"000000000",
  4900=>"000110111",
  4901=>"110101010",
  4902=>"000000000",
  4903=>"111101100",
  4904=>"111111111",
  4905=>"000000001",
  4906=>"000000000",
  4907=>"000000000",
  4908=>"111111000",
  4909=>"000000000",
  4910=>"111011000",
  4911=>"100000000",
  4912=>"110100000",
  4913=>"111100100",
  4914=>"001001101",
  4915=>"101000000",
  4916=>"111111111",
  4917=>"111101111",
  4918=>"111011000",
  4919=>"111111101",
  4920=>"010010000",
  4921=>"011111111",
  4922=>"000101111",
  4923=>"100100111",
  4924=>"100000001",
  4925=>"110100001",
  4926=>"000111111",
  4927=>"111101101",
  4928=>"110111111",
  4929=>"111001101",
  4930=>"001111111",
  4931=>"010010010",
  4932=>"000001111",
  4933=>"000000000",
  4934=>"000010000",
  4935=>"000111111",
  4936=>"111111001",
  4937=>"000000000",
  4938=>"000000000",
  4939=>"011011111",
  4940=>"110000000",
  4941=>"001000000",
  4942=>"111111101",
  4943=>"111010111",
  4944=>"000000000",
  4945=>"000000000",
  4946=>"001000000",
  4947=>"010111011",
  4948=>"000000001",
  4949=>"011011000",
  4950=>"000000000",
  4951=>"111100000",
  4952=>"111111110",
  4953=>"011111000",
  4954=>"110110100",
  4955=>"000000111",
  4956=>"000000001",
  4957=>"001001100",
  4958=>"111101001",
  4959=>"110110101",
  4960=>"111111111",
  4961=>"100000000",
  4962=>"111111011",
  4963=>"000001000",
  4964=>"001111111",
  4965=>"000001100",
  4966=>"000010011",
  4967=>"110110011",
  4968=>"000010011",
  4969=>"000000110",
  4970=>"111111000",
  4971=>"111111111",
  4972=>"001001101",
  4973=>"000000000",
  4974=>"111001001",
  4975=>"111111111",
  4976=>"111111111",
  4977=>"001001101",
  4978=>"000000000",
  4979=>"100100111",
  4980=>"111111111",
  4981=>"111101111",
  4982=>"111111111",
  4983=>"000000000",
  4984=>"001111111",
  4985=>"000001010",
  4986=>"111111111",
  4987=>"110110000",
  4988=>"000101101",
  4989=>"000000000",
  4990=>"010000000",
  4991=>"000000101",
  4992=>"000000001",
  4993=>"110100000",
  4994=>"000000000",
  4995=>"101101111",
  4996=>"001001100",
  4997=>"000010010",
  4998=>"100101101",
  4999=>"111000000",
  5000=>"111111110",
  5001=>"000000111",
  5002=>"100100000",
  5003=>"010010000",
  5004=>"110110000",
  5005=>"001010110",
  5006=>"100110010",
  5007=>"111000000",
  5008=>"111111111",
  5009=>"111011011",
  5010=>"001001101",
  5011=>"000000100",
  5012=>"111111010",
  5013=>"010010010",
  5014=>"001000111",
  5015=>"100100001",
  5016=>"111001000",
  5017=>"000000111",
  5018=>"001000101",
  5019=>"000001111",
  5020=>"000011001",
  5021=>"011111010",
  5022=>"100100100",
  5023=>"000000000",
  5024=>"000001111",
  5025=>"100100000",
  5026=>"000110111",
  5027=>"000000000",
  5028=>"000000101",
  5029=>"000000000",
  5030=>"100100000",
  5031=>"000000000",
  5032=>"100101000",
  5033=>"111110000",
  5034=>"111101110",
  5035=>"111111111",
  5036=>"111101000",
  5037=>"100110100",
  5038=>"000001111",
  5039=>"010110011",
  5040=>"000111111",
  5041=>"000000000",
  5042=>"000000000",
  5043=>"001000001",
  5044=>"011110000",
  5045=>"001000111",
  5046=>"111111111",
  5047=>"010110000",
  5048=>"001001011",
  5049=>"110111111",
  5050=>"100100000",
  5051=>"100100111",
  5052=>"001001000",
  5053=>"111111100",
  5054=>"111111111",
  5055=>"100100101",
  5056=>"100000000",
  5057=>"111111111",
  5058=>"111111111",
  5059=>"111111110",
  5060=>"110110011",
  5061=>"000110011",
  5062=>"010010111",
  5063=>"001111111",
  5064=>"000001001",
  5065=>"100100111",
  5066=>"000001110",
  5067=>"000000000",
  5068=>"100001100",
  5069=>"000000000",
  5070=>"111111111",
  5071=>"111111000",
  5072=>"100101111",
  5073=>"100100100",
  5074=>"000000000",
  5075=>"111101000",
  5076=>"000110110",
  5077=>"100000000",
  5078=>"110111010",
  5079=>"000110101",
  5080=>"111111110",
  5081=>"100110001",
  5082=>"000000000",
  5083=>"111111111",
  5084=>"001000000",
  5085=>"111101110",
  5086=>"011011000",
  5087=>"000000111",
  5088=>"001111111",
  5089=>"110100111",
  5090=>"000000000",
  5091=>"100111111",
  5092=>"110110111",
  5093=>"000111111",
  5094=>"001011000",
  5095=>"000000000",
  5096=>"110110110",
  5097=>"100110000",
  5098=>"000010000",
  5099=>"001001001",
  5100=>"000000101",
  5101=>"011011000",
  5102=>"000000110",
  5103=>"100111111",
  5104=>"101000000",
  5105=>"111111111",
  5106=>"110000000",
  5107=>"001111111",
  5108=>"000000101",
  5109=>"001000000",
  5110=>"111101101",
  5111=>"010010001",
  5112=>"011011111",
  5113=>"111100110",
  5114=>"110110110",
  5115=>"000000000",
  5116=>"001111111",
  5117=>"110010010",
  5118=>"110100101",
  5119=>"101100001",
  5120=>"111100111",
  5121=>"000000011",
  5122=>"111111000",
  5123=>"100000000",
  5124=>"000111111",
  5125=>"111000000",
  5126=>"110000000",
  5127=>"111111111",
  5128=>"011000000",
  5129=>"000000111",
  5130=>"000000000",
  5131=>"000000111",
  5132=>"110100100",
  5133=>"100110111",
  5134=>"000000011",
  5135=>"111000010",
  5136=>"111111111",
  5137=>"000000000",
  5138=>"111111111",
  5139=>"111000000",
  5140=>"000000000",
  5141=>"000000111",
  5142=>"110000110",
  5143=>"111111111",
  5144=>"000000001",
  5145=>"001010000",
  5146=>"001000001",
  5147=>"011000000",
  5148=>"000000000",
  5149=>"000110110",
  5150=>"111100001",
  5151=>"111010000",
  5152=>"110000000",
  5153=>"111111111",
  5154=>"011111100",
  5155=>"101011011",
  5156=>"111010010",
  5157=>"111111011",
  5158=>"000111111",
  5159=>"011110100",
  5160=>"011010000",
  5161=>"000000000",
  5162=>"011010111",
  5163=>"000000000",
  5164=>"001111111",
  5165=>"111111111",
  5166=>"100111101",
  5167=>"000000000",
  5168=>"111111111",
  5169=>"111110001",
  5170=>"000000001",
  5171=>"000100111",
  5172=>"011100000",
  5173=>"110110000",
  5174=>"001000110",
  5175=>"000000111",
  5176=>"000011111",
  5177=>"000100000",
  5178=>"110000000",
  5179=>"000000000",
  5180=>"000000000",
  5181=>"000000000",
  5182=>"011011000",
  5183=>"001000110",
  5184=>"110111000",
  5185=>"011011011",
  5186=>"001111111",
  5187=>"111011111",
  5188=>"000000001",
  5189=>"000001001",
  5190=>"001011111",
  5191=>"111111000",
  5192=>"001011011",
  5193=>"000000001",
  5194=>"011000000",
  5195=>"000000110",
  5196=>"111111111",
  5197=>"000010111",
  5198=>"111110000",
  5199=>"000011001",
  5200=>"000000111",
  5201=>"111000011",
  5202=>"001000000",
  5203=>"111110000",
  5204=>"000010000",
  5205=>"011000000",
  5206=>"111000111",
  5207=>"000001111",
  5208=>"111000100",
  5209=>"000000000",
  5210=>"000000111",
  5211=>"111011000",
  5212=>"000000000",
  5213=>"111111110",
  5214=>"001100110",
  5215=>"111011001",
  5216=>"111000000",
  5217=>"001000011",
  5218=>"000000000",
  5219=>"000000000",
  5220=>"001000000",
  5221=>"111011000",
  5222=>"000100111",
  5223=>"000000000",
  5224=>"000001000",
  5225=>"000000001",
  5226=>"111111110",
  5227=>"011000111",
  5228=>"000000000",
  5229=>"111001000",
  5230=>"111111111",
  5231=>"111001000",
  5232=>"000000011",
  5233=>"000001111",
  5234=>"001011111",
  5235=>"111111111",
  5236=>"000000111",
  5237=>"111111110",
  5238=>"000000000",
  5239=>"000000000",
  5240=>"101111111",
  5241=>"011111011",
  5242=>"000000000",
  5243=>"000000010",
  5244=>"110100011",
  5245=>"000000000",
  5246=>"001000000",
  5247=>"000001111",
  5248=>"011001000",
  5249=>"111111111",
  5250=>"111100000",
  5251=>"000000001",
  5252=>"111110000",
  5253=>"000000000",
  5254=>"111111100",
  5255=>"110111110",
  5256=>"000010000",
  5257=>"000000111",
  5258=>"000000000",
  5259=>"001111111",
  5260=>"000000000",
  5261=>"000000000",
  5262=>"111111011",
  5263=>"110110100",
  5264=>"000000111",
  5265=>"000111111",
  5266=>"000000111",
  5267=>"110111111",
  5268=>"000100000",
  5269=>"000000001",
  5270=>"000000000",
  5271=>"011000001",
  5272=>"001001001",
  5273=>"000001011",
  5274=>"011000111",
  5275=>"000111111",
  5276=>"111001110",
  5277=>"000000000",
  5278=>"110000110",
  5279=>"100000000",
  5280=>"111110000",
  5281=>"011001000",
  5282=>"000000001",
  5283=>"110110111",
  5284=>"000000001",
  5285=>"111000000",
  5286=>"100111111",
  5287=>"001101101",
  5288=>"011000111",
  5289=>"000000000",
  5290=>"000111111",
  5291=>"110111001",
  5292=>"000100111",
  5293=>"011111001",
  5294=>"010010010",
  5295=>"010000010",
  5296=>"010110111",
  5297=>"000001011",
  5298=>"111111111",
  5299=>"111000000",
  5300=>"111000001",
  5301=>"000000000",
  5302=>"111111000",
  5303=>"111111000",
  5304=>"111111110",
  5305=>"000000101",
  5306=>"100000000",
  5307=>"111111111",
  5308=>"100111110",
  5309=>"101001000",
  5310=>"111000001",
  5311=>"000111111",
  5312=>"000000000",
  5313=>"000000000",
  5314=>"111011111",
  5315=>"000100000",
  5316=>"000000000",
  5317=>"111111000",
  5318=>"000000000",
  5319=>"000111111",
  5320=>"000000110",
  5321=>"001000001",
  5322=>"001000000",
  5323=>"000111111",
  5324=>"000000111",
  5325=>"000000111",
  5326=>"000000111",
  5327=>"000000010",
  5328=>"000000000",
  5329=>"000010111",
  5330=>"000001000",
  5331=>"110000000",
  5332=>"100100111",
  5333=>"001001011",
  5334=>"101111000",
  5335=>"000000000",
  5336=>"111011111",
  5337=>"000000100",
  5338=>"000000000",
  5339=>"011000000",
  5340=>"111111000",
  5341=>"101101111",
  5342=>"111111111",
  5343=>"111000000",
  5344=>"001001111",
  5345=>"000001000",
  5346=>"100100000",
  5347=>"111111111",
  5348=>"110110000",
  5349=>"111000000",
  5350=>"001000111",
  5351=>"001011111",
  5352=>"111111000",
  5353=>"000000010",
  5354=>"110111000",
  5355=>"000000001",
  5356=>"111110011",
  5357=>"111000000",
  5358=>"100100001",
  5359=>"000000011",
  5360=>"000000000",
  5361=>"111000000",
  5362=>"111111001",
  5363=>"000000111",
  5364=>"111111000",
  5365=>"111110000",
  5366=>"001111111",
  5367=>"001101000",
  5368=>"111111011",
  5369=>"000111000",
  5370=>"000101111",
  5371=>"000111000",
  5372=>"111011001",
  5373=>"001000000",
  5374=>"010000100",
  5375=>"110111111",
  5376=>"111111110",
  5377=>"111001101",
  5378=>"000000000",
  5379=>"111111111",
  5380=>"101000001",
  5381=>"000011000",
  5382=>"000000000",
  5383=>"111110111",
  5384=>"111111000",
  5385=>"000000000",
  5386=>"000001100",
  5387=>"011000010",
  5388=>"111001101",
  5389=>"101111111",
  5390=>"000000110",
  5391=>"000101111",
  5392=>"111000001",
  5393=>"111110111",
  5394=>"001000000",
  5395=>"001001000",
  5396=>"110111100",
  5397=>"111100000",
  5398=>"001111110",
  5399=>"111111111",
  5400=>"111011011",
  5401=>"000000000",
  5402=>"111000110",
  5403=>"010010000",
  5404=>"111001000",
  5405=>"000000000",
  5406=>"000000011",
  5407=>"111111111",
  5408=>"100111000",
  5409=>"000000011",
  5410=>"000000000",
  5411=>"000011111",
  5412=>"111010000",
  5413=>"000000000",
  5414=>"100110111",
  5415=>"000000100",
  5416=>"111000000",
  5417=>"001000001",
  5418=>"111000000",
  5419=>"111100000",
  5420=>"000000100",
  5421=>"000111111",
  5422=>"000000111",
  5423=>"001000100",
  5424=>"110111111",
  5425=>"000000110",
  5426=>"001011111",
  5427=>"101111000",
  5428=>"000000000",
  5429=>"000110111",
  5430=>"110000010",
  5431=>"000000011",
  5432=>"000000011",
  5433=>"000000000",
  5434=>"000000110",
  5435=>"111111000",
  5436=>"001111111",
  5437=>"100000000",
  5438=>"110000001",
  5439=>"111111010",
  5440=>"000000000",
  5441=>"000111111",
  5442=>"111000000",
  5443=>"000111111",
  5444=>"000000110",
  5445=>"110000000",
  5446=>"011000000",
  5447=>"111000000",
  5448=>"111100000",
  5449=>"000000001",
  5450=>"000000000",
  5451=>"001111000",
  5452=>"000000000",
  5453=>"011000001",
  5454=>"111000000",
  5455=>"001001001",
  5456=>"111100000",
  5457=>"000001111",
  5458=>"111111111",
  5459=>"111000000",
  5460=>"011011111",
  5461=>"011011011",
  5462=>"110100111",
  5463=>"011011011",
  5464=>"111111111",
  5465=>"111010000",
  5466=>"111111111",
  5467=>"101001010",
  5468=>"111011011",
  5469=>"000000000",
  5470=>"110000000",
  5471=>"100000000",
  5472=>"011011111",
  5473=>"000000000",
  5474=>"000011011",
  5475=>"111111011",
  5476=>"000010110",
  5477=>"011011111",
  5478=>"111111000",
  5479=>"000000111",
  5480=>"111111000",
  5481=>"000111111",
  5482=>"110100111",
  5483=>"000001111",
  5484=>"000001011",
  5485=>"000001111",
  5486=>"111000000",
  5487=>"111000111",
  5488=>"100001101",
  5489=>"111111001",
  5490=>"000000011",
  5491=>"111111111",
  5492=>"111111111",
  5493=>"001000010",
  5494=>"111110111",
  5495=>"000000110",
  5496=>"111000000",
  5497=>"000000111",
  5498=>"001001000",
  5499=>"000000111",
  5500=>"111111111",
  5501=>"000110111",
  5502=>"000000001",
  5503=>"000000000",
  5504=>"111000000",
  5505=>"111111000",
  5506=>"000100100",
  5507=>"000101111",
  5508=>"111000011",
  5509=>"000000010",
  5510=>"100000000",
  5511=>"000000000",
  5512=>"001001000",
  5513=>"000111111",
  5514=>"111111111",
  5515=>"011000000",
  5516=>"111101111",
  5517=>"011111111",
  5518=>"111111111",
  5519=>"000000111",
  5520=>"000000111",
  5521=>"001111101",
  5522=>"000010110",
  5523=>"111111110",
  5524=>"000000000",
  5525=>"000000000",
  5526=>"011000000",
  5527=>"100001001",
  5528=>"110111111",
  5529=>"100110111",
  5530=>"000000001",
  5531=>"111011000",
  5532=>"000000000",
  5533=>"110111000",
  5534=>"110000000",
  5535=>"000000111",
  5536=>"000111111",
  5537=>"110100100",
  5538=>"000000100",
  5539=>"000110111",
  5540=>"111011000",
  5541=>"111111000",
  5542=>"111111001",
  5543=>"101100011",
  5544=>"111000000",
  5545=>"111000000",
  5546=>"110110000",
  5547=>"000000000",
  5548=>"111000101",
  5549=>"111001011",
  5550=>"111100000",
  5551=>"111111110",
  5552=>"000000000",
  5553=>"010000001",
  5554=>"010000000",
  5555=>"000000000",
  5556=>"011111111",
  5557=>"111010111",
  5558=>"000000111",
  5559=>"000000000",
  5560=>"001101100",
  5561=>"000111111",
  5562=>"100110001",
  5563=>"001010011",
  5564=>"100100100",
  5565=>"111110000",
  5566=>"110000000",
  5567=>"001011111",
  5568=>"111111110",
  5569=>"001011110",
  5570=>"000000001",
  5571=>"001000000",
  5572=>"111111010",
  5573=>"111001001",
  5574=>"000110111",
  5575=>"000100000",
  5576=>"111111110",
  5577=>"111011000",
  5578=>"111001000",
  5579=>"000000000",
  5580=>"111111000",
  5581=>"111010011",
  5582=>"111110010",
  5583=>"000000000",
  5584=>"000000000",
  5585=>"111000101",
  5586=>"000111111",
  5587=>"111111111",
  5588=>"111110111",
  5589=>"110010000",
  5590=>"111000010",
  5591=>"001001001",
  5592=>"101001000",
  5593=>"000000000",
  5594=>"101111111",
  5595=>"101110110",
  5596=>"111111111",
  5597=>"111010000",
  5598=>"111100111",
  5599=>"101001101",
  5600=>"000001001",
  5601=>"000001000",
  5602=>"111111111",
  5603=>"111111001",
  5604=>"100000000",
  5605=>"000001111",
  5606=>"110000000",
  5607=>"000011111",
  5608=>"000000011",
  5609=>"111111000",
  5610=>"000000000",
  5611=>"000000000",
  5612=>"000000000",
  5613=>"010111110",
  5614=>"000001011",
  5615=>"111111111",
  5616=>"000000111",
  5617=>"011111111",
  5618=>"111111100",
  5619=>"000011111",
  5620=>"111111111",
  5621=>"000000100",
  5622=>"111111011",
  5623=>"111111111",
  5624=>"101111000",
  5625=>"101000000",
  5626=>"000000000",
  5627=>"111011011",
  5628=>"110000000",
  5629=>"111101011",
  5630=>"000000000",
  5631=>"110110010",
  5632=>"111101100",
  5633=>"000000000",
  5634=>"000000000",
  5635=>"111111111",
  5636=>"000000000",
  5637=>"111111101",
  5638=>"001001111",
  5639=>"111111111",
  5640=>"000000001",
  5641=>"000000010",
  5642=>"000000000",
  5643=>"110111111",
  5644=>"001000100",
  5645=>"110000000",
  5646=>"101100101",
  5647=>"000000000",
  5648=>"000000000",
  5649=>"111111011",
  5650=>"011011001",
  5651=>"111111100",
  5652=>"000100111",
  5653=>"000000111",
  5654=>"000000000",
  5655=>"111111110",
  5656=>"000000000",
  5657=>"001000110",
  5658=>"100100100",
  5659=>"000000000",
  5660=>"101111011",
  5661=>"000000100",
  5662=>"111101101",
  5663=>"011000000",
  5664=>"111000000",
  5665=>"011001111",
  5666=>"111111111",
  5667=>"111000000",
  5668=>"111111000",
  5669=>"111111111",
  5670=>"011111100",
  5671=>"000000000",
  5672=>"001000000",
  5673=>"111111000",
  5674=>"101100111",
  5675=>"111111111",
  5676=>"111000111",
  5677=>"111101000",
  5678=>"011000001",
  5679=>"111111111",
  5680=>"111011000",
  5681=>"000000000",
  5682=>"000000000",
  5683=>"011001011",
  5684=>"111101101",
  5685=>"000000000",
  5686=>"111111001",
  5687=>"110111110",
  5688=>"000111011",
  5689=>"100000110",
  5690=>"111101000",
  5691=>"000000100",
  5692=>"101000001",
  5693=>"000000011",
  5694=>"000000000",
  5695=>"100000101",
  5696=>"110100110",
  5697=>"000000100",
  5698=>"111001000",
  5699=>"111111110",
  5700=>"000000000",
  5701=>"110111111",
  5702=>"000000000",
  5703=>"111110000",
  5704=>"101111100",
  5705=>"111111110",
  5706=>"111111111",
  5707=>"110010111",
  5708=>"100000000",
  5709=>"011111111",
  5710=>"001011111",
  5711=>"001111111",
  5712=>"100111111",
  5713=>"000000000",
  5714=>"101111111",
  5715=>"001011000",
  5716=>"000000011",
  5717=>"000000000",
  5718=>"100000000",
  5719=>"111111001",
  5720=>"110111111",
  5721=>"111111111",
  5722=>"111111111",
  5723=>"000111111",
  5724=>"000100100",
  5725=>"000000111",
  5726=>"000000000",
  5727=>"001001000",
  5728=>"000000000",
  5729=>"110100000",
  5730=>"111111111",
  5731=>"100000111",
  5732=>"000010111",
  5733=>"000000000",
  5734=>"111101111",
  5735=>"100111111",
  5736=>"000000111",
  5737=>"001101000",
  5738=>"000000010",
  5739=>"100101111",
  5740=>"000000000",
  5741=>"111111111",
  5742=>"111111001",
  5743=>"000000000",
  5744=>"111111111",
  5745=>"011011111",
  5746=>"001000000",
  5747=>"000000000",
  5748=>"000011011",
  5749=>"101110110",
  5750=>"111111111",
  5751=>"000000011",
  5752=>"000000000",
  5753=>"100110111",
  5754=>"111111111",
  5755=>"111000110",
  5756=>"110110110",
  5757=>"000000000",
  5758=>"011001111",
  5759=>"000110100",
  5760=>"000000000",
  5761=>"000000101",
  5762=>"110110111",
  5763=>"011001000",
  5764=>"111111111",
  5765=>"111111101",
  5766=>"111110110",
  5767=>"000000111",
  5768=>"111111111",
  5769=>"000000000",
  5770=>"000000000",
  5771=>"000000111",
  5772=>"000001001",
  5773=>"001001000",
  5774=>"010010111",
  5775=>"000000000",
  5776=>"111100111",
  5777=>"010011001",
  5778=>"111111100",
  5779=>"000000111",
  5780=>"110110111",
  5781=>"000100000",
  5782=>"111111111",
  5783=>"111110111",
  5784=>"000000000",
  5785=>"111111111",
  5786=>"000000000",
  5787=>"111111110",
  5788=>"110000000",
  5789=>"000000000",
  5790=>"110100100",
  5791=>"000000000",
  5792=>"111111111",
  5793=>"000000000",
  5794=>"011011011",
  5795=>"000000000",
  5796=>"000010110",
  5797=>"111111111",
  5798=>"000101101",
  5799=>"001001001",
  5800=>"000111111",
  5801=>"000000000",
  5802=>"100000000",
  5803=>"111011111",
  5804=>"000000000",
  5805=>"111111111",
  5806=>"111001111",
  5807=>"111111111",
  5808=>"110110010",
  5809=>"000100000",
  5810=>"111111111",
  5811=>"111111101",
  5812=>"110110001",
  5813=>"111111000",
  5814=>"010001000",
  5815=>"111111111",
  5816=>"111000000",
  5817=>"000000111",
  5818=>"000000000",
  5819=>"100000001",
  5820=>"100100110",
  5821=>"111111110",
  5822=>"000111000",
  5823=>"000000000",
  5824=>"111111111",
  5825=>"000000000",
  5826=>"111011100",
  5827=>"000001111",
  5828=>"000000000",
  5829=>"110100000",
  5830=>"000000000",
  5831=>"000000000",
  5832=>"111110110",
  5833=>"000011000",
  5834=>"010011101",
  5835=>"000000000",
  5836=>"000100000",
  5837=>"000000000",
  5838=>"111111111",
  5839=>"111111101",
  5840=>"000000000",
  5841=>"000000001",
  5842=>"000000100",
  5843=>"000000000",
  5844=>"111011110",
  5845=>"110000000",
  5846=>"000111111",
  5847=>"000000110",
  5848=>"111111110",
  5849=>"100100110",
  5850=>"000111110",
  5851=>"000000000",
  5852=>"100000000",
  5853=>"000000011",
  5854=>"000110110",
  5855=>"100000100",
  5856=>"100000000",
  5857=>"000111111",
  5858=>"111111111",
  5859=>"111110000",
  5860=>"000000000",
  5861=>"011001000",
  5862=>"000000111",
  5863=>"001111111",
  5864=>"011111000",
  5865=>"100100111",
  5866=>"000001001",
  5867=>"110111111",
  5868=>"101111111",
  5869=>"111111111",
  5870=>"000100111",
  5871=>"000000000",
  5872=>"000101011",
  5873=>"000000000",
  5874=>"001000000",
  5875=>"000011011",
  5876=>"111000000",
  5877=>"111111111",
  5878=>"000000000",
  5879=>"001101111",
  5880=>"111011011",
  5881=>"111100000",
  5882=>"001000000",
  5883=>"000000000",
  5884=>"000000000",
  5885=>"110110110",
  5886=>"001010111",
  5887=>"111111111",
  5888=>"011111000",
  5889=>"000000000",
  5890=>"111001000",
  5891=>"111111111",
  5892=>"001000000",
  5893=>"000000000",
  5894=>"000000111",
  5895=>"110000101",
  5896=>"001001001",
  5897=>"000000000",
  5898=>"111111111",
  5899=>"111111111",
  5900=>"000000111",
  5901=>"000000010",
  5902=>"111111111",
  5903=>"100000000",
  5904=>"111101111",
  5905=>"000011011",
  5906=>"111111000",
  5907=>"010110110",
  5908=>"010111010",
  5909=>"010000011",
  5910=>"111111101",
  5911=>"111011011",
  5912=>"111111110",
  5913=>"100110110",
  5914=>"111111111",
  5915=>"010010000",
  5916=>"000000010",
  5917=>"011111110",
  5918=>"000000000",
  5919=>"111111101",
  5920=>"100100000",
  5921=>"000000000",
  5922=>"111111110",
  5923=>"001111011",
  5924=>"100100101",
  5925=>"000000111",
  5926=>"110100100",
  5927=>"111111000",
  5928=>"100000000",
  5929=>"111001000",
  5930=>"111000100",
  5931=>"111101111",
  5932=>"000000000",
  5933=>"000000000",
  5934=>"000000001",
  5935=>"000100000",
  5936=>"100111100",
  5937=>"111111000",
  5938=>"111111011",
  5939=>"000000000",
  5940=>"000000111",
  5941=>"111111111",
  5942=>"000000000",
  5943=>"111000000",
  5944=>"000000000",
  5945=>"111111111",
  5946=>"000000011",
  5947=>"000000100",
  5948=>"000000000",
  5949=>"111111111",
  5950=>"000000000",
  5951=>"000000000",
  5952=>"000000000",
  5953=>"111111111",
  5954=>"011011000",
  5955=>"010000000",
  5956=>"000000010",
  5957=>"111111111",
  5958=>"000000000",
  5959=>"000000000",
  5960=>"001111111",
  5961=>"111111111",
  5962=>"000001011",
  5963=>"000100000",
  5964=>"111111111",
  5965=>"000000000",
  5966=>"110110111",
  5967=>"110000000",
  5968=>"100100000",
  5969=>"111111111",
  5970=>"110100010",
  5971=>"101111000",
  5972=>"000000110",
  5973=>"111111011",
  5974=>"100000000",
  5975=>"111011111",
  5976=>"100101000",
  5977=>"000000000",
  5978=>"110100000",
  5979=>"101100110",
  5980=>"111111011",
  5981=>"111000000",
  5982=>"001001000",
  5983=>"011001111",
  5984=>"000000000",
  5985=>"001000000",
  5986=>"010010000",
  5987=>"000001111",
  5988=>"000000000",
  5989=>"010111111",
  5990=>"000000000",
  5991=>"111111111",
  5992=>"101101101",
  5993=>"111111011",
  5994=>"101101000",
  5995=>"100111111",
  5996=>"111111111",
  5997=>"110000010",
  5998=>"010000000",
  5999=>"111111111",
  6000=>"010000000",
  6001=>"111000000",
  6002=>"111111111",
  6003=>"001001000",
  6004=>"000000010",
  6005=>"111111111",
  6006=>"000000000",
  6007=>"000110000",
  6008=>"000000000",
  6009=>"000000000",
  6010=>"111111000",
  6011=>"111101000",
  6012=>"101110000",
  6013=>"111111111",
  6014=>"000000100",
  6015=>"110111111",
  6016=>"111110111",
  6017=>"110000001",
  6018=>"111111111",
  6019=>"010010000",
  6020=>"100111011",
  6021=>"111111111",
  6022=>"000000100",
  6023=>"000111111",
  6024=>"010010000",
  6025=>"011111100",
  6026=>"011111111",
  6027=>"111111011",
  6028=>"111111111",
  6029=>"111100000",
  6030=>"011111110",
  6031=>"001001000",
  6032=>"111111111",
  6033=>"000000000",
  6034=>"000000110",
  6035=>"000000000",
  6036=>"111001000",
  6037=>"000000000",
  6038=>"110111111",
  6039=>"000000000",
  6040=>"000110000",
  6041=>"101000001",
  6042=>"000000100",
  6043=>"000000111",
  6044=>"000000001",
  6045=>"000000000",
  6046=>"000000000",
  6047=>"000100000",
  6048=>"001000000",
  6049=>"100110110",
  6050=>"111111111",
  6051=>"101011010",
  6052=>"011000001",
  6053=>"000000000",
  6054=>"101101111",
  6055=>"000000000",
  6056=>"001000000",
  6057=>"100111111",
  6058=>"101010111",
  6059=>"111111111",
  6060=>"011011000",
  6061=>"110100111",
  6062=>"001011111",
  6063=>"000000000",
  6064=>"000000000",
  6065=>"111111111",
  6066=>"000111111",
  6067=>"111111000",
  6068=>"111100000",
  6069=>"000000000",
  6070=>"111111111",
  6071=>"000000000",
  6072=>"000000111",
  6073=>"111111100",
  6074=>"010000000",
  6075=>"111111111",
  6076=>"111111111",
  6077=>"001111110",
  6078=>"000000000",
  6079=>"111111111",
  6080=>"111001111",
  6081=>"000000000",
  6082=>"000000000",
  6083=>"111111111",
  6084=>"010001001",
  6085=>"000000111",
  6086=>"000000000",
  6087=>"000000111",
  6088=>"011111111",
  6089=>"111111011",
  6090=>"000000100",
  6091=>"111111111",
  6092=>"011111111",
  6093=>"101001000",
  6094=>"100000000",
  6095=>"111111100",
  6096=>"000000100",
  6097=>"111111111",
  6098=>"001001111",
  6099=>"000000000",
  6100=>"100000101",
  6101=>"011111111",
  6102=>"000000110",
  6103=>"000000000",
  6104=>"000000000",
  6105=>"110000000",
  6106=>"001111111",
  6107=>"110111111",
  6108=>"000011111",
  6109=>"000000000",
  6110=>"111011000",
  6111=>"000000000",
  6112=>"000000000",
  6113=>"000000000",
  6114=>"111111111",
  6115=>"111111111",
  6116=>"110111111",
  6117=>"111111111",
  6118=>"000000000",
  6119=>"001111111",
  6120=>"000000100",
  6121=>"000000000",
  6122=>"000000000",
  6123=>"000000000",
  6124=>"111000100",
  6125=>"001000000",
  6126=>"000000000",
  6127=>"100111111",
  6128=>"001011011",
  6129=>"000000000",
  6130=>"000000000",
  6131=>"111110000",
  6132=>"100000000",
  6133=>"111111111",
  6134=>"000001000",
  6135=>"111111111",
  6136=>"001000111",
  6137=>"110100000",
  6138=>"000000000",
  6139=>"111111111",
  6140=>"111111111",
  6141=>"110000000",
  6142=>"100111111",
  6143=>"100111111",
  6144=>"001111111",
  6145=>"001000000",
  6146=>"000000001",
  6147=>"000000000",
  6148=>"111011111",
  6149=>"001000000",
  6150=>"100111111",
  6151=>"111111111",
  6152=>"111011000",
  6153=>"000000111",
  6154=>"100000000",
  6155=>"111100110",
  6156=>"001001011",
  6157=>"000111011",
  6158=>"000100100",
  6159=>"101111100",
  6160=>"111111111",
  6161=>"100000000",
  6162=>"001000110",
  6163=>"111111111",
  6164=>"000000001",
  6165=>"000000111",
  6166=>"000000011",
  6167=>"000000111",
  6168=>"000011111",
  6169=>"000000000",
  6170=>"001111011",
  6171=>"111111010",
  6172=>"000000000",
  6173=>"110000000",
  6174=>"001111111",
  6175=>"000001001",
  6176=>"111111001",
  6177=>"110111111",
  6178=>"000001111",
  6179=>"000000001",
  6180=>"100000000",
  6181=>"111111111",
  6182=>"111000000",
  6183=>"111011000",
  6184=>"001001000",
  6185=>"100111000",
  6186=>"000000000",
  6187=>"100100100",
  6188=>"111110110",
  6189=>"000000000",
  6190=>"111111001",
  6191=>"000010000",
  6192=>"001001111",
  6193=>"000001001",
  6194=>"111111001",
  6195=>"110010000",
  6196=>"110110000",
  6197=>"000000110",
  6198=>"111111111",
  6199=>"000000111",
  6200=>"000110100",
  6201=>"111111111",
  6202=>"000001001",
  6203=>"010000000",
  6204=>"111111000",
  6205=>"101000000",
  6206=>"111100000",
  6207=>"001111111",
  6208=>"111111000",
  6209=>"110000000",
  6210=>"000000000",
  6211=>"000000000",
  6212=>"000011011",
  6213=>"000000000",
  6214=>"001001000",
  6215=>"111111111",
  6216=>"001111000",
  6217=>"111111100",
  6218=>"000100110",
  6219=>"100000110",
  6220=>"010000000",
  6221=>"110000011",
  6222=>"011000000",
  6223=>"111000000",
  6224=>"111111001",
  6225=>"111111111",
  6226=>"000000000",
  6227=>"011011011",
  6228=>"000000000",
  6229=>"110111001",
  6230=>"111000000",
  6231=>"101101000",
  6232=>"001001000",
  6233=>"000000100",
  6234=>"000000000",
  6235=>"001000000",
  6236=>"000000000",
  6237=>"111111111",
  6238=>"100110000",
  6239=>"000000000",
  6240=>"111010000",
  6241=>"000000010",
  6242=>"111111111",
  6243=>"000000110",
  6244=>"000000001",
  6245=>"010010111",
  6246=>"000000000",
  6247=>"100111111",
  6248=>"000000111",
  6249=>"111000001",
  6250=>"111110111",
  6251=>"111111111",
  6252=>"010111110",
  6253=>"000000000",
  6254=>"111000110",
  6255=>"000000111",
  6256=>"000111111",
  6257=>"010000000",
  6258=>"000000011",
  6259=>"100111100",
  6260=>"101101111",
  6261=>"010111111",
  6262=>"011001011",
  6263=>"001000000",
  6264=>"101110000",
  6265=>"101111111",
  6266=>"111101100",
  6267=>"000001001",
  6268=>"011000010",
  6269=>"000000000",
  6270=>"000111110",
  6271=>"000000011",
  6272=>"100000000",
  6273=>"000010111",
  6274=>"111100111",
  6275=>"001101000",
  6276=>"111111111",
  6277=>"111000000",
  6278=>"111111111",
  6279=>"000010111",
  6280=>"111111000",
  6281=>"001100111",
  6282=>"000000000",
  6283=>"111111111",
  6284=>"111111111",
  6285=>"101000111",
  6286=>"010000100",
  6287=>"000111111",
  6288=>"100000000",
  6289=>"000101111",
  6290=>"000000111",
  6291=>"001000010",
  6292=>"111111111",
  6293=>"100111001",
  6294=>"111111000",
  6295=>"000100000",
  6296=>"101111111",
  6297=>"111110111",
  6298=>"111111111",
  6299=>"000010000",
  6300=>"100101101",
  6301=>"000011001",
  6302=>"111110101",
  6303=>"000000000",
  6304=>"000010010",
  6305=>"101101000",
  6306=>"000100111",
  6307=>"101000010",
  6308=>"011111001",
  6309=>"000000111",
  6310=>"000011010",
  6311=>"001011011",
  6312=>"111111111",
  6313=>"000101000",
  6314=>"000000100",
  6315=>"000100111",
  6316=>"000000100",
  6317=>"000000000",
  6318=>"100111110",
  6319=>"000000100",
  6320=>"000000111",
  6321=>"000011010",
  6322=>"111111111",
  6323=>"111101101",
  6324=>"111111110",
  6325=>"000000000",
  6326=>"001001000",
  6327=>"110110000",
  6328=>"001111000",
  6329=>"001000000",
  6330=>"000000000",
  6331=>"011111111",
  6332=>"000000000",
  6333=>"111111000",
  6334=>"000000111",
  6335=>"111111111",
  6336=>"000000111",
  6337=>"111111000",
  6338=>"111111111",
  6339=>"111111000",
  6340=>"000000111",
  6341=>"000111111",
  6342=>"101111100",
  6343=>"000110000",
  6344=>"101111011",
  6345=>"111111110",
  6346=>"111111111",
  6347=>"111111000",
  6348=>"000000110",
  6349=>"100110000",
  6350=>"111111000",
  6351=>"111000000",
  6352=>"000000000",
  6353=>"001000000",
  6354=>"001000000",
  6355=>"100000000",
  6356=>"000000111",
  6357=>"111111000",
  6358=>"111001011",
  6359=>"000000100",
  6360=>"100111111",
  6361=>"000111110",
  6362=>"000111111",
  6363=>"000000111",
  6364=>"000111011",
  6365=>"111111001",
  6366=>"101001111",
  6367=>"111111111",
  6368=>"000000000",
  6369=>"001000000",
  6370=>"000000011",
  6371=>"111111111",
  6372=>"000101101",
  6373=>"110110001",
  6374=>"000000110",
  6375=>"110101000",
  6376=>"000111000",
  6377=>"111001001",
  6378=>"111111110",
  6379=>"000000000",
  6380=>"011000000",
  6381=>"111110000",
  6382=>"111111000",
  6383=>"111000000",
  6384=>"000010000",
  6385=>"100100111",
  6386=>"111111000",
  6387=>"111111111",
  6388=>"000000000",
  6389=>"000000000",
  6390=>"101110111",
  6391=>"101111000",
  6392=>"100111000",
  6393=>"000000000",
  6394=>"011011011",
  6395=>"000000110",
  6396=>"000000000",
  6397=>"011011001",
  6398=>"000000101",
  6399=>"000000000",
  6400=>"111011000",
  6401=>"111011000",
  6402=>"010000100",
  6403=>"000000100",
  6404=>"000000000",
  6405=>"000000000",
  6406=>"001000000",
  6407=>"010000000",
  6408=>"111011001",
  6409=>"111010011",
  6410=>"111101001",
  6411=>"010100110",
  6412=>"110110111",
  6413=>"000000011",
  6414=>"010010111",
  6415=>"111111000",
  6416=>"000111111",
  6417=>"000111111",
  6418=>"011011000",
  6419=>"111111011",
  6420=>"111001001",
  6421=>"100100111",
  6422=>"000011011",
  6423=>"000010000",
  6424=>"010001111",
  6425=>"000100100",
  6426=>"111111110",
  6427=>"000000000",
  6428=>"111110000",
  6429=>"111000000",
  6430=>"000111111",
  6431=>"111111111",
  6432=>"000100100",
  6433=>"000100111",
  6434=>"000111110",
  6435=>"111111111",
  6436=>"111000000",
  6437=>"001001111",
  6438=>"111101100",
  6439=>"100000000",
  6440=>"111111111",
  6441=>"000011111",
  6442=>"111110000",
  6443=>"000000101",
  6444=>"111111111",
  6445=>"011001001",
  6446=>"000111000",
  6447=>"100101000",
  6448=>"000100100",
  6449=>"111111000",
  6450=>"000111111",
  6451=>"001101111",
  6452=>"110101000",
  6453=>"111111111",
  6454=>"000011111",
  6455=>"111101111",
  6456=>"000000000",
  6457=>"000000000",
  6458=>"000000000",
  6459=>"111001000",
  6460=>"000110111",
  6461=>"000110110",
  6462=>"000111000",
  6463=>"111000001",
  6464=>"111111100",
  6465=>"000000111",
  6466=>"111111000",
  6467=>"111001000",
  6468=>"000111001",
  6469=>"111001011",
  6470=>"000000000",
  6471=>"111110110",
  6472=>"111001111",
  6473=>"100000000",
  6474=>"001111111",
  6475=>"111100110",
  6476=>"111000000",
  6477=>"000110111",
  6478=>"111000000",
  6479=>"011001001",
  6480=>"000000001",
  6481=>"100000000",
  6482=>"111011111",
  6483=>"000000000",
  6484=>"111111011",
  6485=>"111010010",
  6486=>"111000111",
  6487=>"000111111",
  6488=>"111111111",
  6489=>"000111000",
  6490=>"111100000",
  6491=>"000000110",
  6492=>"111001000",
  6493=>"001100110",
  6494=>"000000000",
  6495=>"000000011",
  6496=>"000111111",
  6497=>"000000111",
  6498=>"100111111",
  6499=>"100111111",
  6500=>"000110110",
  6501=>"011011000",
  6502=>"000101111",
  6503=>"000100000",
  6504=>"010011000",
  6505=>"110111111",
  6506=>"111111000",
  6507=>"111110111",
  6508=>"011001001",
  6509=>"111011000",
  6510=>"100000000",
  6511=>"000000111",
  6512=>"110000000",
  6513=>"111100000",
  6514=>"000000000",
  6515=>"000011111",
  6516=>"111100100",
  6517=>"000000100",
  6518=>"100000000",
  6519=>"000111111",
  6520=>"110100000",
  6521=>"000110111",
  6522=>"011111111",
  6523=>"000000000",
  6524=>"000000001",
  6525=>"001001111",
  6526=>"000100111",
  6527=>"000000111",
  6528=>"111011011",
  6529=>"000000110",
  6530=>"000000000",
  6531=>"100111111",
  6532=>"010000111",
  6533=>"111111100",
  6534=>"000110100",
  6535=>"101100000",
  6536=>"111110000",
  6537=>"010000100",
  6538=>"111110000",
  6539=>"100101000",
  6540=>"010000111",
  6541=>"000000111",
  6542=>"000000100",
  6543=>"000111111",
  6544=>"000011111",
  6545=>"100000000",
  6546=>"000000000",
  6547=>"000011011",
  6548=>"100000000",
  6549=>"000000000",
  6550=>"111111111",
  6551=>"110010010",
  6552=>"000011111",
  6553=>"000011000",
  6554=>"000110000",
  6555=>"000000000",
  6556=>"111111101",
  6557=>"011010000",
  6558=>"111111001",
  6559=>"000001001",
  6560=>"111111000",
  6561=>"111110100",
  6562=>"000000000",
  6563=>"000000000",
  6564=>"000111111",
  6565=>"000000000",
  6566=>"000101000",
  6567=>"011001000",
  6568=>"000000000",
  6569=>"111111110",
  6570=>"111111100",
  6571=>"000000111",
  6572=>"100000000",
  6573=>"110111101",
  6574=>"111000100",
  6575=>"111011000",
  6576=>"000000111",
  6577=>"100100110",
  6578=>"000000001",
  6579=>"111011010",
  6580=>"000000000",
  6581=>"000111111",
  6582=>"000111000",
  6583=>"111111111",
  6584=>"000000000",
  6585=>"111011001",
  6586=>"110000000",
  6587=>"111111001",
  6588=>"000011001",
  6589=>"000000000",
  6590=>"000010111",
  6591=>"000011110",
  6592=>"001011010",
  6593=>"111111111",
  6594=>"000000111",
  6595=>"000000001",
  6596=>"111011111",
  6597=>"111111111",
  6598=>"111000001",
  6599=>"000000000",
  6600=>"111000000",
  6601=>"000000101",
  6602=>"100000000",
  6603=>"000000000",
  6604=>"000000010",
  6605=>"000000000",
  6606=>"000000000",
  6607=>"111111111",
  6608=>"111110000",
  6609=>"000000000",
  6610=>"010000111",
  6611=>"111101100",
  6612=>"000000000",
  6613=>"111111111",
  6614=>"000011111",
  6615=>"111111111",
  6616=>"000111111",
  6617=>"000000011",
  6618=>"111111111",
  6619=>"000000100",
  6620=>"000011111",
  6621=>"110110111",
  6622=>"000000000",
  6623=>"000001001",
  6624=>"110110111",
  6625=>"111111000",
  6626=>"000000000",
  6627=>"000000010",
  6628=>"111111111",
  6629=>"000000000",
  6630=>"010111111",
  6631=>"110110111",
  6632=>"101111010",
  6633=>"000000000",
  6634=>"111111111",
  6635=>"110000000",
  6636=>"001001000",
  6637=>"101000000",
  6638=>"101101000",
  6639=>"000000000",
  6640=>"000111111",
  6641=>"111100000",
  6642=>"111011000",
  6643=>"000011000",
  6644=>"011010110",
  6645=>"100110011",
  6646=>"000010111",
  6647=>"110111011",
  6648=>"111111001",
  6649=>"000111100",
  6650=>"000000000",
  6651=>"110111011",
  6652=>"111000000",
  6653=>"111111000",
  6654=>"011000000",
  6655=>"000000000",
  6656=>"000100100",
  6657=>"000000000",
  6658=>"000000000",
  6659=>"111111110",
  6660=>"111100100",
  6661=>"111111000",
  6662=>"100100110",
  6663=>"000000100",
  6664=>"110111111",
  6665=>"111111111",
  6666=>"100000100",
  6667=>"111111000",
  6668=>"001111110",
  6669=>"000100111",
  6670=>"000001000",
  6671=>"111111111",
  6672=>"000101100",
  6673=>"110000000",
  6674=>"111001100",
  6675=>"000000000",
  6676=>"101111111",
  6677=>"000000000",
  6678=>"111110110",
  6679=>"111110110",
  6680=>"000000000",
  6681=>"100100111",
  6682=>"000000000",
  6683=>"000011011",
  6684=>"001000001",
  6685=>"000000000",
  6686=>"111111111",
  6687=>"000010111",
  6688=>"100100000",
  6689=>"000111111",
  6690=>"111111110",
  6691=>"101111111",
  6692=>"000001001",
  6693=>"111000000",
  6694=>"111000000",
  6695=>"000010111",
  6696=>"111111111",
  6697=>"000000000",
  6698=>"100000111",
  6699=>"000000000",
  6700=>"000000111",
  6701=>"000000000",
  6702=>"000111111",
  6703=>"111111101",
  6704=>"000100000",
  6705=>"111111111",
  6706=>"111011010",
  6707=>"000000000",
  6708=>"111111101",
  6709=>"111001000",
  6710=>"111111011",
  6711=>"101101000",
  6712=>"000010010",
  6713=>"000000000",
  6714=>"111111111",
  6715=>"001000001",
  6716=>"000010111",
  6717=>"000000101",
  6718=>"111111001",
  6719=>"000000000",
  6720=>"111111011",
  6721=>"111111111",
  6722=>"000000001",
  6723=>"000010111",
  6724=>"111011000",
  6725=>"000010000",
  6726=>"101000000",
  6727=>"110111111",
  6728=>"001001000",
  6729=>"111001000",
  6730=>"010111111",
  6731=>"111111111",
  6732=>"111111111",
  6733=>"110110000",
  6734=>"000000000",
  6735=>"001111111",
  6736=>"000000000",
  6737=>"000000101",
  6738=>"110111101",
  6739=>"000000000",
  6740=>"000000000",
  6741=>"011111111",
  6742=>"000000111",
  6743=>"110000000",
  6744=>"111111111",
  6745=>"111001001",
  6746=>"010010000",
  6747=>"100100000",
  6748=>"000000000",
  6749=>"111110110",
  6750=>"000010111",
  6751=>"111111011",
  6752=>"000000000",
  6753=>"101000000",
  6754=>"001001111",
  6755=>"000000100",
  6756=>"000100110",
  6757=>"111111000",
  6758=>"111000111",
  6759=>"000000000",
  6760=>"000000000",
  6761=>"111111000",
  6762=>"000000100",
  6763=>"001000000",
  6764=>"110110100",
  6765=>"000000110",
  6766=>"111111011",
  6767=>"111010110",
  6768=>"000000000",
  6769=>"111111101",
  6770=>"101111111",
  6771=>"000000101",
  6772=>"000000110",
  6773=>"110100000",
  6774=>"111110000",
  6775=>"111111000",
  6776=>"011001000",
  6777=>"111111111",
  6778=>"100000100",
  6779=>"000001000",
  6780=>"100010110",
  6781=>"111111111",
  6782=>"111111111",
  6783=>"000000000",
  6784=>"000000000",
  6785=>"111111111",
  6786=>"000000000",
  6787=>"001000001",
  6788=>"000000110",
  6789=>"000000111",
  6790=>"101100000",
  6791=>"111011011",
  6792=>"111111111",
  6793=>"010111111",
  6794=>"000000000",
  6795=>"111111111",
  6796=>"000011011",
  6797=>"101000110",
  6798=>"111111111",
  6799=>"000110110",
  6800=>"000000000",
  6801=>"111001001",
  6802=>"111111111",
  6803=>"010111111",
  6804=>"000000000",
  6805=>"111110110",
  6806=>"000000110",
  6807=>"111111000",
  6808=>"000000000",
  6809=>"111111111",
  6810=>"111111111",
  6811=>"111111000",
  6812=>"000000000",
  6813=>"100110100",
  6814=>"110100000",
  6815=>"000000000",
  6816=>"000000111",
  6817=>"111111101",
  6818=>"000000000",
  6819=>"111011010",
  6820=>"111111111",
  6821=>"000000001",
  6822=>"000000000",
  6823=>"111011000",
  6824=>"111111111",
  6825=>"000000000",
  6826=>"000000000",
  6827=>"000100111",
  6828=>"000000101",
  6829=>"101110110",
  6830=>"111110110",
  6831=>"111111111",
  6832=>"000000000",
  6833=>"111001011",
  6834=>"000000010",
  6835=>"000000000",
  6836=>"000101111",
  6837=>"100000000",
  6838=>"111111011",
  6839=>"000001000",
  6840=>"101011001",
  6841=>"111111011",
  6842=>"111111111",
  6843=>"000000000",
  6844=>"000000000",
  6845=>"000000000",
  6846=>"111111111",
  6847=>"111111000",
  6848=>"100100110",
  6849=>"000000000",
  6850=>"001000000",
  6851=>"111111111",
  6852=>"110000000",
  6853=>"111111111",
  6854=>"000000100",
  6855=>"111111111",
  6856=>"010010010",
  6857=>"000000110",
  6858=>"111111111",
  6859=>"111111111",
  6860=>"111111011",
  6861=>"111000000",
  6862=>"000000000",
  6863=>"111110100",
  6864=>"000000101",
  6865=>"111111011",
  6866=>"000000000",
  6867=>"000000000",
  6868=>"000100011",
  6869=>"011111111",
  6870=>"000000000",
  6871=>"111111011",
  6872=>"000011000",
  6873=>"000100111",
  6874=>"000000111",
  6875=>"111111111",
  6876=>"101000000",
  6877=>"111001001",
  6878=>"000000000",
  6879=>"100100100",
  6880=>"000000000",
  6881=>"011111110",
  6882=>"111111111",
  6883=>"000111111",
  6884=>"111110110",
  6885=>"011000000",
  6886=>"110110111",
  6887=>"110000000",
  6888=>"000111001",
  6889=>"000000110",
  6890=>"000010110",
  6891=>"000000000",
  6892=>"111111111",
  6893=>"011111111",
  6894=>"000000101",
  6895=>"111111000",
  6896=>"001001111",
  6897=>"111111111",
  6898=>"111000000",
  6899=>"001000000",
  6900=>"000111111",
  6901=>"100110100",
  6902=>"111111011",
  6903=>"101111111",
  6904=>"000001011",
  6905=>"000000100",
  6906=>"000000000",
  6907=>"011001000",
  6908=>"110100100",
  6909=>"000010011",
  6910=>"000110111",
  6911=>"110111011",
  6912=>"000000100",
  6913=>"011001001",
  6914=>"000000000",
  6915=>"111101111",
  6916=>"000101111",
  6917=>"101000000",
  6918=>"000100100",
  6919=>"000101001",
  6920=>"000000000",
  6921=>"111111011",
  6922=>"001000111",
  6923=>"000101001",
  6924=>"111111111",
  6925=>"000000011",
  6926=>"111111111",
  6927=>"111011011",
  6928=>"111000000",
  6929=>"000000000",
  6930=>"010110111",
  6931=>"110000000",
  6932=>"101011000",
  6933=>"000111111",
  6934=>"000000000",
  6935=>"000000000",
  6936=>"000000110",
  6937=>"111111100",
  6938=>"111111000",
  6939=>"100111110",
  6940=>"000100100",
  6941=>"000000000",
  6942=>"111111011",
  6943=>"111111111",
  6944=>"011001111",
  6945=>"001000000",
  6946=>"000111110",
  6947=>"101111110",
  6948=>"000000000",
  6949=>"101000000",
  6950=>"001001001",
  6951=>"111001000",
  6952=>"000000111",
  6953=>"111111111",
  6954=>"111101111",
  6955=>"100000001",
  6956=>"100111111",
  6957=>"001001011",
  6958=>"000000000",
  6959=>"000000011",
  6960=>"000000000",
  6961=>"000000001",
  6962=>"111111110",
  6963=>"011000000",
  6964=>"000001001",
  6965=>"111101110",
  6966=>"000000000",
  6967=>"000000000",
  6968=>"000000000",
  6969=>"000010000",
  6970=>"111111111",
  6971=>"001111111",
  6972=>"000000000",
  6973=>"000000000",
  6974=>"110111111",
  6975=>"111111100",
  6976=>"100101111",
  6977=>"000000010",
  6978=>"000000001",
  6979=>"110110011",
  6980=>"001000000",
  6981=>"111111111",
  6982=>"000001000",
  6983=>"111111011",
  6984=>"000011111",
  6985=>"000000000",
  6986=>"000000000",
  6987=>"000000011",
  6988=>"111110110",
  6989=>"100011001",
  6990=>"000000000",
  6991=>"111110100",
  6992=>"100000000",
  6993=>"111001111",
  6994=>"111110111",
  6995=>"000111111",
  6996=>"111111111",
  6997=>"000000001",
  6998=>"110110011",
  6999=>"111111111",
  7000=>"100100111",
  7001=>"011011011",
  7002=>"000111111",
  7003=>"000000000",
  7004=>"100110100",
  7005=>"111111111",
  7006=>"000000000",
  7007=>"000000000",
  7008=>"111111000",
  7009=>"100100111",
  7010=>"000000000",
  7011=>"000000010",
  7012=>"001000000",
  7013=>"111011111",
  7014=>"111111111",
  7015=>"110100011",
  7016=>"001000000",
  7017=>"110111011",
  7018=>"000000000",
  7019=>"111000010",
  7020=>"000000110",
  7021=>"000000000",
  7022=>"111111111",
  7023=>"000010101",
  7024=>"000000000",
  7025=>"100110110",
  7026=>"100000110",
  7027=>"000000000",
  7028=>"111111001",
  7029=>"111011000",
  7030=>"111111000",
  7031=>"001011011",
  7032=>"111111111",
  7033=>"001001111",
  7034=>"111111111",
  7035=>"110110000",
  7036=>"000000110",
  7037=>"000000000",
  7038=>"110000000",
  7039=>"100111110",
  7040=>"111111111",
  7041=>"111111111",
  7042=>"110110000",
  7043=>"100101110",
  7044=>"000100000",
  7045=>"001111100",
  7046=>"001000110",
  7047=>"111000111",
  7048=>"000000100",
  7049=>"100100001",
  7050=>"000000000",
  7051=>"111111111",
  7052=>"111010110",
  7053=>"001000001",
  7054=>"100000000",
  7055=>"000000000",
  7056=>"000111011",
  7057=>"000100100",
  7058=>"101011000",
  7059=>"001100100",
  7060=>"001001011",
  7061=>"111010000",
  7062=>"000000000",
  7063=>"001000101",
  7064=>"000000110",
  7065=>"111110000",
  7066=>"100111111",
  7067=>"000000000",
  7068=>"000000000",
  7069=>"100000000",
  7070=>"110110111",
  7071=>"111111111",
  7072=>"100110110",
  7073=>"011011000",
  7074=>"111101111",
  7075=>"000000000",
  7076=>"000000111",
  7077=>"110110100",
  7078=>"111111001",
  7079=>"100100000",
  7080=>"111000000",
  7081=>"000000001",
  7082=>"111000000",
  7083=>"111111111",
  7084=>"111111111",
  7085=>"000000011",
  7086=>"001111001",
  7087=>"000000000",
  7088=>"111111101",
  7089=>"111111111",
  7090=>"001001001",
  7091=>"111111111",
  7092=>"111111111",
  7093=>"001111111",
  7094=>"000101110",
  7095=>"000000100",
  7096=>"000000010",
  7097=>"111111111",
  7098=>"000000000",
  7099=>"111100110",
  7100=>"000000000",
  7101=>"111111001",
  7102=>"000000111",
  7103=>"111111011",
  7104=>"111111111",
  7105=>"110110000",
  7106=>"111111011",
  7107=>"111111111",
  7108=>"000000000",
  7109=>"100001001",
  7110=>"110110110",
  7111=>"000000000",
  7112=>"001001000",
  7113=>"000110110",
  7114=>"100000000",
  7115=>"111111111",
  7116=>"001001011",
  7117=>"000000000",
  7118=>"111111000",
  7119=>"010010000",
  7120=>"111110010",
  7121=>"001101011",
  7122=>"110110110",
  7123=>"011111111",
  7124=>"111111111",
  7125=>"111111111",
  7126=>"010110111",
  7127=>"010000000",
  7128=>"000000100",
  7129=>"111000000",
  7130=>"110010010",
  7131=>"000000000",
  7132=>"001000000",
  7133=>"111111000",
  7134=>"000000000",
  7135=>"010011111",
  7136=>"000000000",
  7137=>"111111111",
  7138=>"001000111",
  7139=>"000000000",
  7140=>"110110111",
  7141=>"100101111",
  7142=>"111011000",
  7143=>"000000000",
  7144=>"111011111",
  7145=>"110100000",
  7146=>"000000000",
  7147=>"000111111",
  7148=>"101001001",
  7149=>"011110110",
  7150=>"001111001",
  7151=>"000001001",
  7152=>"111111111",
  7153=>"111111111",
  7154=>"011011011",
  7155=>"011011001",
  7156=>"111111111",
  7157=>"000000000",
  7158=>"110010000",
  7159=>"110111111",
  7160=>"111111000",
  7161=>"000000000",
  7162=>"000000000",
  7163=>"110111111",
  7164=>"111111100",
  7165=>"101100000",
  7166=>"111111000",
  7167=>"000000000",
  7168=>"100100111",
  7169=>"010110000",
  7170=>"000000111",
  7171=>"000010110",
  7172=>"000000000",
  7173=>"111000000",
  7174=>"010010000",
  7175=>"111111111",
  7176=>"111010000",
  7177=>"000000000",
  7178=>"000000001",
  7179=>"011111110",
  7180=>"000000000",
  7181=>"000000000",
  7182=>"000000000",
  7183=>"000110111",
  7184=>"010000000",
  7185=>"000110110",
  7186=>"001001111",
  7187=>"000000000",
  7188=>"000000000",
  7189=>"111111000",
  7190=>"000000000",
  7191=>"111001001",
  7192=>"101100000",
  7193=>"000000000",
  7194=>"010000000",
  7195=>"100001000",
  7196=>"111111111",
  7197=>"000000000",
  7198=>"111100101",
  7199=>"000000000",
  7200=>"000000000",
  7201=>"100100000",
  7202=>"111000110",
  7203=>"000000110",
  7204=>"000000100",
  7205=>"111111111",
  7206=>"101101000",
  7207=>"100000000",
  7208=>"111111101",
  7209=>"111111111",
  7210=>"110000110",
  7211=>"000011011",
  7212=>"000000010",
  7213=>"011011001",
  7214=>"111111110",
  7215=>"110000000",
  7216=>"001000101",
  7217=>"111101000",
  7218=>"001001111",
  7219=>"001000000",
  7220=>"000010111",
  7221=>"001111111",
  7222=>"000100111",
  7223=>"100000000",
  7224=>"111111111",
  7225=>"000000000",
  7226=>"010111110",
  7227=>"010010000",
  7228=>"000000000",
  7229=>"001111111",
  7230=>"000000100",
  7231=>"011001000",
  7232=>"001001001",
  7233=>"000101111",
  7234=>"111111111",
  7235=>"011111000",
  7236=>"011001000",
  7237=>"111011000",
  7238=>"000000000",
  7239=>"000111111",
  7240=>"111011001",
  7241=>"000000000",
  7242=>"010011111",
  7243=>"000000000",
  7244=>"000000000",
  7245=>"000000000",
  7246=>"111100111",
  7247=>"000010011",
  7248=>"000000000",
  7249=>"111111000",
  7250=>"111100000",
  7251=>"001001111",
  7252=>"000000010",
  7253=>"011011101",
  7254=>"100111111",
  7255=>"101111111",
  7256=>"000000100",
  7257=>"000101111",
  7258=>"000011110",
  7259=>"000000000",
  7260=>"100000000",
  7261=>"111001011",
  7262=>"100110001",
  7263=>"000000000",
  7264=>"101100000",
  7265=>"111111111",
  7266=>"111111111",
  7267=>"000010111",
  7268=>"111101000",
  7269=>"000000000",
  7270=>"000110111",
  7271=>"110000111",
  7272=>"100110011",
  7273=>"010000001",
  7274=>"000000000",
  7275=>"100111111",
  7276=>"111011011",
  7277=>"100000000",
  7278=>"000000000",
  7279=>"000000111",
  7280=>"000000000",
  7281=>"000000000",
  7282=>"000100111",
  7283=>"111100100",
  7284=>"001000001",
  7285=>"110110110",
  7286=>"111111011",
  7287=>"111111111",
  7288=>"010000000",
  7289=>"000000000",
  7290=>"100110000",
  7291=>"000000000",
  7292=>"011010010",
  7293=>"011111111",
  7294=>"110100000",
  7295=>"111111110",
  7296=>"111000000",
  7297=>"111111111",
  7298=>"000000100",
  7299=>"111111111",
  7300=>"111010100",
  7301=>"111000000",
  7302=>"000001111",
  7303=>"000000000",
  7304=>"000010110",
  7305=>"100111000",
  7306=>"000000000",
  7307=>"001111100",
  7308=>"111111111",
  7309=>"111111111",
  7310=>"000000100",
  7311=>"011010111",
  7312=>"000010111",
  7313=>"111111111",
  7314=>"000010111",
  7315=>"111000000",
  7316=>"000000000",
  7317=>"000000000",
  7318=>"111001111",
  7319=>"000101000",
  7320=>"000000000",
  7321=>"111111111",
  7322=>"111011111",
  7323=>"000000000",
  7324=>"000000000",
  7325=>"110110000",
  7326=>"000101111",
  7327=>"000000000",
  7328=>"001001000",
  7329=>"000101010",
  7330=>"111111001",
  7331=>"111000000",
  7332=>"000110110",
  7333=>"001000110",
  7334=>"010010010",
  7335=>"111111111",
  7336=>"000110000",
  7337=>"101000111",
  7338=>"000000001",
  7339=>"000000100",
  7340=>"000100111",
  7341=>"001001100",
  7342=>"111111111",
  7343=>"001011000",
  7344=>"000000000",
  7345=>"011001000",
  7346=>"000000010",
  7347=>"111001000",
  7348=>"101111011",
  7349=>"011011001",
  7350=>"111110000",
  7351=>"000000000",
  7352=>"000110110",
  7353=>"110110100",
  7354=>"000100111",
  7355=>"000111100",
  7356=>"000000000",
  7357=>"111111110",
  7358=>"111100100",
  7359=>"111110000",
  7360=>"111111100",
  7361=>"110000000",
  7362=>"000000000",
  7363=>"111101000",
  7364=>"110000000",
  7365=>"000011010",
  7366=>"111111111",
  7367=>"111100000",
  7368=>"111111111",
  7369=>"100000000",
  7370=>"000100110",
  7371=>"111111110",
  7372=>"000101111",
  7373=>"111111011",
  7374=>"001111011",
  7375=>"000000001",
  7376=>"011000000",
  7377=>"111100000",
  7378=>"100000000",
  7379=>"110000000",
  7380=>"000010111",
  7381=>"000111111",
  7382=>"011000000",
  7383=>"111111111",
  7384=>"101111111",
  7385=>"111111111",
  7386=>"101001100",
  7387=>"000111000",
  7388=>"011011000",
  7389=>"000111110",
  7390=>"000000000",
  7391=>"111101001",
  7392=>"000000000",
  7393=>"111100111",
  7394=>"000100000",
  7395=>"011011000",
  7396=>"011000110",
  7397=>"001000000",
  7398=>"000010111",
  7399=>"111100110",
  7400=>"000000000",
  7401=>"111111111",
  7402=>"101001000",
  7403=>"000000000",
  7404=>"111000000",
  7405=>"001000000",
  7406=>"000000000",
  7407=>"000001111",
  7408=>"111011011",
  7409=>"011111111",
  7410=>"000000000",
  7411=>"000001011",
  7412=>"100010000",
  7413=>"000000111",
  7414=>"111111100",
  7415=>"000000000",
  7416=>"111111110",
  7417=>"111111111",
  7418=>"000001111",
  7419=>"000000000",
  7420=>"111100100",
  7421=>"111010000",
  7422=>"101111110",
  7423=>"100000000",
  7424=>"000111111",
  7425=>"110110110",
  7426=>"111111011",
  7427=>"100111000",
  7428=>"111111111",
  7429=>"000010110",
  7430=>"000000000",
  7431=>"000001101",
  7432=>"110001111",
  7433=>"011111111",
  7434=>"000110000",
  7435=>"000000000",
  7436=>"110000010",
  7437=>"011111111",
  7438=>"001100001",
  7439=>"110110111",
  7440=>"001011011",
  7441=>"000000000",
  7442=>"111111111",
  7443=>"000010000",
  7444=>"000000110",
  7445=>"000000111",
  7446=>"110110110",
  7447=>"110110110",
  7448=>"111111111",
  7449=>"111111111",
  7450=>"000110110",
  7451=>"100111111",
  7452=>"111111111",
  7453=>"000000000",
  7454=>"111111111",
  7455=>"000111001",
  7456=>"011101001",
  7457=>"000000000",
  7458=>"000000011",
  7459=>"000001001",
  7460=>"111111111",
  7461=>"000000000",
  7462=>"000011011",
  7463=>"000000000",
  7464=>"100111111",
  7465=>"000000000",
  7466=>"000000001",
  7467=>"010000001",
  7468=>"000000000",
  7469=>"111111111",
  7470=>"000000000",
  7471=>"100010111",
  7472=>"101011001",
  7473=>"001011111",
  7474=>"101000000",
  7475=>"111100000",
  7476=>"111111111",
  7477=>"000010110",
  7478=>"000100101",
  7479=>"111111000",
  7480=>"011111110",
  7481=>"000100000",
  7482=>"111111111",
  7483=>"110000000",
  7484=>"010110110",
  7485=>"001111001",
  7486=>"111111000",
  7487=>"111111111",
  7488=>"000000000",
  7489=>"010111011",
  7490=>"000100100",
  7491=>"111010010",
  7492=>"000000000",
  7493=>"111111111",
  7494=>"111111111",
  7495=>"000000000",
  7496=>"110110000",
  7497=>"000000000",
  7498=>"000101111",
  7499=>"111011111",
  7500=>"000000010",
  7501=>"110000001",
  7502=>"001000000",
  7503=>"111111101",
  7504=>"001011111",
  7505=>"000000000",
  7506=>"010010110",
  7507=>"111000001",
  7508=>"000000001",
  7509=>"010000000",
  7510=>"000011111",
  7511=>"011111101",
  7512=>"111001000",
  7513=>"000000000",
  7514=>"000000011",
  7515=>"000000111",
  7516=>"111110001",
  7517=>"100110110",
  7518=>"000110011",
  7519=>"100100111",
  7520=>"000000000",
  7521=>"111111111",
  7522=>"010011000",
  7523=>"000000110",
  7524=>"000000000",
  7525=>"000000000",
  7526=>"000000000",
  7527=>"111111011",
  7528=>"000000110",
  7529=>"100100000",
  7530=>"110111000",
  7531=>"111111010",
  7532=>"111001000",
  7533=>"000111110",
  7534=>"111111111",
  7535=>"000111011",
  7536=>"111111111",
  7537=>"111101111",
  7538=>"111111001",
  7539=>"111001001",
  7540=>"111111111",
  7541=>"111111111",
  7542=>"000000000",
  7543=>"111111111",
  7544=>"111111111",
  7545=>"111111111",
  7546=>"110110111",
  7547=>"001001001",
  7548=>"100110010",
  7549=>"000000000",
  7550=>"111111001",
  7551=>"111111000",
  7552=>"111111110",
  7553=>"111110000",
  7554=>"111110000",
  7555=>"000000000",
  7556=>"011000000",
  7557=>"000000000",
  7558=>"101000000",
  7559=>"110111000",
  7560=>"111111111",
  7561=>"001001011",
  7562=>"111110100",
  7563=>"000000100",
  7564=>"000000000",
  7565=>"000001101",
  7566=>"100000010",
  7567=>"111111111",
  7568=>"001111111",
  7569=>"110001000",
  7570=>"111111111",
  7571=>"011111011",
  7572=>"111110110",
  7573=>"001110000",
  7574=>"001010111",
  7575=>"000100111",
  7576=>"111110000",
  7577=>"111010010",
  7578=>"111110111",
  7579=>"111111100",
  7580=>"111111111",
  7581=>"000000011",
  7582=>"000000111",
  7583=>"000000100",
  7584=>"111011000",
  7585=>"111111111",
  7586=>"000110110",
  7587=>"011111111",
  7588=>"111111100",
  7589=>"111011001",
  7590=>"000100110",
  7591=>"011000110",
  7592=>"000000000",
  7593=>"001000111",
  7594=>"001000000",
  7595=>"000111111",
  7596=>"011000000",
  7597=>"000000000",
  7598=>"000000111",
  7599=>"000000000",
  7600=>"000000001",
  7601=>"000110111",
  7602=>"000001111",
  7603=>"000000101",
  7604=>"100000000",
  7605=>"011000000",
  7606=>"111111101",
  7607=>"001000000",
  7608=>"000111000",
  7609=>"001111000",
  7610=>"000001111",
  7611=>"001011010",
  7612=>"111001000",
  7613=>"111111001",
  7614=>"110111110",
  7615=>"000011011",
  7616=>"111110111",
  7617=>"011011010",
  7618=>"000000000",
  7619=>"110011000",
  7620=>"000111001",
  7621=>"011011001",
  7622=>"000111111",
  7623=>"000111111",
  7624=>"000001111",
  7625=>"000111111",
  7626=>"000000000",
  7627=>"111110000",
  7628=>"000000000",
  7629=>"111111111",
  7630=>"000000000",
  7631=>"000000011",
  7632=>"001001111",
  7633=>"101111001",
  7634=>"000000000",
  7635=>"111110010",
  7636=>"000100100",
  7637=>"000000000",
  7638=>"000000111",
  7639=>"000001001",
  7640=>"000000000",
  7641=>"000000100",
  7642=>"001111111",
  7643=>"011000101",
  7644=>"101011001",
  7645=>"000000000",
  7646=>"100000000",
  7647=>"000000001",
  7648=>"111111111",
  7649=>"111111000",
  7650=>"011111000",
  7651=>"000000000",
  7652=>"000011000",
  7653=>"000000000",
  7654=>"000000010",
  7655=>"111001010",
  7656=>"111100000",
  7657=>"000000000",
  7658=>"111100100",
  7659=>"000001011",
  7660=>"111111000",
  7661=>"000000001",
  7662=>"111111111",
  7663=>"100010000",
  7664=>"000100111",
  7665=>"000000111",
  7666=>"111111001",
  7667=>"111101101",
  7668=>"000111111",
  7669=>"001010011",
  7670=>"000000000",
  7671=>"011111111",
  7672=>"000000000",
  7673=>"101101111",
  7674=>"001000000",
  7675=>"111111111",
  7676=>"110111111",
  7677=>"111111111",
  7678=>"000111111",
  7679=>"111111111",
  7680=>"001101000",
  7681=>"111111100",
  7682=>"111111001",
  7683=>"100100000",
  7684=>"111110111",
  7685=>"000000000",
  7686=>"100000100",
  7687=>"111111111",
  7688=>"111111111",
  7689=>"111111111",
  7690=>"001000000",
  7691=>"101100100",
  7692=>"111111111",
  7693=>"000011011",
  7694=>"000000000",
  7695=>"000000000",
  7696=>"111111001",
  7697=>"010110000",
  7698=>"111101111",
  7699=>"011011011",
  7700=>"000011111",
  7701=>"101101001",
  7702=>"111011100",
  7703=>"111111110",
  7704=>"000000000",
  7705=>"110100000",
  7706=>"000000111",
  7707=>"110111011",
  7708=>"111111111",
  7709=>"000000000",
  7710=>"111000000",
  7711=>"111111111",
  7712=>"000000111",
  7713=>"111111100",
  7714=>"000000101",
  7715=>"000000000",
  7716=>"111110100",
  7717=>"000001001",
  7718=>"111010111",
  7719=>"111111100",
  7720=>"111111111",
  7721=>"000000000",
  7722=>"000000000",
  7723=>"110100000",
  7724=>"000000000",
  7725=>"000000011",
  7726=>"111111101",
  7727=>"111100000",
  7728=>"001000000",
  7729=>"111111111",
  7730=>"101001000",
  7731=>"111111111",
  7732=>"111011001",
  7733=>"111001001",
  7734=>"000000000",
  7735=>"111111111",
  7736=>"100100111",
  7737=>"000000000",
  7738=>"000000000",
  7739=>"010111111",
  7740=>"000001011",
  7741=>"000000000",
  7742=>"111111111",
  7743=>"000000000",
  7744=>"010100111",
  7745=>"000111001",
  7746=>"000000000",
  7747=>"000100100",
  7748=>"110110000",
  7749=>"001001001",
  7750=>"001001111",
  7751=>"111111111",
  7752=>"000000000",
  7753=>"000000000",
  7754=>"001001001",
  7755=>"111000011",
  7756=>"000000000",
  7757=>"000111111",
  7758=>"000000000",
  7759=>"110100111",
  7760=>"000010000",
  7761=>"011011011",
  7762=>"000100110",
  7763=>"111111111",
  7764=>"111111111",
  7765=>"111111000",
  7766=>"000100100",
  7767=>"111111111",
  7768=>"000000000",
  7769=>"001000000",
  7770=>"001000000",
  7771=>"111011001",
  7772=>"110111111",
  7773=>"001011111",
  7774=>"010010000",
  7775=>"111110111",
  7776=>"111111001",
  7777=>"000000000",
  7778=>"111101100",
  7779=>"111111111",
  7780=>"100110000",
  7781=>"000000000",
  7782=>"000000100",
  7783=>"111000001",
  7784=>"110010111",
  7785=>"100000111",
  7786=>"111111110",
  7787=>"011001000",
  7788=>"111111111",
  7789=>"000000111",
  7790=>"111111011",
  7791=>"011000000",
  7792=>"101111111",
  7793=>"111111111",
  7794=>"011000001",
  7795=>"000000010",
  7796=>"111111111",
  7797=>"011111000",
  7798=>"000000000",
  7799=>"001000000",
  7800=>"000000100",
  7801=>"000001000",
  7802=>"110010011",
  7803=>"000000000",
  7804=>"111111111",
  7805=>"111111110",
  7806=>"110111110",
  7807=>"101101001",
  7808=>"000000000",
  7809=>"111110111",
  7810=>"000000000",
  7811=>"100111111",
  7812=>"000111111",
  7813=>"111011111",
  7814=>"111111001",
  7815=>"111000001",
  7816=>"100100111",
  7817=>"000111100",
  7818=>"000000111",
  7819=>"000100000",
  7820=>"101111110",
  7821=>"001000001",
  7822=>"011110111",
  7823=>"111011001",
  7824=>"000000110",
  7825=>"110100111",
  7826=>"000110111",
  7827=>"111111110",
  7828=>"011000000",
  7829=>"111001000",
  7830=>"011011011",
  7831=>"111111111",
  7832=>"111100111",
  7833=>"111110110",
  7834=>"000000000",
  7835=>"000001000",
  7836=>"000000000",
  7837=>"100110000",
  7838=>"111001111",
  7839=>"000000000",
  7840=>"111001111",
  7841=>"000000000",
  7842=>"101101111",
  7843=>"011000000",
  7844=>"111111111",
  7845=>"111111111",
  7846=>"111001110",
  7847=>"011011000",
  7848=>"111111111",
  7849=>"000000100",
  7850=>"000000000",
  7851=>"000000001",
  7852=>"011111000",
  7853=>"110101011",
  7854=>"111111111",
  7855=>"101001011",
  7856=>"111000000",
  7857=>"001110000",
  7858=>"111001111",
  7859=>"000000100",
  7860=>"111111111",
  7861=>"000000000",
  7862=>"000000000",
  7863=>"000010111",
  7864=>"000000001",
  7865=>"011001000",
  7866=>"000000000",
  7867=>"110110110",
  7868=>"001001001",
  7869=>"000110110",
  7870=>"000111111",
  7871=>"100100111",
  7872=>"111111111",
  7873=>"110000111",
  7874=>"000000000",
  7875=>"000000000",
  7876=>"100100001",
  7877=>"000000000",
  7878=>"011011000",
  7879=>"000101111",
  7880=>"000011001",
  7881=>"111101101",
  7882=>"000000111",
  7883=>"111001111",
  7884=>"111111011",
  7885=>"111000000",
  7886=>"110000000",
  7887=>"111111111",
  7888=>"000000000",
  7889=>"011111011",
  7890=>"110111110",
  7891=>"000001000",
  7892=>"000101111",
  7893=>"111111111",
  7894=>"000000000",
  7895=>"000110000",
  7896=>"001001011",
  7897=>"100000000",
  7898=>"000001011",
  7899=>"011010000",
  7900=>"111111000",
  7901=>"111001001",
  7902=>"000001111",
  7903=>"000000111",
  7904=>"000111111",
  7905=>"001000000",
  7906=>"000000000",
  7907=>"000000000",
  7908=>"000010111",
  7909=>"011010111",
  7910=>"111111110",
  7911=>"100110110",
  7912=>"100100111",
  7913=>"100101111",
  7914=>"110000000",
  7915=>"111111111",
  7916=>"111111111",
  7917=>"000001000",
  7918=>"000000000",
  7919=>"111001000",
  7920=>"010100000",
  7921=>"111111111",
  7922=>"000000000",
  7923=>"100100111",
  7924=>"111111111",
  7925=>"011011011",
  7926=>"000000001",
  7927=>"111101111",
  7928=>"111111110",
  7929=>"000000000",
  7930=>"111111111",
  7931=>"000000000",
  7932=>"111111111",
  7933=>"011001000",
  7934=>"001001100",
  7935=>"000000010",
  7936=>"111110110",
  7937=>"011000000",
  7938=>"111111000",
  7939=>"111111111",
  7940=>"000010111",
  7941=>"111000000",
  7942=>"011111111",
  7943=>"100100100",
  7944=>"000000100",
  7945=>"111111111",
  7946=>"111111111",
  7947=>"100000000",
  7948=>"111001001",
  7949=>"011011001",
  7950=>"110111111",
  7951=>"000111011",
  7952=>"111111000",
  7953=>"110110111",
  7954=>"000000000",
  7955=>"110110100",
  7956=>"000000000",
  7957=>"101101011",
  7958=>"011011001",
  7959=>"111000000",
  7960=>"001000111",
  7961=>"110110110",
  7962=>"111001000",
  7963=>"000000000",
  7964=>"100000000",
  7965=>"111111111",
  7966=>"000010000",
  7967=>"110110011",
  7968=>"111111101",
  7969=>"111110110",
  7970=>"100110110",
  7971=>"000000000",
  7972=>"001001001",
  7973=>"111101000",
  7974=>"111111111",
  7975=>"000001101",
  7976=>"000000010",
  7977=>"111111111",
  7978=>"100110111",
  7979=>"000010010",
  7980=>"001001001",
  7981=>"100100100",
  7982=>"000000000",
  7983=>"000000000",
  7984=>"111111111",
  7985=>"111011001",
  7986=>"011011000",
  7987=>"001001100",
  7988=>"000000000",
  7989=>"111111101",
  7990=>"111001011",
  7991=>"111110000",
  7992=>"000000011",
  7993=>"111111111",
  7994=>"011000000",
  7995=>"111110000",
  7996=>"000000000",
  7997=>"101100100",
  7998=>"110111111",
  7999=>"000000011",
  8000=>"000000000",
  8001=>"011111000",
  8002=>"110110000",
  8003=>"110100001",
  8004=>"011111101",
  8005=>"011011111",
  8006=>"111111111",
  8007=>"100000000",
  8008=>"111011111",
  8009=>"111111011",
  8010=>"000000000",
  8011=>"000111111",
  8012=>"111111011",
  8013=>"000100000",
  8014=>"111111111",
  8015=>"001001011",
  8016=>"001001001",
  8017=>"000110111",
  8018=>"110111111",
  8019=>"110111111",
  8020=>"000000000",
  8021=>"011111111",
  8022=>"000000001",
  8023=>"111111111",
  8024=>"000101110",
  8025=>"111001001",
  8026=>"100110111",
  8027=>"000001011",
  8028=>"000010111",
  8029=>"001101111",
  8030=>"000100100",
  8031=>"000000000",
  8032=>"000000000",
  8033=>"000000000",
  8034=>"111111101",
  8035=>"011101011",
  8036=>"111110110",
  8037=>"111111111",
  8038=>"000000111",
  8039=>"111111111",
  8040=>"001001001",
  8041=>"111111110",
  8042=>"000000001",
  8043=>"000110111",
  8044=>"111111001",
  8045=>"000110110",
  8046=>"000111111",
  8047=>"000000111",
  8048=>"111111011",
  8049=>"000000000",
  8050=>"111111111",
  8051=>"100111110",
  8052=>"001000000",
  8053=>"011000000",
  8054=>"000000000",
  8055=>"110000011",
  8056=>"000100110",
  8057=>"001000001",
  8058=>"111111111",
  8059=>"011000001",
  8060=>"111111111",
  8061=>"111011111",
  8062=>"111011111",
  8063=>"111111111",
  8064=>"000000000",
  8065=>"111111101",
  8066=>"110110111",
  8067=>"111111111",
  8068=>"000000100",
  8069=>"110110110",
  8070=>"001001000",
  8071=>"000011000",
  8072=>"111011000",
  8073=>"011001000",
  8074=>"011111000",
  8075=>"011011000",
  8076=>"000000000",
  8077=>"111010010",
  8078=>"001000010",
  8079=>"000000000",
  8080=>"111111000",
  8081=>"111111000",
  8082=>"000000000",
  8083=>"111110110",
  8084=>"100111111",
  8085=>"000000000",
  8086=>"111111111",
  8087=>"111101111",
  8088=>"111110111",
  8089=>"010111011",
  8090=>"111111111",
  8091=>"000000111",
  8092=>"110100111",
  8093=>"000000000",
  8094=>"000000000",
  8095=>"000000111",
  8096=>"111000000",
  8097=>"111011011",
  8098=>"011111111",
  8099=>"000000000",
  8100=>"111001111",
  8101=>"011111111",
  8102=>"111000000",
  8103=>"000000000",
  8104=>"000000000",
  8105=>"001001111",
  8106=>"000000110",
  8107=>"111111101",
  8108=>"100001001",
  8109=>"111110110",
  8110=>"000000000",
  8111=>"000000000",
  8112=>"000000000",
  8113=>"000000000",
  8114=>"111100000",
  8115=>"001000001",
  8116=>"010111111",
  8117=>"011000000",
  8118=>"000110110",
  8119=>"110000000",
  8120=>"111000000",
  8121=>"111111101",
  8122=>"101100011",
  8123=>"100100110",
  8124=>"001001001",
  8125=>"111100100",
  8126=>"000000000",
  8127=>"001011011",
  8128=>"100110000",
  8129=>"001000000",
  8130=>"001000000",
  8131=>"000000000",
  8132=>"000000000",
  8133=>"000000100",
  8134=>"111111111",
  8135=>"000001000",
  8136=>"011000000",
  8137=>"000000100",
  8138=>"011000101",
  8139=>"000000000",
  8140=>"000000111",
  8141=>"111111111",
  8142=>"001110111",
  8143=>"000001001",
  8144=>"000000000",
  8145=>"111111111",
  8146=>"011000001",
  8147=>"111111111",
  8148=>"111111111",
  8149=>"011111000",
  8150=>"111111111",
  8151=>"110110001",
  8152=>"110000000",
  8153=>"000010000",
  8154=>"000000000",
  8155=>"000000000",
  8156=>"011000000",
  8157=>"000100100",
  8158=>"001010000",
  8159=>"110010110",
  8160=>"111101000",
  8161=>"011001000",
  8162=>"000111111",
  8163=>"000000000",
  8164=>"111111111",
  8165=>"000001101",
  8166=>"000001000",
  8167=>"000000001",
  8168=>"100000000",
  8169=>"011011000",
  8170=>"111111100",
  8171=>"000000000",
  8172=>"111101100",
  8173=>"111011011",
  8174=>"000000000",
  8175=>"010010010",
  8176=>"011000111",
  8177=>"011001001",
  8178=>"000000000",
  8179=>"011111011",
  8180=>"111111001",
  8181=>"000000000",
  8182=>"101111111",
  8183=>"000000100",
  8184=>"011011011",
  8185=>"001101111",
  8186=>"000000000",
  8187=>"001001001",
  8188=>"000011011",
  8189=>"111101101",
  8190=>"011111000",
  8191=>"000011010",
  8192=>"001001001",
  8193=>"111011011",
  8194=>"001001111",
  8195=>"101100100",
  8196=>"011011000",
  8197=>"101111000",
  8198=>"010110010",
  8199=>"111111111",
  8200=>"111111000",
  8201=>"011000000",
  8202=>"000000101",
  8203=>"000000000",
  8204=>"000000101",
  8205=>"111111101",
  8206=>"100100000",
  8207=>"111111110",
  8208=>"110111010",
  8209=>"000111111",
  8210=>"001000000",
  8211=>"110000000",
  8212=>"101001111",
  8213=>"111100100",
  8214=>"111111010",
  8215=>"110000000",
  8216=>"111111111",
  8217=>"111111000",
  8218=>"101100111",
  8219=>"101111100",
  8220=>"001000111",
  8221=>"101111000",
  8222=>"000000000",
  8223=>"101001110",
  8224=>"010000000",
  8225=>"000110111",
  8226=>"001001001",
  8227=>"000000111",
  8228=>"001000111",
  8229=>"001011111",
  8230=>"000000001",
  8231=>"000000000",
  8232=>"000000000",
  8233=>"111011111",
  8234=>"000000101",
  8235=>"111111100",
  8236=>"001001101",
  8237=>"100100000",
  8238=>"000000001",
  8239=>"000110010",
  8240=>"110111111",
  8241=>"001001110",
  8242=>"111101000",
  8243=>"000001011",
  8244=>"000000100",
  8245=>"110110000",
  8246=>"000001001",
  8247=>"000000000",
  8248=>"001000000",
  8249=>"110111101",
  8250=>"000001001",
  8251=>"000000000",
  8252=>"001000111",
  8253=>"100100100",
  8254=>"011111100",
  8255=>"110100000",
  8256=>"011001000",
  8257=>"000010000",
  8258=>"010111111",
  8259=>"111111100",
  8260=>"110110110",
  8261=>"000001000",
  8262=>"111111111",
  8263=>"111101101",
  8264=>"011111011",
  8265=>"100101111",
  8266=>"010111000",
  8267=>"111010000",
  8268=>"000000000",
  8269=>"111000101",
  8270=>"000110001",
  8271=>"111000000",
  8272=>"110100100",
  8273=>"000000000",
  8274=>"101001101",
  8275=>"100100110",
  8276=>"111111000",
  8277=>"000000000",
  8278=>"111111011",
  8279=>"010000000",
  8280=>"000000000",
  8281=>"111000100",
  8282=>"010001111",
  8283=>"010000000",
  8284=>"000001000",
  8285=>"111111110",
  8286=>"001000001",
  8287=>"000000000",
  8288=>"111110010",
  8289=>"101010000",
  8290=>"000011111",
  8291=>"000000000",
  8292=>"100000000",
  8293=>"001011111",
  8294=>"001000001",
  8295=>"000000010",
  8296=>"010111110",
  8297=>"000000010",
  8298=>"011001100",
  8299=>"010010011",
  8300=>"111110100",
  8301=>"000000001",
  8302=>"100000000",
  8303=>"111111011",
  8304=>"000000000",
  8305=>"110110100",
  8306=>"111111111",
  8307=>"000000000",
  8308=>"111011000",
  8309=>"110111000",
  8310=>"000000000",
  8311=>"111101101",
  8312=>"010111001",
  8313=>"000000000",
  8314=>"111101000",
  8315=>"000100111",
  8316=>"100110110",
  8317=>"000000101",
  8318=>"011011001",
  8319=>"100000000",
  8320=>"000001011",
  8321=>"111111001",
  8322=>"000000000",
  8323=>"111111111",
  8324=>"000000000",
  8325=>"010110000",
  8326=>"110110000",
  8327=>"000110110",
  8328=>"000000000",
  8329=>"100100111",
  8330=>"001111111",
  8331=>"001000000",
  8332=>"110111111",
  8333=>"111110111",
  8334=>"110111010",
  8335=>"000001001",
  8336=>"101000100",
  8337=>"111100000",
  8338=>"000000110",
  8339=>"001010000",
  8340=>"111011111",
  8341=>"000100111",
  8342=>"111000000",
  8343=>"001000000",
  8344=>"001000101",
  8345=>"101000001",
  8346=>"111111111",
  8347=>"011011000",
  8348=>"111010010",
  8349=>"000011000",
  8350=>"100000000",
  8351=>"000010000",
  8352=>"000011110",
  8353=>"000000000",
  8354=>"110111000",
  8355=>"010000000",
  8356=>"011011001",
  8357=>"110111001",
  8358=>"111111000",
  8359=>"000000000",
  8360=>"111111011",
  8361=>"100111111",
  8362=>"001000000",
  8363=>"111111101",
  8364=>"011001001",
  8365=>"100110000",
  8366=>"110111001",
  8367=>"100111111",
  8368=>"100001000",
  8369=>"001000000",
  8370=>"111111000",
  8371=>"110110000",
  8372=>"110110111",
  8373=>"111000000",
  8374=>"111111000",
  8375=>"010000000",
  8376=>"011111011",
  8377=>"001001111",
  8378=>"011011111",
  8379=>"111000100",
  8380=>"111111100",
  8381=>"000000000",
  8382=>"000000111",
  8383=>"001000111",
  8384=>"101000100",
  8385=>"111111001",
  8386=>"000000000",
  8387=>"000001001",
  8388=>"001111111",
  8389=>"011111111",
  8390=>"110100110",
  8391=>"001000001",
  8392=>"110110110",
  8393=>"000000000",
  8394=>"111111111",
  8395=>"000000000",
  8396=>"100001000",
  8397=>"100111101",
  8398=>"000110110",
  8399=>"000000000",
  8400=>"010100100",
  8401=>"000111111",
  8402=>"110111000",
  8403=>"001000001",
  8404=>"000111111",
  8405=>"001011010",
  8406=>"111001000",
  8407=>"110111000",
  8408=>"111111001",
  8409=>"111111111",
  8410=>"111111111",
  8411=>"110000111",
  8412=>"111110000",
  8413=>"000101100",
  8414=>"100100111",
  8415=>"000000000",
  8416=>"000000111",
  8417=>"000011111",
  8418=>"111111111",
  8419=>"111111011",
  8420=>"000110110",
  8421=>"110100000",
  8422=>"111111010",
  8423=>"111111111",
  8424=>"111110001",
  8425=>"000000000",
  8426=>"001101011",
  8427=>"101000011",
  8428=>"011111100",
  8429=>"100000111",
  8430=>"101000000",
  8431=>"110010000",
  8432=>"000111110",
  8433=>"000100100",
  8434=>"000011011",
  8435=>"000000100",
  8436=>"110000000",
  8437=>"010000000",
  8438=>"111111101",
  8439=>"000000001",
  8440=>"000000000",
  8441=>"000000000",
  8442=>"111111000",
  8443=>"111010010",
  8444=>"100100100",
  8445=>"011001001",
  8446=>"010000111",
  8447=>"100100100",
  8448=>"001000000",
  8449=>"011001001",
  8450=>"001001000",
  8451=>"100000000",
  8452=>"000011111",
  8453=>"000000111",
  8454=>"110111000",
  8455=>"111010010",
  8456=>"001000000",
  8457=>"000000100",
  8458=>"010101000",
  8459=>"111111101",
  8460=>"000000100",
  8461=>"111111010",
  8462=>"000000000",
  8463=>"000000000",
  8464=>"100100000",
  8465=>"010111111",
  8466=>"101101111",
  8467=>"000000001",
  8468=>"000000000",
  8469=>"000000000",
  8470=>"001001001",
  8471=>"000110100",
  8472=>"000000000",
  8473=>"111111111",
  8474=>"000000100",
  8475=>"111100000",
  8476=>"110110110",
  8477=>"011001000",
  8478=>"011111111",
  8479=>"111111000",
  8480=>"110100000",
  8481=>"111111111",
  8482=>"111000000",
  8483=>"000000101",
  8484=>"000000111",
  8485=>"111111111",
  8486=>"001000100",
  8487=>"100000110",
  8488=>"011111111",
  8489=>"110110000",
  8490=>"111111111",
  8491=>"111111000",
  8492=>"000000000",
  8493=>"000000000",
  8494=>"010010000",
  8495=>"100101111",
  8496=>"111111111",
  8497=>"000100100",
  8498=>"111001000",
  8499=>"110010011",
  8500=>"000000000",
  8501=>"000000000",
  8502=>"000100110",
  8503=>"010111010",
  8504=>"000000100",
  8505=>"110100110",
  8506=>"111110111",
  8507=>"001000000",
  8508=>"110110000",
  8509=>"111111000",
  8510=>"000111100",
  8511=>"000000000",
  8512=>"101001000",
  8513=>"000100000",
  8514=>"101000111",
  8515=>"100000110",
  8516=>"110010000",
  8517=>"111000100",
  8518=>"111001001",
  8519=>"101100000",
  8520=>"100100000",
  8521=>"011111110",
  8522=>"000100010",
  8523=>"100110110",
  8524=>"100100100",
  8525=>"000000000",
  8526=>"000000101",
  8527=>"000000010",
  8528=>"001000000",
  8529=>"000000011",
  8530=>"111000000",
  8531=>"000000000",
  8532=>"000000000",
  8533=>"011011011",
  8534=>"000110111",
  8535=>"100111111",
  8536=>"000000000",
  8537=>"001100100",
  8538=>"100111000",
  8539=>"111111001",
  8540=>"111010000",
  8541=>"100000000",
  8542=>"111111011",
  8543=>"101001111",
  8544=>"010111010",
  8545=>"101000000",
  8546=>"000000111",
  8547=>"111101100",
  8548=>"110110100",
  8549=>"000000000",
  8550=>"001111111",
  8551=>"111000011",
  8552=>"111111010",
  8553=>"000000000",
  8554=>"101000000",
  8555=>"010111000",
  8556=>"001001000",
  8557=>"001001101",
  8558=>"101111000",
  8559=>"111111000",
  8560=>"000000000",
  8561=>"000000000",
  8562=>"010111111",
  8563=>"000100111",
  8564=>"011011011",
  8565=>"000100100",
  8566=>"000000111",
  8567=>"110010000",
  8568=>"101000000",
  8569=>"111110000",
  8570=>"111011011",
  8571=>"000000100",
  8572=>"111111011",
  8573=>"000000001",
  8574=>"000110111",
  8575=>"101101111",
  8576=>"100000000",
  8577=>"000001011",
  8578=>"000000000",
  8579=>"001001001",
  8580=>"100000111",
  8581=>"000000111",
  8582=>"010010011",
  8583=>"000000001",
  8584=>"001000111",
  8585=>"111111101",
  8586=>"101001001",
  8587=>"110111111",
  8588=>"111111111",
  8589=>"100111000",
  8590=>"000000000",
  8591=>"111111010",
  8592=>"000000010",
  8593=>"111000000",
  8594=>"100111111",
  8595=>"111001000",
  8596=>"010000010",
  8597=>"000010000",
  8598=>"111111001",
  8599=>"110000001",
  8600=>"111111111",
  8601=>"101001000",
  8602=>"111111111",
  8603=>"101000111",
  8604=>"111111011",
  8605=>"111111000",
  8606=>"000000000",
  8607=>"111111111",
  8608=>"000000110",
  8609=>"100100011",
  8610=>"111111010",
  8611=>"111111111",
  8612=>"110111100",
  8613=>"011111000",
  8614=>"001001000",
  8615=>"111111111",
  8616=>"000000000",
  8617=>"111111011",
  8618=>"111111111",
  8619=>"000000000",
  8620=>"000000000",
  8621=>"000001001",
  8622=>"011111111",
  8623=>"111111100",
  8624=>"101000110",
  8625=>"000000000",
  8626=>"000010000",
  8627=>"100000111",
  8628=>"100100110",
  8629=>"001001101",
  8630=>"000001101",
  8631=>"110000000",
  8632=>"111000000",
  8633=>"111001100",
  8634=>"001000011",
  8635=>"110111111",
  8636=>"100000000",
  8637=>"111111111",
  8638=>"000000000",
  8639=>"100100100",
  8640=>"000000000",
  8641=>"101000111",
  8642=>"111110000",
  8643=>"110111000",
  8644=>"111111001",
  8645=>"000101111",
  8646=>"000000000",
  8647=>"110110100",
  8648=>"001000100",
  8649=>"001000111",
  8650=>"000000000",
  8651=>"011000000",
  8652=>"111000000",
  8653=>"111111001",
  8654=>"110001000",
  8655=>"100111110",
  8656=>"000000000",
  8657=>"000000100",
  8658=>"000111111",
  8659=>"000000000",
  8660=>"111111000",
  8661=>"111111000",
  8662=>"100101111",
  8663=>"000000011",
  8664=>"111111111",
  8665=>"111111110",
  8666=>"111000001",
  8667=>"111010100",
  8668=>"000010010",
  8669=>"111111010",
  8670=>"000000000",
  8671=>"100100100",
  8672=>"111111111",
  8673=>"011011000",
  8674=>"011011010",
  8675=>"111111000",
  8676=>"111111111",
  8677=>"100110111",
  8678=>"110000000",
  8679=>"111111011",
  8680=>"001001000",
  8681=>"111110000",
  8682=>"011011111",
  8683=>"100000100",
  8684=>"110111001",
  8685=>"100100100",
  8686=>"111111111",
  8687=>"000011111",
  8688=>"000001111",
  8689=>"010011010",
  8690=>"001001111",
  8691=>"111111000",
  8692=>"111011010",
  8693=>"000000000",
  8694=>"011011111",
  8695=>"110000000",
  8696=>"000000000",
  8697=>"000010000",
  8698=>"000000000",
  8699=>"100100100",
  8700=>"101001111",
  8701=>"101000000",
  8702=>"000101111",
  8703=>"000000111",
  8704=>"000000111",
  8705=>"111011111",
  8706=>"000111111",
  8707=>"111111011",
  8708=>"100000000",
  8709=>"111110100",
  8710=>"000000000",
  8711=>"000000011",
  8712=>"111111000",
  8713=>"010010111",
  8714=>"000001000",
  8715=>"111111111",
  8716=>"110110110",
  8717=>"111000000",
  8718=>"110000101",
  8719=>"001101101",
  8720=>"011110011",
  8721=>"111111111",
  8722=>"111111111",
  8723=>"000111111",
  8724=>"000110111",
  8725=>"000000110",
  8726=>"000000000",
  8727=>"000111111",
  8728=>"110000000",
  8729=>"000111111",
  8730=>"000000100",
  8731=>"001011111",
  8732=>"111000000",
  8733=>"111111111",
  8734=>"000011011",
  8735=>"011001000",
  8736=>"000000010",
  8737=>"100101111",
  8738=>"111110100",
  8739=>"000000000",
  8740=>"000000000",
  8741=>"111111111",
  8742=>"111111111",
  8743=>"010000000",
  8744=>"111111111",
  8745=>"001001111",
  8746=>"000000000",
  8747=>"101000001",
  8748=>"011111000",
  8749=>"000000011",
  8750=>"000000000",
  8751=>"000110111",
  8752=>"001111111",
  8753=>"000000000",
  8754=>"111011000",
  8755=>"111111011",
  8756=>"111011000",
  8757=>"110110100",
  8758=>"000000111",
  8759=>"000001001",
  8760=>"111111000",
  8761=>"000000001",
  8762=>"111100000",
  8763=>"000000000",
  8764=>"000000111",
  8765=>"110110110",
  8766=>"011011011",
  8767=>"001111111",
  8768=>"011001111",
  8769=>"011100000",
  8770=>"000000000",
  8771=>"110100111",
  8772=>"110111100",
  8773=>"000100111",
  8774=>"111101110",
  8775=>"100100000",
  8776=>"000000000",
  8777=>"100110111",
  8778=>"111011101",
  8779=>"111111110",
  8780=>"011111110",
  8781=>"101111111",
  8782=>"000010000",
  8783=>"111110000",
  8784=>"000110111",
  8785=>"000010010",
  8786=>"111111101",
  8787=>"111101100",
  8788=>"110111000",
  8789=>"111000000",
  8790=>"000001111",
  8791=>"111111000",
  8792=>"111111110",
  8793=>"111111000",
  8794=>"111111000",
  8795=>"111001000",
  8796=>"111111111",
  8797=>"110111111",
  8798=>"010001000",
  8799=>"111000000",
  8800=>"000100000",
  8801=>"000000000",
  8802=>"100000000",
  8803=>"111111111",
  8804=>"110000000",
  8805=>"000000100",
  8806=>"011000111",
  8807=>"111111111",
  8808=>"000011110",
  8809=>"001000000",
  8810=>"000000000",
  8811=>"000000000",
  8812=>"000000100",
  8813=>"010000111",
  8814=>"011000000",
  8815=>"001001111",
  8816=>"000111111",
  8817=>"000000111",
  8818=>"001000000",
  8819=>"111001000",
  8820=>"001111111",
  8821=>"111111111",
  8822=>"000000000",
  8823=>"000000000",
  8824=>"110110110",
  8825=>"000000001",
  8826=>"111111111",
  8827=>"111000000",
  8828=>"111111100",
  8829=>"011010011",
  8830=>"100000000",
  8831=>"111110100",
  8832=>"010111111",
  8833=>"111100110",
  8834=>"111111101",
  8835=>"011000000",
  8836=>"000000011",
  8837=>"111000000",
  8838=>"000000110",
  8839=>"000000000",
  8840=>"111011001",
  8841=>"000000000",
  8842=>"111000000",
  8843=>"000111111",
  8844=>"000000000",
  8845=>"000010111",
  8846=>"111100111",
  8847=>"100101111",
  8848=>"001001000",
  8849=>"000000000",
  8850=>"011110010",
  8851=>"111111000",
  8852=>"000000000",
  8853=>"110000000",
  8854=>"000111111",
  8855=>"110010000",
  8856=>"000110111",
  8857=>"000000001",
  8858=>"011000000",
  8859=>"111100000",
  8860=>"111111111",
  8861=>"000000111",
  8862=>"000000011",
  8863=>"110111000",
  8864=>"111111111",
  8865=>"111111111",
  8866=>"110000100",
  8867=>"000010111",
  8868=>"110100110",
  8869=>"010000010",
  8870=>"111111111",
  8871=>"110111001",
  8872=>"000000111",
  8873=>"111111100",
  8874=>"111111111",
  8875=>"000000000",
  8876=>"000000000",
  8877=>"000000000",
  8878=>"111000000",
  8879=>"111111010",
  8880=>"000100000",
  8881=>"000100100",
  8882=>"110111111",
  8883=>"000000000",
  8884=>"001000000",
  8885=>"111001000",
  8886=>"000000000",
  8887=>"101111111",
  8888=>"100100000",
  8889=>"110111010",
  8890=>"000000001",
  8891=>"111111111",
  8892=>"010000000",
  8893=>"100110000",
  8894=>"000000111",
  8895=>"001001111",
  8896=>"111111111",
  8897=>"000000111",
  8898=>"000000000",
  8899=>"111111111",
  8900=>"000000000",
  8901=>"011111111",
  8902=>"000100111",
  8903=>"111111100",
  8904=>"010110111",
  8905=>"000000101",
  8906=>"001000110",
  8907=>"110111111",
  8908=>"000000111",
  8909=>"000000001",
  8910=>"111111111",
  8911=>"000111000",
  8912=>"000011001",
  8913=>"111111111",
  8914=>"000000000",
  8915=>"000000000",
  8916=>"000000000",
  8917=>"111111101",
  8918=>"000000111",
  8919=>"000000101",
  8920=>"111000100",
  8921=>"001000001",
  8922=>"111011011",
  8923=>"000000000",
  8924=>"001000001",
  8925=>"110100000",
  8926=>"111000000",
  8927=>"000000110",
  8928=>"000010000",
  8929=>"100100011",
  8930=>"011111111",
  8931=>"001001000",
  8932=>"001001111",
  8933=>"110000000",
  8934=>"110111111",
  8935=>"111011010",
  8936=>"111011000",
  8937=>"100111011",
  8938=>"111000000",
  8939=>"000000111",
  8940=>"111111000",
  8941=>"111111110",
  8942=>"000111111",
  8943=>"111111111",
  8944=>"000000000",
  8945=>"111111111",
  8946=>"111111111",
  8947=>"101111111",
  8948=>"111111000",
  8949=>"111000011",
  8950=>"111000001",
  8951=>"111000000",
  8952=>"000000111",
  8953=>"000000010",
  8954=>"111000000",
  8955=>"111111000",
  8956=>"101101010",
  8957=>"000100110",
  8958=>"000011000",
  8959=>"000000000",
  8960=>"000000000",
  8961=>"111011011",
  8962=>"000100111",
  8963=>"011000000",
  8964=>"000000000",
  8965=>"111111111",
  8966=>"000000111",
  8967=>"111111000",
  8968=>"000100110",
  8969=>"000000000",
  8970=>"111000000",
  8971=>"001000000",
  8972=>"100000000",
  8973=>"000000111",
  8974=>"000000000",
  8975=>"000000000",
  8976=>"000000000",
  8977=>"000000101",
  8978=>"011000000",
  8979=>"111111000",
  8980=>"100000010",
  8981=>"000110111",
  8982=>"001001001",
  8983=>"000000000",
  8984=>"111001011",
  8985=>"000000000",
  8986=>"000111000",
  8987=>"000000000",
  8988=>"110111111",
  8989=>"111111101",
  8990=>"111011111",
  8991=>"111100000",
  8992=>"000000001",
  8993=>"111000000",
  8994=>"000000000",
  8995=>"001001111",
  8996=>"100101111",
  8997=>"011111111",
  8998=>"010111111",
  8999=>"111111001",
  9000=>"010010011",
  9001=>"110000000",
  9002=>"111000001",
  9003=>"001000000",
  9004=>"111111001",
  9005=>"111111100",
  9006=>"110111000",
  9007=>"111010000",
  9008=>"000000000",
  9009=>"110111111",
  9010=>"000001000",
  9011=>"111111111",
  9012=>"000000000",
  9013=>"111111010",
  9014=>"111111000",
  9015=>"100000111",
  9016=>"000000000",
  9017=>"111010011",
  9018=>"110111111",
  9019=>"000111111",
  9020=>"000000000",
  9021=>"000000000",
  9022=>"011001001",
  9023=>"111111111",
  9024=>"000000111",
  9025=>"011111011",
  9026=>"111111111",
  9027=>"111000000",
  9028=>"000000000",
  9029=>"111110111",
  9030=>"000000000",
  9031=>"000010000",
  9032=>"111111111",
  9033=>"100010111",
  9034=>"001000000",
  9035=>"000000100",
  9036=>"000000000",
  9037=>"101111111",
  9038=>"111111111",
  9039=>"111111111",
  9040=>"000000100",
  9041=>"000000110",
  9042=>"000000000",
  9043=>"000000011",
  9044=>"000011000",
  9045=>"011011011",
  9046=>"011000000",
  9047=>"111111111",
  9048=>"101100000",
  9049=>"001000000",
  9050=>"111111111",
  9051=>"010110111",
  9052=>"110111111",
  9053=>"111111111",
  9054=>"000000101",
  9055=>"000001011",
  9056=>"000000100",
  9057=>"111000000",
  9058=>"000100101",
  9059=>"010000111",
  9060=>"111000000",
  9061=>"000000000",
  9062=>"000001111",
  9063=>"111111111",
  9064=>"001001011",
  9065=>"000000111",
  9066=>"111111000",
  9067=>"010000001",
  9068=>"000001001",
  9069=>"001111111",
  9070=>"000000000",
  9071=>"111011010",
  9072=>"111001000",
  9073=>"000000000",
  9074=>"001000000",
  9075=>"000000000",
  9076=>"000111111",
  9077=>"001000000",
  9078=>"000111111",
  9079=>"111111111",
  9080=>"011000111",
  9081=>"111111001",
  9082=>"000000000",
  9083=>"110000000",
  9084=>"111111111",
  9085=>"000001111",
  9086=>"000000000",
  9087=>"000110000",
  9088=>"000110111",
  9089=>"111100100",
  9090=>"001001011",
  9091=>"100111111",
  9092=>"111111111",
  9093=>"111111010",
  9094=>"111111111",
  9095=>"001001101",
  9096=>"000000000",
  9097=>"001001111",
  9098=>"000000001",
  9099=>"111000000",
  9100=>"111001111",
  9101=>"000100110",
  9102=>"110000000",
  9103=>"111111000",
  9104=>"100000000",
  9105=>"001000000",
  9106=>"000000101",
  9107=>"000100110",
  9108=>"011000000",
  9109=>"000000000",
  9110=>"101101111",
  9111=>"000000100",
  9112=>"111011111",
  9113=>"000000000",
  9114=>"000000111",
  9115=>"111111001",
  9116=>"111111000",
  9117=>"110111000",
  9118=>"100110111",
  9119=>"111111000",
  9120=>"111110000",
  9121=>"110110011",
  9122=>"000000000",
  9123=>"010110111",
  9124=>"001111111",
  9125=>"000100000",
  9126=>"000000000",
  9127=>"111111111",
  9128=>"001000100",
  9129=>"111001111",
  9130=>"111000000",
  9131=>"000000000",
  9132=>"000001111",
  9133=>"111111001",
  9134=>"111111111",
  9135=>"100000000",
  9136=>"000000000",
  9137=>"000000000",
  9138=>"110100100",
  9139=>"000111111",
  9140=>"100100110",
  9141=>"111011011",
  9142=>"111111111",
  9143=>"111100100",
  9144=>"000000000",
  9145=>"111111111",
  9146=>"100000001",
  9147=>"111111011",
  9148=>"000001011",
  9149=>"111000100",
  9150=>"011000000",
  9151=>"010010000",
  9152=>"000000000",
  9153=>"111111110",
  9154=>"111111111",
  9155=>"000000111",
  9156=>"000000111",
  9157=>"000000011",
  9158=>"000000000",
  9159=>"011001000",
  9160=>"000000000",
  9161=>"111111110",
  9162=>"000000000",
  9163=>"111111000",
  9164=>"000000000",
  9165=>"111111111",
  9166=>"000000000",
  9167=>"000111111",
  9168=>"010000000",
  9169=>"000111000",
  9170=>"000000001",
  9171=>"101001001",
  9172=>"010000000",
  9173=>"000000000",
  9174=>"111111011",
  9175=>"111011000",
  9176=>"000000000",
  9177=>"000011111",
  9178=>"101000111",
  9179=>"000000000",
  9180=>"111000001",
  9181=>"001000000",
  9182=>"100000000",
  9183=>"011000000",
  9184=>"000000111",
  9185=>"111000000",
  9186=>"111111010",
  9187=>"111111000",
  9188=>"100010111",
  9189=>"111111100",
  9190=>"000000000",
  9191=>"111101111",
  9192=>"011011111",
  9193=>"001011011",
  9194=>"111000111",
  9195=>"000000111",
  9196=>"111111111",
  9197=>"000000000",
  9198=>"011111000",
  9199=>"000010000",
  9200=>"100000000",
  9201=>"111111111",
  9202=>"000100111",
  9203=>"111111100",
  9204=>"000000000",
  9205=>"100000000",
  9206=>"011111111",
  9207=>"110111111",
  9208=>"000000111",
  9209=>"000100100",
  9210=>"010111110",
  9211=>"000000000",
  9212=>"000000000",
  9213=>"000000111",
  9214=>"000000001",
  9215=>"100000100",
  9216=>"111111111",
  9217=>"000000000",
  9218=>"111111111",
  9219=>"111111000",
  9220=>"000011000",
  9221=>"001000000",
  9222=>"111111111",
  9223=>"111111101",
  9224=>"000110111",
  9225=>"100101111",
  9226=>"000000000",
  9227=>"001000001",
  9228=>"110110110",
  9229=>"111111111",
  9230=>"101000100",
  9231=>"000000111",
  9232=>"000000000",
  9233=>"000011000",
  9234=>"111111111",
  9235=>"000000100",
  9236=>"000000000",
  9237=>"111111101",
  9238=>"111111111",
  9239=>"000000000",
  9240=>"101111011",
  9241=>"000100111",
  9242=>"000000011",
  9243=>"111111011",
  9244=>"111111111",
  9245=>"100011000",
  9246=>"100111111",
  9247=>"000000100",
  9248=>"111111111",
  9249=>"100000000",
  9250=>"000000000",
  9251=>"000000000",
  9252=>"001111111",
  9253=>"000111101",
  9254=>"111100111",
  9255=>"100100001",
  9256=>"001011100",
  9257=>"010010000",
  9258=>"000000101",
  9259=>"000000001",
  9260=>"111111000",
  9261=>"110111111",
  9262=>"000000000",
  9263=>"001000000",
  9264=>"110111111",
  9265=>"000000001",
  9266=>"111101111",
  9267=>"000000000",
  9268=>"000000000",
  9269=>"000000000",
  9270=>"111111111",
  9271=>"111111111",
  9272=>"111111111",
  9273=>"000000001",
  9274=>"000000000",
  9275=>"000000000",
  9276=>"101101111",
  9277=>"000000000",
  9278=>"111111100",
  9279=>"111000000",
  9280=>"111001000",
  9281=>"111111111",
  9282=>"111001000",
  9283=>"100101100",
  9284=>"011011111",
  9285=>"110011001",
  9286=>"111110011",
  9287=>"111111000",
  9288=>"111111111",
  9289=>"000100110",
  9290=>"111111111",
  9291=>"000000000",
  9292=>"000000000",
  9293=>"000001001",
  9294=>"100100000",
  9295=>"111011111",
  9296=>"000000000",
  9297=>"111011000",
  9298=>"000000000",
  9299=>"011001111",
  9300=>"000000000",
  9301=>"000000000",
  9302=>"111111111",
  9303=>"000000000",
  9304=>"110100001",
  9305=>"000000100",
  9306=>"111111111",
  9307=>"000001110",
  9308=>"000000000",
  9309=>"111011011",
  9310=>"110111111",
  9311=>"000000000",
  9312=>"000000000",
  9313=>"000001111",
  9314=>"110110111",
  9315=>"000101111",
  9316=>"001000000",
  9317=>"111111000",
  9318=>"011001111",
  9319=>"111111111",
  9320=>"101111111",
  9321=>"011000000",
  9322=>"000011001",
  9323=>"000000000",
  9324=>"001011011",
  9325=>"000000011",
  9326=>"111111111",
  9327=>"111111101",
  9328=>"111111111",
  9329=>"101111111",
  9330=>"110010000",
  9331=>"100101000",
  9332=>"111111111",
  9333=>"000010000",
  9334=>"000000111",
  9335=>"001001001",
  9336=>"000001101",
  9337=>"111111111",
  9338=>"000011011",
  9339=>"001000001",
  9340=>"111111011",
  9341=>"000000000",
  9342=>"000000100",
  9343=>"000000000",
  9344=>"111111111",
  9345=>"100000000",
  9346=>"111110111",
  9347=>"111110100",
  9348=>"111111111",
  9349=>"100100100",
  9350=>"000100110",
  9351=>"011000000",
  9352=>"000000111",
  9353=>"000000000",
  9354=>"000010110",
  9355=>"000000110",
  9356=>"111011000",
  9357=>"111111111",
  9358=>"111111100",
  9359=>"001001001",
  9360=>"000000101",
  9361=>"000000000",
  9362=>"000000000",
  9363=>"010001111",
  9364=>"110111111",
  9365=>"000000000",
  9366=>"111111111",
  9367=>"111111111",
  9368=>"000010000",
  9369=>"000100110",
  9370=>"000000111",
  9371=>"000000000",
  9372=>"001001001",
  9373=>"001001000",
  9374=>"111000000",
  9375=>"111111111",
  9376=>"001001000",
  9377=>"001111111",
  9378=>"111111111",
  9379=>"000000010",
  9380=>"100110110",
  9381=>"000000000",
  9382=>"111111111",
  9383=>"000000000",
  9384=>"111001000",
  9385=>"001001001",
  9386=>"000000000",
  9387=>"101101100",
  9388=>"001000000",
  9389=>"111111111",
  9390=>"111111111",
  9391=>"000000000",
  9392=>"000001000",
  9393=>"111111000",
  9394=>"111111000",
  9395=>"111101111",
  9396=>"000000000",
  9397=>"100100000",
  9398=>"000000000",
  9399=>"000000000",
  9400=>"111111110",
  9401=>"111111111",
  9402=>"000100000",
  9403=>"000000000",
  9404=>"000000000",
  9405=>"000000000",
  9406=>"110111111",
  9407=>"000000000",
  9408=>"000000000",
  9409=>"000000000",
  9410=>"000100111",
  9411=>"010111111",
  9412=>"001000001",
  9413=>"111111010",
  9414=>"111111000",
  9415=>"010000000",
  9416=>"000110000",
  9417=>"111111101",
  9418=>"101000000",
  9419=>"100100000",
  9420=>"001000000",
  9421=>"000000111",
  9422=>"111111111",
  9423=>"000000100",
  9424=>"000000001",
  9425=>"111111011",
  9426=>"000001001",
  9427=>"111111010",
  9428=>"000000000",
  9429=>"110000000",
  9430=>"111111000",
  9431=>"111111111",
  9432=>"011111111",
  9433=>"110000110",
  9434=>"111101111",
  9435=>"111111011",
  9436=>"000111111",
  9437=>"111111111",
  9438=>"000000000",
  9439=>"001000000",
  9440=>"100000110",
  9441=>"000111111",
  9442=>"111111111",
  9443=>"111111111",
  9444=>"111111111",
  9445=>"000000000",
  9446=>"111000111",
  9447=>"000010010",
  9448=>"000000001",
  9449=>"111111111",
  9450=>"111111111",
  9451=>"101101101",
  9452=>"111111111",
  9453=>"111111111",
  9454=>"111111111",
  9455=>"000000000",
  9456=>"000000000",
  9457=>"000000111",
  9458=>"111111111",
  9459=>"101001111",
  9460=>"000000000",
  9461=>"000000000",
  9462=>"110000001",
  9463=>"011011000",
  9464=>"111111111",
  9465=>"000000000",
  9466=>"000000000",
  9467=>"111010000",
  9468=>"001000000",
  9469=>"111101111",
  9470=>"011001001",
  9471=>"110111111",
  9472=>"000000000",
  9473=>"111111111",
  9474=>"111111111",
  9475=>"001000000",
  9476=>"111101111",
  9477=>"000111100",
  9478=>"111111001",
  9479=>"100000100",
  9480=>"000000011",
  9481=>"011000000",
  9482=>"111111111",
  9483=>"111111111",
  9484=>"000000000",
  9485=>"000000000",
  9486=>"000000000",
  9487=>"000000000",
  9488=>"000000000",
  9489=>"001000000",
  9490=>"101000000",
  9491=>"110010011",
  9492=>"011011011",
  9493=>"010000000",
  9494=>"111111111",
  9495=>"001111111",
  9496=>"111011111",
  9497=>"100100111",
  9498=>"111111111",
  9499=>"000000000",
  9500=>"110100000",
  9501=>"100000101",
  9502=>"000000111",
  9503=>"111111111",
  9504=>"111111111",
  9505=>"100011000",
  9506=>"111111111",
  9507=>"000000101",
  9508=>"111110110",
  9509=>"111000000",
  9510=>"111000000",
  9511=>"100111010",
  9512=>"000000011",
  9513=>"000000110",
  9514=>"111001101",
  9515=>"100000111",
  9516=>"000000000",
  9517=>"001001111",
  9518=>"000000000",
  9519=>"000000000",
  9520=>"111111111",
  9521=>"000000000",
  9522=>"000000000",
  9523=>"000000000",
  9524=>"000000000",
  9525=>"110101110",
  9526=>"010000111",
  9527=>"111000000",
  9528=>"000000000",
  9529=>"111111111",
  9530=>"000000000",
  9531=>"111111001",
  9532=>"111111111",
  9533=>"000000000",
  9534=>"000111000",
  9535=>"000000101",
  9536=>"111101111",
  9537=>"111100000",
  9538=>"111011111",
  9539=>"111101000",
  9540=>"000000001",
  9541=>"000000000",
  9542=>"011011001",
  9543=>"111111101",
  9544=>"000000000",
  9545=>"000000010",
  9546=>"101001111",
  9547=>"100100000",
  9548=>"000000000",
  9549=>"000000000",
  9550=>"110110000",
  9551=>"011011011",
  9552=>"000011011",
  9553=>"001001000",
  9554=>"111111111",
  9555=>"000000000",
  9556=>"000000000",
  9557=>"011011011",
  9558=>"111111000",
  9559=>"100100100",
  9560=>"111111111",
  9561=>"100000000",
  9562=>"101101000",
  9563=>"000000000",
  9564=>"111111111",
  9565=>"000000000",
  9566=>"111111111",
  9567=>"110110111",
  9568=>"000000110",
  9569=>"000000000",
  9570=>"111101101",
  9571=>"000000000",
  9572=>"000000000",
  9573=>"000001000",
  9574=>"111111000",
  9575=>"000000111",
  9576=>"001001000",
  9577=>"000000000",
  9578=>"000000111",
  9579=>"111111001",
  9580=>"111111111",
  9581=>"111111101",
  9582=>"000000000",
  9583=>"000001000",
  9584=>"111111111",
  9585=>"111111111",
  9586=>"000000000",
  9587=>"001000000",
  9588=>"000000000",
  9589=>"000111111",
  9590=>"000000111",
  9591=>"111111111",
  9592=>"111111001",
  9593=>"001111111",
  9594=>"000000000",
  9595=>"111111111",
  9596=>"000000000",
  9597=>"000000001",
  9598=>"000000000",
  9599=>"011011011",
  9600=>"110000110",
  9601=>"000000111",
  9602=>"110000100",
  9603=>"000000000",
  9604=>"110111111",
  9605=>"000000111",
  9606=>"100100101",
  9607=>"111101000",
  9608=>"000110111",
  9609=>"000000111",
  9610=>"001001011",
  9611=>"010111111",
  9612=>"111111111",
  9613=>"000000000",
  9614=>"110000010",
  9615=>"000000000",
  9616=>"000000000",
  9617=>"110010111",
  9618=>"111111110",
  9619=>"111111110",
  9620=>"110111111",
  9621=>"000000000",
  9622=>"000000111",
  9623=>"111000001",
  9624=>"111111111",
  9625=>"000000000",
  9626=>"100000000",
  9627=>"100000111",
  9628=>"000000011",
  9629=>"111111001",
  9630=>"000001000",
  9631=>"000000000",
  9632=>"110111011",
  9633=>"110011011",
  9634=>"101111101",
  9635=>"111111111",
  9636=>"111001100",
  9637=>"000000100",
  9638=>"000000000",
  9639=>"010111001",
  9640=>"111111011",
  9641=>"000000000",
  9642=>"111111111",
  9643=>"000000001",
  9644=>"000000000",
  9645=>"101111100",
  9646=>"110111001",
  9647=>"000000001",
  9648=>"000000100",
  9649=>"000000010",
  9650=>"111111001",
  9651=>"000001011",
  9652=>"001001001",
  9653=>"111100000",
  9654=>"000000000",
  9655=>"000000000",
  9656=>"111111111",
  9657=>"111111000",
  9658=>"110000011",
  9659=>"011000000",
  9660=>"111011111",
  9661=>"100111111",
  9662=>"111001111",
  9663=>"011001000",
  9664=>"000000110",
  9665=>"111111111",
  9666=>"000000001",
  9667=>"000000000",
  9668=>"111001111",
  9669=>"011111101",
  9670=>"000000000",
  9671=>"111011011",
  9672=>"101111111",
  9673=>"000000000",
  9674=>"000000001",
  9675=>"111111111",
  9676=>"011001111",
  9677=>"111111101",
  9678=>"111111111",
  9679=>"000000000",
  9680=>"111111111",
  9681=>"001001001",
  9682=>"000000000",
  9683=>"111011000",
  9684=>"000000101",
  9685=>"111111111",
  9686=>"111111000",
  9687=>"001011011",
  9688=>"000000000",
  9689=>"000000000",
  9690=>"000010111",
  9691=>"111111111",
  9692=>"111111111",
  9693=>"000000101",
  9694=>"000111111",
  9695=>"000000100",
  9696=>"111111000",
  9697=>"000000000",
  9698=>"000000000",
  9699=>"000001000",
  9700=>"000000001",
  9701=>"111111011",
  9702=>"100000000",
  9703=>"000000000",
  9704=>"111111111",
  9705=>"011010000",
  9706=>"000000000",
  9707=>"011010111",
  9708=>"000001001",
  9709=>"101000000",
  9710=>"010011111",
  9711=>"001101101",
  9712=>"000001000",
  9713=>"011000001",
  9714=>"111111111",
  9715=>"000000000",
  9716=>"001011000",
  9717=>"000000000",
  9718=>"000000000",
  9719=>"000100000",
  9720=>"000000000",
  9721=>"000000000",
  9722=>"111111111",
  9723=>"001001111",
  9724=>"111111111",
  9725=>"111111111",
  9726=>"000000000",
  9727=>"000000000",
  9728=>"010111011",
  9729=>"111001000",
  9730=>"000111111",
  9731=>"000000001",
  9732=>"100111111",
  9733=>"000111111",
  9734=>"100000100",
  9735=>"111100000",
  9736=>"111111111",
  9737=>"111111111",
  9738=>"000000000",
  9739=>"011011000",
  9740=>"000000000",
  9741=>"111111111",
  9742=>"000000000",
  9743=>"010000000",
  9744=>"111110001",
  9745=>"101111111",
  9746=>"000000001",
  9747=>"010010111",
  9748=>"001101000",
  9749=>"000101111",
  9750=>"111011000",
  9751=>"110110000",
  9752=>"011111111",
  9753=>"111011000",
  9754=>"011011111",
  9755=>"010010000",
  9756=>"111111111",
  9757=>"000000010",
  9758=>"111011011",
  9759=>"111111111",
  9760=>"000000111",
  9761=>"111111111",
  9762=>"110111111",
  9763=>"100100111",
  9764=>"110100000",
  9765=>"111111000",
  9766=>"010010111",
  9767=>"000100111",
  9768=>"010111111",
  9769=>"000000000",
  9770=>"011011010",
  9771=>"000101111",
  9772=>"111111111",
  9773=>"000000111",
  9774=>"111111111",
  9775=>"000000000",
  9776=>"111111111",
  9777=>"000000000",
  9778=>"111010000",
  9779=>"110011011",
  9780=>"000000000",
  9781=>"000000000",
  9782=>"001100100",
  9783=>"000000110",
  9784=>"111100111",
  9785=>"000000000",
  9786=>"000000000",
  9787=>"000000111",
  9788=>"001001000",
  9789=>"111011001",
  9790=>"111110000",
  9791=>"000000000",
  9792=>"000001111",
  9793=>"001110000",
  9794=>"100111111",
  9795=>"111111001",
  9796=>"000000000",
  9797=>"000000011",
  9798=>"111111111",
  9799=>"111111010",
  9800=>"111111110",
  9801=>"101101111",
  9802=>"000000000",
  9803=>"000010010",
  9804=>"111001101",
  9805=>"111110000",
  9806=>"000110111",
  9807=>"110000111",
  9808=>"000000000",
  9809=>"000000000",
  9810=>"111111111",
  9811=>"110111000",
  9812=>"000000000",
  9813=>"000000000",
  9814=>"011000110",
  9815=>"000000000",
  9816=>"000000000",
  9817=>"001001001",
  9818=>"000000101",
  9819=>"111111111",
  9820=>"000000000",
  9821=>"000011000",
  9822=>"001111111",
  9823=>"111100000",
  9824=>"000000110",
  9825=>"000000111",
  9826=>"000000000",
  9827=>"000001111",
  9828=>"111111111",
  9829=>"000000000",
  9830=>"000000000",
  9831=>"000000000",
  9832=>"110111000",
  9833=>"000000010",
  9834=>"011000000",
  9835=>"000000000",
  9836=>"001011000",
  9837=>"111111100",
  9838=>"000000011",
  9839=>"111111000",
  9840=>"000000111",
  9841=>"111010001",
  9842=>"111111000",
  9843=>"000000110",
  9844=>"111111000",
  9845=>"000111111",
  9846=>"000000001",
  9847=>"000000111",
  9848=>"000011111",
  9849=>"000000000",
  9850=>"000000111",
  9851=>"000000000",
  9852=>"111110000",
  9853=>"011111111",
  9854=>"100100111",
  9855=>"111111010",
  9856=>"000100111",
  9857=>"111000111",
  9858=>"011011111",
  9859=>"110111000",
  9860=>"000000000",
  9861=>"001000000",
  9862=>"011111000",
  9863=>"010110111",
  9864=>"010000010",
  9865=>"000000111",
  9866=>"000000000",
  9867=>"000111111",
  9868=>"110000000",
  9869=>"000000010",
  9870=>"000000111",
  9871=>"111111000",
  9872=>"111000000",
  9873=>"101100111",
  9874=>"110000010",
  9875=>"111111010",
  9876=>"000000000",
  9877=>"000000000",
  9878=>"000000000",
  9879=>"000111111",
  9880=>"000000100",
  9881=>"111111000",
  9882=>"100000000",
  9883=>"000010011",
  9884=>"000000010",
  9885=>"000000010",
  9886=>"011011001",
  9887=>"000000100",
  9888=>"110000000",
  9889=>"001000010",
  9890=>"100000010",
  9891=>"110010000",
  9892=>"000000001",
  9893=>"110111111",
  9894=>"111111000",
  9895=>"000000000",
  9896=>"111111111",
  9897=>"111111111",
  9898=>"111111111",
  9899=>"100000010",
  9900=>"000000000",
  9901=>"110010000",
  9902=>"111111111",
  9903=>"110110000",
  9904=>"000000111",
  9905=>"111010010",
  9906=>"111111111",
  9907=>"111111000",
  9908=>"110000000",
  9909=>"000001111",
  9910=>"000000000",
  9911=>"111111111",
  9912=>"110110011",
  9913=>"000000000",
  9914=>"000000000",
  9915=>"000000111",
  9916=>"111000010",
  9917=>"000111111",
  9918=>"001100111",
  9919=>"000111110",
  9920=>"111111110",
  9921=>"111110111",
  9922=>"111111111",
  9923=>"111101111",
  9924=>"000111110",
  9925=>"111111111",
  9926=>"000010111",
  9927=>"000011111",
  9928=>"000000000",
  9929=>"111111000",
  9930=>"000100000",
  9931=>"000000111",
  9932=>"111111101",
  9933=>"111111111",
  9934=>"000000110",
  9935=>"111111111",
  9936=>"000000000",
  9937=>"001001111",
  9938=>"111101000",
  9939=>"000000000",
  9940=>"110101000",
  9941=>"111111111",
  9942=>"000000010",
  9943=>"000000000",
  9944=>"000000000",
  9945=>"011011011",
  9946=>"000000000",
  9947=>"000100100",
  9948=>"000000000",
  9949=>"111111111",
  9950=>"000000000",
  9951=>"000000011",
  9952=>"000000000",
  9953=>"011111111",
  9954=>"000000000",
  9955=>"101111111",
  9956=>"111110000",
  9957=>"111101100",
  9958=>"011000000",
  9959=>"111011011",
  9960=>"000000000",
  9961=>"011111111",
  9962=>"000100111",
  9963=>"000000000",
  9964=>"000000000",
  9965=>"000010111",
  9966=>"000000111",
  9967=>"111111111",
  9968=>"000111000",
  9969=>"000010010",
  9970=>"000100111",
  9971=>"011010011",
  9972=>"111111111",
  9973=>"110011001",
  9974=>"111111111",
  9975=>"000000001",
  9976=>"000000010",
  9977=>"111100000",
  9978=>"111111010",
  9979=>"000111111",
  9980=>"111110000",
  9981=>"111001011",
  9982=>"111111111",
  9983=>"111111111",
  9984=>"010000000",
  9985=>"111111000",
  9986=>"111000000",
  9987=>"100111111",
  9988=>"100101111",
  9989=>"111111111",
  9990=>"000111111",
  9991=>"111111000",
  9992=>"111110100",
  9993=>"000010111",
  9994=>"000000000",
  9995=>"100000000",
  9996=>"001001111",
  9997=>"111111110",
  9998=>"111111000",
  9999=>"111111110",
  10000=>"110000000",
  10001=>"000000000",
  10002=>"000000111",
  10003=>"000000000",
  10004=>"111000000",
  10005=>"000000000",
  10006=>"100000000",
  10007=>"000000000",
  10008=>"000001011",
  10009=>"000000101",
  10010=>"000000110",
  10011=>"100101111",
  10012=>"101111110",
  10013=>"000000000",
  10014=>"111111000",
  10015=>"110100000",
  10016=>"010000000",
  10017=>"100111111",
  10018=>"111111000",
  10019=>"100101000",
  10020=>"000000000",
  10021=>"101000000",
  10022=>"011111111",
  10023=>"111111111",
  10024=>"000000110",
  10025=>"011111111",
  10026=>"111111111",
  10027=>"011011111",
  10028=>"000000100",
  10029=>"000011111",
  10030=>"000100100",
  10031=>"000000000",
  10032=>"000011111",
  10033=>"011111111",
  10034=>"111001001",
  10035=>"000110111",
  10036=>"111111110",
  10037=>"110111111",
  10038=>"000000000",
  10039=>"000000000",
  10040=>"000000100",
  10041=>"111111100",
  10042=>"000001011",
  10043=>"001001111",
  10044=>"000011011",
  10045=>"111111000",
  10046=>"111110000",
  10047=>"000010111",
  10048=>"000000000",
  10049=>"110111111",
  10050=>"000111100",
  10051=>"111000000",
  10052=>"000011111",
  10053=>"101000000",
  10054=>"111111000",
  10055=>"000001111",
  10056=>"000110110",
  10057=>"000000000",
  10058=>"001000000",
  10059=>"111000000",
  10060=>"000000000",
  10061=>"000000000",
  10062=>"000000001",
  10063=>"000000000",
  10064=>"000000000",
  10065=>"111100111",
  10066=>"111100000",
  10067=>"110010000",
  10068=>"010111110",
  10069=>"111011000",
  10070=>"111111000",
  10071=>"000000000",
  10072=>"110111111",
  10073=>"000000100",
  10074=>"111011011",
  10075=>"110111111",
  10076=>"111111101",
  10077=>"000000000",
  10078=>"001000010",
  10079=>"110000000",
  10080=>"000000000",
  10081=>"111111001",
  10082=>"111100000",
  10083=>"000000000",
  10084=>"000000000",
  10085=>"010000000",
  10086=>"000000010",
  10087=>"110111111",
  10088=>"000000000",
  10089=>"000000000",
  10090=>"111111111",
  10091=>"111101111",
  10092=>"111011000",
  10093=>"000010010",
  10094=>"000111111",
  10095=>"000000100",
  10096=>"000000000",
  10097=>"000000000",
  10098=>"111111111",
  10099=>"000100001",
  10100=>"111111111",
  10101=>"111110000",
  10102=>"000000100",
  10103=>"100000000",
  10104=>"111111111",
  10105=>"110111111",
  10106=>"000000000",
  10107=>"111111110",
  10108=>"111000000",
  10109=>"111101111",
  10110=>"000000000",
  10111=>"001001111",
  10112=>"110111001",
  10113=>"111111111",
  10114=>"100000000",
  10115=>"011000110",
  10116=>"000000000",
  10117=>"000001111",
  10118=>"100000100",
  10119=>"111111010",
  10120=>"000000000",
  10121=>"000010100",
  10122=>"000000101",
  10123=>"111001111",
  10124=>"111111111",
  10125=>"011111011",
  10126=>"111111000",
  10127=>"011011000",
  10128=>"111101000",
  10129=>"000000000",
  10130=>"110110111",
  10131=>"110110110",
  10132=>"111000000",
  10133=>"000000000",
  10134=>"111111100",
  10135=>"011010000",
  10136=>"000011111",
  10137=>"111111111",
  10138=>"111111000",
  10139=>"111111011",
  10140=>"001000101",
  10141=>"111111111",
  10142=>"111001001",
  10143=>"111011111",
  10144=>"000000000",
  10145=>"111111000",
  10146=>"000000111",
  10147=>"000011111",
  10148=>"111111111",
  10149=>"110100000",
  10150=>"100101111",
  10151=>"111111111",
  10152=>"000000000",
  10153=>"100000000",
  10154=>"000000000",
  10155=>"110001001",
  10156=>"000000000",
  10157=>"100101111",
  10158=>"000001111",
  10159=>"000000000",
  10160=>"011111010",
  10161=>"111011011",
  10162=>"111100001",
  10163=>"000000000",
  10164=>"000000000",
  10165=>"000000001",
  10166=>"000000001",
  10167=>"100100000",
  10168=>"111111000",
  10169=>"001111111",
  10170=>"111001100",
  10171=>"100010001",
  10172=>"111111111",
  10173=>"100100000",
  10174=>"000001111",
  10175=>"000000000",
  10176=>"001111111",
  10177=>"000000000",
  10178=>"111111000",
  10179=>"000000000",
  10180=>"111111111",
  10181=>"110110000",
  10182=>"000011111",
  10183=>"000111011",
  10184=>"000000000",
  10185=>"111000111",
  10186=>"000000110",
  10187=>"111110000",
  10188=>"111001100",
  10189=>"111111000",
  10190=>"000011111",
  10191=>"100100000",
  10192=>"000000111",
  10193=>"000000000",
  10194=>"000100111",
  10195=>"111100110",
  10196=>"111010011",
  10197=>"111111100",
  10198=>"000000111",
  10199=>"000000010",
  10200=>"000110111",
  10201=>"110000000",
  10202=>"000000000",
  10203=>"111111111",
  10204=>"111111100",
  10205=>"010010000",
  10206=>"110111110",
  10207=>"000001000",
  10208=>"111101111",
  10209=>"000000011",
  10210=>"111111111",
  10211=>"111110000",
  10212=>"111111111",
  10213=>"000000001",
  10214=>"111111100",
  10215=>"000000000",
  10216=>"111011011",
  10217=>"111111111",
  10218=>"111111111",
  10219=>"100100100",
  10220=>"000011111",
  10221=>"000000000",
  10222=>"000000000",
  10223=>"100000001",
  10224=>"111100000",
  10225=>"111111111",
  10226=>"110110111",
  10227=>"000000111",
  10228=>"000111111",
  10229=>"000000000",
  10230=>"000000101",
  10231=>"001000000",
  10232=>"111111111",
  10233=>"011001000",
  10234=>"101000000",
  10235=>"111011111",
  10236=>"111111111",
  10237=>"100000000",
  10238=>"111111111",
  10239=>"000000101",
  10240=>"110000000",
  10241=>"111110110",
  10242=>"111011111",
  10243=>"110000000",
  10244=>"000000000",
  10245=>"111000000",
  10246=>"101100100",
  10247=>"000011111",
  10248=>"001011000",
  10249=>"000001111",
  10250=>"011010000",
  10251=>"000111110",
  10252=>"000000110",
  10253=>"111000000",
  10254=>"110111011",
  10255=>"000000100",
  10256=>"000000010",
  10257=>"111111111",
  10258=>"000000100",
  10259=>"011111111",
  10260=>"111000000",
  10261=>"000000111",
  10262=>"000000111",
  10263=>"110100000",
  10264=>"111111000",
  10265=>"011011111",
  10266=>"011011000",
  10267=>"111011111",
  10268=>"000000111",
  10269=>"000000000",
  10270=>"001111101",
  10271=>"111000011",
  10272=>"110110110",
  10273=>"111100000",
  10274=>"000001000",
  10275=>"000101100",
  10276=>"110011011",
  10277=>"010111110",
  10278=>"010111111",
  10279=>"111000111",
  10280=>"111111111",
  10281=>"000111000",
  10282=>"001000000",
  10283=>"000100100",
  10284=>"100111000",
  10285=>"000101111",
  10286=>"101100111",
  10287=>"100110110",
  10288=>"000000000",
  10289=>"111001001",
  10290=>"000111111",
  10291=>"111111000",
  10292=>"000010000",
  10293=>"110111101",
  10294=>"000000111",
  10295=>"000011111",
  10296=>"110110111",
  10297=>"000110010",
  10298=>"000000101",
  10299=>"000000111",
  10300=>"111110000",
  10301=>"010111111",
  10302=>"001000000",
  10303=>"100100101",
  10304=>"000000101",
  10305=>"000000000",
  10306=>"100100101",
  10307=>"100000000",
  10308=>"000001000",
  10309=>"000000111",
  10310=>"111110000",
  10311=>"111111000",
  10312=>"000000001",
  10313=>"111111111",
  10314=>"100110000",
  10315=>"110100110",
  10316=>"111000000",
  10317=>"111111000",
  10318=>"111011001",
  10319=>"000000111",
  10320=>"000000110",
  10321=>"000000000",
  10322=>"110100000",
  10323=>"111100100",
  10324=>"011000000",
  10325=>"001000000",
  10326=>"000000101",
  10327=>"000111111",
  10328=>"000001000",
  10329=>"111000000",
  10330=>"100000001",
  10331=>"111111100",
  10332=>"111111000",
  10333=>"000001100",
  10334=>"000100100",
  10335=>"110110000",
  10336=>"100110000",
  10337=>"100000000",
  10338=>"011111011",
  10339=>"111111111",
  10340=>"000001000",
  10341=>"111111000",
  10342=>"000000111",
  10343=>"111111111",
  10344=>"101111111",
  10345=>"000000110",
  10346=>"111010111",
  10347=>"000000001",
  10348=>"100000000",
  10349=>"100110111",
  10350=>"000000111",
  10351=>"000111111",
  10352=>"000111111",
  10353=>"111001000",
  10354=>"000111111",
  10355=>"000110011",
  10356=>"010000001",
  10357=>"111111111",
  10358=>"000000000",
  10359=>"100110100",
  10360=>"110110000",
  10361=>"111111111",
  10362=>"111000000",
  10363=>"000000000",
  10364=>"110111000",
  10365=>"111111111",
  10366=>"010000000",
  10367=>"000000000",
  10368=>"000100111",
  10369=>"100000110",
  10370=>"111000111",
  10371=>"011111000",
  10372=>"111110110",
  10373=>"111111001",
  10374=>"111111111",
  10375=>"111111000",
  10376=>"001101111",
  10377=>"100000111",
  10378=>"111010010",
  10379=>"100000101",
  10380=>"000000010",
  10381=>"000111111",
  10382=>"000001101",
  10383=>"000000000",
  10384=>"000111001",
  10385=>"111111001",
  10386=>"000100111",
  10387=>"111000111",
  10388=>"111110000",
  10389=>"111000111",
  10390=>"111111111",
  10391=>"111111000",
  10392=>"000000101",
  10393=>"100111111",
  10394=>"010111110",
  10395=>"101011000",
  10396=>"111111111",
  10397=>"110111100",
  10398=>"111110000",
  10399=>"100100100",
  10400=>"111111110",
  10401=>"000000011",
  10402=>"000000111",
  10403=>"110111001",
  10404=>"111000000",
  10405=>"111000000",
  10406=>"000111000",
  10407=>"000110010",
  10408=>"000011111",
  10409=>"100000000",
  10410=>"110000001",
  10411=>"111001001",
  10412=>"000111111",
  10413=>"111111000",
  10414=>"101000000",
  10415=>"110110000",
  10416=>"110000000",
  10417=>"110111111",
  10418=>"111111000",
  10419=>"111111000",
  10420=>"000000000",
  10421=>"111111010",
  10422=>"000101100",
  10423=>"111110000",
  10424=>"111010000",
  10425=>"000000111",
  10426=>"111100000",
  10427=>"000011111",
  10428=>"000111111",
  10429=>"111111011",
  10430=>"111111111",
  10431=>"000011011",
  10432=>"000000000",
  10433=>"000110110",
  10434=>"000000111",
  10435=>"010111010",
  10436=>"111111110",
  10437=>"000110011",
  10438=>"111111111",
  10439=>"111110000",
  10440=>"000000111",
  10441=>"000101111",
  10442=>"101101100",
  10443=>"000000000",
  10444=>"100000100",
  10445=>"000000111",
  10446=>"111100111",
  10447=>"000101111",
  10448=>"111111111",
  10449=>"010110110",
  10450=>"000000100",
  10451=>"110000000",
  10452=>"000000011",
  10453=>"111000001",
  10454=>"000111111",
  10455=>"100101110",
  10456=>"110110111",
  10457=>"000111111",
  10458=>"111101101",
  10459=>"000111111",
  10460=>"000011111",
  10461=>"111101000",
  10462=>"000000111",
  10463=>"100000000",
  10464=>"111111111",
  10465=>"111111000",
  10466=>"000001001",
  10467=>"000000001",
  10468=>"111101000",
  10469=>"111111111",
  10470=>"111111110",
  10471=>"000000000",
  10472=>"111111000",
  10473=>"000010010",
  10474=>"011000001",
  10475=>"100111111",
  10476=>"000000111",
  10477=>"111111111",
  10478=>"000000000",
  10479=>"000000100",
  10480=>"101001000",
  10481=>"100100111",
  10482=>"111111101",
  10483=>"111000000",
  10484=>"001011011",
  10485=>"000111111",
  10486=>"000100000",
  10487=>"010000000",
  10488=>"111101101",
  10489=>"000111111",
  10490=>"111111111",
  10491=>"010111010",
  10492=>"000001111",
  10493=>"101111111",
  10494=>"000100110",
  10495=>"100000101",
  10496=>"000000000",
  10497=>"000000111",
  10498=>"100111111",
  10499=>"000011111",
  10500=>"000100111",
  10501=>"000000000",
  10502=>"100000110",
  10503=>"000111000",
  10504=>"011000000",
  10505=>"011000010",
  10506=>"100000000",
  10507=>"111000111",
  10508=>"101000111",
  10509=>"100100100",
  10510=>"110110000",
  10511=>"000111111",
  10512=>"000101000",
  10513=>"000101101",
  10514=>"111000000",
  10515=>"110101000",
  10516=>"001000000",
  10517=>"100111001",
  10518=>"001111111",
  10519=>"111111000",
  10520=>"011001111",
  10521=>"111111001",
  10522=>"000111111",
  10523=>"000111111",
  10524=>"001000110",
  10525=>"000000111",
  10526=>"111111111",
  10527=>"110000000",
  10528=>"110100000",
  10529=>"011000000",
  10530=>"000111110",
  10531=>"001000001",
  10532=>"111111000",
  10533=>"010110000",
  10534=>"000000101",
  10535=>"110100100",
  10536=>"111100110",
  10537=>"000000111",
  10538=>"000011011",
  10539=>"011011001",
  10540=>"111111111",
  10541=>"110011010",
  10542=>"111111000",
  10543=>"000000000",
  10544=>"111111110",
  10545=>"111101111",
  10546=>"111000000",
  10547=>"000001111",
  10548=>"111001000",
  10549=>"000000000",
  10550=>"000011111",
  10551=>"011001000",
  10552=>"111111000",
  10553=>"111001111",
  10554=>"111110101",
  10555=>"000000111",
  10556=>"001011001",
  10557=>"101001000",
  10558=>"000000000",
  10559=>"000000000",
  10560=>"111011000",
  10561=>"111000000",
  10562=>"111111011",
  10563=>"111000010",
  10564=>"000110111",
  10565=>"111111111",
  10566=>"111111111",
  10567=>"001111000",
  10568=>"110101000",
  10569=>"111100000",
  10570=>"100000110",
  10571=>"010000010",
  10572=>"000111111",
  10573=>"000011111",
  10574=>"100000000",
  10575=>"000111111",
  10576=>"000111000",
  10577=>"111111000",
  10578=>"000110110",
  10579=>"000111110",
  10580=>"000011000",
  10581=>"111011000",
  10582=>"100000010",
  10583=>"000000111",
  10584=>"110000000",
  10585=>"001001000",
  10586=>"111111000",
  10587=>"111111100",
  10588=>"000011111",
  10589=>"000100110",
  10590=>"000000000",
  10591=>"011111111",
  10592=>"111000001",
  10593=>"000000111",
  10594=>"011111111",
  10595=>"101111111",
  10596=>"000011111",
  10597=>"000000110",
  10598=>"000100000",
  10599=>"001110100",
  10600=>"001000110",
  10601=>"010111111",
  10602=>"001010010",
  10603=>"000001001",
  10604=>"110000000",
  10605=>"111011000",
  10606=>"110100100",
  10607=>"000000000",
  10608=>"000000000",
  10609=>"111001000",
  10610=>"110000000",
  10611=>"011000000",
  10612=>"000000111",
  10613=>"101000000",
  10614=>"000000001",
  10615=>"000011011",
  10616=>"111111111",
  10617=>"011000000",
  10618=>"111000000",
  10619=>"001111111",
  10620=>"111111111",
  10621=>"110110111",
  10622=>"000000000",
  10623=>"000000100",
  10624=>"000010110",
  10625=>"100100000",
  10626=>"000000111",
  10627=>"000000000",
  10628=>"000011001",
  10629=>"111111111",
  10630=>"000000000",
  10631=>"111000000",
  10632=>"000000000",
  10633=>"011011011",
  10634=>"000000000",
  10635=>"001111111",
  10636=>"101000001",
  10637=>"011010000",
  10638=>"011111011",
  10639=>"111111111",
  10640=>"110000000",
  10641=>"111111111",
  10642=>"000001111",
  10643=>"000000000",
  10644=>"111001111",
  10645=>"000110000",
  10646=>"011000000",
  10647=>"111111000",
  10648=>"111001111",
  10649=>"000001100",
  10650=>"000000111",
  10651=>"111111111",
  10652=>"101111111",
  10653=>"111111110",
  10654=>"000011111",
  10655=>"111110010",
  10656=>"000000101",
  10657=>"011111111",
  10658=>"010000100",
  10659=>"011111011",
  10660=>"100000111",
  10661=>"100110000",
  10662=>"111111000",
  10663=>"111111000",
  10664=>"010000100",
  10665=>"000000011",
  10666=>"000000010",
  10667=>"111111000",
  10668=>"000110111",
  10669=>"100110000",
  10670=>"000111111",
  10671=>"011111001",
  10672=>"101111111",
  10673=>"000000011",
  10674=>"000000000",
  10675=>"000000000",
  10676=>"111111000",
  10677=>"111110111",
  10678=>"100000111",
  10679=>"001011011",
  10680=>"100001111",
  10681=>"101000000",
  10682=>"100000111",
  10683=>"010001011",
  10684=>"011000000",
  10685=>"111111011",
  10686=>"000111111",
  10687=>"111111001",
  10688=>"100110000",
  10689=>"010110000",
  10690=>"000111010",
  10691=>"000110000",
  10692=>"100000000",
  10693=>"000011111",
  10694=>"111110000",
  10695=>"000111111",
  10696=>"001000111",
  10697=>"111100001",
  10698=>"000000111",
  10699=>"111000000",
  10700=>"111111010",
  10701=>"000000000",
  10702=>"110110100",
  10703=>"100111111",
  10704=>"011000000",
  10705=>"010000000",
  10706=>"000111111",
  10707=>"001111111",
  10708=>"010110110",
  10709=>"111000000",
  10710=>"000010000",
  10711=>"000110001",
  10712=>"001111111",
  10713=>"111111000",
  10714=>"111000011",
  10715=>"000000111",
  10716=>"000111111",
  10717=>"110100000",
  10718=>"111111000",
  10719=>"000111111",
  10720=>"000001111",
  10721=>"111111000",
  10722=>"111000000",
  10723=>"111111111",
  10724=>"100000110",
  10725=>"100000011",
  10726=>"110111000",
  10727=>"000101111",
  10728=>"000000111",
  10729=>"000001001",
  10730=>"100111111",
  10731=>"100100111",
  10732=>"111000000",
  10733=>"111111000",
  10734=>"000010111",
  10735=>"111111111",
  10736=>"111111001",
  10737=>"110001000",
  10738=>"101100100",
  10739=>"000000000",
  10740=>"111000000",
  10741=>"000000111",
  10742=>"100000000",
  10743=>"111111000",
  10744=>"111111111",
  10745=>"010110000",
  10746=>"110000001",
  10747=>"110111000",
  10748=>"000000101",
  10749=>"111111000",
  10750=>"000000111",
  10751=>"000000011",
  10752=>"111111110",
  10753=>"111111101",
  10754=>"111111111",
  10755=>"111111100",
  10756=>"111110110",
  10757=>"001111111",
  10758=>"111001000",
  10759=>"000000000",
  10760=>"000000010",
  10761=>"100000000",
  10762=>"110000000",
  10763=>"111111111",
  10764=>"111100100",
  10765=>"111111111",
  10766=>"000000000",
  10767=>"101000100",
  10768=>"011011011",
  10769=>"000010000",
  10770=>"100111000",
  10771=>"000000111",
  10772=>"001001111",
  10773=>"000000000",
  10774=>"001000000",
  10775=>"111111111",
  10776=>"100001001",
  10777=>"111111110",
  10778=>"111111111",
  10779=>"001011001",
  10780=>"000011111",
  10781=>"011010101",
  10782=>"111111111",
  10783=>"100101111",
  10784=>"111000111",
  10785=>"110110100",
  10786=>"100000100",
  10787=>"110000110",
  10788=>"000000000",
  10789=>"111111011",
  10790=>"110110110",
  10791=>"111001000",
  10792=>"111111100",
  10793=>"000000000",
  10794=>"000001000",
  10795=>"110100111",
  10796=>"000101111",
  10797=>"000000110",
  10798=>"000000000",
  10799=>"000100011",
  10800=>"111111101",
  10801=>"001000000",
  10802=>"011011000",
  10803=>"111011011",
  10804=>"100110110",
  10805=>"111111110",
  10806=>"000000000",
  10807=>"011001000",
  10808=>"000000000",
  10809=>"111111100",
  10810=>"000000000",
  10811=>"000001001",
  10812=>"111111111",
  10813=>"000111111",
  10814=>"000000011",
  10815=>"000000001",
  10816=>"000000110",
  10817=>"010000000",
  10818=>"111111111",
  10819=>"111111110",
  10820=>"001001111",
  10821=>"000000000",
  10822=>"000000001",
  10823=>"111111111",
  10824=>"111111111",
  10825=>"111000111",
  10826=>"000010011",
  10827=>"111111111",
  10828=>"111111000",
  10829=>"111111111",
  10830=>"000100100",
  10831=>"011011000",
  10832=>"000011000",
  10833=>"111001111",
  10834=>"011011011",
  10835=>"100100000",
  10836=>"111111010",
  10837=>"111010000",
  10838=>"111110110",
  10839=>"000000000",
  10840=>"111111111",
  10841=>"111000001",
  10842=>"000010011",
  10843=>"000000100",
  10844=>"111111111",
  10845=>"101111111",
  10846=>"000000000",
  10847=>"000000000",
  10848=>"000000000",
  10849=>"100100100",
  10850=>"111000110",
  10851=>"000101000",
  10852=>"111101100",
  10853=>"111000000",
  10854=>"000010000",
  10855=>"010000000",
  10856=>"000000000",
  10857=>"000000111",
  10858=>"010000000",
  10859=>"010010011",
  10860=>"111111111",
  10861=>"000000000",
  10862=>"101000000",
  10863=>"000000000",
  10864=>"111111111",
  10865=>"111010110",
  10866=>"110110111",
  10867=>"110111111",
  10868=>"111101101",
  10869=>"000000000",
  10870=>"000000000",
  10871=>"011011000",
  10872=>"111111111",
  10873=>"110101111",
  10874=>"010011000",
  10875=>"000000100",
  10876=>"110101100",
  10877=>"000000000",
  10878=>"111110000",
  10879=>"000000000",
  10880=>"111101001",
  10881=>"000111011",
  10882=>"100111111",
  10883=>"111111111",
  10884=>"101110000",
  10885=>"100100111",
  10886=>"111110000",
  10887=>"111001000",
  10888=>"111111111",
  10889=>"000000000",
  10890=>"011000000",
  10891=>"011011111",
  10892=>"000000000",
  10893=>"000000111",
  10894=>"100110000",
  10895=>"011110110",
  10896=>"101111110",
  10897=>"000000000",
  10898=>"000100000",
  10899=>"111001001",
  10900=>"111000000",
  10901=>"111111111",
  10902=>"000000111",
  10903=>"000000011",
  10904=>"000000000",
  10905=>"010011110",
  10906=>"111111111",
  10907=>"000000000",
  10908=>"111111111",
  10909=>"111000000",
  10910=>"111111111",
  10911=>"111111111",
  10912=>"100110000",
  10913=>"000001001",
  10914=>"000000000",
  10915=>"000000000",
  10916=>"000000000",
  10917=>"000010000",
  10918=>"000001111",
  10919=>"000000000",
  10920=>"111011111",
  10921=>"111111111",
  10922=>"000000000",
  10923=>"111110000",
  10924=>"100000100",
  10925=>"001001100",
  10926=>"000100111",
  10927=>"111011111",
  10928=>"111111100",
  10929=>"001100100",
  10930=>"100000000",
  10931=>"111001111",
  10932=>"001101101",
  10933=>"011111111",
  10934=>"000000000",
  10935=>"000011111",
  10936=>"111110101",
  10937=>"000000011",
  10938=>"000000000",
  10939=>"010010000",
  10940=>"111101111",
  10941=>"111010000",
  10942=>"010110110",
  10943=>"000000110",
  10944=>"000000000",
  10945=>"000000111",
  10946=>"000000000",
  10947=>"111111111",
  10948=>"111111000",
  10949=>"000000000",
  10950=>"110000100",
  10951=>"111111111",
  10952=>"111111111",
  10953=>"001001000",
  10954=>"110000000",
  10955=>"000010011",
  10956=>"000100111",
  10957=>"000000000",
  10958=>"111111111",
  10959=>"001001000",
  10960=>"000000000",
  10961=>"001001000",
  10962=>"111111111",
  10963=>"000000000",
  10964=>"101001000",
  10965=>"000011111",
  10966=>"000000000",
  10967=>"000110111",
  10968=>"111111111",
  10969=>"000000110",
  10970=>"000000000",
  10971=>"100000000",
  10972=>"000000000",
  10973=>"000010000",
  10974=>"000000000",
  10975=>"000000000",
  10976=>"000000000",
  10977=>"000000000",
  10978=>"111111100",
  10979=>"100100101",
  10980=>"110110000",
  10981=>"000000000",
  10982=>"011011011",
  10983=>"010000000",
  10984=>"001001000",
  10985=>"000000000",
  10986=>"001110110",
  10987=>"000000101",
  10988=>"000000000",
  10989=>"000000000",
  10990=>"001111111",
  10991=>"111000111",
  10992=>"100111110",
  10993=>"000010011",
  10994=>"010000110",
  10995=>"001011111",
  10996=>"011111111",
  10997=>"000000100",
  10998=>"001110000",
  10999=>"100001001",
  11000=>"111111111",
  11001=>"111111111",
  11002=>"000000000",
  11003=>"111111111",
  11004=>"001101001",
  11005=>"111011111",
  11006=>"000100000",
  11007=>"111111101",
  11008=>"000000000",
  11009=>"110111100",
  11010=>"000111111",
  11011=>"000000000",
  11012=>"111000000",
  11013=>"001000000",
  11014=>"011000000",
  11015=>"000111111",
  11016=>"000000000",
  11017=>"000000000",
  11018=>"000000000",
  11019=>"111110110",
  11020=>"101001000",
  11021=>"111011001",
  11022=>"000000111",
  11023=>"001000000",
  11024=>"000010110",
  11025=>"000000101",
  11026=>"111000000",
  11027=>"100001001",
  11028=>"000000001",
  11029=>"000000000",
  11030=>"111111111",
  11031=>"110000000",
  11032=>"000000100",
  11033=>"001010011",
  11034=>"000111111",
  11035=>"000000000",
  11036=>"101100100",
  11037=>"000000000",
  11038=>"000000000",
  11039=>"000000000",
  11040=>"000000001",
  11041=>"100000001",
  11042=>"111111000",
  11043=>"110110111",
  11044=>"001001100",
  11045=>"000000000",
  11046=>"111101101",
  11047=>"000000001",
  11048=>"000000000",
  11049=>"000000000",
  11050=>"000000000",
  11051=>"111011111",
  11052=>"000000000",
  11053=>"000100100",
  11054=>"111111010",
  11055=>"110111111",
  11056=>"111111111",
  11057=>"000000000",
  11058=>"111111111",
  11059=>"000000000",
  11060=>"011111111",
  11061=>"111111111",
  11062=>"000000000",
  11063=>"000000011",
  11064=>"000000000",
  11065=>"000001000",
  11066=>"111111110",
  11067=>"000000000",
  11068=>"111111111",
  11069=>"000001111",
  11070=>"111101001",
  11071=>"111110111",
  11072=>"000000100",
  11073=>"000000001",
  11074=>"110100111",
  11075=>"011000000",
  11076=>"111111111",
  11077=>"000000000",
  11078=>"000000100",
  11079=>"000000111",
  11080=>"111000100",
  11081=>"000000000",
  11082=>"100000000",
  11083=>"000000110",
  11084=>"000000000",
  11085=>"010000000",
  11086=>"110111111",
  11087=>"111001101",
  11088=>"000001010",
  11089=>"111111111",
  11090=>"100111110",
  11091=>"111111111",
  11092=>"000100000",
  11093=>"011011011",
  11094=>"110100000",
  11095=>"000000000",
  11096=>"011100000",
  11097=>"111111000",
  11098=>"111110000",
  11099=>"111111111",
  11100=>"000000111",
  11101=>"111000000",
  11102=>"000000000",
  11103=>"000000111",
  11104=>"111111111",
  11105=>"110100100",
  11106=>"111111111",
  11107=>"111111111",
  11108=>"001001000",
  11109=>"000000000",
  11110=>"011010111",
  11111=>"000000000",
  11112=>"001001011",
  11113=>"001011111",
  11114=>"000000000",
  11115=>"101101110",
  11116=>"100000000",
  11117=>"000000000",
  11118=>"000000000",
  11119=>"000000000",
  11120=>"000000000",
  11121=>"000000000",
  11122=>"100100100",
  11123=>"000100111",
  11124=>"000000000",
  11125=>"111111111",
  11126=>"111011111",
  11127=>"110110000",
  11128=>"101100100",
  11129=>"000000000",
  11130=>"000000001",
  11131=>"001111100",
  11132=>"000000011",
  11133=>"000000001",
  11134=>"111000000",
  11135=>"110111111",
  11136=>"000000000",
  11137=>"000010000",
  11138=>"000000000",
  11139=>"000000000",
  11140=>"111100100",
  11141=>"000000000",
  11142=>"001111101",
  11143=>"111111111",
  11144=>"000000000",
  11145=>"100110010",
  11146=>"000000000",
  11147=>"000000000",
  11148=>"111111111",
  11149=>"111111111",
  11150=>"110010111",
  11151=>"010111111",
  11152=>"000000000",
  11153=>"011111111",
  11154=>"000000000",
  11155=>"111111110",
  11156=>"000000000",
  11157=>"000000000",
  11158=>"111111111",
  11159=>"000000000",
  11160=>"001000000",
  11161=>"000000000",
  11162=>"010000000",
  11163=>"111000000",
  11164=>"000000000",
  11165=>"111111111",
  11166=>"001000000",
  11167=>"000000100",
  11168=>"100111111",
  11169=>"111111111",
  11170=>"011000000",
  11171=>"011001000",
  11172=>"110110110",
  11173=>"111111111",
  11174=>"111111011",
  11175=>"000000100",
  11176=>"111111111",
  11177=>"110100100",
  11178=>"000000010",
  11179=>"000001000",
  11180=>"000000000",
  11181=>"110110000",
  11182=>"000000000",
  11183=>"011011111",
  11184=>"111111111",
  11185=>"100011111",
  11186=>"011011100",
  11187=>"000000000",
  11188=>"001111111",
  11189=>"111111011",
  11190=>"110110111",
  11191=>"101111111",
  11192=>"011011110",
  11193=>"000000000",
  11194=>"111111010",
  11195=>"011011011",
  11196=>"000000110",
  11197=>"000000000",
  11198=>"000000000",
  11199=>"011111111",
  11200=>"111111111",
  11201=>"100101111",
  11202=>"001111111",
  11203=>"111111011",
  11204=>"111011100",
  11205=>"001111111",
  11206=>"000111110",
  11207=>"000000000",
  11208=>"011000100",
  11209=>"100111111",
  11210=>"000000111",
  11211=>"100000111",
  11212=>"000000000",
  11213=>"111111111",
  11214=>"100111111",
  11215=>"010000000",
  11216=>"100100111",
  11217=>"110101101",
  11218=>"111111100",
  11219=>"111111111",
  11220=>"100110111",
  11221=>"111111111",
  11222=>"000000000",
  11223=>"011011001",
  11224=>"110111111",
  11225=>"111111111",
  11226=>"111111011",
  11227=>"111111001",
  11228=>"011011010",
  11229=>"111011000",
  11230=>"111111111",
  11231=>"001000000",
  11232=>"100000010",
  11233=>"000000000",
  11234=>"111111111",
  11235=>"111111111",
  11236=>"111000111",
  11237=>"000000000",
  11238=>"000000000",
  11239=>"110111100",
  11240=>"111000000",
  11241=>"111110000",
  11242=>"000000000",
  11243=>"000000011",
  11244=>"000000000",
  11245=>"110010000",
  11246=>"100100100",
  11247=>"001000100",
  11248=>"000000000",
  11249=>"111111011",
  11250=>"111111111",
  11251=>"000000000",
  11252=>"000000000",
  11253=>"110110100",
  11254=>"101111111",
  11255=>"011010101",
  11256=>"000000011",
  11257=>"111111111",
  11258=>"111110101",
  11259=>"000000111",
  11260=>"111000000",
  11261=>"001111111",
  11262=>"110000000",
  11263=>"000000000",
  11264=>"000000100",
  11265=>"000000000",
  11266=>"111111111",
  11267=>"010111110",
  11268=>"000000101",
  11269=>"110011011",
  11270=>"101001101",
  11271=>"111111111",
  11272=>"010000000",
  11273=>"000000000",
  11274=>"000000000",
  11275=>"111110111",
  11276=>"100110110",
  11277=>"100000000",
  11278=>"100001001",
  11279=>"111000000",
  11280=>"000000110",
  11281=>"000111111",
  11282=>"111111101",
  11283=>"011000001",
  11284=>"000000100",
  11285=>"001000001",
  11286=>"001010000",
  11287=>"111111111",
  11288=>"110110110",
  11289=>"001000000",
  11290=>"111111111",
  11291=>"111001011",
  11292=>"111101111",
  11293=>"111110111",
  11294=>"111011001",
  11295=>"000000000",
  11296=>"111000000",
  11297=>"000000110",
  11298=>"110110100",
  11299=>"000000000",
  11300=>"110000000",
  11301=>"111110101",
  11302=>"111111000",
  11303=>"100000100",
  11304=>"101111111",
  11305=>"101000000",
  11306=>"000000001",
  11307=>"011001000",
  11308=>"011011011",
  11309=>"000000000",
  11310=>"101001000",
  11311=>"001001000",
  11312=>"100100000",
  11313=>"000000001",
  11314=>"000000000",
  11315=>"000000000",
  11316=>"100100111",
  11317=>"100111111",
  11318=>"001101101",
  11319=>"000000100",
  11320=>"000000000",
  11321=>"111110101",
  11322=>"000000001",
  11323=>"010000000",
  11324=>"111101111",
  11325=>"000000000",
  11326=>"000000000",
  11327=>"001000001",
  11328=>"011011010",
  11329=>"001001000",
  11330=>"000000000",
  11331=>"000000000",
  11332=>"000010110",
  11333=>"110010000",
  11334=>"110000000",
  11335=>"111111111",
  11336=>"111111011",
  11337=>"001000001",
  11338=>"000000001",
  11339=>"000001001",
  11340=>"110110010",
  11341=>"000000000",
  11342=>"000100000",
  11343=>"001001101",
  11344=>"000000000",
  11345=>"111011000",
  11346=>"111101111",
  11347=>"000000001",
  11348=>"000000101",
  11349=>"111001110",
  11350=>"111111111",
  11351=>"110110010",
  11352=>"000000011",
  11353=>"101101101",
  11354=>"111101111",
  11355=>"000000000",
  11356=>"000000001",
  11357=>"111101111",
  11358=>"111000101",
  11359=>"111111000",
  11360=>"111000100",
  11361=>"110111011",
  11362=>"001111111",
  11363=>"001001001",
  11364=>"111110010",
  11365=>"000000000",
  11366=>"111111000",
  11367=>"000001010",
  11368=>"111111111",
  11369=>"001111111",
  11370=>"110010110",
  11371=>"000000000",
  11372=>"001001011",
  11373=>"111101111",
  11374=>"110110111",
  11375=>"111111110",
  11376=>"111111111",
  11377=>"000001111",
  11378=>"100111111",
  11379=>"110111111",
  11380=>"000000000",
  11381=>"110110111",
  11382=>"111111111",
  11383=>"001001001",
  11384=>"000000010",
  11385=>"010111111",
  11386=>"000000000",
  11387=>"000000000",
  11388=>"111110100",
  11389=>"111111111",
  11390=>"000111100",
  11391=>"010000001",
  11392=>"000000000",
  11393=>"000000001",
  11394=>"000000111",
  11395=>"001001001",
  11396=>"101011000",
  11397=>"000110100",
  11398=>"110110100",
  11399=>"111011010",
  11400=>"111001001",
  11401=>"110110000",
  11402=>"000000000",
  11403=>"111111111",
  11404=>"111011111",
  11405=>"000000000",
  11406=>"111111101",
  11407=>"110110110",
  11408=>"000111110",
  11409=>"000000000",
  11410=>"011011111",
  11411=>"011111111",
  11412=>"000000111",
  11413=>"011010000",
  11414=>"000001101",
  11415=>"100111110",
  11416=>"001000001",
  11417=>"111111111",
  11418=>"111111010",
  11419=>"101000001",
  11420=>"000100111",
  11421=>"111111000",
  11422=>"111111000",
  11423=>"111111010",
  11424=>"011000000",
  11425=>"000111111",
  11426=>"010011000",
  11427=>"000000000",
  11428=>"001001111",
  11429=>"101000000",
  11430=>"111101111",
  11431=>"011010000",
  11432=>"101001101",
  11433=>"001000000",
  11434=>"101101101",
  11435=>"011010011",
  11436=>"110111111",
  11437=>"101000001",
  11438=>"000001000",
  11439=>"000000101",
  11440=>"011010000",
  11441=>"100000000",
  11442=>"110111111",
  11443=>"000000000",
  11444=>"111111111",
  11445=>"111001001",
  11446=>"000000100",
  11447=>"111111111",
  11448=>"111111111",
  11449=>"000000000",
  11450=>"001000000",
  11451=>"101001000",
  11452=>"111111100",
  11453=>"001001101",
  11454=>"001000000",
  11455=>"000010110",
  11456=>"111111111",
  11457=>"111111111",
  11458=>"111101100",
  11459=>"000101100",
  11460=>"111100111",
  11461=>"111001001",
  11462=>"111011011",
  11463=>"111111011",
  11464=>"111010000",
  11465=>"110111111",
  11466=>"000000000",
  11467=>"111111111",
  11468=>"100101111",
  11469=>"000000000",
  11470=>"111111111",
  11471=>"111111111",
  11472=>"111111011",
  11473=>"001111111",
  11474=>"000000110",
  11475=>"111101001",
  11476=>"110000000",
  11477=>"110110000",
  11478=>"111111111",
  11479=>"111001000",
  11480=>"000111111",
  11481=>"100111111",
  11482=>"101000000",
  11483=>"101001001",
  11484=>"000000000",
  11485=>"111000001",
  11486=>"000000000",
  11487=>"000000001",
  11488=>"111000000",
  11489=>"000000000",
  11490=>"011111111",
  11491=>"111001111",
  11492=>"000000111",
  11493=>"101001001",
  11494=>"000000101",
  11495=>"101000100",
  11496=>"010010010",
  11497=>"101000000",
  11498=>"100111111",
  11499=>"110111000",
  11500=>"100100100",
  11501=>"000000000",
  11502=>"000000111",
  11503=>"111011000",
  11504=>"111111111",
  11505=>"111111111",
  11506=>"001000001",
  11507=>"100001001",
  11508=>"001001111",
  11509=>"111111000",
  11510=>"000001011",
  11511=>"110100000",
  11512=>"001101110",
  11513=>"000011011",
  11514=>"001000000",
  11515=>"000000000",
  11516=>"111101001",
  11517=>"101001100",
  11518=>"000010000",
  11519=>"001001111",
  11520=>"000000001",
  11521=>"001001111",
  11522=>"001001111",
  11523=>"000000000",
  11524=>"101000000",
  11525=>"000101111",
  11526=>"101101111",
  11527=>"110010000",
  11528=>"000100000",
  11529=>"101000101",
  11530=>"111101000",
  11531=>"000000111",
  11532=>"101000101",
  11533=>"011000000",
  11534=>"111111111",
  11535=>"111000110",
  11536=>"011111100",
  11537=>"000100111",
  11538=>"101000101",
  11539=>"000000010",
  11540=>"100111111",
  11541=>"111000000",
  11542=>"001101111",
  11543=>"001111001",
  11544=>"111111011",
  11545=>"000000111",
  11546=>"111111010",
  11547=>"110110110",
  11548=>"000000100",
  11549=>"001000000",
  11550=>"000000000",
  11551=>"110100000",
  11552=>"010111001",
  11553=>"100111111",
  11554=>"111111111",
  11555=>"101001000",
  11556=>"111000001",
  11557=>"000001001",
  11558=>"000000000",
  11559=>"111100001",
  11560=>"111111001",
  11561=>"111111010",
  11562=>"111000000",
  11563=>"000000111",
  11564=>"110100000",
  11565=>"100000000",
  11566=>"000000000",
  11567=>"000000000",
  11568=>"111111110",
  11569=>"000010000",
  11570=>"111101101",
  11571=>"111001000",
  11572=>"010000010",
  11573=>"111000000",
  11574=>"111111111",
  11575=>"111101001",
  11576=>"001001101",
  11577=>"001000000",
  11578=>"000100101",
  11579=>"000000111",
  11580=>"000000000",
  11581=>"000111110",
  11582=>"000000100",
  11583=>"110100000",
  11584=>"001101111",
  11585=>"110111110",
  11586=>"111011011",
  11587=>"001000000",
  11588=>"001000000",
  11589=>"001111000",
  11590=>"011111001",
  11591=>"000000000",
  11592=>"001000000",
  11593=>"111001011",
  11594=>"111000000",
  11595=>"111001011",
  11596=>"110110110",
  11597=>"111111110",
  11598=>"100000001",
  11599=>"010110110",
  11600=>"000000100",
  11601=>"001000101",
  11602=>"111001111",
  11603=>"000000111",
  11604=>"000000011",
  11605=>"011011011",
  11606=>"111111111",
  11607=>"110111110",
  11608=>"000000101",
  11609=>"000000000",
  11610=>"111010000",
  11611=>"100000000",
  11612=>"111111111",
  11613=>"110111110",
  11614=>"101001101",
  11615=>"100110111",
  11616=>"101111111",
  11617=>"111111111",
  11618=>"100100111",
  11619=>"101000000",
  11620=>"000000001",
  11621=>"100000000",
  11622=>"000000000",
  11623=>"110110110",
  11624=>"110100100",
  11625=>"101101111",
  11626=>"000000001",
  11627=>"010110111",
  11628=>"110110111",
  11629=>"000001001",
  11630=>"001000001",
  11631=>"000000000",
  11632=>"111000000",
  11633=>"000000010",
  11634=>"111000000",
  11635=>"111111000",
  11636=>"010111111",
  11637=>"110111111",
  11638=>"000000100",
  11639=>"111111111",
  11640=>"101000000",
  11641=>"111000110",
  11642=>"000000010",
  11643=>"000000000",
  11644=>"110110110",
  11645=>"111000000",
  11646=>"111111111",
  11647=>"000000000",
  11648=>"000000000",
  11649=>"110010000",
  11650=>"110011011",
  11651=>"000000000",
  11652=>"111000100",
  11653=>"000111000",
  11654=>"111111110",
  11655=>"000000000",
  11656=>"000001101",
  11657=>"000000100",
  11658=>"111011111",
  11659=>"100100100",
  11660=>"111000000",
  11661=>"111111111",
  11662=>"000000000",
  11663=>"000101101",
  11664=>"000000000",
  11665=>"111111111",
  11666=>"111011111",
  11667=>"000100011",
  11668=>"001000000",
  11669=>"000000000",
  11670=>"110111111",
  11671=>"101111111",
  11672=>"001000110",
  11673=>"111010000",
  11674=>"000000001",
  11675=>"101101101",
  11676=>"111111010",
  11677=>"000000111",
  11678=>"111111111",
  11679=>"111010000",
  11680=>"000111011",
  11681=>"000011111",
  11682=>"101000001",
  11683=>"111110110",
  11684=>"101101101",
  11685=>"000001001",
  11686=>"000001001",
  11687=>"010110111",
  11688=>"100000000",
  11689=>"001000000",
  11690=>"000000001",
  11691=>"111001000",
  11692=>"111100000",
  11693=>"111110100",
  11694=>"000111101",
  11695=>"000000000",
  11696=>"000000001",
  11697=>"111000001",
  11698=>"101100100",
  11699=>"000000000",
  11700=>"001001001",
  11701=>"111110110",
  11702=>"000000101",
  11703=>"000100110",
  11704=>"111011111",
  11705=>"010010011",
  11706=>"111111010",
  11707=>"000000000",
  11708=>"111111111",
  11709=>"111111110",
  11710=>"101000000",
  11711=>"011110111",
  11712=>"111011000",
  11713=>"000000111",
  11714=>"011001001",
  11715=>"111000000",
  11716=>"101101001",
  11717=>"111111000",
  11718=>"001001001",
  11719=>"001000110",
  11720=>"001001000",
  11721=>"000000000",
  11722=>"101001001",
  11723=>"110010000",
  11724=>"001011111",
  11725=>"111111111",
  11726=>"110110010",
  11727=>"010111111",
  11728=>"011111010",
  11729=>"001001011",
  11730=>"000000000",
  11731=>"111011111",
  11732=>"111000000",
  11733=>"111110000",
  11734=>"111111000",
  11735=>"011011011",
  11736=>"000000000",
  11737=>"000000000",
  11738=>"001000000",
  11739=>"111111111",
  11740=>"111111111",
  11741=>"111101101",
  11742=>"011111111",
  11743=>"000000001",
  11744=>"111000000",
  11745=>"000011011",
  11746=>"111100111",
  11747=>"001000100",
  11748=>"111000110",
  11749=>"000000001",
  11750=>"101111111",
  11751=>"010010000",
  11752=>"100000000",
  11753=>"000001111",
  11754=>"111111111",
  11755=>"010111011",
  11756=>"111111101",
  11757=>"110000100",
  11758=>"001001000",
  11759=>"101111111",
  11760=>"000000101",
  11761=>"110110000",
  11762=>"010011010",
  11763=>"000001111",
  11764=>"000001111",
  11765=>"100000000",
  11766=>"110110111",
  11767=>"101000000",
  11768=>"111111111",
  11769=>"011001001",
  11770=>"110111001",
  11771=>"001000000",
  11772=>"111111011",
  11773=>"110110110",
  11774=>"100100100",
  11775=>"111111110",
  11776=>"010110110",
  11777=>"000000000",
  11778=>"111111111",
  11779=>"111111111",
  11780=>"000010000",
  11781=>"111111111",
  11782=>"001000100",
  11783=>"000000000",
  11784=>"111011111",
  11785=>"100111111",
  11786=>"110111111",
  11787=>"000111011",
  11788=>"111011000",
  11789=>"001101111",
  11790=>"000000000",
  11791=>"110111111",
  11792=>"000000000",
  11793=>"111101101",
  11794=>"111111111",
  11795=>"011011011",
  11796=>"000000110",
  11797=>"101100111",
  11798=>"001101111",
  11799=>"111111110",
  11800=>"111110111",
  11801=>"011011011",
  11802=>"101111111",
  11803=>"111111111",
  11804=>"111101111",
  11805=>"000010000",
  11806=>"001001001",
  11807=>"000000000",
  11808=>"111111111",
  11809=>"011111110",
  11810=>"001000111",
  11811=>"000000100",
  11812=>"111111111",
  11813=>"000111111",
  11814=>"111111011",
  11815=>"001111011",
  11816=>"000000011",
  11817=>"101000000",
  11818=>"100000011",
  11819=>"000000111",
  11820=>"000000100",
  11821=>"110100000",
  11822=>"001001000",
  11823=>"000111000",
  11824=>"110010010",
  11825=>"000000000",
  11826=>"000000000",
  11827=>"000000000",
  11828=>"001000111",
  11829=>"110101100",
  11830=>"000000000",
  11831=>"010011001",
  11832=>"010110110",
  11833=>"000000000",
  11834=>"000101111",
  11835=>"111000000",
  11836=>"111111100",
  11837=>"000000000",
  11838=>"000000011",
  11839=>"000000111",
  11840=>"000000000",
  11841=>"011000000",
  11842=>"111111111",
  11843=>"100110111",
  11844=>"000000000",
  11845=>"010011011",
  11846=>"000000111",
  11847=>"111111111",
  11848=>"111000111",
  11849=>"000000000",
  11850=>"111111111",
  11851=>"000111111",
  11852=>"110111111",
  11853=>"111010000",
  11854=>"010000000",
  11855=>"100111111",
  11856=>"001001000",
  11857=>"111001000",
  11858=>"010111111",
  11859=>"111111000",
  11860=>"000110010",
  11861=>"011111111",
  11862=>"000010011",
  11863=>"101111111",
  11864=>"111111111",
  11865=>"100000100",
  11866=>"110000111",
  11867=>"001111110",
  11868=>"110000000",
  11869=>"111111111",
  11870=>"000000000",
  11871=>"111111110",
  11872=>"111111111",
  11873=>"111011000",
  11874=>"001001000",
  11875=>"000000000",
  11876=>"000000000",
  11877=>"110110111",
  11878=>"111111110",
  11879=>"111111110",
  11880=>"010110110",
  11881=>"000000000",
  11882=>"000000111",
  11883=>"000000000",
  11884=>"000110111",
  11885=>"000100111",
  11886=>"111001000",
  11887=>"001000000",
  11888=>"000000000",
  11889=>"110010010",
  11890=>"101100100",
  11891=>"001001000",
  11892=>"000000000",
  11893=>"000001111",
  11894=>"000000111",
  11895=>"111111111",
  11896=>"101111110",
  11897=>"000000000",
  11898=>"111111000",
  11899=>"111111111",
  11900=>"100100110",
  11901=>"110111111",
  11902=>"111111011",
  11903=>"000011010",
  11904=>"111111111",
  11905=>"000001000",
  11906=>"001000000",
  11907=>"000000000",
  11908=>"000111101",
  11909=>"110000101",
  11910=>"110111111",
  11911=>"111111011",
  11912=>"000000000",
  11913=>"001101111",
  11914=>"000000000",
  11915=>"111011110",
  11916=>"000000000",
  11917=>"001001000",
  11918=>"111111111",
  11919=>"000000111",
  11920=>"000000111",
  11921=>"000000000",
  11922=>"111111000",
  11923=>"000000111",
  11924=>"000000000",
  11925=>"011011010",
  11926=>"000001111",
  11927=>"000000000",
  11928=>"111111100",
  11929=>"010010010",
  11930=>"111111111",
  11931=>"111111111",
  11932=>"000001111",
  11933=>"111011111",
  11934=>"010000011",
  11935=>"000000000",
  11936=>"111110111",
  11937=>"111100100",
  11938=>"110010111",
  11939=>"111111110",
  11940=>"111001001",
  11941=>"010010000",
  11942=>"111111111",
  11943=>"011111011",
  11944=>"000000000",
  11945=>"111011010",
  11946=>"111111111",
  11947=>"111111111",
  11948=>"111111000",
  11949=>"000110111",
  11950=>"110110111",
  11951=>"111110100",
  11952=>"000000000",
  11953=>"111111111",
  11954=>"111111111",
  11955=>"011100111",
  11956=>"011111111",
  11957=>"111111110",
  11958=>"111111111",
  11959=>"110110111",
  11960=>"000001001",
  11961=>"000000000",
  11962=>"111010000",
  11963=>"111111111",
  11964=>"111111000",
  11965=>"001111111",
  11966=>"111111111",
  11967=>"000000000",
  11968=>"001000000",
  11969=>"111111010",
  11970=>"111111111",
  11971=>"000000000",
  11972=>"111111111",
  11973=>"111111111",
  11974=>"111000000",
  11975=>"000110110",
  11976=>"001111111",
  11977=>"001000101",
  11978=>"000000000",
  11979=>"111101101",
  11980=>"001000100",
  11981=>"000010100",
  11982=>"111111111",
  11983=>"000000000",
  11984=>"111111001",
  11985=>"111111111",
  11986=>"101111111",
  11987=>"111000000",
  11988=>"110111111",
  11989=>"110110111",
  11990=>"111101100",
  11991=>"000000000",
  11992=>"111111111",
  11993=>"000011111",
  11994=>"000000000",
  11995=>"000010000",
  11996=>"111001000",
  11997=>"000000000",
  11998=>"000000000",
  11999=>"000000000",
  12000=>"000010000",
  12001=>"010000000",
  12002=>"111111111",
  12003=>"111111111",
  12004=>"111111111",
  12005=>"111111111",
  12006=>"000000001",
  12007=>"111101101",
  12008=>"111111111",
  12009=>"100010010",
  12010=>"000000001",
  12011=>"000000000",
  12012=>"011101111",
  12013=>"111111111",
  12014=>"000000000",
  12015=>"000000111",
  12016=>"111111011",
  12017=>"000000000",
  12018=>"010111111",
  12019=>"000000110",
  12020=>"000100111",
  12021=>"111111110",
  12022=>"000000000",
  12023=>"010010000",
  12024=>"111111101",
  12025=>"000000001",
  12026=>"111111111",
  12027=>"011111111",
  12028=>"000100100",
  12029=>"000000000",
  12030=>"010111111",
  12031=>"111111100",
  12032=>"111111110",
  12033=>"000100100",
  12034=>"010010000",
  12035=>"111111000",
  12036=>"111111111",
  12037=>"000000100",
  12038=>"000111111",
  12039=>"001111111",
  12040=>"010000000",
  12041=>"000000000",
  12042=>"001000100",
  12043=>"000101111",
  12044=>"001001111",
  12045=>"000000000",
  12046=>"000000010",
  12047=>"000000000",
  12048=>"111111111",
  12049=>"100100100",
  12050=>"001000101",
  12051=>"001111111",
  12052=>"000000110",
  12053=>"111111100",
  12054=>"000000111",
  12055=>"111110100",
  12056=>"111111111",
  12057=>"111111111",
  12058=>"111111111",
  12059=>"011011111",
  12060=>"110111100",
  12061=>"111011001",
  12062=>"000000111",
  12063=>"111000100",
  12064=>"000000000",
  12065=>"000000111",
  12066=>"111111111",
  12067=>"000100110",
  12068=>"111100000",
  12069=>"110110110",
  12070=>"000000110",
  12071=>"000000010",
  12072=>"000000110",
  12073=>"000000000",
  12074=>"111111111",
  12075=>"100101111",
  12076=>"111101100",
  12077=>"110111111",
  12078=>"111111111",
  12079=>"000000000",
  12080=>"001001001",
  12081=>"000000000",
  12082=>"000001000",
  12083=>"000000000",
  12084=>"111111001",
  12085=>"001001011",
  12086=>"000001011",
  12087=>"111011111",
  12088=>"001001001",
  12089=>"000000111",
  12090=>"001111111",
  12091=>"010010000",
  12092=>"111111111",
  12093=>"000001101",
  12094=>"000000010",
  12095=>"111111111",
  12096=>"000000000",
  12097=>"000000000",
  12098=>"000111111",
  12099=>"000000110",
  12100=>"000000000",
  12101=>"000010111",
  12102=>"111111111",
  12103=>"111111111",
  12104=>"111100101",
  12105=>"000000111",
  12106=>"000000111",
  12107=>"100110100",
  12108=>"100000111",
  12109=>"111011000",
  12110=>"000011111",
  12111=>"010011011",
  12112=>"111111111",
  12113=>"111111110",
  12114=>"001111111",
  12115=>"000000000",
  12116=>"101000001",
  12117=>"011011011",
  12118=>"100000000",
  12119=>"111111111",
  12120=>"000111111",
  12121=>"111111111",
  12122=>"000000000",
  12123=>"111111111",
  12124=>"000000000",
  12125=>"100110111",
  12126=>"001001001",
  12127=>"000000000",
  12128=>"000000000",
  12129=>"110111111",
  12130=>"100100000",
  12131=>"000100000",
  12132=>"111111111",
  12133=>"111111000",
  12134=>"111111111",
  12135=>"000000000",
  12136=>"111100001",
  12137=>"001001001",
  12138=>"111001111",
  12139=>"111111110",
  12140=>"010111111",
  12141=>"110110110",
  12142=>"111111111",
  12143=>"100101100",
  12144=>"001000111",
  12145=>"000000000",
  12146=>"110101101",
  12147=>"100111111",
  12148=>"000100100",
  12149=>"111110111",
  12150=>"011011000",
  12151=>"101111010",
  12152=>"111111111",
  12153=>"011011001",
  12154=>"000000000",
  12155=>"000000111",
  12156=>"001000000",
  12157=>"111110111",
  12158=>"111111101",
  12159=>"100000100",
  12160=>"000111011",
  12161=>"100100000",
  12162=>"000000100",
  12163=>"000000000",
  12164=>"111111111",
  12165=>"111101000",
  12166=>"111111001",
  12167=>"111000000",
  12168=>"111111111",
  12169=>"100100100",
  12170=>"111111111",
  12171=>"111111111",
  12172=>"000000111",
  12173=>"011011001",
  12174=>"000010000",
  12175=>"000000000",
  12176=>"111011000",
  12177=>"111011100",
  12178=>"000000000",
  12179=>"111111110",
  12180=>"000110111",
  12181=>"011011000",
  12182=>"000000010",
  12183=>"000000000",
  12184=>"111111111",
  12185=>"001001001",
  12186=>"000100110",
  12187=>"010011000",
  12188=>"000000000",
  12189=>"000000111",
  12190=>"000000101",
  12191=>"111111011",
  12192=>"001011000",
  12193=>"100110111",
  12194=>"000000111",
  12195=>"011111111",
  12196=>"111110000",
  12197=>"111101101",
  12198=>"111111111",
  12199=>"000110111",
  12200=>"111101000",
  12201=>"001111010",
  12202=>"011111100",
  12203=>"000111111",
  12204=>"100111111",
  12205=>"111111111",
  12206=>"000000000",
  12207=>"001001000",
  12208=>"000000000",
  12209=>"111111111",
  12210=>"100100111",
  12211=>"000000000",
  12212=>"000000000",
  12213=>"111111111",
  12214=>"000111111",
  12215=>"111111111",
  12216=>"000000000",
  12217=>"110110111",
  12218=>"111111111",
  12219=>"111111111",
  12220=>"000000111",
  12221=>"111111111",
  12222=>"000101111",
  12223=>"000100100",
  12224=>"010111111",
  12225=>"111111111",
  12226=>"000000101",
  12227=>"000000100",
  12228=>"000000110",
  12229=>"010010000",
  12230=>"000000010",
  12231=>"000000011",
  12232=>"111000111",
  12233=>"110010011",
  12234=>"000000000",
  12235=>"100000000",
  12236=>"111111000",
  12237=>"001111000",
  12238=>"000000000",
  12239=>"010001001",
  12240=>"000010000",
  12241=>"000000111",
  12242=>"000000111",
  12243=>"111111011",
  12244=>"000000000",
  12245=>"111111111",
  12246=>"011010010",
  12247=>"111111100",
  12248=>"000100111",
  12249=>"000000000",
  12250=>"000000000",
  12251=>"000000110",
  12252=>"010000010",
  12253=>"000000001",
  12254=>"111111111",
  12255=>"010010011",
  12256=>"000000100",
  12257=>"000000001",
  12258=>"001101110",
  12259=>"000000000",
  12260=>"000000000",
  12261=>"001111111",
  12262=>"000100111",
  12263=>"110010010",
  12264=>"001101111",
  12265=>"000110011",
  12266=>"111111010",
  12267=>"000000000",
  12268=>"000000101",
  12269=>"011011001",
  12270=>"111111111",
  12271=>"000000000",
  12272=>"000000111",
  12273=>"000110110",
  12274=>"111111111",
  12275=>"000000000",
  12276=>"111111111",
  12277=>"111111111",
  12278=>"000000000",
  12279=>"000000000",
  12280=>"111111111",
  12281=>"110001001",
  12282=>"000000111",
  12283=>"000000000",
  12284=>"000000000",
  12285=>"000000000",
  12286=>"000100000",
  12287=>"001111111",
  12288=>"101111111",
  12289=>"000000000",
  12290=>"111000000",
  12291=>"110100000",
  12292=>"110111111",
  12293=>"111000001",
  12294=>"000000001",
  12295=>"111111111",
  12296=>"111010111",
  12297=>"111111000",
  12298=>"000000000",
  12299=>"111110110",
  12300=>"000000111",
  12301=>"000001001",
  12302=>"011000000",
  12303=>"000000000",
  12304=>"011001000",
  12305=>"111111111",
  12306=>"111111111",
  12307=>"111111111",
  12308=>"111111111",
  12309=>"000001000",
  12310=>"011111000",
  12311=>"111000000",
  12312=>"000000000",
  12313=>"111101111",
  12314=>"000000001",
  12315=>"000000000",
  12316=>"111111111",
  12317=>"000000000",
  12318=>"001000001",
  12319=>"111110111",
  12320=>"000000000",
  12321=>"111110111",
  12322=>"111111111",
  12323=>"000000000",
  12324=>"011111111",
  12325=>"111101000",
  12326=>"000000000",
  12327=>"000000000",
  12328=>"000000000",
  12329=>"000000000",
  12330=>"111111111",
  12331=>"110100000",
  12332=>"000110111",
  12333=>"111111111",
  12334=>"000000111",
  12335=>"010000000",
  12336=>"000001000",
  12337=>"000100101",
  12338=>"111110110",
  12339=>"000000000",
  12340=>"111111111",
  12341=>"011000000",
  12342=>"000000000",
  12343=>"010110100",
  12344=>"010000001",
  12345=>"000000000",
  12346=>"011111111",
  12347=>"001000000",
  12348=>"111111111",
  12349=>"111111000",
  12350=>"001011011",
  12351=>"111111111",
  12352=>"111111111",
  12353=>"010111111",
  12354=>"000000000",
  12355=>"000000010",
  12356=>"100110011",
  12357=>"000000000",
  12358=>"101000000",
  12359=>"100100000",
  12360=>"111111111",
  12361=>"100101111",
  12362=>"111110100",
  12363=>"001001111",
  12364=>"111101111",
  12365=>"000000000",
  12366=>"000000000",
  12367=>"000000000",
  12368=>"000000000",
  12369=>"111111111",
  12370=>"000000000",
  12371=>"000000000",
  12372=>"001000000",
  12373=>"111111101",
  12374=>"000000000",
  12375=>"000000000",
  12376=>"000000001",
  12377=>"111101111",
  12378=>"011000000",
  12379=>"000101111",
  12380=>"111111111",
  12381=>"000111000",
  12382=>"111111000",
  12383=>"110110111",
  12384=>"000111111",
  12385=>"111111111",
  12386=>"000000110",
  12387=>"100000110",
  12388=>"000000000",
  12389=>"011111111",
  12390=>"000000000",
  12391=>"111111111",
  12392=>"111111111",
  12393=>"111000000",
  12394=>"000000000",
  12395=>"110111010",
  12396=>"100000111",
  12397=>"000000011",
  12398=>"000000000",
  12399=>"111111111",
  12400=>"000000001",
  12401=>"000000001",
  12402=>"000000000",
  12403=>"000000001",
  12404=>"011000000",
  12405=>"111111111",
  12406=>"111111111",
  12407=>"000000100",
  12408=>"111111010",
  12409=>"111111001",
  12410=>"001000000",
  12411=>"111111111",
  12412=>"110110110",
  12413=>"000000000",
  12414=>"000001000",
  12415=>"001101111",
  12416=>"011000000",
  12417=>"000000000",
  12418=>"000000011",
  12419=>"000111111",
  12420=>"111111101",
  12421=>"001111111",
  12422=>"111111111",
  12423=>"000000000",
  12424=>"001000001",
  12425=>"111110000",
  12426=>"000000000",
  12427=>"000000100",
  12428=>"001011000",
  12429=>"011000000",
  12430=>"000000000",
  12431=>"000000000",
  12432=>"000101111",
  12433=>"000000001",
  12434=>"000001000",
  12435=>"000000000",
  12436=>"111101111",
  12437=>"000000001",
  12438=>"000011000",
  12439=>"000000000",
  12440=>"111011001",
  12441=>"110100001",
  12442=>"100000001",
  12443=>"111111111",
  12444=>"111111111",
  12445=>"101000001",
  12446=>"111111111",
  12447=>"001100000",
  12448=>"001001100",
  12449=>"000000000",
  12450=>"111111111",
  12451=>"010010000",
  12452=>"011001000",
  12453=>"110110110",
  12454=>"000010000",
  12455=>"001001001",
  12456=>"000110000",
  12457=>"111111011",
  12458=>"000000000",
  12459=>"111111111",
  12460=>"000000000",
  12461=>"111111110",
  12462=>"100101111",
  12463=>"011000001",
  12464=>"000110110",
  12465=>"111111110",
  12466=>"111111111",
  12467=>"000001000",
  12468=>"000000000",
  12469=>"111111000",
  12470=>"000000000",
  12471=>"000000000",
  12472=>"100000111",
  12473=>"111111000",
  12474=>"000000000",
  12475=>"001000000",
  12476=>"111010111",
  12477=>"101101001",
  12478=>"111110011",
  12479=>"000000000",
  12480=>"111111111",
  12481=>"000000000",
  12482=>"111111111",
  12483=>"000001000",
  12484=>"000000000",
  12485=>"011110010",
  12486=>"000000000",
  12487=>"000000000",
  12488=>"111111111",
  12489=>"111110111",
  12490=>"001111111",
  12491=>"000100111",
  12492=>"111111111",
  12493=>"101101001",
  12494=>"000000001",
  12495=>"000000000",
  12496=>"000000000",
  12497=>"000000111",
  12498=>"000001101",
  12499=>"110111111",
  12500=>"111111111",
  12501=>"100110111",
  12502=>"000000000",
  12503=>"000000000",
  12504=>"111111111",
  12505=>"110000101",
  12506=>"000000000",
  12507=>"111111111",
  12508=>"100000000",
  12509=>"000000111",
  12510=>"000011000",
  12511=>"111001000",
  12512=>"111000000",
  12513=>"000110000",
  12514=>"111111000",
  12515=>"001000000",
  12516=>"111111111",
  12517=>"000000000",
  12518=>"000000111",
  12519=>"000000000",
  12520=>"111111000",
  12521=>"111111111",
  12522=>"011000000",
  12523=>"111111100",
  12524=>"000000111",
  12525=>"000000000",
  12526=>"111100111",
  12527=>"000000000",
  12528=>"000110111",
  12529=>"111111100",
  12530=>"111000000",
  12531=>"111111001",
  12532=>"001001001",
  12533=>"011111111",
  12534=>"000000000",
  12535=>"111111111",
  12536=>"000000000",
  12537=>"111100000",
  12538=>"111110000",
  12539=>"000010111",
  12540=>"110110110",
  12541=>"111110110",
  12542=>"011011111",
  12543=>"000000000",
  12544=>"111111101",
  12545=>"111111101",
  12546=>"111111111",
  12547=>"001001111",
  12548=>"000000101",
  12549=>"111101000",
  12550=>"000001111",
  12551=>"000001001",
  12552=>"000000000",
  12553=>"111111111",
  12554=>"000000001",
  12555=>"111111001",
  12556=>"000000111",
  12557=>"111111111",
  12558=>"110000001",
  12559=>"011000000",
  12560=>"000000000",
  12561=>"001000001",
  12562=>"111111111",
  12563=>"010011000",
  12564=>"111000000",
  12565=>"111101001",
  12566=>"110111111",
  12567=>"111111111",
  12568=>"111101001",
  12569=>"000111111",
  12570=>"000000000",
  12571=>"000000000",
  12572=>"001001101",
  12573=>"000000011",
  12574=>"111111111",
  12575=>"000000111",
  12576=>"111111111",
  12577=>"000000001",
  12578=>"111001000",
  12579=>"000110000",
  12580=>"111111010",
  12581=>"100100101",
  12582=>"001011111",
  12583=>"111110110",
  12584=>"011001001",
  12585=>"111111111",
  12586=>"111110000",
  12587=>"000000000",
  12588=>"000111111",
  12589=>"000000000",
  12590=>"111000000",
  12591=>"000001000",
  12592=>"110110110",
  12593=>"000001000",
  12594=>"111111111",
  12595=>"000001000",
  12596=>"111000000",
  12597=>"110111111",
  12598=>"110001111",
  12599=>"100100111",
  12600=>"111010110",
  12601=>"001000000",
  12602=>"111111111",
  12603=>"111100000",
  12604=>"011001000",
  12605=>"000000011",
  12606=>"001001111",
  12607=>"000000000",
  12608=>"000000000",
  12609=>"000000000",
  12610=>"001001111",
  12611=>"000000000",
  12612=>"000001001",
  12613=>"111001111",
  12614=>"111111010",
  12615=>"111111001",
  12616=>"111111111",
  12617=>"000000000",
  12618=>"111111111",
  12619=>"100111111",
  12620=>"001111111",
  12621=>"111111001",
  12622=>"000000000",
  12623=>"010011011",
  12624=>"111111101",
  12625=>"000000000",
  12626=>"000000101",
  12627=>"110100110",
  12628=>"001000000",
  12629=>"011011011",
  12630=>"001111101",
  12631=>"000000000",
  12632=>"000011001",
  12633=>"000000000",
  12634=>"111011011",
  12635=>"100000000",
  12636=>"111111111",
  12637=>"000000111",
  12638=>"000100000",
  12639=>"111111110",
  12640=>"111100101",
  12641=>"111111111",
  12642=>"000100111",
  12643=>"111000000",
  12644=>"000001001",
  12645=>"000000000",
  12646=>"100000011",
  12647=>"111111011",
  12648=>"111111111",
  12649=>"011011000",
  12650=>"100110111",
  12651=>"011000000",
  12652=>"001100111",
  12653=>"111111001",
  12654=>"000000000",
  12655=>"000000000",
  12656=>"111111111",
  12657=>"111111111",
  12658=>"100100110",
  12659=>"111101001",
  12660=>"000000000",
  12661=>"000000000",
  12662=>"111101111",
  12663=>"100111000",
  12664=>"000000000",
  12665=>"111001011",
  12666=>"001000000",
  12667=>"011011000",
  12668=>"011001111",
  12669=>"110000111",
  12670=>"000000001",
  12671=>"001111111",
  12672=>"010000010",
  12673=>"111111111",
  12674=>"111000000",
  12675=>"110000000",
  12676=>"010000000",
  12677=>"000000000",
  12678=>"000000000",
  12679=>"000000000",
  12680=>"000000000",
  12681=>"000000000",
  12682=>"110111111",
  12683=>"000000000",
  12684=>"111111111",
  12685=>"101000111",
  12686=>"100000001",
  12687=>"000111111",
  12688=>"000000000",
  12689=>"010110111",
  12690=>"000011101",
  12691=>"100100001",
  12692=>"011001000",
  12693=>"000000000",
  12694=>"000011011",
  12695=>"111000000",
  12696=>"010011000",
  12697=>"000000000",
  12698=>"110000000",
  12699=>"111111111",
  12700=>"010111111",
  12701=>"010100000",
  12702=>"111111111",
  12703=>"000000000",
  12704=>"000000000",
  12705=>"000000000",
  12706=>"111111111",
  12707=>"000000000",
  12708=>"000111111",
  12709=>"001111010",
  12710=>"111111000",
  12711=>"110100110",
  12712=>"011000000",
  12713=>"100100000",
  12714=>"000000000",
  12715=>"111111001",
  12716=>"111001000",
  12717=>"000100000",
  12718=>"111111111",
  12719=>"111111111",
  12720=>"111001000",
  12721=>"111001000",
  12722=>"000000000",
  12723=>"000000110",
  12724=>"000001111",
  12725=>"000000000",
  12726=>"000111111",
  12727=>"111101111",
  12728=>"111111111",
  12729=>"111111110",
  12730=>"000000000",
  12731=>"111110100",
  12732=>"011111111",
  12733=>"100111111",
  12734=>"000000000",
  12735=>"001011011",
  12736=>"111111111",
  12737=>"101000000",
  12738=>"000111111",
  12739=>"111011000",
  12740=>"000000111",
  12741=>"000001001",
  12742=>"110000101",
  12743=>"000000000",
  12744=>"111011001",
  12745=>"110111111",
  12746=>"000101111",
  12747=>"000110111",
  12748=>"111111000",
  12749=>"111111111",
  12750=>"111101111",
  12751=>"000001111",
  12752=>"000111111",
  12753=>"011011111",
  12754=>"101000101",
  12755=>"001000000",
  12756=>"011111010",
  12757=>"000000001",
  12758=>"000000100",
  12759=>"000000100",
  12760=>"111101111",
  12761=>"111111111",
  12762=>"110110000",
  12763=>"001000000",
  12764=>"011101111",
  12765=>"000011011",
  12766=>"000000000",
  12767=>"000100000",
  12768=>"111111111",
  12769=>"000000111",
  12770=>"000000000",
  12771=>"000000000",
  12772=>"001101111",
  12773=>"111111111",
  12774=>"000110111",
  12775=>"010000000",
  12776=>"111111001",
  12777=>"011111011",
  12778=>"000000000",
  12779=>"111001001",
  12780=>"001111111",
  12781=>"111100001",
  12782=>"000000000",
  12783=>"111111110",
  12784=>"111100111",
  12785=>"001011101",
  12786=>"000000111",
  12787=>"111111111",
  12788=>"111111111",
  12789=>"100000000",
  12790=>"101001001",
  12791=>"001011011",
  12792=>"000001111",
  12793=>"001001101",
  12794=>"000000000",
  12795=>"111001000",
  12796=>"000000111",
  12797=>"000011111",
  12798=>"111110000",
  12799=>"111110001",
  12800=>"001001101",
  12801=>"000111111",
  12802=>"111111111",
  12803=>"000111111",
  12804=>"100100111",
  12805=>"000100110",
  12806=>"001000000",
  12807=>"000000100",
  12808=>"000000011",
  12809=>"111111111",
  12810=>"011000000",
  12811=>"100111111",
  12812=>"100100100",
  12813=>"101100100",
  12814=>"110111111",
  12815=>"011111100",
  12816=>"111111111",
  12817=>"000111100",
  12818=>"010011011",
  12819=>"000000000",
  12820=>"000000111",
  12821=>"111111111",
  12822=>"101111111",
  12823=>"100100110",
  12824=>"100100100",
  12825=>"000010000",
  12826=>"000000001",
  12827=>"000000000",
  12828=>"111111111",
  12829=>"111011001",
  12830=>"000000000",
  12831=>"000000000",
  12832=>"101000001",
  12833=>"011000000",
  12834=>"110100111",
  12835=>"111111111",
  12836=>"000000000",
  12837=>"111111111",
  12838=>"110110110",
  12839=>"001000000",
  12840=>"111101111",
  12841=>"111111111",
  12842=>"011111111",
  12843=>"111111110",
  12844=>"000000000",
  12845=>"111111111",
  12846=>"000000001",
  12847=>"000010000",
  12848=>"111000100",
  12849=>"111001000",
  12850=>"000000000",
  12851=>"000000000",
  12852=>"110011000",
  12853=>"001001001",
  12854=>"011000000",
  12855=>"111111111",
  12856=>"000000110",
  12857=>"000000100",
  12858=>"111111111",
  12859=>"111111111",
  12860=>"000000000",
  12861=>"111011000",
  12862=>"000000000",
  12863=>"000110110",
  12864=>"000000000",
  12865=>"000100000",
  12866=>"011000000",
  12867=>"001001000",
  12868=>"111000001",
  12869=>"111110111",
  12870=>"000000000",
  12871=>"000100000",
  12872=>"110000000",
  12873=>"110000000",
  12874=>"000000000",
  12875=>"000000000",
  12876=>"000000011",
  12877=>"011011000",
  12878=>"111000000",
  12879=>"000110110",
  12880=>"000000101",
  12881=>"111111111",
  12882=>"000000000",
  12883=>"101101111",
  12884=>"111111001",
  12885=>"111100000",
  12886=>"111111100",
  12887=>"111011001",
  12888=>"000000111",
  12889=>"111111010",
  12890=>"111100000",
  12891=>"011011011",
  12892=>"000000111",
  12893=>"110100111",
  12894=>"000001000",
  12895=>"111000000",
  12896=>"111111111",
  12897=>"111111111",
  12898=>"000000000",
  12899=>"000000000",
  12900=>"111111111",
  12901=>"111100100",
  12902=>"000000011",
  12903=>"110111100",
  12904=>"111111111",
  12905=>"000000000",
  12906=>"000000000",
  12907=>"000000000",
  12908=>"110110110",
  12909=>"000000000",
  12910=>"000000000",
  12911=>"000011111",
  12912=>"000000000",
  12913=>"000000101",
  12914=>"000110110",
  12915=>"111111111",
  12916=>"000010000",
  12917=>"010001111",
  12918=>"000111111",
  12919=>"000000000",
  12920=>"000001001",
  12921=>"000100100",
  12922=>"000010000",
  12923=>"111110100",
  12924=>"001001011",
  12925=>"111100111",
  12926=>"000100111",
  12927=>"000010011",
  12928=>"010111111",
  12929=>"111101111",
  12930=>"000000000",
  12931=>"000000000",
  12932=>"000000100",
  12933=>"000000111",
  12934=>"111111111",
  12935=>"000101111",
  12936=>"000000000",
  12937=>"000000011",
  12938=>"111111111",
  12939=>"111111000",
  12940=>"111101111",
  12941=>"000000000",
  12942=>"000000000",
  12943=>"111111111",
  12944=>"000110110",
  12945=>"000000000",
  12946=>"000000000",
  12947=>"000010110",
  12948=>"010010000",
  12949=>"001000100",
  12950=>"000001111",
  12951=>"000000001",
  12952=>"000000000",
  12953=>"111111111",
  12954=>"111001000",
  12955=>"111100000",
  12956=>"111111111",
  12957=>"000000100",
  12958=>"001000000",
  12959=>"000000111",
  12960=>"011010100",
  12961=>"111001001",
  12962=>"111111111",
  12963=>"000111111",
  12964=>"000010000",
  12965=>"000011111",
  12966=>"111000000",
  12967=>"100000000",
  12968=>"000000000",
  12969=>"000011010",
  12970=>"111111111",
  12971=>"111100100",
  12972=>"011111111",
  12973=>"000000000",
  12974=>"111001111",
  12975=>"100101111",
  12976=>"010111111",
  12977=>"001001000",
  12978=>"111111111",
  12979=>"101000101",
  12980=>"000000101",
  12981=>"010111111",
  12982=>"001001001",
  12983=>"111110110",
  12984=>"101100000",
  12985=>"111111111",
  12986=>"000110000",
  12987=>"011000001",
  12988=>"111111111",
  12989=>"111111111",
  12990=>"110111000",
  12991=>"000010110",
  12992=>"111101111",
  12993=>"110110001",
  12994=>"000000111",
  12995=>"000000000",
  12996=>"000111111",
  12997=>"000000001",
  12998=>"000000011",
  12999=>"111111111",
  13000=>"011111111",
  13001=>"100001101",
  13002=>"101000000",
  13003=>"000001001",
  13004=>"110000110",
  13005=>"110010000",
  13006=>"000000000",
  13007=>"000000000",
  13008=>"000000110",
  13009=>"011011011",
  13010=>"101101111",
  13011=>"000000000",
  13012=>"111111111",
  13013=>"110110111",
  13014=>"001111011",
  13015=>"111111000",
  13016=>"110000000",
  13017=>"000000100",
  13018=>"111111111",
  13019=>"000111111",
  13020=>"111111111",
  13021=>"000000000",
  13022=>"000100111",
  13023=>"000000000",
  13024=>"111111000",
  13025=>"010010000",
  13026=>"000000000",
  13027=>"011011000",
  13028=>"111111111",
  13029=>"100110100",
  13030=>"000011111",
  13031=>"111111111",
  13032=>"100100111",
  13033=>"000000000",
  13034=>"111111111",
  13035=>"001000100",
  13036=>"000000100",
  13037=>"000000000",
  13038=>"000000011",
  13039=>"000000000",
  13040=>"000000000",
  13041=>"000111111",
  13042=>"011011111",
  13043=>"000100000",
  13044=>"111111111",
  13045=>"010001001",
  13046=>"100000000",
  13047=>"111111111",
  13048=>"010010000",
  13049=>"111111111",
  13050=>"000000000",
  13051=>"110111111",
  13052=>"001001001",
  13053=>"000000000",
  13054=>"000000000",
  13055=>"000000000",
  13056=>"011111001",
  13057=>"000001001",
  13058=>"000000000",
  13059=>"111100000",
  13060=>"000001111",
  13061=>"000000001",
  13062=>"111111111",
  13063=>"111100111",
  13064=>"111111111",
  13065=>"000000000",
  13066=>"111111111",
  13067=>"111100001",
  13068=>"111000000",
  13069=>"111111000",
  13070=>"001000000",
  13071=>"000000000",
  13072=>"000000000",
  13073=>"000110111",
  13074=>"111111111",
  13075=>"000011011",
  13076=>"000000000",
  13077=>"010010000",
  13078=>"000000110",
  13079=>"111100000",
  13080=>"011011111",
  13081=>"111111100",
  13082=>"111111111",
  13083=>"000000010",
  13084=>"100000001",
  13085=>"000000001",
  13086=>"000000000",
  13087=>"111101111",
  13088=>"000000000",
  13089=>"000000101",
  13090=>"100000000",
  13091=>"111100101",
  13092=>"001001111",
  13093=>"000100000",
  13094=>"011001011",
  13095=>"110000111",
  13096=>"110111111",
  13097=>"111110000",
  13098=>"111111111",
  13099=>"111110100",
  13100=>"101100100",
  13101=>"011001011",
  13102=>"000000111",
  13103=>"111111010",
  13104=>"111010010",
  13105=>"111000000",
  13106=>"001000000",
  13107=>"000000000",
  13108=>"101000000",
  13109=>"000000001",
  13110=>"111101100",
  13111=>"000000000",
  13112=>"000000011",
  13113=>"000000111",
  13114=>"111111111",
  13115=>"000000111",
  13116=>"100000000",
  13117=>"111110111",
  13118=>"000111111",
  13119=>"000000000",
  13120=>"000000000",
  13121=>"111111111",
  13122=>"100100100",
  13123=>"111111111",
  13124=>"000000000",
  13125=>"000000000",
  13126=>"111111111",
  13127=>"110111111",
  13128=>"110110000",
  13129=>"000000011",
  13130=>"000000111",
  13131=>"110110000",
  13132=>"011111111",
  13133=>"101101111",
  13134=>"001001100",
  13135=>"000111110",
  13136=>"000000000",
  13137=>"001010000",
  13138=>"111100000",
  13139=>"000000000",
  13140=>"111111111",
  13141=>"011011011",
  13142=>"111000100",
  13143=>"111100100",
  13144=>"111111101",
  13145=>"000000100",
  13146=>"000000000",
  13147=>"000000000",
  13148=>"000111111",
  13149=>"111111111",
  13150=>"011110111",
  13151=>"011001101",
  13152=>"111111110",
  13153=>"111111111",
  13154=>"000000100",
  13155=>"101000001",
  13156=>"011111111",
  13157=>"000000100",
  13158=>"000000100",
  13159=>"110111111",
  13160=>"011011000",
  13161=>"010010010",
  13162=>"000000000",
  13163=>"111000010",
  13164=>"100000000",
  13165=>"011111000",
  13166=>"001001000",
  13167=>"000000111",
  13168=>"000000000",
  13169=>"111111000",
  13170=>"000000000",
  13171=>"100100111",
  13172=>"000110110",
  13173=>"111110111",
  13174=>"000100110",
  13175=>"111111000",
  13176=>"000001000",
  13177=>"000000000",
  13178=>"111000100",
  13179=>"000000000",
  13180=>"111111111",
  13181=>"000000000",
  13182=>"000100100",
  13183=>"000000000",
  13184=>"001000000",
  13185=>"000000000",
  13186=>"011011011",
  13187=>"101101110",
  13188=>"000000000",
  13189=>"110110001",
  13190=>"000000100",
  13191=>"010010010",
  13192=>"111111111",
  13193=>"111111000",
  13194=>"000000000",
  13195=>"000000000",
  13196=>"000000000",
  13197=>"001001001",
  13198=>"000001000",
  13199=>"100111111",
  13200=>"000000000",
  13201=>"111001000",
  13202=>"111000000",
  13203=>"001000000",
  13204=>"001001011",
  13205=>"011001001",
  13206=>"111101111",
  13207=>"000000000",
  13208=>"011011011",
  13209=>"000000000",
  13210=>"000000100",
  13211=>"000000000",
  13212=>"011111011",
  13213=>"000000000",
  13214=>"000001111",
  13215=>"000000111",
  13216=>"000111111",
  13217=>"010000010",
  13218=>"111111111",
  13219=>"111000000",
  13220=>"111111111",
  13221=>"010010010",
  13222=>"000000000",
  13223=>"111111001",
  13224=>"100110111",
  13225=>"010000000",
  13226=>"000000001",
  13227=>"000001001",
  13228=>"000000000",
  13229=>"001000000",
  13230=>"000101101",
  13231=>"000000110",
  13232=>"111111111",
  13233=>"011111111",
  13234=>"000100110",
  13235=>"000000000",
  13236=>"111011000",
  13237=>"110111111",
  13238=>"100111111",
  13239=>"100000000",
  13240=>"000000000",
  13241=>"000000101",
  13242=>"100110111",
  13243=>"111111111",
  13244=>"000000000",
  13245=>"111111000",
  13246=>"000000000",
  13247=>"001001000",
  13248=>"000000100",
  13249=>"010010111",
  13250=>"000000011",
  13251=>"000000000",
  13252=>"111111111",
  13253=>"000010000",
  13254=>"000000000",
  13255=>"100110000",
  13256=>"000111110",
  13257=>"000000000",
  13258=>"001000000",
  13259=>"000000111",
  13260=>"000000001",
  13261=>"000000000",
  13262=>"011111111",
  13263=>"000000111",
  13264=>"000000010",
  13265=>"110000110",
  13266=>"000000101",
  13267=>"000000100",
  13268=>"000000000",
  13269=>"100100000",
  13270=>"100100000",
  13271=>"000000001",
  13272=>"001000000",
  13273=>"001001000",
  13274=>"001000000",
  13275=>"000000000",
  13276=>"111111111",
  13277=>"100000000",
  13278=>"000000000",
  13279=>"000001001",
  13280=>"111001000",
  13281=>"000110111",
  13282=>"000000111",
  13283=>"100000110",
  13284=>"000000000",
  13285=>"001001011",
  13286=>"111101111",
  13287=>"000110111",
  13288=>"000000000",
  13289=>"011011111",
  13290=>"000111111",
  13291=>"000000000",
  13292=>"111111111",
  13293=>"000000000",
  13294=>"000110100",
  13295=>"001001111",
  13296=>"000000000",
  13297=>"000000000",
  13298=>"111111111",
  13299=>"000000000",
  13300=>"000000000",
  13301=>"111111111",
  13302=>"111011001",
  13303=>"010010000",
  13304=>"111110010",
  13305=>"000000000",
  13306=>"000010010",
  13307=>"111111111",
  13308=>"000000110",
  13309=>"110111111",
  13310=>"000000000",
  13311=>"000000000",
  13312=>"001001001",
  13313=>"000100000",
  13314=>"000000000",
  13315=>"100100101",
  13316=>"111111111",
  13317=>"000000110",
  13318=>"000011011",
  13319=>"000000000",
  13320=>"100110100",
  13321=>"000001001",
  13322=>"111111111",
  13323=>"111111100",
  13324=>"000000000",
  13325=>"111101100",
  13326=>"000001001",
  13327=>"100100110",
  13328=>"100101111",
  13329=>"110110100",
  13330=>"100010000",
  13331=>"111111001",
  13332=>"000010000",
  13333=>"000000110",
  13334=>"000000000",
  13335=>"000000000",
  13336=>"111111111",
  13337=>"100000000",
  13338=>"000000111",
  13339=>"001101111",
  13340=>"111111111",
  13341=>"001000000",
  13342=>"100110111",
  13343=>"111111111",
  13344=>"111111111",
  13345=>"000000000",
  13346=>"011001000",
  13347=>"000110111",
  13348=>"110110000",
  13349=>"000001111",
  13350=>"100100110",
  13351=>"111110111",
  13352=>"110110000",
  13353=>"000000000",
  13354=>"111000000",
  13355=>"000000000",
  13356=>"111011000",
  13357=>"000000000",
  13358=>"010011011",
  13359=>"111100111",
  13360=>"100111101",
  13361=>"000110000",
  13362=>"111111110",
  13363=>"000100110",
  13364=>"011000010",
  13365=>"101011110",
  13366=>"001111111",
  13367=>"000000001",
  13368=>"111100000",
  13369=>"100100001",
  13370=>"101000000",
  13371=>"110110111",
  13372=>"111000000",
  13373=>"111111100",
  13374=>"111111111",
  13375=>"000000100",
  13376=>"100100000",
  13377=>"111111111",
  13378=>"000110110",
  13379=>"111001000",
  13380=>"001000000",
  13381=>"111111111",
  13382=>"011011011",
  13383=>"000000000",
  13384=>"000000001",
  13385=>"111000000",
  13386=>"111100000",
  13387=>"000000000",
  13388=>"010101111",
  13389=>"111111001",
  13390=>"100000000",
  13391=>"111111110",
  13392=>"100110111",
  13393=>"000110111",
  13394=>"001011000",
  13395=>"011000000",
  13396=>"110110000",
  13397=>"000011111",
  13398=>"000000001",
  13399=>"111111111",
  13400=>"110111101",
  13401=>"011001001",
  13402=>"111111111",
  13403=>"000000001",
  13404=>"000000000",
  13405=>"111111111",
  13406=>"001100111",
  13407=>"000000000",
  13408=>"110111110",
  13409=>"011011001",
  13410=>"000000000",
  13411=>"110000000",
  13412=>"010000000",
  13413=>"101110111",
  13414=>"011111111",
  13415=>"111111111",
  13416=>"111111000",
  13417=>"000000110",
  13418=>"001011111",
  13419=>"001001000",
  13420=>"000000110",
  13421=>"001000000",
  13422=>"001001111",
  13423=>"011010000",
  13424=>"000000011",
  13425=>"000000010",
  13426=>"111111111",
  13427=>"100100000",
  13428=>"100000000",
  13429=>"000000000",
  13430=>"011000010",
  13431=>"000000000",
  13432=>"111100100",
  13433=>"000100101",
  13434=>"000000000",
  13435=>"000000011",
  13436=>"000000110",
  13437=>"111111111",
  13438=>"000000000",
  13439=>"000000111",
  13440=>"111000000",
  13441=>"111111111",
  13442=>"000011111",
  13443=>"000000100",
  13444=>"111111111",
  13445=>"000000101",
  13446=>"111111110",
  13447=>"111000000",
  13448=>"000000010",
  13449=>"000000110",
  13450=>"111111000",
  13451=>"000000111",
  13452=>"000011011",
  13453=>"000100100",
  13454=>"000010000",
  13455=>"111001001",
  13456=>"011011011",
  13457=>"111111111",
  13458=>"111100000",
  13459=>"000000000",
  13460=>"111111101",
  13461=>"000001011",
  13462=>"110110000",
  13463=>"000000110",
  13464=>"000000000",
  13465=>"000000000",
  13466=>"111111111",
  13467=>"000000000",
  13468=>"111101000",
  13469=>"111101100",
  13470=>"100000000",
  13471=>"111110111",
  13472=>"000110111",
  13473=>"000000001",
  13474=>"000000011",
  13475=>"111111111",
  13476=>"100100101",
  13477=>"110000000",
  13478=>"011000000",
  13479=>"110100111",
  13480=>"000000100",
  13481=>"100101111",
  13482=>"011011110",
  13483=>"111000000",
  13484=>"100100110",
  13485=>"001001111",
  13486=>"100000111",
  13487=>"110110111",
  13488=>"111111111",
  13489=>"110110000",
  13490=>"110110010",
  13491=>"000000000",
  13492=>"111111111",
  13493=>"100001011",
  13494=>"110111111",
  13495=>"000100100",
  13496=>"111101111",
  13497=>"010111111",
  13498=>"000000000",
  13499=>"111111111",
  13500=>"111111111",
  13501=>"110100000",
  13502=>"000111111",
  13503=>"110000000",
  13504=>"111111111",
  13505=>"000000000",
  13506=>"000000000",
  13507=>"101111111",
  13508=>"111100111",
  13509=>"111111111",
  13510=>"100101101",
  13511=>"100101011",
  13512=>"100100000",
  13513=>"111111111",
  13514=>"111000000",
  13515=>"111111111",
  13516=>"000001111",
  13517=>"000011001",
  13518=>"110000100",
  13519=>"000000100",
  13520=>"000101111",
  13521=>"000000000",
  13522=>"110000000",
  13523=>"000000000",
  13524=>"000000000",
  13525=>"100001001",
  13526=>"000111111",
  13527=>"001111011",
  13528=>"000000000",
  13529=>"010011111",
  13530=>"111010000",
  13531=>"111111111",
  13532=>"111001000",
  13533=>"111111111",
  13534=>"111111000",
  13535=>"100100101",
  13536=>"111111111",
  13537=>"011111011",
  13538=>"000011111",
  13539=>"000000010",
  13540=>"111111001",
  13541=>"000000000",
  13542=>"111110110",
  13543=>"111111000",
  13544=>"000010001",
  13545=>"001111111",
  13546=>"000011111",
  13547=>"100100111",
  13548=>"111111000",
  13549=>"011010000",
  13550=>"100110000",
  13551=>"110000000",
  13552=>"111111101",
  13553=>"110010000",
  13554=>"111111111",
  13555=>"000011010",
  13556=>"000000000",
  13557=>"110111111",
  13558=>"011011011",
  13559=>"111111001",
  13560=>"000011111",
  13561=>"100100100",
  13562=>"000000000",
  13563=>"111011011",
  13564=>"001001111",
  13565=>"100000100",
  13566=>"100110100",
  13567=>"100111111",
  13568=>"110111111",
  13569=>"101001001",
  13570=>"000000000",
  13571=>"000111111",
  13572=>"000000000",
  13573=>"000110000",
  13574=>"111111111",
  13575=>"000000000",
  13576=>"000000000",
  13577=>"000111111",
  13578=>"000000000",
  13579=>"111111110",
  13580=>"111000000",
  13581=>"000010111",
  13582=>"111111111",
  13583=>"111111000",
  13584=>"100100101",
  13585=>"100000000",
  13586=>"000000000",
  13587=>"111111101",
  13588=>"111111000",
  13589=>"111111111",
  13590=>"001110100",
  13591=>"111111111",
  13592=>"010110110",
  13593=>"000000000",
  13594=>"000000110",
  13595=>"111110110",
  13596=>"100100111",
  13597=>"011000000",
  13598=>"000000110",
  13599=>"000000000",
  13600=>"001000000",
  13601=>"111000000",
  13602=>"111111100",
  13603=>"111111100",
  13604=>"111101000",
  13605=>"001111111",
  13606=>"000000000",
  13607=>"000000011",
  13608=>"111111000",
  13609=>"110000000",
  13610=>"010011111",
  13611=>"000101000",
  13612=>"000000100",
  13613=>"001011011",
  13614=>"000011000",
  13615=>"000000100",
  13616=>"011011110",
  13617=>"101000001",
  13618=>"000011000",
  13619=>"011110000",
  13620=>"000011111",
  13621=>"100111110",
  13622=>"100000000",
  13623=>"100100000",
  13624=>"000000111",
  13625=>"000000011",
  13626=>"000000000",
  13627=>"100000000",
  13628=>"101001000",
  13629=>"000000110",
  13630=>"100100100",
  13631=>"000000000",
  13632=>"101111111",
  13633=>"100111110",
  13634=>"110001001",
  13635=>"111111111",
  13636=>"101101111",
  13637=>"110111111",
  13638=>"100000000",
  13639=>"000000000",
  13640=>"000000001",
  13641=>"011010000",
  13642=>"100110110",
  13643=>"010110110",
  13644=>"000000000",
  13645=>"000000111",
  13646=>"000001001",
  13647=>"001001111",
  13648=>"111111111",
  13649=>"001001011",
  13650=>"001111111",
  13651=>"001001111",
  13652=>"100000000",
  13653=>"011011111",
  13654=>"110000110",
  13655=>"110110111",
  13656=>"000000000",
  13657=>"111111111",
  13658=>"111101000",
  13659=>"000000010",
  13660=>"000000000",
  13661=>"000000001",
  13662=>"101001111",
  13663=>"000000000",
  13664=>"000000011",
  13665=>"000000000",
  13666=>"001001001",
  13667=>"000000011",
  13668=>"111011011",
  13669=>"111000000",
  13670=>"011111111",
  13671=>"000000000",
  13672=>"001101101",
  13673=>"000010010",
  13674=>"110000000",
  13675=>"111111111",
  13676=>"000000000",
  13677=>"000000000",
  13678=>"111100000",
  13679=>"110111011",
  13680=>"111011000",
  13681=>"000000000",
  13682=>"100000000",
  13683=>"111111001",
  13684=>"000011001",
  13685=>"001010010",
  13686=>"110111111",
  13687=>"000000000",
  13688=>"001001011",
  13689=>"000000000",
  13690=>"100000100",
  13691=>"111100110",
  13692=>"000000000",
  13693=>"111111111",
  13694=>"111111111",
  13695=>"111110000",
  13696=>"111111111",
  13697=>"111111111",
  13698=>"000110110",
  13699=>"111111111",
  13700=>"111100100",
  13701=>"000000111",
  13702=>"000000001",
  13703=>"111011111",
  13704=>"000000000",
  13705=>"101100111",
  13706=>"110000000",
  13707=>"111111011",
  13708=>"111111111",
  13709=>"000000000",
  13710=>"010010000",
  13711=>"000000000",
  13712=>"111111000",
  13713=>"000000000",
  13714=>"011011001",
  13715=>"110110000",
  13716=>"011000000",
  13717=>"000110010",
  13718=>"111101111",
  13719=>"011011111",
  13720=>"101011111",
  13721=>"100000000",
  13722=>"000001001",
  13723=>"000000000",
  13724=>"000000100",
  13725=>"000000000",
  13726=>"100000000",
  13727=>"110110000",
  13728=>"000000000",
  13729=>"100000000",
  13730=>"000000110",
  13731=>"000010000",
  13732=>"000000101",
  13733=>"111111110",
  13734=>"000011011",
  13735=>"111111111",
  13736=>"000110111",
  13737=>"001000000",
  13738=>"111110100",
  13739=>"111001000",
  13740=>"110111010",
  13741=>"011011111",
  13742=>"000110000",
  13743=>"110110000",
  13744=>"000000010",
  13745=>"111111111",
  13746=>"110000000",
  13747=>"111011110",
  13748=>"000010110",
  13749=>"000000101",
  13750=>"101111100",
  13751=>"110110100",
  13752=>"000000100",
  13753=>"110100100",
  13754=>"110110000",
  13755=>"110111000",
  13756=>"011010110",
  13757=>"111011111",
  13758=>"111111111",
  13759=>"000101101",
  13760=>"000110000",
  13761=>"110010110",
  13762=>"000000000",
  13763=>"011111111",
  13764=>"000000110",
  13765=>"000000100",
  13766=>"001111111",
  13767=>"111111111",
  13768=>"100000000",
  13769=>"111111111",
  13770=>"011011011",
  13771=>"000000000",
  13772=>"000000100",
  13773=>"111111011",
  13774=>"111111111",
  13775=>"111100101",
  13776=>"111110000",
  13777=>"101111111",
  13778=>"111111000",
  13779=>"001100111",
  13780=>"001001111",
  13781=>"011001111",
  13782=>"100101000",
  13783=>"010000000",
  13784=>"000000000",
  13785=>"100111111",
  13786=>"000000000",
  13787=>"000100000",
  13788=>"111010011",
  13789=>"001001001",
  13790=>"111111111",
  13791=>"100100111",
  13792=>"010010011",
  13793=>"001001100",
  13794=>"111000000",
  13795=>"000000001",
  13796=>"000100111",
  13797=>"000000100",
  13798=>"111111111",
  13799=>"010011000",
  13800=>"001001000",
  13801=>"111111111",
  13802=>"011111110",
  13803=>"101111111",
  13804=>"110110100",
  13805=>"110100100",
  13806=>"111111000",
  13807=>"000100100",
  13808=>"000000000",
  13809=>"000100111",
  13810=>"000000110",
  13811=>"111111011",
  13812=>"000000000",
  13813=>"000000000",
  13814=>"111111111",
  13815=>"111011001",
  13816=>"000000000",
  13817=>"000100110",
  13818=>"000010111",
  13819=>"110010000",
  13820=>"100010010",
  13821=>"101011111",
  13822=>"111111111",
  13823=>"110111011",
  13824=>"111111111",
  13825=>"000000001",
  13826=>"111111111",
  13827=>"111111000",
  13828=>"111111111",
  13829=>"111000000",
  13830=>"111111111",
  13831=>"111001000",
  13832=>"000001111",
  13833=>"111111000",
  13834=>"100100111",
  13835=>"000000000",
  13836=>"110110110",
  13837=>"000000100",
  13838=>"110001110",
  13839=>"111111111",
  13840=>"000100100",
  13841=>"000000000",
  13842=>"000000000",
  13843=>"000000000",
  13844=>"100000000",
  13845=>"111111000",
  13846=>"000011001",
  13847=>"001000000",
  13848=>"000000000",
  13849=>"000001001",
  13850=>"000000000",
  13851=>"111111001",
  13852=>"111111111",
  13853=>"110000000",
  13854=>"100000000",
  13855=>"000001001",
  13856=>"001000000",
  13857=>"111111111",
  13858=>"110100000",
  13859=>"111111111",
  13860=>"011011011",
  13861=>"101001000",
  13862=>"111010111",
  13863=>"011111110",
  13864=>"000100100",
  13865=>"111111010",
  13866=>"000000001",
  13867=>"111111111",
  13868=>"100001000",
  13869=>"111111000",
  13870=>"111111111",
  13871=>"100000000",
  13872=>"111111111",
  13873=>"111111111",
  13874=>"001101001",
  13875=>"000100100",
  13876=>"000100100",
  13877=>"000011001",
  13878=>"000001000",
  13879=>"111000010",
  13880=>"111101100",
  13881=>"001000000",
  13882=>"110000000",
  13883=>"000000111",
  13884=>"101101000",
  13885=>"011011111",
  13886=>"111110100",
  13887=>"000000000",
  13888=>"111111111",
  13889=>"101111111",
  13890=>"000001001",
  13891=>"000010010",
  13892=>"111011001",
  13893=>"001001001",
  13894=>"110000000",
  13895=>"111111111",
  13896=>"000011111",
  13897=>"000000000",
  13898=>"011011011",
  13899=>"000011011",
  13900=>"111111111",
  13901=>"011011111",
  13902=>"000000000",
  13903=>"111111111",
  13904=>"110100000",
  13905=>"111110000",
  13906=>"001000000",
  13907=>"000000001",
  13908=>"111111111",
  13909=>"000000000",
  13910=>"011011111",
  13911=>"000000000",
  13912=>"000000000",
  13913=>"100000000",
  13914=>"100111000",
  13915=>"111100000",
  13916=>"111111111",
  13917=>"000000000",
  13918=>"110001111",
  13919=>"010000101",
  13920=>"000111111",
  13921=>"000000000",
  13922=>"011111101",
  13923=>"000000000",
  13924=>"111111000",
  13925=>"111111001",
  13926=>"111111011",
  13927=>"000000000",
  13928=>"111101101",
  13929=>"000100111",
  13930=>"000000000",
  13931=>"101111111",
  13932=>"111111111",
  13933=>"111111111",
  13934=>"111111111",
  13935=>"110110110",
  13936=>"000000001",
  13937=>"100000000",
  13938=>"111111111",
  13939=>"111111111",
  13940=>"000000100",
  13941=>"111111111",
  13942=>"111111000",
  13943=>"000000000",
  13944=>"001101001",
  13945=>"111111111",
  13946=>"100100100",
  13947=>"111111110",
  13948=>"110011110",
  13949=>"000000100",
  13950=>"100111101",
  13951=>"000000000",
  13952=>"000000000",
  13953=>"111111111",
  13954=>"000000001",
  13955=>"000101100",
  13956=>"011000000",
  13957=>"000000000",
  13958=>"111111111",
  13959=>"000000000",
  13960=>"000000000",
  13961=>"111111111",
  13962=>"000000111",
  13963=>"000000000",
  13964=>"111111000",
  13965=>"000000000",
  13966=>"111111010",
  13967=>"000001000",
  13968=>"000000000",
  13969=>"111111111",
  13970=>"000000110",
  13971=>"000000110",
  13972=>"111111111",
  13973=>"111001011",
  13974=>"000000000",
  13975=>"000000111",
  13976=>"000000111",
  13977=>"111111111",
  13978=>"000000000",
  13979=>"000001001",
  13980=>"100111111",
  13981=>"111001001",
  13982=>"111111111",
  13983=>"111111011",
  13984=>"011010011",
  13985=>"000000000",
  13986=>"111101101",
  13987=>"000000111",
  13988=>"000110000",
  13989=>"100101111",
  13990=>"101111000",
  13991=>"000001001",
  13992=>"100000100",
  13993=>"000000000",
  13994=>"111111111",
  13995=>"111111111",
  13996=>"111111111",
  13997=>"111011011",
  13998=>"111111111",
  13999=>"111001001",
  14000=>"100111111",
  14001=>"000001001",
  14002=>"110111110",
  14003=>"111111111",
  14004=>"001001001",
  14005=>"000110000",
  14006=>"000000000",
  14007=>"110111111",
  14008=>"000000001",
  14009=>"111000000",
  14010=>"000000000",
  14011=>"111000011",
  14012=>"001000111",
  14013=>"111010000",
  14014=>"111000111",
  14015=>"111111111",
  14016=>"000000001",
  14017=>"000100100",
  14018=>"000000000",
  14019=>"000000011",
  14020=>"000100000",
  14021=>"000100111",
  14022=>"111111111",
  14023=>"000000000",
  14024=>"111111111",
  14025=>"000000000",
  14026=>"001101111",
  14027=>"100000100",
  14028=>"000000000",
  14029=>"111111111",
  14030=>"111001101",
  14031=>"000000111",
  14032=>"110111111",
  14033=>"101000111",
  14034=>"111011111",
  14035=>"111111100",
  14036=>"111111111",
  14037=>"000000000",
  14038=>"000100111",
  14039=>"000000000",
  14040=>"111101100",
  14041=>"101111110",
  14042=>"111111011",
  14043=>"000111111",
  14044=>"001111111",
  14045=>"000100000",
  14046=>"000111000",
  14047=>"000000000",
  14048=>"111111111",
  14049=>"000000000",
  14050=>"000011000",
  14051=>"000000000",
  14052=>"101101111",
  14053=>"111001001",
  14054=>"100000000",
  14055=>"111111111",
  14056=>"111111100",
  14057=>"111101111",
  14058=>"001000100",
  14059=>"111111000",
  14060=>"111111111",
  14061=>"110010000",
  14062=>"000000100",
  14063=>"000000000",
  14064=>"111111000",
  14065=>"000000011",
  14066=>"011011011",
  14067=>"000001011",
  14068=>"000000000",
  14069=>"000001001",
  14070=>"000000000",
  14071=>"000000100",
  14072=>"100111100",
  14073=>"111111111",
  14074=>"111111111",
  14075=>"111111111",
  14076=>"000111101",
  14077=>"001001001",
  14078=>"110111111",
  14079=>"000000000",
  14080=>"100000000",
  14081=>"111100100",
  14082=>"000000010",
  14083=>"000000001",
  14084=>"000001111",
  14085=>"000000000",
  14086=>"000000110",
  14087=>"000000111",
  14088=>"000111111",
  14089=>"100100110",
  14090=>"000000111",
  14091=>"000100100",
  14092=>"001000110",
  14093=>"100110111",
  14094=>"111111111",
  14095=>"111111001",
  14096=>"000000000",
  14097=>"101000100",
  14098=>"000000000",
  14099=>"111000000",
  14100=>"000000110",
  14101=>"010010110",
  14102=>"000100110",
  14103=>"000111111",
  14104=>"101111111",
  14105=>"111111111",
  14106=>"111111001",
  14107=>"100000110",
  14108=>"000000000",
  14109=>"000000000",
  14110=>"111111001",
  14111=>"111111111",
  14112=>"000110110",
  14113=>"000000001",
  14114=>"000111110",
  14115=>"111101111",
  14116=>"111011000",
  14117=>"110110000",
  14118=>"111111000",
  14119=>"001101111",
  14120=>"111111111",
  14121=>"111111111",
  14122=>"101001011",
  14123=>"110111111",
  14124=>"111111111",
  14125=>"000000011",
  14126=>"111111111",
  14127=>"000000000",
  14128=>"000000000",
  14129=>"110000000",
  14130=>"000001100",
  14131=>"111111110",
  14132=>"111100100",
  14133=>"111001001",
  14134=>"111111100",
  14135=>"111111011",
  14136=>"000000000",
  14137=>"101111111",
  14138=>"101000101",
  14139=>"111111100",
  14140=>"101001000",
  14141=>"110110000",
  14142=>"111111000",
  14143=>"111111111",
  14144=>"000000111",
  14145=>"000000000",
  14146=>"111101101",
  14147=>"100100111",
  14148=>"011000000",
  14149=>"000000000",
  14150=>"011111111",
  14151=>"001001111",
  14152=>"000000000",
  14153=>"011111111",
  14154=>"000100001",
  14155=>"110111111",
  14156=>"110100100",
  14157=>"000000000",
  14158=>"000011111",
  14159=>"000001001",
  14160=>"011010000",
  14161=>"000101111",
  14162=>"000001001",
  14163=>"000000000",
  14164=>"000000000",
  14165=>"011011011",
  14166=>"000000000",
  14167=>"111111111",
  14168=>"111111111",
  14169=>"000111111",
  14170=>"011011000",
  14171=>"000000100",
  14172=>"000000111",
  14173=>"000000000",
  14174=>"000000001",
  14175=>"011111111",
  14176=>"111110110",
  14177=>"000000111",
  14178=>"000000000",
  14179=>"100000000",
  14180=>"011010000",
  14181=>"000000000",
  14182=>"111111111",
  14183=>"111011111",
  14184=>"001001111",
  14185=>"111111111",
  14186=>"010011111",
  14187=>"111001000",
  14188=>"100011001",
  14189=>"000000111",
  14190=>"000000000",
  14191=>"101000000",
  14192=>"111111111",
  14193=>"000000000",
  14194=>"111000011",
  14195=>"100010000",
  14196=>"000000000",
  14197=>"000100111",
  14198=>"011011100",
  14199=>"111111111",
  14200=>"111000000",
  14201=>"111000000",
  14202=>"000000000",
  14203=>"000000000",
  14204=>"111110110",
  14205=>"111000000",
  14206=>"011100000",
  14207=>"100000011",
  14208=>"000000100",
  14209=>"000000000",
  14210=>"110100100",
  14211=>"111111111",
  14212=>"000000000",
  14213=>"111111111",
  14214=>"000001010",
  14215=>"110100000",
  14216=>"000000000",
  14217=>"010100100",
  14218=>"000111111",
  14219=>"110000100",
  14220=>"101001011",
  14221=>"111110100",
  14222=>"111111111",
  14223=>"111111111",
  14224=>"000000000",
  14225=>"111111111",
  14226=>"000000000",
  14227=>"000000000",
  14228=>"111111110",
  14229=>"000000000",
  14230=>"111111111",
  14231=>"001011011",
  14232=>"000000000",
  14233=>"000000101",
  14234=>"111111111",
  14235=>"110101001",
  14236=>"000011011",
  14237=>"111000000",
  14238=>"001011001",
  14239=>"000000000",
  14240=>"101111001",
  14241=>"011000101",
  14242=>"101000000",
  14243=>"111111111",
  14244=>"000000000",
  14245=>"011000000",
  14246=>"111111111",
  14247=>"000001111",
  14248=>"000000001",
  14249=>"001000101",
  14250=>"011111100",
  14251=>"001111111",
  14252=>"000000000",
  14253=>"111111111",
  14254=>"000110100",
  14255=>"110100001",
  14256=>"000111111",
  14257=>"111111110",
  14258=>"011101000",
  14259=>"000000111",
  14260=>"000000000",
  14261=>"111111111",
  14262=>"110111111",
  14263=>"100111001",
  14264=>"000000000",
  14265=>"100110110",
  14266=>"111101001",
  14267=>"001000000",
  14268=>"111111101",
  14269=>"000000000",
  14270=>"111111111",
  14271=>"100100100",
  14272=>"111111111",
  14273=>"101001001",
  14274=>"000000000",
  14275=>"111111100",
  14276=>"000000101",
  14277=>"011010110",
  14278=>"001000000",
  14279=>"001000000",
  14280=>"111011111",
  14281=>"111000000",
  14282=>"000000000",
  14283=>"111111111",
  14284=>"111111110",
  14285=>"111111111",
  14286=>"010000100",
  14287=>"000000000",
  14288=>"000000000",
  14289=>"000000011",
  14290=>"111111111",
  14291=>"100000000",
  14292=>"111111111",
  14293=>"001111001",
  14294=>"000000000",
  14295=>"111111001",
  14296=>"011111111",
  14297=>"000000001",
  14298=>"111111111",
  14299=>"111101111",
  14300=>"000100100",
  14301=>"001011111",
  14302=>"011011111",
  14303=>"000000000",
  14304=>"000000000",
  14305=>"111111111",
  14306=>"011011000",
  14307=>"000011111",
  14308=>"000000000",
  14309=>"001001011",
  14310=>"000000000",
  14311=>"000000000",
  14312=>"101100100",
  14313=>"000011011",
  14314=>"011000000",
  14315=>"100000000",
  14316=>"111111111",
  14317=>"111001001",
  14318=>"000011111",
  14319=>"000000000",
  14320=>"111111111",
  14321=>"111111011",
  14322=>"000000100",
  14323=>"111000101",
  14324=>"001001001",
  14325=>"111000011",
  14326=>"111100000",
  14327=>"100100100",
  14328=>"110110111",
  14329=>"011011001",
  14330=>"000000000",
  14331=>"000000000",
  14332=>"000000011",
  14333=>"110100110",
  14334=>"111111001",
  14335=>"000000000",
  14336=>"111000000",
  14337=>"111111000",
  14338=>"000000000",
  14339=>"000000000",
  14340=>"100001001",
  14341=>"011111111",
  14342=>"001001001",
  14343=>"100101101",
  14344=>"111111011",
  14345=>"000000011",
  14346=>"111011011",
  14347=>"001000000",
  14348=>"100100111",
  14349=>"111101100",
  14350=>"000000000",
  14351=>"000001001",
  14352=>"111000100",
  14353=>"000000111",
  14354=>"111001001",
  14355=>"111111111",
  14356=>"000000000",
  14357=>"111111111",
  14358=>"110110111",
  14359=>"001100100",
  14360=>"001011111",
  14361=>"111101001",
  14362=>"000000111",
  14363=>"111010100",
  14364=>"000000000",
  14365=>"001001000",
  14366=>"000000110",
  14367=>"111110110",
  14368=>"000001001",
  14369=>"100110110",
  14370=>"000000000",
  14371=>"110111001",
  14372=>"011000000",
  14373=>"111111111",
  14374=>"001111111",
  14375=>"111101001",
  14376=>"111101100",
  14377=>"000000000",
  14378=>"111101111",
  14379=>"000011000",
  14380=>"010110110",
  14381=>"001111011",
  14382=>"001001011",
  14383=>"001001011",
  14384=>"000000000",
  14385=>"101001111",
  14386=>"000001001",
  14387=>"000111100",
  14388=>"111111001",
  14389=>"001000001",
  14390=>"111111111",
  14391=>"011110110",
  14392=>"001000000",
  14393=>"000000000",
  14394=>"111111111",
  14395=>"111000000",
  14396=>"100001111",
  14397=>"000110110",
  14398=>"101001011",
  14399=>"000000000",
  14400=>"111111111",
  14401=>"110110000",
  14402=>"011011101",
  14403=>"000000010",
  14404=>"110100100",
  14405=>"001001001",
  14406=>"000000000",
  14407=>"000100100",
  14408=>"001000011",
  14409=>"100000000",
  14410=>"000000111",
  14411=>"000111000",
  14412=>"101101000",
  14413=>"000000111",
  14414=>"000001011",
  14415=>"000111111",
  14416=>"000000000",
  14417=>"000111111",
  14418=>"000000000",
  14419=>"111010001",
  14420=>"001000000",
  14421=>"011000111",
  14422=>"000111000",
  14423=>"111101101",
  14424=>"111111010",
  14425=>"100000000",
  14426=>"110111111",
  14427=>"001000000",
  14428=>"000000000",
  14429=>"110100111",
  14430=>"000000000",
  14431=>"111111011",
  14432=>"101101001",
  14433=>"111111010",
  14434=>"100111111",
  14435=>"100100000",
  14436=>"111111111",
  14437=>"000111111",
  14438=>"000000011",
  14439=>"111110111",
  14440=>"111111111",
  14441=>"111101000",
  14442=>"000000000",
  14443=>"111110011",
  14444=>"000000000",
  14445=>"001011111",
  14446=>"000000001",
  14447=>"010111110",
  14448=>"100111010",
  14449=>"000000000",
  14450=>"111111111",
  14451=>"000000011",
  14452=>"011111001",
  14453=>"111111111",
  14454=>"111001000",
  14455=>"111011011",
  14456=>"000000000",
  14457=>"111111110",
  14458=>"111111111",
  14459=>"000000000",
  14460=>"111111110",
  14461=>"100001101",
  14462=>"000110111",
  14463=>"111111111",
  14464=>"000000010",
  14465=>"111111111",
  14466=>"000000000",
  14467=>"010111111",
  14468=>"001000001",
  14469=>"110000000",
  14470=>"111001001",
  14471=>"000000000",
  14472=>"000010010",
  14473=>"111111111",
  14474=>"000101111",
  14475=>"010111111",
  14476=>"000000000",
  14477=>"001101111",
  14478=>"001001101",
  14479=>"111100110",
  14480=>"110110000",
  14481=>"100000000",
  14482=>"000111000",
  14483=>"100000100",
  14484=>"111111000",
  14485=>"111111111",
  14486=>"000000000",
  14487=>"000000000",
  14488=>"000000000",
  14489=>"110111110",
  14490=>"111100111",
  14491=>"111100000",
  14492=>"110111111",
  14493=>"111011011",
  14494=>"000000000",
  14495=>"000010011",
  14496=>"011010000",
  14497=>"001000010",
  14498=>"000001001",
  14499=>"111111111",
  14500=>"000000100",
  14501=>"011001001",
  14502=>"000000000",
  14503=>"100100110",
  14504=>"000111000",
  14505=>"000001111",
  14506=>"001000101",
  14507=>"100000000",
  14508=>"111111111",
  14509=>"000000000",
  14510=>"111111111",
  14511=>"111011111",
  14512=>"000111000",
  14513=>"011011111",
  14514=>"100110110",
  14515=>"000000000",
  14516=>"101001111",
  14517=>"011111111",
  14518=>"111100100",
  14519=>"001000000",
  14520=>"000000000",
  14521=>"010000000",
  14522=>"110100111",
  14523=>"000110100",
  14524=>"000000000",
  14525=>"000000000",
  14526=>"111111011",
  14527=>"000010000",
  14528=>"111001001",
  14529=>"001011111",
  14530=>"111111111",
  14531=>"000000000",
  14532=>"100100000",
  14533=>"000000000",
  14534=>"111000000",
  14535=>"000000000",
  14536=>"000000111",
  14537=>"000010000",
  14538=>"100100101",
  14539=>"111011011",
  14540=>"000000000",
  14541=>"001011111",
  14542=>"011011011",
  14543=>"111101000",
  14544=>"111111111",
  14545=>"111110110",
  14546=>"000000110",
  14547=>"111111111",
  14548=>"000000000",
  14549=>"000101000",
  14550=>"000000000",
  14551=>"100110010",
  14552=>"000001111",
  14553=>"000111000",
  14554=>"000000000",
  14555=>"000000000",
  14556=>"111111111",
  14557=>"000111111",
  14558=>"000000000",
  14559=>"011111111",
  14560=>"100111001",
  14561=>"000100010",
  14562=>"010100000",
  14563=>"000000000",
  14564=>"111000000",
  14565=>"000100000",
  14566=>"111111111",
  14567=>"000000000",
  14568=>"000111111",
  14569=>"111111010",
  14570=>"011000111",
  14571=>"011111111",
  14572=>"111011010",
  14573=>"111110000",
  14574=>"111111111",
  14575=>"000000000",
  14576=>"111100100",
  14577=>"000000100",
  14578=>"110001000",
  14579=>"000000000",
  14580=>"000000100",
  14581=>"110110000",
  14582=>"111111111",
  14583=>"111110111",
  14584=>"111110010",
  14585=>"000000000",
  14586=>"000110001",
  14587=>"000111111",
  14588=>"011001010",
  14589=>"110111111",
  14590=>"001111110",
  14591=>"011011111",
  14592=>"000001001",
  14593=>"111110110",
  14594=>"000000000",
  14595=>"000000111",
  14596=>"000010000",
  14597=>"000000111",
  14598=>"000000001",
  14599=>"111011011",
  14600=>"000111111",
  14601=>"000000111",
  14602=>"000000100",
  14603=>"000000000",
  14604=>"100000000",
  14605=>"001001000",
  14606=>"111111111",
  14607=>"001011111",
  14608=>"100100000",
  14609=>"000000000",
  14610=>"101101111",
  14611=>"000111010",
  14612=>"111111111",
  14613=>"100000000",
  14614=>"100000000",
  14615=>"001100101",
  14616=>"000000000",
  14617=>"110110111",
  14618=>"000000000",
  14619=>"111111000",
  14620=>"000100000",
  14621=>"000000000",
  14622=>"101000000",
  14623=>"000000000",
  14624=>"111111011",
  14625=>"000011111",
  14626=>"001000000",
  14627=>"111111000",
  14628=>"000001001",
  14629=>"101101101",
  14630=>"111111111",
  14631=>"000000010",
  14632=>"101001100",
  14633=>"111111111",
  14634=>"000011011",
  14635=>"111111001",
  14636=>"111111101",
  14637=>"001111111",
  14638=>"000000000",
  14639=>"110110100",
  14640=>"111000000",
  14641=>"000000000",
  14642=>"101000000",
  14643=>"010011011",
  14644=>"000000000",
  14645=>"110111111",
  14646=>"000111111",
  14647=>"111111000",
  14648=>"111110110",
  14649=>"000000111",
  14650=>"001011011",
  14651=>"101001000",
  14652=>"000000001",
  14653=>"011111111",
  14654=>"000100110",
  14655=>"111111111",
  14656=>"100111111",
  14657=>"100100000",
  14658=>"000000000",
  14659=>"111101111",
  14660=>"111111000",
  14661=>"000110100",
  14662=>"111000111",
  14663=>"000000100",
  14664=>"000000000",
  14665=>"111111000",
  14666=>"000000110",
  14667=>"001111111",
  14668=>"111011001",
  14669=>"110000100",
  14670=>"111111100",
  14671=>"111101101",
  14672=>"001001111",
  14673=>"011011011",
  14674=>"000000000",
  14675=>"000000000",
  14676=>"100100000",
  14677=>"011011011",
  14678=>"111111111",
  14679=>"000001111",
  14680=>"001111111",
  14681=>"000000000",
  14682=>"000001111",
  14683=>"000000000",
  14684=>"000000010",
  14685=>"001000000",
  14686=>"110000010",
  14687=>"111111110",
  14688=>"001011011",
  14689=>"110111001",
  14690=>"000000001",
  14691=>"011111111",
  14692=>"000000101",
  14693=>"111011011",
  14694=>"001000000",
  14695=>"000110100",
  14696=>"111011101",
  14697=>"111000000",
  14698=>"101000000",
  14699=>"000100000",
  14700=>"001000000",
  14701=>"000000011",
  14702=>"000001000",
  14703=>"100111111",
  14704=>"000000000",
  14705=>"001001001",
  14706=>"011111111",
  14707=>"001001100",
  14708=>"000011011",
  14709=>"010010110",
  14710=>"000011001",
  14711=>"000000111",
  14712=>"000010000",
  14713=>"000000000",
  14714=>"110110000",
  14715=>"000000000",
  14716=>"111111111",
  14717=>"111111111",
  14718=>"001011011",
  14719=>"111111101",
  14720=>"110100100",
  14721=>"111110111",
  14722=>"011000001",
  14723=>"010111001",
  14724=>"111111111",
  14725=>"000001001",
  14726=>"010000000",
  14727=>"000001111",
  14728=>"000000010",
  14729=>"000000000",
  14730=>"001000000",
  14731=>"110000000",
  14732=>"111111111",
  14733=>"100000100",
  14734=>"111111101",
  14735=>"100111100",
  14736=>"000000100",
  14737=>"000000000",
  14738=>"111111111",
  14739=>"000000000",
  14740=>"111000000",
  14741=>"011001011",
  14742=>"101000000",
  14743=>"010011011",
  14744=>"111101111",
  14745=>"000111111",
  14746=>"000101011",
  14747=>"111111111",
  14748=>"000101111",
  14749=>"000000000",
  14750=>"100000000",
  14751=>"000000000",
  14752=>"111111111",
  14753=>"011001111",
  14754=>"000100000",
  14755=>"000111111",
  14756=>"000000100",
  14757=>"111111111",
  14758=>"111111000",
  14759=>"100111101",
  14760=>"100110000",
  14761=>"110111111",
  14762=>"000110100",
  14763=>"001001100",
  14764=>"111111111",
  14765=>"011001000",
  14766=>"111111111",
  14767=>"000001011",
  14768=>"000100100",
  14769=>"111111001",
  14770=>"100000100",
  14771=>"000110110",
  14772=>"011111000",
  14773=>"000000111",
  14774=>"100110111",
  14775=>"000110110",
  14776=>"000000000",
  14777=>"000111111",
  14778=>"000000000",
  14779=>"101001000",
  14780=>"100100000",
  14781=>"001101100",
  14782=>"100100111",
  14783=>"100110110",
  14784=>"000000001",
  14785=>"000000000",
  14786=>"110110000",
  14787=>"000000000",
  14788=>"000000000",
  14789=>"001111110",
  14790=>"000000000",
  14791=>"000000111",
  14792=>"000010000",
  14793=>"111011011",
  14794=>"111111000",
  14795=>"100100111",
  14796=>"100111111",
  14797=>"000000000",
  14798=>"110001000",
  14799=>"111110111",
  14800=>"000000110",
  14801=>"111111111",
  14802=>"110111111",
  14803=>"000000101",
  14804=>"110110110",
  14805=>"000000000",
  14806=>"111111101",
  14807=>"000000001",
  14808=>"000111001",
  14809=>"111111111",
  14810=>"111111111",
  14811=>"000100111",
  14812=>"111000100",
  14813=>"111111011",
  14814=>"000000000",
  14815=>"100100100",
  14816=>"000000001",
  14817=>"000001000",
  14818=>"000000100",
  14819=>"111111111",
  14820=>"000111111",
  14821=>"111111111",
  14822=>"111111111",
  14823=>"000000000",
  14824=>"000011011",
  14825=>"001001001",
  14826=>"000000011",
  14827=>"101101100",
  14828=>"100000000",
  14829=>"011001001",
  14830=>"000000110",
  14831=>"000001000",
  14832=>"100101111",
  14833=>"001111101",
  14834=>"111100101",
  14835=>"100111000",
  14836=>"000000001",
  14837=>"101100111",
  14838=>"000000000",
  14839=>"111001000",
  14840=>"111111000",
  14841=>"101111101",
  14842=>"000111111",
  14843=>"001001101",
  14844=>"100000111",
  14845=>"000000000",
  14846=>"001000000",
  14847=>"111111111",
  14848=>"000000000",
  14849=>"000000100",
  14850=>"000100111",
  14851=>"101000000",
  14852=>"111011000",
  14853=>"000100000",
  14854=>"111000000",
  14855=>"111011011",
  14856=>"000100111",
  14857=>"111111110",
  14858=>"111111111",
  14859=>"000111000",
  14860=>"111111000",
  14861=>"000000000",
  14862=>"011011111",
  14863=>"111001001",
  14864=>"000000000",
  14865=>"111111111",
  14866=>"000000000",
  14867=>"000111111",
  14868=>"000000000",
  14869=>"000111111",
  14870=>"111110110",
  14871=>"111111101",
  14872=>"011011111",
  14873=>"011011000",
  14874=>"100111111",
  14875=>"000000000",
  14876=>"111110100",
  14877=>"110111011",
  14878=>"000100001",
  14879=>"110111111",
  14880=>"000100101",
  14881=>"001111111",
  14882=>"000011111",
  14883=>"000000000",
  14884=>"000111111",
  14885=>"000000000",
  14886=>"101001111",
  14887=>"000000111",
  14888=>"000000000",
  14889=>"001100100",
  14890=>"000111111",
  14891=>"000110110",
  14892=>"011010000",
  14893=>"001111111",
  14894=>"011000000",
  14895=>"000110111",
  14896=>"000000000",
  14897=>"111001000",
  14898=>"110000000",
  14899=>"111011000",
  14900=>"001001111",
  14901=>"000000000",
  14902=>"000110110",
  14903=>"111011001",
  14904=>"011110110",
  14905=>"110111111",
  14906=>"101001000",
  14907=>"000000000",
  14908=>"111110000",
  14909=>"001100000",
  14910=>"110110000",
  14911=>"000110000",
  14912=>"010010110",
  14913=>"101111111",
  14914=>"111000000",
  14915=>"000000000",
  14916=>"111111111",
  14917=>"111000000",
  14918=>"111000000",
  14919=>"101000000",
  14920=>"001011000",
  14921=>"000000111",
  14922=>"000100000",
  14923=>"111011111",
  14924=>"000000000",
  14925=>"111100111",
  14926=>"111110111",
  14927=>"111011000",
  14928=>"000100111",
  14929=>"111110000",
  14930=>"000100111",
  14931=>"111011001",
  14932=>"111001000",
  14933=>"000000000",
  14934=>"100110000",
  14935=>"000000000",
  14936=>"000111111",
  14937=>"000000111",
  14938=>"100000100",
  14939=>"011111111",
  14940=>"000000111",
  14941=>"000111111",
  14942=>"000111111",
  14943=>"111111110",
  14944=>"000000000",
  14945=>"100000000",
  14946=>"110110100",
  14947=>"111100001",
  14948=>"100000000",
  14949=>"101101111",
  14950=>"111111000",
  14951=>"111000111",
  14952=>"000000000",
  14953=>"101100101",
  14954=>"111111111",
  14955=>"011011111",
  14956=>"111000001",
  14957=>"000000000",
  14958=>"110000000",
  14959=>"111100111",
  14960=>"000000000",
  14961=>"101100000",
  14962=>"000000000",
  14963=>"000000000",
  14964=>"000000000",
  14965=>"000111111",
  14966=>"000000001",
  14967=>"000111000",
  14968=>"000111111",
  14969=>"111111101",
  14970=>"111000000",
  14971=>"000000110",
  14972=>"011011110",
  14973=>"011111110",
  14974=>"000000000",
  14975=>"000001111",
  14976=>"000000000",
  14977=>"000011111",
  14978=>"110110111",
  14979=>"100100000",
  14980=>"000000111",
  14981=>"110000000",
  14982=>"000000001",
  14983=>"111111011",
  14984=>"111000000",
  14985=>"111111001",
  14986=>"000000111",
  14987=>"111110000",
  14988=>"000011111",
  14989=>"000000000",
  14990=>"111000000",
  14991=>"000000001",
  14992=>"111000000",
  14993=>"111001000",
  14994=>"000000000",
  14995=>"111111110",
  14996=>"010000011",
  14997=>"111011001",
  14998=>"000001000",
  14999=>"000000110",
  15000=>"111101111",
  15001=>"000000010",
  15002=>"111111111",
  15003=>"111111111",
  15004=>"000011111",
  15005=>"111100000",
  15006=>"000111111",
  15007=>"000000000",
  15008=>"111001000",
  15009=>"110110110",
  15010=>"111111111",
  15011=>"000110110",
  15012=>"101000101",
  15013=>"000000000",
  15014=>"111111111",
  15015=>"000111000",
  15016=>"111111111",
  15017=>"100011011",
  15018=>"001111111",
  15019=>"111111111",
  15020=>"000000000",
  15021=>"000000011",
  15022=>"000000000",
  15023=>"101000000",
  15024=>"111011011",
  15025=>"100000000",
  15026=>"111111011",
  15027=>"111001000",
  15028=>"000010110",
  15029=>"000011111",
  15030=>"110111111",
  15031=>"100100110",
  15032=>"000000000",
  15033=>"000000000",
  15034=>"111000000",
  15035=>"111000011",
  15036=>"000000110",
  15037=>"000000000",
  15038=>"000000000",
  15039=>"111111111",
  15040=>"111110000",
  15041=>"000100111",
  15042=>"111111111",
  15043=>"000000001",
  15044=>"000001111",
  15045=>"000000001",
  15046=>"000000001",
  15047=>"000111111",
  15048=>"000000000",
  15049=>"100111111",
  15050=>"010000000",
  15051=>"111111001",
  15052=>"000000000",
  15053=>"110110000",
  15054=>"010010111",
  15055=>"111100100",
  15056=>"000000001",
  15057=>"111001000",
  15058=>"111000000",
  15059=>"000000011",
  15060=>"110110000",
  15061=>"000000000",
  15062=>"000000101",
  15063=>"110110100",
  15064=>"011000111",
  15065=>"111000100",
  15066=>"000000111",
  15067=>"110011000",
  15068=>"000010001",
  15069=>"001001001",
  15070=>"000111111",
  15071=>"000010000",
  15072=>"000000001",
  15073=>"001111111",
  15074=>"111111100",
  15075=>"110111110",
  15076=>"000000000",
  15077=>"010110111",
  15078=>"000110111",
  15079=>"111110010",
  15080=>"010000100",
  15081=>"111100000",
  15082=>"000110100",
  15083=>"110000000",
  15084=>"111000000",
  15085=>"110111111",
  15086=>"111110000",
  15087=>"111001001",
  15088=>"000011111",
  15089=>"111010111",
  15090=>"000000111",
  15091=>"000100000",
  15092=>"111011000",
  15093=>"001111000",
  15094=>"011111110",
  15095=>"101000000",
  15096=>"111111000",
  15097=>"111111111",
  15098=>"111111000",
  15099=>"000000000",
  15100=>"100110001",
  15101=>"111110100",
  15102=>"000010001",
  15103=>"000000000",
  15104=>"000000000",
  15105=>"000011011",
  15106=>"111101001",
  15107=>"000000111",
  15108=>"000010110",
  15109=>"011001001",
  15110=>"001000101",
  15111=>"000100000",
  15112=>"100101110",
  15113=>"111111111",
  15114=>"000111111",
  15115=>"001001000",
  15116=>"000000000",
  15117=>"111111111",
  15118=>"111111000",
  15119=>"111111001",
  15120=>"101111110",
  15121=>"011001001",
  15122=>"000100000",
  15123=>"100110100",
  15124=>"011000000",
  15125=>"111000000",
  15126=>"011001001",
  15127=>"111001001",
  15128=>"111111000",
  15129=>"111111111",
  15130=>"000000111",
  15131=>"010000001",
  15132=>"111111110",
  15133=>"001011111",
  15134=>"011111111",
  15135=>"000001111",
  15136=>"110110001",
  15137=>"111111111",
  15138=>"000111111",
  15139=>"110000000",
  15140=>"011111111",
  15141=>"001000000",
  15142=>"111111100",
  15143=>"111111111",
  15144=>"110000001",
  15145=>"100100001",
  15146=>"000001001",
  15147=>"000111111",
  15148=>"000101101",
  15149=>"000100111",
  15150=>"101111111",
  15151=>"111000000",
  15152=>"110111010",
  15153=>"111111100",
  15154=>"111001000",
  15155=>"111100000",
  15156=>"000011000",
  15157=>"101000000",
  15158=>"000000001",
  15159=>"110011111",
  15160=>"011011000",
  15161=>"111000000",
  15162=>"111001000",
  15163=>"111111111",
  15164=>"001001001",
  15165=>"000000011",
  15166=>"110100100",
  15167=>"100000001",
  15168=>"000010000",
  15169=>"111000000",
  15170=>"011111111",
  15171=>"111001011",
  15172=>"111001000",
  15173=>"000000000",
  15174=>"000000000",
  15175=>"111011000",
  15176=>"000000000",
  15177=>"000001111",
  15178=>"000001011",
  15179=>"000110000",
  15180=>"000000000",
  15181=>"001111111",
  15182=>"000000110",
  15183=>"010110110",
  15184=>"010111110",
  15185=>"110000000",
  15186=>"000011111",
  15187=>"101000101",
  15188=>"000000100",
  15189=>"111100001",
  15190=>"011111111",
  15191=>"111111101",
  15192=>"000000000",
  15193=>"000010001",
  15194=>"111111111",
  15195=>"110111100",
  15196=>"000010100",
  15197=>"111101000",
  15198=>"000100000",
  15199=>"111011000",
  15200=>"001001101",
  15201=>"000111111",
  15202=>"010000000",
  15203=>"000000000",
  15204=>"000111100",
  15205=>"000000000",
  15206=>"000000000",
  15207=>"100000111",
  15208=>"001001011",
  15209=>"000111111",
  15210=>"111101111",
  15211=>"100111111",
  15212=>"000111111",
  15213=>"111000000",
  15214=>"111111111",
  15215=>"001000000",
  15216=>"011000000",
  15217=>"111110110",
  15218=>"000000111",
  15219=>"111111101",
  15220=>"111111000",
  15221=>"111000111",
  15222=>"011111111",
  15223=>"001000001",
  15224=>"000111100",
  15225=>"111111111",
  15226=>"011000000",
  15227=>"111100000",
  15228=>"000000001",
  15229=>"111100111",
  15230=>"111000000",
  15231=>"100000111",
  15232=>"000000000",
  15233=>"100110111",
  15234=>"110100000",
  15235=>"000000111",
  15236=>"000010111",
  15237=>"010000000",
  15238=>"000011011",
  15239=>"011000000",
  15240=>"000000000",
  15241=>"111101001",
  15242=>"010000000",
  15243=>"111111111",
  15244=>"111111111",
  15245=>"111000001",
  15246=>"000001000",
  15247=>"111111001",
  15248=>"100111111",
  15249=>"001011111",
  15250=>"111111111",
  15251=>"000100110",
  15252=>"111001101",
  15253=>"010000000",
  15254=>"010000000",
  15255=>"100001001",
  15256=>"110000000",
  15257=>"110111111",
  15258=>"000000000",
  15259=>"111111111",
  15260=>"000000000",
  15261=>"101111000",
  15262=>"100000101",
  15263=>"000111111",
  15264=>"000100000",
  15265=>"100011011",
  15266=>"011111111",
  15267=>"000000000",
  15268=>"000000000",
  15269=>"000111111",
  15270=>"000000000",
  15271=>"011011000",
  15272=>"010000000",
  15273=>"111111111",
  15274=>"011111001",
  15275=>"111111001",
  15276=>"111101100",
  15277=>"011001000",
  15278=>"000010010",
  15279=>"000111111",
  15280=>"000000000",
  15281=>"111101101",
  15282=>"001000000",
  15283=>"111100110",
  15284=>"000000000",
  15285=>"001001001",
  15286=>"000000011",
  15287=>"000000000",
  15288=>"000000000",
  15289=>"001111111",
  15290=>"111111100",
  15291=>"110111111",
  15292=>"011000000",
  15293=>"010010000",
  15294=>"011000000",
  15295=>"001001000",
  15296=>"110111000",
  15297=>"100000000",
  15298=>"000000000",
  15299=>"001000111",
  15300=>"111000000",
  15301=>"100100000",
  15302=>"000000000",
  15303=>"111110010",
  15304=>"000100010",
  15305=>"000000000",
  15306=>"110111001",
  15307=>"000000110",
  15308=>"100000000",
  15309=>"000010110",
  15310=>"000000001",
  15311=>"000010111",
  15312=>"000010111",
  15313=>"111000011",
  15314=>"101000000",
  15315=>"111100101",
  15316=>"000011111",
  15317=>"100111110",
  15318=>"100100110",
  15319=>"000000000",
  15320=>"100000000",
  15321=>"001111101",
  15322=>"111111111",
  15323=>"100100111",
  15324=>"111111000",
  15325=>"001111000",
  15326=>"111111111",
  15327=>"110110010",
  15328=>"111000000",
  15329=>"001000000",
  15330=>"111000000",
  15331=>"000000111",
  15332=>"000100111",
  15333=>"101000000",
  15334=>"001001000",
  15335=>"000000000",
  15336=>"000000000",
  15337=>"011111111",
  15338=>"000010111",
  15339=>"111101000",
  15340=>"001011111",
  15341=>"011010000",
  15342=>"000000000",
  15343=>"010000010",
  15344=>"111000000",
  15345=>"010000000",
  15346=>"001000111",
  15347=>"001000000",
  15348=>"000000000",
  15349=>"100000000",
  15350=>"111010000",
  15351=>"100010111",
  15352=>"000000111",
  15353=>"010010010",
  15354=>"011001111",
  15355=>"000111111",
  15356=>"000000000",
  15357=>"000111111",
  15358=>"000000111",
  15359=>"001011011",
  15360=>"011111111",
  15361=>"000000000",
  15362=>"000000110",
  15363=>"111000000",
  15364=>"000000110",
  15365=>"110110000",
  15366=>"100111111",
  15367=>"111111111",
  15368=>"111111001",
  15369=>"000000111",
  15370=>"000000001",
  15371=>"000000100",
  15372=>"100110110",
  15373=>"100000101",
  15374=>"100000000",
  15375=>"111001000",
  15376=>"111111111",
  15377=>"000000111",
  15378=>"000101111",
  15379=>"111110111",
  15380=>"000000011",
  15381=>"111000000",
  15382=>"111001000",
  15383=>"000011111",
  15384=>"100111111",
  15385=>"000110111",
  15386=>"100000111",
  15387=>"111100000",
  15388=>"000000010",
  15389=>"110111111",
  15390=>"000011111",
  15391=>"111111011",
  15392=>"000000000",
  15393=>"000000110",
  15394=>"111111000",
  15395=>"100110111",
  15396=>"000000110",
  15397=>"000101000",
  15398=>"000100001",
  15399=>"000000000",
  15400=>"000100010",
  15401=>"111111111",
  15402=>"001000001",
  15403=>"100100111",
  15404=>"111000000",
  15405=>"111111111",
  15406=>"100110111",
  15407=>"000101111",
  15408=>"111111111",
  15409=>"000000000",
  15410=>"011010011",
  15411=>"100100110",
  15412=>"001011011",
  15413=>"000011001",
  15414=>"000000000",
  15415=>"110110101",
  15416=>"000000111",
  15417=>"000000111",
  15418=>"111111111",
  15419=>"111000000",
  15420=>"000000000",
  15421=>"001000000",
  15422=>"000000111",
  15423=>"111111111",
  15424=>"011000000",
  15425=>"111001001",
  15426=>"000000001",
  15427=>"011111001",
  15428=>"110110110",
  15429=>"000000000",
  15430=>"000000100",
  15431=>"000001001",
  15432=>"011111011",
  15433=>"000000111",
  15434=>"100111010",
  15435=>"111101111",
  15436=>"000000110",
  15437=>"100110100",
  15438=>"110111110",
  15439=>"000000111",
  15440=>"111111111",
  15441=>"000000000",
  15442=>"110110010",
  15443=>"000110110",
  15444=>"000011111",
  15445=>"100000000",
  15446=>"000000000",
  15447=>"000000000",
  15448=>"000001111",
  15449=>"111111111",
  15450=>"010110100",
  15451=>"100011011",
  15452=>"100011111",
  15453=>"111110111",
  15454=>"001000001",
  15455=>"111111011",
  15456=>"000011000",
  15457=>"100110000",
  15458=>"000000000",
  15459=>"000000000",
  15460=>"000110000",
  15461=>"111111111",
  15462=>"000110110",
  15463=>"011111111",
  15464=>"111000000",
  15465=>"111001000",
  15466=>"001000100",
  15467=>"001001001",
  15468=>"001101111",
  15469=>"111111010",
  15470=>"110100000",
  15471=>"000000000",
  15472=>"000001011",
  15473=>"000000111",
  15474=>"001011011",
  15475=>"000001001",
  15476=>"001000111",
  15477=>"000111011",
  15478=>"110000000",
  15479=>"000000111",
  15480=>"000000000",
  15481=>"001101111",
  15482=>"111101100",
  15483=>"110110100",
  15484=>"100100100",
  15485=>"110111111",
  15486=>"000000001",
  15487=>"000000000",
  15488=>"000000110",
  15489=>"000000000",
  15490=>"001111111",
  15491=>"111111000",
  15492=>"000000001",
  15493=>"111000000",
  15494=>"111111001",
  15495=>"111111000",
  15496=>"000000111",
  15497=>"111111101",
  15498=>"111111111",
  15499=>"001001111",
  15500=>"111111000",
  15501=>"000000001",
  15502=>"100100111",
  15503=>"000111111",
  15504=>"001000011",
  15505=>"100001011",
  15506=>"010000000",
  15507=>"110011001",
  15508=>"000001011",
  15509=>"000100100",
  15510=>"000000000",
  15511=>"000000000",
  15512=>"111000001",
  15513=>"000000110",
  15514=>"111111100",
  15515=>"010100001",
  15516=>"000000001",
  15517=>"100000000",
  15518=>"000111111",
  15519=>"111111110",
  15520=>"111011111",
  15521=>"010111111",
  15522=>"000000000",
  15523=>"000000000",
  15524=>"111101111",
  15525=>"101111110",
  15526=>"111111111",
  15527=>"000101000",
  15528=>"000010111",
  15529=>"000000000",
  15530=>"000000111",
  15531=>"111111111",
  15532=>"000000000",
  15533=>"000011111",
  15534=>"100110101",
  15535=>"110011001",
  15536=>"000000001",
  15537=>"101111101",
  15538=>"111111011",
  15539=>"010000000",
  15540=>"100100000",
  15541=>"111111000",
  15542=>"000010000",
  15543=>"100111111",
  15544=>"011000000",
  15545=>"111111111",
  15546=>"000000000",
  15547=>"111101000",
  15548=>"000000000",
  15549=>"000001101",
  15550=>"111111111",
  15551=>"111000111",
  15552=>"111110000",
  15553=>"111111111",
  15554=>"000000110",
  15555=>"000000000",
  15556=>"000000111",
  15557=>"111111111",
  15558=>"000111000",
  15559=>"100000000",
  15560=>"111011000",
  15561=>"100111111",
  15562=>"110111011",
  15563=>"111111111",
  15564=>"111111011",
  15565=>"010011000",
  15566=>"111111000",
  15567=>"000001111",
  15568=>"000000000",
  15569=>"001001000",
  15570=>"000000000",
  15571=>"100100111",
  15572=>"010010000",
  15573=>"000100111",
  15574=>"000000000",
  15575=>"000111111",
  15576=>"000001000",
  15577=>"000000111",
  15578=>"100000000",
  15579=>"000000000",
  15580=>"000000000",
  15581=>"000000101",
  15582=>"111011000",
  15583=>"000100101",
  15584=>"110100000",
  15585=>"000110000",
  15586=>"111111111",
  15587=>"111111111",
  15588=>"110111111",
  15589=>"111110000",
  15590=>"000000001",
  15591=>"111111000",
  15592=>"111010000",
  15593=>"000000111",
  15594=>"111111000",
  15595=>"001000101",
  15596=>"111111000",
  15597=>"111001000",
  15598=>"000100111",
  15599=>"111111110",
  15600=>"100000000",
  15601=>"000000000",
  15602=>"000011001",
  15603=>"000010000",
  15604=>"111111111",
  15605=>"110100010",
  15606=>"000001111",
  15607=>"111000000",
  15608=>"111111111",
  15609=>"001000000",
  15610=>"111111111",
  15611=>"110100000",
  15612=>"100101111",
  15613=>"100001111",
  15614=>"000000000",
  15615=>"000000000",
  15616=>"111111111",
  15617=>"000000000",
  15618=>"111111011",
  15619=>"111101111",
  15620=>"000000110",
  15621=>"001000000",
  15622=>"001111111",
  15623=>"000000000",
  15624=>"111111010",
  15625=>"100101101",
  15626=>"111111111",
  15627=>"111111010",
  15628=>"100101111",
  15629=>"111000000",
  15630=>"000000111",
  15631=>"000000000",
  15632=>"111101111",
  15633=>"100111101",
  15634=>"111111111",
  15635=>"111100111",
  15636=>"010111111",
  15637=>"100111111",
  15638=>"100111011",
  15639=>"100100100",
  15640=>"111111011",
  15641=>"000000111",
  15642=>"100000000",
  15643=>"010011000",
  15644=>"100000111",
  15645=>"111100111",
  15646=>"000000111",
  15647=>"000010010",
  15648=>"000001000",
  15649=>"111111111",
  15650=>"010000100",
  15651=>"111111110",
  15652=>"110100100",
  15653=>"111111111",
  15654=>"000011111",
  15655=>"111111110",
  15656=>"110101111",
  15657=>"000000011",
  15658=>"111111001",
  15659=>"101101101",
  15660=>"110000000",
  15661=>"100110110",
  15662=>"100000011",
  15663=>"000000001",
  15664=>"000001111",
  15665=>"110110111",
  15666=>"000000111",
  15667=>"000000000",
  15668=>"000010110",
  15669=>"111111111",
  15670=>"000001111",
  15671=>"000000000",
  15672=>"110111111",
  15673=>"111100110",
  15674=>"000000001",
  15675=>"111110111",
  15676=>"000000000",
  15677=>"000010010",
  15678=>"110100000",
  15679=>"100000000",
  15680=>"101111111",
  15681=>"111111000",
  15682=>"111111000",
  15683=>"111111111",
  15684=>"000011111",
  15685=>"111100111",
  15686=>"101111111",
  15687=>"000000000",
  15688=>"000000000",
  15689=>"010110100",
  15690=>"000111010",
  15691=>"000000111",
  15692=>"111111101",
  15693=>"111111000",
  15694=>"000110000",
  15695=>"001001000",
  15696=>"011011011",
  15697=>"000000000",
  15698=>"000111111",
  15699=>"111111111",
  15700=>"000111111",
  15701=>"011001001",
  15702=>"000000000",
  15703=>"010001111",
  15704=>"100100111",
  15705=>"000000000",
  15706=>"000000000",
  15707=>"001000100",
  15708=>"000000001",
  15709=>"000000000",
  15710=>"000011011",
  15711=>"111111111",
  15712=>"111111111",
  15713=>"111000001",
  15714=>"000111111",
  15715=>"000000000",
  15716=>"000000000",
  15717=>"000000000",
  15718=>"000000000",
  15719=>"000000000",
  15720=>"111011011",
  15721=>"001001001",
  15722=>"111111111",
  15723=>"011111111",
  15724=>"111111000",
  15725=>"000000111",
  15726=>"111111000",
  15727=>"000001001",
  15728=>"000001111",
  15729=>"000000001",
  15730=>"000000000",
  15731=>"111111000",
  15732=>"000011001",
  15733=>"000000000",
  15734=>"111111110",
  15735=>"000000000",
  15736=>"000010001",
  15737=>"000000100",
  15738=>"000000000",
  15739=>"011001111",
  15740=>"000000110",
  15741=>"101001001",
  15742=>"011001000",
  15743=>"111111111",
  15744=>"110111100",
  15745=>"111111111",
  15746=>"000000000",
  15747=>"000000101",
  15748=>"000010000",
  15749=>"000000000",
  15750=>"111110000",
  15751=>"011111111",
  15752=>"000000000",
  15753=>"111011111",
  15754=>"000000000",
  15755=>"011011011",
  15756=>"111111111",
  15757=>"100110000",
  15758=>"111111110",
  15759=>"111111111",
  15760=>"000000000",
  15761=>"000000011",
  15762=>"111011011",
  15763=>"100000111",
  15764=>"111010000",
  15765=>"000011000",
  15766=>"111000100",
  15767=>"000000110",
  15768=>"100111111",
  15769=>"110000000",
  15770=>"111110110",
  15771=>"100111011",
  15772=>"100000001",
  15773=>"011000000",
  15774=>"000000100",
  15775=>"110111001",
  15776=>"111111111",
  15777=>"000000000",
  15778=>"111111001",
  15779=>"000100100",
  15780=>"111111101",
  15781=>"000110110",
  15782=>"000000111",
  15783=>"011000011",
  15784=>"111111001",
  15785=>"000000100",
  15786=>"111111011",
  15787=>"000011010",
  15788=>"000000000",
  15789=>"100100100",
  15790=>"000000111",
  15791=>"000000010",
  15792=>"111000000",
  15793=>"000000000",
  15794=>"000000000",
  15795=>"000000000",
  15796=>"101000000",
  15797=>"001000000",
  15798=>"000000011",
  15799=>"011001111",
  15800=>"000000000",
  15801=>"000000000",
  15802=>"110010000",
  15803=>"111000000",
  15804=>"000000100",
  15805=>"000000000",
  15806=>"110111111",
  15807=>"111111001",
  15808=>"111111011",
  15809=>"111111011",
  15810=>"111111111",
  15811=>"000000000",
  15812=>"110110000",
  15813=>"000000000",
  15814=>"101101111",
  15815=>"111111001",
  15816=>"001001001",
  15817=>"101100111",
  15818=>"000101111",
  15819=>"000000000",
  15820=>"010111110",
  15821=>"011001000",
  15822=>"101001001",
  15823=>"000000000",
  15824=>"000111011",
  15825=>"111111101",
  15826=>"001101111",
  15827=>"011000000",
  15828=>"000000000",
  15829=>"111111111",
  15830=>"000000110",
  15831=>"111111011",
  15832=>"000000001",
  15833=>"111010000",
  15834=>"011001000",
  15835=>"000000001",
  15836=>"100110111",
  15837=>"001011000",
  15838=>"110111011",
  15839=>"111000000",
  15840=>"001101001",
  15841=>"111111101",
  15842=>"001000000",
  15843=>"100111010",
  15844=>"000000000",
  15845=>"111111001",
  15846=>"000000111",
  15847=>"100000000",
  15848=>"000000000",
  15849=>"111010000",
  15850=>"111111111",
  15851=>"100101101",
  15852=>"100101000",
  15853=>"001000110",
  15854=>"111001001",
  15855=>"100100111",
  15856=>"000000100",
  15857=>"000000000",
  15858=>"110111111",
  15859=>"001000011",
  15860=>"111111010",
  15861=>"111100110",
  15862=>"111111111",
  15863=>"110000000",
  15864=>"010000001",
  15865=>"001001111",
  15866=>"000000000",
  15867=>"101100110",
  15868=>"010010011",
  15869=>"110111100",
  15870=>"001111111",
  15871=>"001001011",
  15872=>"000000000",
  15873=>"001001011",
  15874=>"111111101",
  15875=>"001011011",
  15876=>"000000000",
  15877=>"111111010",
  15878=>"000000000",
  15879=>"000000000",
  15880=>"111111111",
  15881=>"000000110",
  15882=>"111111001",
  15883=>"100000100",
  15884=>"000000000",
  15885=>"011001000",
  15886=>"000000000",
  15887=>"000100111",
  15888=>"000000100",
  15889=>"000000000",
  15890=>"111111111",
  15891=>"111111101",
  15892=>"111101111",
  15893=>"111111111",
  15894=>"110110000",
  15895=>"111111111",
  15896=>"111111011",
  15897=>"000000000",
  15898=>"100000000",
  15899=>"111101000",
  15900=>"111000001",
  15901=>"111111100",
  15902=>"111110000",
  15903=>"110110111",
  15904=>"111111111",
  15905=>"111111001",
  15906=>"001111100",
  15907=>"000100100",
  15908=>"000000000",
  15909=>"000001001",
  15910=>"011011000",
  15911=>"111111111",
  15912=>"111111111",
  15913=>"101000111",
  15914=>"011001000",
  15915=>"000000000",
  15916=>"111111111",
  15917=>"000000111",
  15918=>"000000000",
  15919=>"111000001",
  15920=>"000000100",
  15921=>"000000100",
  15922=>"100100000",
  15923=>"111111111",
  15924=>"000000000",
  15925=>"011011000",
  15926=>"000000000",
  15927=>"000100111",
  15928=>"111111111",
  15929=>"011000110",
  15930=>"000000000",
  15931=>"000000111",
  15932=>"100000000",
  15933=>"110111000",
  15934=>"000011011",
  15935=>"001111111",
  15936=>"011000101",
  15937=>"110110111",
  15938=>"000000000",
  15939=>"000000111",
  15940=>"110100000",
  15941=>"011011111",
  15942=>"000000111",
  15943=>"111111111",
  15944=>"000000000",
  15945=>"000000000",
  15946=>"001111000",
  15947=>"000000000",
  15948=>"000000011",
  15949=>"100000111",
  15950=>"000000000",
  15951=>"111111111",
  15952=>"111111111",
  15953=>"111111101",
  15954=>"000011011",
  15955=>"000000100",
  15956=>"000010000",
  15957=>"111111100",
  15958=>"101001000",
  15959=>"111110101",
  15960=>"111111111",
  15961=>"000001011",
  15962=>"010111111",
  15963=>"111111110",
  15964=>"000000000",
  15965=>"111111111",
  15966=>"110110111",
  15967=>"000000000",
  15968=>"000000000",
  15969=>"000000000",
  15970=>"111111111",
  15971=>"111111111",
  15972=>"000001000",
  15973=>"000000101",
  15974=>"000000011",
  15975=>"001000000",
  15976=>"111111111",
  15977=>"101000000",
  15978=>"100101000",
  15979=>"010110010",
  15980=>"000100110",
  15981=>"001001000",
  15982=>"000000001",
  15983=>"101001101",
  15984=>"111000000",
  15985=>"000111111",
  15986=>"111111111",
  15987=>"011011110",
  15988=>"011111111",
  15989=>"011011011",
  15990=>"001001011",
  15991=>"111011000",
  15992=>"111111111",
  15993=>"000000000",
  15994=>"000000000",
  15995=>"011000000",
  15996=>"000100100",
  15997=>"111111111",
  15998=>"000000000",
  15999=>"111000000",
  16000=>"111111011",
  16001=>"111100000",
  16002=>"000000000",
  16003=>"011011011",
  16004=>"110100100",
  16005=>"000001111",
  16006=>"000000000",
  16007=>"100111111",
  16008=>"000000000",
  16009=>"011111111",
  16010=>"011000000",
  16011=>"111011000",
  16012=>"111111111",
  16013=>"000000000",
  16014=>"000100110",
  16015=>"100111111",
  16016=>"000000011",
  16017=>"011110011",
  16018=>"111000000",
  16019=>"000011011",
  16020=>"000000000",
  16021=>"001001000",
  16022=>"111111111",
  16023=>"000111111",
  16024=>"001111111",
  16025=>"111111111",
  16026=>"111000100",
  16027=>"000100000",
  16028=>"100100111",
  16029=>"000001011",
  16030=>"000110000",
  16031=>"000000000",
  16032=>"111111111",
  16033=>"001111000",
  16034=>"111111000",
  16035=>"111111111",
  16036=>"000000100",
  16037=>"111111100",
  16038=>"111011011",
  16039=>"000010011",
  16040=>"000110111",
  16041=>"111111111",
  16042=>"011000000",
  16043=>"000000000",
  16044=>"111111111",
  16045=>"001001011",
  16046=>"000100000",
  16047=>"000000011",
  16048=>"000000000",
  16049=>"000010111",
  16050=>"111100111",
  16051=>"000000000",
  16052=>"111111000",
  16053=>"000000000",
  16054=>"000000000",
  16055=>"000000000",
  16056=>"000101001",
  16057=>"000000000",
  16058=>"010111000",
  16059=>"011110010",
  16060=>"111111101",
  16061=>"001000000",
  16062=>"000000000",
  16063=>"000000000",
  16064=>"111111111",
  16065=>"111001000",
  16066=>"000000000",
  16067=>"001011010",
  16068=>"111000000",
  16069=>"110100100",
  16070=>"000100001",
  16071=>"000000000",
  16072=>"000000000",
  16073=>"111111111",
  16074=>"111111110",
  16075=>"111111111",
  16076=>"000000000",
  16077=>"000001000",
  16078=>"111111111",
  16079=>"000000000",
  16080=>"000000000",
  16081=>"000000000",
  16082=>"000000000",
  16083=>"111111111",
  16084=>"000000001",
  16085=>"111111111",
  16086=>"000000000",
  16087=>"001101111",
  16088=>"001001000",
  16089=>"011111001",
  16090=>"111111111",
  16091=>"111111111",
  16092=>"001101000",
  16093=>"111011001",
  16094=>"110111111",
  16095=>"000111111",
  16096=>"000000001",
  16097=>"000000111",
  16098=>"111111111",
  16099=>"000110000",
  16100=>"000000000",
  16101=>"111111111",
  16102=>"111111111",
  16103=>"000000000",
  16104=>"111011011",
  16105=>"001000111",
  16106=>"111110110",
  16107=>"100000000",
  16108=>"001010011",
  16109=>"111111111",
  16110=>"111011000",
  16111=>"111111000",
  16112=>"111110111",
  16113=>"111111111",
  16114=>"111110111",
  16115=>"101000101",
  16116=>"000000101",
  16117=>"001001000",
  16118=>"000000000",
  16119=>"111111111",
  16120=>"111111000",
  16121=>"000000000",
  16122=>"110111110",
  16123=>"000111101",
  16124=>"111111011",
  16125=>"111011001",
  16126=>"101111111",
  16127=>"000000000",
  16128=>"000010111",
  16129=>"111110111",
  16130=>"011110111",
  16131=>"111001101",
  16132=>"111111111",
  16133=>"111101000",
  16134=>"101111111",
  16135=>"001111111",
  16136=>"111111001",
  16137=>"000000000",
  16138=>"001000011",
  16139=>"111111100",
  16140=>"001000100",
  16141=>"000001001",
  16142=>"111111010",
  16143=>"100111111",
  16144=>"000001111",
  16145=>"111111111",
  16146=>"011000100",
  16147=>"111111000",
  16148=>"101000000",
  16149=>"000000111",
  16150=>"000000001",
  16151=>"111111111",
  16152=>"000000011",
  16153=>"000000000",
  16154=>"000000100",
  16155=>"110111111",
  16156=>"110110000",
  16157=>"000000000",
  16158=>"000000001",
  16159=>"111111111",
  16160=>"000001110",
  16161=>"000000000",
  16162=>"111111111",
  16163=>"110000001",
  16164=>"001111111",
  16165=>"111111111",
  16166=>"000000100",
  16167=>"111111111",
  16168=>"011111110",
  16169=>"101100111",
  16170=>"011110000",
  16171=>"111111111",
  16172=>"000000000",
  16173=>"011011011",
  16174=>"000000000",
  16175=>"000000000",
  16176=>"000000000",
  16177=>"000000000",
  16178=>"111110000",
  16179=>"000001111",
  16180=>"000000000",
  16181=>"000000110",
  16182=>"000000111",
  16183=>"000000111",
  16184=>"000000000",
  16185=>"111111000",
  16186=>"000000000",
  16187=>"000001001",
  16188=>"000001001",
  16189=>"111001001",
  16190=>"000000110",
  16191=>"111111000",
  16192=>"111111000",
  16193=>"010010001",
  16194=>"000000000",
  16195=>"000000000",
  16196=>"000000001",
  16197=>"000111111",
  16198=>"000100110",
  16199=>"000000000",
  16200=>"111111000",
  16201=>"111111111",
  16202=>"111111011",
  16203=>"111111011",
  16204=>"011111010",
  16205=>"100000000",
  16206=>"111111110",
  16207=>"011111111",
  16208=>"011000111",
  16209=>"111111001",
  16210=>"111111111",
  16211=>"111111111",
  16212=>"111011111",
  16213=>"011011011",
  16214=>"011001111",
  16215=>"111111111",
  16216=>"001001011",
  16217=>"111000001",
  16218=>"000000000",
  16219=>"111111111",
  16220=>"001000101",
  16221=>"000000111",
  16222=>"101100111",
  16223=>"000000001",
  16224=>"000000000",
  16225=>"000000111",
  16226=>"111111000",
  16227=>"100111111",
  16228=>"011001001",
  16229=>"000000000",
  16230=>"000000111",
  16231=>"111111011",
  16232=>"111111100",
  16233=>"000000000",
  16234=>"000000000",
  16235=>"000001001",
  16236=>"110000000",
  16237=>"010001001",
  16238=>"100000000",
  16239=>"011011000",
  16240=>"000000000",
  16241=>"111111001",
  16242=>"111111110",
  16243=>"001011011",
  16244=>"100101001",
  16245=>"001000001",
  16246=>"100011000",
  16247=>"100100100",
  16248=>"111111111",
  16249=>"011000111",
  16250=>"100000111",
  16251=>"000000000",
  16252=>"000000000",
  16253=>"000000000",
  16254=>"111111111",
  16255=>"000000111",
  16256=>"111111011",
  16257=>"111101000",
  16258=>"111111111",
  16259=>"111111111",
  16260=>"001001000",
  16261=>"000000011",
  16262=>"000110100",
  16263=>"111111111",
  16264=>"111010000",
  16265=>"100000000",
  16266=>"111111111",
  16267=>"010110111",
  16268=>"000000000",
  16269=>"011011001",
  16270=>"000000000",
  16271=>"000000001",
  16272=>"000000000",
  16273=>"111111000",
  16274=>"111111011",
  16275=>"000110000",
  16276=>"111111111",
  16277=>"000010110",
  16278=>"111111000",
  16279=>"000000000",
  16280=>"111001001",
  16281=>"011111111",
  16282=>"111111111",
  16283=>"101111111",
  16284=>"000111111",
  16285=>"000000001",
  16286=>"000000000",
  16287=>"101101111",
  16288=>"110010000",
  16289=>"100111111",
  16290=>"100111111",
  16291=>"011001100",
  16292=>"000111000",
  16293=>"100111111",
  16294=>"111001000",
  16295=>"111111000",
  16296=>"011011011",
  16297=>"001000111",
  16298=>"000110000",
  16299=>"000000000",
  16300=>"000000000",
  16301=>"111111000",
  16302=>"000000111",
  16303=>"000001001",
  16304=>"000000000",
  16305=>"000000000",
  16306=>"111100000",
  16307=>"111111111",
  16308=>"111111111",
  16309=>"100100100",
  16310=>"111111001",
  16311=>"000001111",
  16312=>"111001000",
  16313=>"111111000",
  16314=>"111011111",
  16315=>"101100100",
  16316=>"101111111",
  16317=>"110111101",
  16318=>"111100000",
  16319=>"000000000",
  16320=>"010110000",
  16321=>"111111111",
  16322=>"000000000",
  16323=>"001001000",
  16324=>"000001000",
  16325=>"010000000",
  16326=>"000000001",
  16327=>"000000000",
  16328=>"000000000",
  16329=>"000000111",
  16330=>"000000000",
  16331=>"000000000",
  16332=>"000000000",
  16333=>"100001111",
  16334=>"100000000",
  16335=>"110100000",
  16336=>"100000000",
  16337=>"011111111",
  16338=>"111111111",
  16339=>"000000001",
  16340=>"000000001",
  16341=>"000001001",
  16342=>"000000111",
  16343=>"010000000",
  16344=>"001000000",
  16345=>"111111000",
  16346=>"101000111",
  16347=>"000000000",
  16348=>"100001001",
  16349=>"000111111",
  16350=>"000100000",
  16351=>"011001001",
  16352=>"011011010",
  16353=>"001001000",
  16354=>"001000001",
  16355=>"111111110",
  16356=>"011001000",
  16357=>"000101101",
  16358=>"111010111",
  16359=>"000000100",
  16360=>"101000000",
  16361=>"001001111",
  16362=>"111000100",
  16363=>"111111111",
  16364=>"111111111",
  16365=>"110000110",
  16366=>"111000000",
  16367=>"000001101",
  16368=>"000000000",
  16369=>"100100111",
  16370=>"101001000",
  16371=>"111111111",
  16372=>"101111100",
  16373=>"000000000",
  16374=>"111111111",
  16375=>"111011011",
  16376=>"111111000",
  16377=>"000110110",
  16378=>"000000000",
  16379=>"000000000",
  16380=>"000000000",
  16381=>"111111111",
  16382=>"111111111",
  16383=>"000000000",
  16384=>"111111000",
  16385=>"000000000",
  16386=>"000100100",
  16387=>"111111111",
  16388=>"100111111",
  16389=>"010010010",
  16390=>"000000010",
  16391=>"001001000",
  16392=>"111101101",
  16393=>"000000000",
  16394=>"111000111",
  16395=>"011110111",
  16396=>"000000110",
  16397=>"001011111",
  16398=>"111111111",
  16399=>"001000000",
  16400=>"011000000",
  16401=>"001111111",
  16402=>"000000000",
  16403=>"000000000",
  16404=>"000000101",
  16405=>"001001111",
  16406=>"000000000",
  16407=>"100100111",
  16408=>"111111111",
  16409=>"100100001",
  16410=>"000000001",
  16411=>"110000001",
  16412=>"011111111",
  16413=>"111110111",
  16414=>"111111101",
  16415=>"011111111",
  16416=>"011000100",
  16417=>"001001011",
  16418=>"110000000",
  16419=>"011000000",
  16420=>"111011011",
  16421=>"000000000",
  16422=>"110100111",
  16423=>"000001001",
  16424=>"111111111",
  16425=>"000000000",
  16426=>"111110111",
  16427=>"111100000",
  16428=>"000000011",
  16429=>"000100100",
  16430=>"110110010",
  16431=>"111111111",
  16432=>"111111111",
  16433=>"000110010",
  16434=>"001000000",
  16435=>"000110101",
  16436=>"011010000",
  16437=>"000000100",
  16438=>"010000000",
  16439=>"000000000",
  16440=>"000000000",
  16441=>"111001000",
  16442=>"000000011",
  16443=>"100000000",
  16444=>"111111111",
  16445=>"011000100",
  16446=>"000010110",
  16447=>"000000000",
  16448=>"110110111",
  16449=>"000101111",
  16450=>"001000000",
  16451=>"010010111",
  16452=>"000001000",
  16453=>"000111111",
  16454=>"000000100",
  16455=>"000000000",
  16456=>"000000100",
  16457=>"001111111",
  16458=>"000000000",
  16459=>"001001111",
  16460=>"000011111",
  16461=>"001000000",
  16462=>"000000000",
  16463=>"000000000",
  16464=>"000000000",
  16465=>"000000000",
  16466=>"000000000",
  16467=>"001000100",
  16468=>"111111110",
  16469=>"110000000",
  16470=>"000110111",
  16471=>"110111111",
  16472=>"111111111",
  16473=>"000000000",
  16474=>"010111110",
  16475=>"000011011",
  16476=>"111001111",
  16477=>"000000000",
  16478=>"001000001",
  16479=>"111111111",
  16480=>"111101111",
  16481=>"111110110",
  16482=>"000100110",
  16483=>"011011111",
  16484=>"111111111",
  16485=>"111111111",
  16486=>"100111111",
  16487=>"000000110",
  16488=>"101001000",
  16489=>"000000100",
  16490=>"111111111",
  16491=>"000000000",
  16492=>"111111011",
  16493=>"000110111",
  16494=>"000001111",
  16495=>"111111100",
  16496=>"000111111",
  16497=>"000000000",
  16498=>"111011001",
  16499=>"111111111",
  16500=>"011011001",
  16501=>"111000000",
  16502=>"111111111",
  16503=>"111111111",
  16504=>"111111111",
  16505=>"000000000",
  16506=>"000000000",
  16507=>"111111111",
  16508=>"011010000",
  16509=>"111111111",
  16510=>"000000000",
  16511=>"110001111",
  16512=>"111111011",
  16513=>"111111100",
  16514=>"000000000",
  16515=>"111111111",
  16516=>"000001000",
  16517=>"000000000",
  16518=>"100100110",
  16519=>"000000000",
  16520=>"111111100",
  16521=>"000000000",
  16522=>"110100000",
  16523=>"011111111",
  16524=>"011111111",
  16525=>"111100110",
  16526=>"010000000",
  16527=>"000000000",
  16528=>"111111111",
  16529=>"111111111",
  16530=>"100111111",
  16531=>"111100000",
  16532=>"111011111",
  16533=>"101111110",
  16534=>"000000000",
  16535=>"010000010",
  16536=>"111000000",
  16537=>"111111111",
  16538=>"111111111",
  16539=>"111111111",
  16540=>"111111111",
  16541=>"111111100",
  16542=>"000000000",
  16543=>"000000000",
  16544=>"000000000",
  16545=>"001000000",
  16546=>"111111011",
  16547=>"101111011",
  16548=>"000010110",
  16549=>"111111000",
  16550=>"111111111",
  16551=>"111110000",
  16552=>"000001011",
  16553=>"111111001",
  16554=>"111101111",
  16555=>"101101000",
  16556=>"110100111",
  16557=>"011011011",
  16558=>"000001111",
  16559=>"110010000",
  16560=>"111000000",
  16561=>"001000000",
  16562=>"011011011",
  16563=>"011001000",
  16564=>"111111111",
  16565=>"110110010",
  16566=>"111111011",
  16567=>"111001000",
  16568=>"001111111",
  16569=>"000110000",
  16570=>"000010000",
  16571=>"111011011",
  16572=>"000000000",
  16573=>"111000000",
  16574=>"000000000",
  16575=>"000000000",
  16576=>"100100111",
  16577=>"101111001",
  16578=>"111111111",
  16579=>"111111111",
  16580=>"111001001",
  16581=>"111111000",
  16582=>"100110101",
  16583=>"000000001",
  16584=>"111111111",
  16585=>"000000001",
  16586=>"000000000",
  16587=>"000000000",
  16588=>"100000000",
  16589=>"111111100",
  16590=>"000000000",
  16591=>"000001100",
  16592=>"001000000",
  16593=>"000000000",
  16594=>"001111110",
  16595=>"000000000",
  16596=>"011111111",
  16597=>"000000110",
  16598=>"111011111",
  16599=>"100100100",
  16600=>"000110111",
  16601=>"000000000",
  16602=>"111011001",
  16603=>"101000001",
  16604=>"111111111",
  16605=>"111111111",
  16606=>"000000111",
  16607=>"111111000",
  16608=>"111111111",
  16609=>"000000100",
  16610=>"000010010",
  16611=>"110000000",
  16612=>"111001111",
  16613=>"110100100",
  16614=>"000000000",
  16615=>"111111011",
  16616=>"000000000",
  16617=>"011001001",
  16618=>"011000000",
  16619=>"000000000",
  16620=>"011001000",
  16621=>"001111111",
  16622=>"101111000",
  16623=>"001101000",
  16624=>"011001111",
  16625=>"000001001",
  16626=>"111111111",
  16627=>"000000000",
  16628=>"000000000",
  16629=>"111111111",
  16630=>"011000111",
  16631=>"000000000",
  16632=>"000000000",
  16633=>"111111000",
  16634=>"110000111",
  16635=>"101000000",
  16636=>"111000100",
  16637=>"000111011",
  16638=>"111001001",
  16639=>"111111111",
  16640=>"000000000",
  16641=>"011011011",
  16642=>"000000000",
  16643=>"110111111",
  16644=>"000100111",
  16645=>"111110111",
  16646=>"110111111",
  16647=>"000000111",
  16648=>"111101001",
  16649=>"110110110",
  16650=>"100100110",
  16651=>"111111111",
  16652=>"111110000",
  16653=>"100100100",
  16654=>"111011111",
  16655=>"000000000",
  16656=>"111111111",
  16657=>"000100101",
  16658=>"101100110",
  16659=>"000000000",
  16660=>"000000000",
  16661=>"000000111",
  16662=>"000000000",
  16663=>"011111011",
  16664=>"111111111",
  16665=>"000000000",
  16666=>"101101111",
  16667=>"000000000",
  16668=>"111011011",
  16669=>"000000000",
  16670=>"111111111",
  16671=>"000001101",
  16672=>"000100101",
  16673=>"000110110",
  16674=>"110111111",
  16675=>"100000000",
  16676=>"111000000",
  16677=>"000000111",
  16678=>"000000000",
  16679=>"000000000",
  16680=>"111111111",
  16681=>"000011000",
  16682=>"111111001",
  16683=>"000000100",
  16684=>"110100001",
  16685=>"000000100",
  16686=>"111111111",
  16687=>"000000000",
  16688=>"011011011",
  16689=>"000000000",
  16690=>"111000000",
  16691=>"000000000",
  16692=>"111111111",
  16693=>"000000000",
  16694=>"000000000",
  16695=>"111111111",
  16696=>"000111111",
  16697=>"000000000",
  16698=>"000111000",
  16699=>"111111110",
  16700=>"011001001",
  16701=>"000000111",
  16702=>"000000000",
  16703=>"100101111",
  16704=>"100000000",
  16705=>"111111111",
  16706=>"000001111",
  16707=>"000000111",
  16708=>"111000111",
  16709=>"100110110",
  16710=>"111001000",
  16711=>"000000011",
  16712=>"111000000",
  16713=>"000000000",
  16714=>"111000000",
  16715=>"011111111",
  16716=>"000000000",
  16717=>"111111111",
  16718=>"111010111",
  16719=>"111111111",
  16720=>"011011011",
  16721=>"111111110",
  16722=>"000000000",
  16723=>"111111111",
  16724=>"000000000",
  16725=>"000001110",
  16726=>"111100000",
  16727=>"000000000",
  16728=>"111111111",
  16729=>"111011011",
  16730=>"100000000",
  16731=>"111111111",
  16732=>"010000000",
  16733=>"000000000",
  16734=>"111111111",
  16735=>"000000000",
  16736=>"111111111",
  16737=>"000000000",
  16738=>"111111110",
  16739=>"111111110",
  16740=>"111100000",
  16741=>"000000000",
  16742=>"000000000",
  16743=>"111111111",
  16744=>"000001101",
  16745=>"111111111",
  16746=>"000000000",
  16747=>"001011111",
  16748=>"011111111",
  16749=>"000000000",
  16750=>"001001011",
  16751=>"000000000",
  16752=>"000001111",
  16753=>"111111111",
  16754=>"101100101",
  16755=>"000000000",
  16756=>"000000001",
  16757=>"100000011",
  16758=>"001000000",
  16759=>"000000000",
  16760=>"111000111",
  16761=>"000000000",
  16762=>"111111111",
  16763=>"000000011",
  16764=>"010000100",
  16765=>"100100001",
  16766=>"100101101",
  16767=>"000000011",
  16768=>"111111101",
  16769=>"000000000",
  16770=>"011011011",
  16771=>"000000000",
  16772=>"111100111",
  16773=>"111111111",
  16774=>"111101001",
  16775=>"000000000",
  16776=>"001011111",
  16777=>"110000000",
  16778=>"111111000",
  16779=>"111111110",
  16780=>"111111111",
  16781=>"111111111",
  16782=>"111111111",
  16783=>"110110111",
  16784=>"111111111",
  16785=>"111111110",
  16786=>"101001101",
  16787=>"100000001",
  16788=>"111111111",
  16789=>"101000000",
  16790=>"101100001",
  16791=>"011011101",
  16792=>"001111111",
  16793=>"111001001",
  16794=>"000000000",
  16795=>"000000101",
  16796=>"000000111",
  16797=>"000100000",
  16798=>"000000000",
  16799=>"011110000",
  16800=>"000100110",
  16801=>"001111111",
  16802=>"000001100",
  16803=>"111111111",
  16804=>"110100100",
  16805=>"100111111",
  16806=>"011111111",
  16807=>"000000110",
  16808=>"000011010",
  16809=>"010011000",
  16810=>"000000000",
  16811=>"000000000",
  16812=>"111101101",
  16813=>"100101011",
  16814=>"111111111",
  16815=>"000000000",
  16816=>"111111001",
  16817=>"111110110",
  16818=>"011011001",
  16819=>"110111111",
  16820=>"000000000",
  16821=>"000010011",
  16822=>"000000000",
  16823=>"111111000",
  16824=>"001000000",
  16825=>"000000111",
  16826=>"100000000",
  16827=>"001001000",
  16828=>"110000110",
  16829=>"101000000",
  16830=>"000000000",
  16831=>"011011000",
  16832=>"000000000",
  16833=>"111111111",
  16834=>"000010000",
  16835=>"111111010",
  16836=>"110111111",
  16837=>"011011111",
  16838=>"000000100",
  16839=>"111111111",
  16840=>"000000000",
  16841=>"100000000",
  16842=>"000000000",
  16843=>"011110110",
  16844=>"111111111",
  16845=>"111111100",
  16846=>"100101001",
  16847=>"111111111",
  16848=>"001000000",
  16849=>"000000000",
  16850=>"001111111",
  16851=>"111111111",
  16852=>"111011111",
  16853=>"111111111",
  16854=>"111111111",
  16855=>"001011011",
  16856=>"111111011",
  16857=>"111111110",
  16858=>"011111111",
  16859=>"111001001",
  16860=>"111111111",
  16861=>"000000000",
  16862=>"000000111",
  16863=>"011111101",
  16864=>"000000000",
  16865=>"111101101",
  16866=>"000000000",
  16867=>"111111000",
  16868=>"111000111",
  16869=>"111111001",
  16870=>"111111111",
  16871=>"000100110",
  16872=>"010010000",
  16873=>"000000000",
  16874=>"001111111",
  16875=>"000010000",
  16876=>"011000000",
  16877=>"110111011",
  16878=>"010000000",
  16879=>"000000111",
  16880=>"000000000",
  16881=>"000010111",
  16882=>"111111111",
  16883=>"000000000",
  16884=>"110000000",
  16885=>"111111111",
  16886=>"111110110",
  16887=>"101100000",
  16888=>"011111111",
  16889=>"100000000",
  16890=>"111111111",
  16891=>"000000000",
  16892=>"100000000",
  16893=>"000101111",
  16894=>"000001001",
  16895=>"000110110",
  16896=>"000000000",
  16897=>"000000000",
  16898=>"000000111",
  16899=>"101111111",
  16900=>"100111111",
  16901=>"111110000",
  16902=>"110010111",
  16903=>"111111111",
  16904=>"111111111",
  16905=>"111110111",
  16906=>"100111111",
  16907=>"111111111",
  16908=>"100100100",
  16909=>"111000000",
  16910=>"111001011",
  16911=>"111001000",
  16912=>"110111110",
  16913=>"111111111",
  16914=>"100000000",
  16915=>"000000000",
  16916=>"111111000",
  16917=>"111100110",
  16918=>"000000010",
  16919=>"111000000",
  16920=>"111000000",
  16921=>"111001111",
  16922=>"100111111",
  16923=>"100100100",
  16924=>"111100110",
  16925=>"111111111",
  16926=>"010010011",
  16927=>"000111111",
  16928=>"111111100",
  16929=>"010111110",
  16930=>"011000111",
  16931=>"000110000",
  16932=>"101111011",
  16933=>"000100101",
  16934=>"000111110",
  16935=>"001111111",
  16936=>"110111111",
  16937=>"100111111",
  16938=>"011111111",
  16939=>"000000000",
  16940=>"000000000",
  16941=>"111111111",
  16942=>"111111111",
  16943=>"111000010",
  16944=>"111111111",
  16945=>"000001001",
  16946=>"001001001",
  16947=>"000101000",
  16948=>"000100111",
  16949=>"001111110",
  16950=>"000000000",
  16951=>"000000000",
  16952=>"111111110",
  16953=>"000001001",
  16954=>"000000000",
  16955=>"110100000",
  16956=>"001000000",
  16957=>"000000111",
  16958=>"110000000",
  16959=>"111111000",
  16960=>"100000111",
  16961=>"000000110",
  16962=>"000000000",
  16963=>"001000000",
  16964=>"000000000",
  16965=>"111111111",
  16966=>"000000000",
  16967=>"111101111",
  16968=>"011111011",
  16969=>"001101111",
  16970=>"000000000",
  16971=>"100100101",
  16972=>"011000100",
  16973=>"110000000",
  16974=>"000000000",
  16975=>"011001001",
  16976=>"101101011",
  16977=>"011010001",
  16978=>"101111110",
  16979=>"000000000",
  16980=>"000000111",
  16981=>"000000000",
  16982=>"001101111",
  16983=>"000000000",
  16984=>"111111110",
  16985=>"000000000",
  16986=>"000000011",
  16987=>"110110111",
  16988=>"100000111",
  16989=>"000100111",
  16990=>"111111111",
  16991=>"011111111",
  16992=>"000000111",
  16993=>"111000000",
  16994=>"001001001",
  16995=>"000000000",
  16996=>"111110000",
  16997=>"111111011",
  16998=>"000000000",
  16999=>"111100000",
  17000=>"111111111",
  17001=>"000110110",
  17002=>"000000000",
  17003=>"111111110",
  17004=>"000000000",
  17005=>"111111111",
  17006=>"000000000",
  17007=>"000000110",
  17008=>"000000001",
  17009=>"000000111",
  17010=>"000001111",
  17011=>"001001000",
  17012=>"000001111",
  17013=>"000000000",
  17014=>"000000000",
  17015=>"101111111",
  17016=>"000000000",
  17017=>"000000000",
  17018=>"111100100",
  17019=>"000000000",
  17020=>"000000000",
  17021=>"000000000",
  17022=>"101000110",
  17023=>"000000000",
  17024=>"111110000",
  17025=>"111111110",
  17026=>"111110111",
  17027=>"001001001",
  17028=>"111000000",
  17029=>"111111111",
  17030=>"110110000",
  17031=>"000011000",
  17032=>"111111000",
  17033=>"111000000",
  17034=>"011001111",
  17035=>"000000000",
  17036=>"111111111",
  17037=>"000000000",
  17038=>"111111110",
  17039=>"000001001",
  17040=>"000111010",
  17041=>"000000000",
  17042=>"111111000",
  17043=>"001000000",
  17044=>"000000000",
  17045=>"000000000",
  17046=>"000111111",
  17047=>"010000000",
  17048=>"000000110",
  17049=>"000000000",
  17050=>"000111111",
  17051=>"111111111",
  17052=>"000000000",
  17053=>"101100110",
  17054=>"000000101",
  17055=>"010010100",
  17056=>"000000001",
  17057=>"000000000",
  17058=>"111111000",
  17059=>"110000111",
  17060=>"100000001",
  17061=>"111111110",
  17062=>"111000000",
  17063=>"000001011",
  17064=>"011000000",
  17065=>"000000000",
  17066=>"110000000",
  17067=>"111110111",
  17068=>"001000001",
  17069=>"111010000",
  17070=>"000000111",
  17071=>"110111001",
  17072=>"000000000",
  17073=>"111111110",
  17074=>"111111000",
  17075=>"011000000",
  17076=>"111111110",
  17077=>"111000111",
  17078=>"101111011",
  17079=>"100000000",
  17080=>"000100111",
  17081=>"000000001",
  17082=>"111000110",
  17083=>"111111110",
  17084=>"000000001",
  17085=>"000000010",
  17086=>"000000000",
  17087=>"101111111",
  17088=>"000010000",
  17089=>"000100000",
  17090=>"000000000",
  17091=>"000001000",
  17092=>"000100000",
  17093=>"000111111",
  17094=>"111100000",
  17095=>"000000111",
  17096=>"101111111",
  17097=>"111111111",
  17098=>"111110100",
  17099=>"011111111",
  17100=>"000000111",
  17101=>"000111101",
  17102=>"111111010",
  17103=>"000000000",
  17104=>"110111110",
  17105=>"001000111",
  17106=>"100000000",
  17107=>"000000000",
  17108=>"111111111",
  17109=>"111111111",
  17110=>"000000000",
  17111=>"000001001",
  17112=>"000000000",
  17113=>"000000001",
  17114=>"001001011",
  17115=>"000001000",
  17116=>"110111111",
  17117=>"111100111",
  17118=>"111111110",
  17119=>"111110000",
  17120=>"000000000",
  17121=>"111111110",
  17122=>"000111111",
  17123=>"000000000",
  17124=>"110000000",
  17125=>"111111111",
  17126=>"000000110",
  17127=>"000000010",
  17128=>"001111111",
  17129=>"001111110",
  17130=>"000001111",
  17131=>"111100000",
  17132=>"000000000",
  17133=>"000010010",
  17134=>"111000000",
  17135=>"000000000",
  17136=>"111111011",
  17137=>"111000000",
  17138=>"111000011",
  17139=>"110111111",
  17140=>"111111111",
  17141=>"111110111",
  17142=>"100100000",
  17143=>"110101100",
  17144=>"000000010",
  17145=>"000000000",
  17146=>"000000110",
  17147=>"000000000",
  17148=>"101111001",
  17149=>"000000000",
  17150=>"101111111",
  17151=>"000000000",
  17152=>"100000000",
  17153=>"010011011",
  17154=>"111111000",
  17155=>"111100000",
  17156=>"111011111",
  17157=>"001000000",
  17158=>"000000000",
  17159=>"000000000",
  17160=>"100000100",
  17161=>"111000000",
  17162=>"000000000",
  17163=>"111111111",
  17164=>"001001001",
  17165=>"000000001",
  17166=>"000000000",
  17167=>"000010111",
  17168=>"001011000",
  17169=>"100001001",
  17170=>"000100000",
  17171=>"110111111",
  17172=>"000000000",
  17173=>"000111111",
  17174=>"110110110",
  17175=>"000000100",
  17176=>"000001111",
  17177=>"101101000",
  17178=>"000001000",
  17179=>"001000000",
  17180=>"000001000",
  17181=>"000000000",
  17182=>"000000000",
  17183=>"110000000",
  17184=>"000010000",
  17185=>"111111111",
  17186=>"000000000",
  17187=>"001000000",
  17188=>"111111110",
  17189=>"000000000",
  17190=>"011111000",
  17191=>"111011000",
  17192=>"000000111",
  17193=>"111111000",
  17194=>"111110111",
  17195=>"111111110",
  17196=>"000011110",
  17197=>"000000000",
  17198=>"000000010",
  17199=>"000000000",
  17200=>"110111001",
  17201=>"000000110",
  17202=>"111111111",
  17203=>"000000000",
  17204=>"111111111",
  17205=>"000000000",
  17206=>"000000010",
  17207=>"111100000",
  17208=>"000000110",
  17209=>"000000000",
  17210=>"111101111",
  17211=>"000010000",
  17212=>"000000000",
  17213=>"000000000",
  17214=>"111111111",
  17215=>"011111000",
  17216=>"000100000",
  17217=>"111111111",
  17218=>"111111111",
  17219=>"000111111",
  17220=>"000000000",
  17221=>"000000000",
  17222=>"001111111",
  17223=>"000000000",
  17224=>"111001000",
  17225=>"100111100",
  17226=>"101000010",
  17227=>"001100100",
  17228=>"100000010",
  17229=>"000000000",
  17230=>"110111110",
  17231=>"011000101",
  17232=>"000000001",
  17233=>"111111011",
  17234=>"111011011",
  17235=>"110110100",
  17236=>"000111111",
  17237=>"011001001",
  17238=>"111011011",
  17239=>"111101101",
  17240=>"000000000",
  17241=>"111111000",
  17242=>"000000000",
  17243=>"111011111",
  17244=>"000000000",
  17245=>"111111001",
  17246=>"000000000",
  17247=>"111111111",
  17248=>"100000000",
  17249=>"111111111",
  17250=>"101101101",
  17251=>"000000111",
  17252=>"000100110",
  17253=>"011111000",
  17254=>"111110000",
  17255=>"111001110",
  17256=>"000000001",
  17257=>"110111000",
  17258=>"111000100",
  17259=>"110100101",
  17260=>"000010000",
  17261=>"110000000",
  17262=>"011111110",
  17263=>"000000000",
  17264=>"000000111",
  17265=>"011000000",
  17266=>"000000001",
  17267=>"011001001",
  17268=>"000000000",
  17269=>"111000111",
  17270=>"110111111",
  17271=>"111111110",
  17272=>"001011011",
  17273=>"111111111",
  17274=>"111111000",
  17275=>"110111111",
  17276=>"011110111",
  17277=>"000000111",
  17278=>"000000000",
  17279=>"000000000",
  17280=>"000000000",
  17281=>"000001101",
  17282=>"111011011",
  17283=>"111111111",
  17284=>"000111111",
  17285=>"000000000",
  17286=>"011000000",
  17287=>"000000001",
  17288=>"000000001",
  17289=>"000100100",
  17290=>"101000000",
  17291=>"111111000",
  17292=>"000000000",
  17293=>"100100110",
  17294=>"000000000",
  17295=>"000101000",
  17296=>"000000000",
  17297=>"000000000",
  17298=>"000101000",
  17299=>"100000000",
  17300=>"111110111",
  17301=>"000000000",
  17302=>"111100110",
  17303=>"110100000",
  17304=>"001000000",
  17305=>"111111111",
  17306=>"000000011",
  17307=>"111001000",
  17308=>"100100110",
  17309=>"100110000",
  17310=>"001111111",
  17311=>"000000000",
  17312=>"000000100",
  17313=>"100000010",
  17314=>"100110111",
  17315=>"110110000",
  17316=>"000000110",
  17317=>"110111111",
  17318=>"111011000",
  17319=>"111111000",
  17320=>"000100111",
  17321=>"000000000",
  17322=>"000000000",
  17323=>"111000011",
  17324=>"000000000",
  17325=>"111111110",
  17326=>"111111111",
  17327=>"001011100",
  17328=>"111000001",
  17329=>"111111111",
  17330=>"111110000",
  17331=>"000000000",
  17332=>"100100111",
  17333=>"000000000",
  17334=>"000000000",
  17335=>"001001010",
  17336=>"111111000",
  17337=>"111111111",
  17338=>"000110010",
  17339=>"110110111",
  17340=>"000000000",
  17341=>"000000000",
  17342=>"010001001",
  17343=>"000011000",
  17344=>"111111011",
  17345=>"111111111",
  17346=>"000000000",
  17347=>"111111111",
  17348=>"001111111",
  17349=>"111001001",
  17350=>"000111111",
  17351=>"000000000",
  17352=>"100000111",
  17353=>"011001011",
  17354=>"000000000",
  17355=>"000100000",
  17356=>"000000000",
  17357=>"010010000",
  17358=>"000000000",
  17359=>"000011010",
  17360=>"011111111",
  17361=>"010100000",
  17362=>"100110111",
  17363=>"011011000",
  17364=>"001001011",
  17365=>"000000010",
  17366=>"000111110",
  17367=>"001000001",
  17368=>"001101000",
  17369=>"100100111",
  17370=>"111011110",
  17371=>"110100001",
  17372=>"111111111",
  17373=>"100110100",
  17374=>"000000000",
  17375=>"110010011",
  17376=>"111111111",
  17377=>"000000000",
  17378=>"110110110",
  17379=>"110111111",
  17380=>"111010010",
  17381=>"111111111",
  17382=>"111111110",
  17383=>"110111111",
  17384=>"110000000",
  17385=>"000000000",
  17386=>"000001011",
  17387=>"111111111",
  17388=>"001001111",
  17389=>"111111111",
  17390=>"001001001",
  17391=>"000000000",
  17392=>"011001001",
  17393=>"010000000",
  17394=>"111111111",
  17395=>"001111011",
  17396=>"000000010",
  17397=>"000000000",
  17398=>"111111111",
  17399=>"011001000",
  17400=>"111011001",
  17401=>"101101001",
  17402=>"111111000",
  17403=>"110000000",
  17404=>"000000000",
  17405=>"111001111",
  17406=>"000011000",
  17407=>"000000010",
  17408=>"111111001",
  17409=>"111000000",
  17410=>"111111101",
  17411=>"100000111",
  17412=>"000000010",
  17413=>"111000000",
  17414=>"011000000",
  17415=>"100000000",
  17416=>"011000000",
  17417=>"000001111",
  17418=>"111111011",
  17419=>"000000111",
  17420=>"100110111",
  17421=>"110110111",
  17422=>"111111111",
  17423=>"000000000",
  17424=>"001000000",
  17425=>"111001000",
  17426=>"100000010",
  17427=>"000001111",
  17428=>"000111111",
  17429=>"110000000",
  17430=>"000100000",
  17431=>"010110110",
  17432=>"000000111",
  17433=>"111111111",
  17434=>"100000000",
  17435=>"001000000",
  17436=>"111110000",
  17437=>"000110111",
  17438=>"001000000",
  17439=>"111111111",
  17440=>"001011000",
  17441=>"111000110",
  17442=>"000110111",
  17443=>"011000000",
  17444=>"011111111",
  17445=>"000100101",
  17446=>"010000001",
  17447=>"101110100",
  17448=>"000000001",
  17449=>"000000000",
  17450=>"111111011",
  17451=>"111111110",
  17452=>"111100000",
  17453=>"111111111",
  17454=>"111111111",
  17455=>"111100000",
  17456=>"111111111",
  17457=>"000000000",
  17458=>"100000000",
  17459=>"000000111",
  17460=>"111111100",
  17461=>"010000000",
  17462=>"111000001",
  17463=>"000000011",
  17464=>"000000000",
  17465=>"111001011",
  17466=>"000000111",
  17467=>"111001111",
  17468=>"011111000",
  17469=>"011000000",
  17470=>"111111011",
  17471=>"011000000",
  17472=>"000001111",
  17473=>"111111111",
  17474=>"000110111",
  17475=>"111111101",
  17476=>"000001000",
  17477=>"000000111",
  17478=>"100000110",
  17479=>"111111110",
  17480=>"101101001",
  17481=>"000000010",
  17482=>"111111111",
  17483=>"000000100",
  17484=>"000000000",
  17485=>"111111011",
  17486=>"101001000",
  17487=>"111111000",
  17488=>"000111111",
  17489=>"111111000",
  17490=>"111111111",
  17491=>"011011001",
  17492=>"111000000",
  17493=>"000000000",
  17494=>"111111000",
  17495=>"000100000",
  17496=>"000110111",
  17497=>"111001000",
  17498=>"111001000",
  17499=>"111000110",
  17500=>"000000011",
  17501=>"001111100",
  17502=>"000100000",
  17503=>"001001001",
  17504=>"111011010",
  17505=>"100000000",
  17506=>"000111111",
  17507=>"000000111",
  17508=>"000000000",
  17509=>"111111101",
  17510=>"111111000",
  17511=>"111000000",
  17512=>"111111111",
  17513=>"000000001",
  17514=>"111111100",
  17515=>"011011001",
  17516=>"111110100",
  17517=>"111111111",
  17518=>"101001000",
  17519=>"111111101",
  17520=>"000111111",
  17521=>"110111000",
  17522=>"001111100",
  17523=>"000000000",
  17524=>"000000001",
  17525=>"111110000",
  17526=>"000011000",
  17527=>"111000000",
  17528=>"000000111",
  17529=>"111000111",
  17530=>"011000000",
  17531=>"111001000",
  17532=>"110101101",
  17533=>"111111111",
  17534=>"000111000",
  17535=>"001000000",
  17536=>"000000000",
  17537=>"000000110",
  17538=>"111111000",
  17539=>"000110110",
  17540=>"110100000",
  17541=>"000000000",
  17542=>"111111111",
  17543=>"110111111",
  17544=>"111111110",
  17545=>"000000100",
  17546=>"000010111",
  17547=>"000000110",
  17548=>"011111100",
  17549=>"011111111",
  17550=>"100000111",
  17551=>"111111111",
  17552=>"100100000",
  17553=>"000000111",
  17554=>"111110000",
  17555=>"100110111",
  17556=>"000111000",
  17557=>"111111111",
  17558=>"000110110",
  17559=>"000000000",
  17560=>"110000000",
  17561=>"111111111",
  17562=>"111111111",
  17563=>"000110110",
  17564=>"000011011",
  17565=>"111111010",
  17566=>"000011111",
  17567=>"010110111",
  17568=>"000000000",
  17569=>"000000000",
  17570=>"000011111",
  17571=>"000000000",
  17572=>"000000000",
  17573=>"000100110",
  17574=>"001111111",
  17575=>"000000011",
  17576=>"111000000",
  17577=>"000001111",
  17578=>"111000000",
  17579=>"000000000",
  17580=>"111000000",
  17581=>"011111111",
  17582=>"111000000",
  17583=>"100000000",
  17584=>"000000000",
  17585=>"110110011",
  17586=>"010111111",
  17587=>"111101000",
  17588=>"000000000",
  17589=>"111111001",
  17590=>"000111111",
  17591=>"111110000",
  17592=>"111111111",
  17593=>"000000000",
  17594=>"111011000",
  17595=>"111111000",
  17596=>"000000000",
  17597=>"000010110",
  17598=>"000000000",
  17599=>"000000000",
  17600=>"011011100",
  17601=>"011000100",
  17602=>"001111111",
  17603=>"111111000",
  17604=>"000001110",
  17605=>"111111100",
  17606=>"100000011",
  17607=>"100100000",
  17608=>"100000000",
  17609=>"000000010",
  17610=>"011001000",
  17611=>"111011000",
  17612=>"000100111",
  17613=>"111010101",
  17614=>"001111111",
  17615=>"111000000",
  17616=>"111111111",
  17617=>"111000000",
  17618=>"000101111",
  17619=>"111110000",
  17620=>"011111001",
  17621=>"000111111",
  17622=>"000000000",
  17623=>"111011111",
  17624=>"000000111",
  17625=>"111111111",
  17626=>"000000000",
  17627=>"101111110",
  17628=>"001011111",
  17629=>"011111111",
  17630=>"000000000",
  17631=>"001111111",
  17632=>"001001011",
  17633=>"011001000",
  17634=>"110111110",
  17635=>"000111111",
  17636=>"011011011",
  17637=>"100100000",
  17638=>"111000000",
  17639=>"110111001",
  17640=>"101000000",
  17641=>"001101111",
  17642=>"111111111",
  17643=>"111000000",
  17644=>"000011111",
  17645=>"001100110",
  17646=>"000000111",
  17647=>"111111111",
  17648=>"000000000",
  17649=>"100111111",
  17650=>"000111111",
  17651=>"000110000",
  17652=>"111000000",
  17653=>"110110110",
  17654=>"110000000",
  17655=>"110000000",
  17656=>"111111111",
  17657=>"111111111",
  17658=>"000111000",
  17659=>"111110000",
  17660=>"011010110",
  17661=>"000010111",
  17662=>"110000000",
  17663=>"110110000",
  17664=>"001000000",
  17665=>"011001011",
  17666=>"111011000",
  17667=>"000000010",
  17668=>"111000000",
  17669=>"000000000",
  17670=>"000000000",
  17671=>"000111111",
  17672=>"000000110",
  17673=>"000000000",
  17674=>"101101000",
  17675=>"111111000",
  17676=>"011000111",
  17677=>"000000000",
  17678=>"100100100",
  17679=>"011111111",
  17680=>"000000111",
  17681=>"011111111",
  17682=>"000000100",
  17683=>"001000000",
  17684=>"111111111",
  17685=>"000000000",
  17686=>"100100010",
  17687=>"111110000",
  17688=>"111111111",
  17689=>"011111111",
  17690=>"000000111",
  17691=>"000000100",
  17692=>"111110000",
  17693=>"000011000",
  17694=>"000110111",
  17695=>"000111111",
  17696=>"011111111",
  17697=>"110000000",
  17698=>"000000000",
  17699=>"110100000",
  17700=>"110110111",
  17701=>"111111111",
  17702=>"000000000",
  17703=>"111111000",
  17704=>"111111111",
  17705=>"111011000",
  17706=>"000001111",
  17707=>"000111000",
  17708=>"111111111",
  17709=>"011011001",
  17710=>"111000111",
  17711=>"000000000",
  17712=>"001011111",
  17713=>"011101000",
  17714=>"000000000",
  17715=>"000110110",
  17716=>"111111100",
  17717=>"111111010",
  17718=>"001100000",
  17719=>"110110110",
  17720=>"011001111",
  17721=>"100111111",
  17722=>"111111000",
  17723=>"000000111",
  17724=>"011011011",
  17725=>"000000100",
  17726=>"010111111",
  17727=>"111011111",
  17728=>"000000000",
  17729=>"000000000",
  17730=>"000110111",
  17731=>"110000000",
  17732=>"110000111",
  17733=>"111111101",
  17734=>"001000000",
  17735=>"110111111",
  17736=>"111111000",
  17737=>"110111111",
  17738=>"001001001",
  17739=>"111111011",
  17740=>"011000100",
  17741=>"111100111",
  17742=>"000100111",
  17743=>"100110111",
  17744=>"101101101",
  17745=>"111001000",
  17746=>"110111111",
  17747=>"000000111",
  17748=>"000000010",
  17749=>"011011001",
  17750=>"111100100",
  17751=>"100100101",
  17752=>"000110001",
  17753=>"000000100",
  17754=>"011111111",
  17755=>"001011111",
  17756=>"000000000",
  17757=>"000111111",
  17758=>"000100001",
  17759=>"111111111",
  17760=>"011001000",
  17761=>"111111001",
  17762=>"100100000",
  17763=>"111000000",
  17764=>"110110111",
  17765=>"111111000",
  17766=>"110000000",
  17767=>"000000011",
  17768=>"110100111",
  17769=>"001110100",
  17770=>"111001000",
  17771=>"000000111",
  17772=>"111111000",
  17773=>"111011111",
  17774=>"000000000",
  17775=>"000000000",
  17776=>"111111111",
  17777=>"111111011",
  17778=>"111111111",
  17779=>"000011111",
  17780=>"000000001",
  17781=>"100100100",
  17782=>"000000000",
  17783=>"000000000",
  17784=>"000000100",
  17785=>"111110000",
  17786=>"000000001",
  17787=>"101101000",
  17788=>"001001000",
  17789=>"001011100",
  17790=>"000000000",
  17791=>"000000011",
  17792=>"000001100",
  17793=>"000100100",
  17794=>"001001111",
  17795=>"000000000",
  17796=>"011111111",
  17797=>"000111000",
  17798=>"111111111",
  17799=>"100100111",
  17800=>"000000001",
  17801=>"111111111",
  17802=>"100111111",
  17803=>"111111111",
  17804=>"001001111",
  17805=>"000001011",
  17806=>"111100000",
  17807=>"111000000",
  17808=>"111000000",
  17809=>"111111000",
  17810=>"111111000",
  17811=>"000111111",
  17812=>"000000100",
  17813=>"000000000",
  17814=>"000010010",
  17815=>"111001100",
  17816=>"100000000",
  17817=>"000111111",
  17818=>"111110000",
  17819=>"100000100",
  17820=>"000000000",
  17821=>"011111000",
  17822=>"000000000",
  17823=>"000000000",
  17824=>"001011111",
  17825=>"101100111",
  17826=>"000010010",
  17827=>"111111001",
  17828=>"111111000",
  17829=>"000001111",
  17830=>"100100110",
  17831=>"001000111",
  17832=>"110111001",
  17833=>"111111111",
  17834=>"000000000",
  17835=>"000000000",
  17836=>"101000000",
  17837=>"111101000",
  17838=>"100101000",
  17839=>"001011111",
  17840=>"000111111",
  17841=>"000000000",
  17842=>"000100111",
  17843=>"111100000",
  17844=>"111110111",
  17845=>"111111000",
  17846=>"111111110",
  17847=>"110111111",
  17848=>"000000000",
  17849=>"110000000",
  17850=>"001000000",
  17851=>"001101111",
  17852=>"000000111",
  17853=>"100111111",
  17854=>"111000011",
  17855=>"110000000",
  17856=>"010010111",
  17857=>"000000000",
  17858=>"111000000",
  17859=>"111111111",
  17860=>"010010110",
  17861=>"000001011",
  17862=>"001101000",
  17863=>"111000000",
  17864=>"010010111",
  17865=>"000000000",
  17866=>"000000000",
  17867=>"111111111",
  17868=>"111111000",
  17869=>"011110000",
  17870=>"111100001",
  17871=>"000000111",
  17872=>"110110111",
  17873=>"001000111",
  17874=>"000101100",
  17875=>"100011000",
  17876=>"101101001",
  17877=>"111110010",
  17878=>"101111000",
  17879=>"010011010",
  17880=>"000000000",
  17881=>"000001111",
  17882=>"111111111",
  17883=>"000000000",
  17884=>"110111011",
  17885=>"111111000",
  17886=>"100001111",
  17887=>"100000000",
  17888=>"100000000",
  17889=>"000100110",
  17890=>"001000000",
  17891=>"000110111",
  17892=>"111111111",
  17893=>"111111000",
  17894=>"001100111",
  17895=>"000001111",
  17896=>"000000000",
  17897=>"000111111",
  17898=>"000000000",
  17899=>"111111000",
  17900=>"000000110",
  17901=>"111111111",
  17902=>"000000000",
  17903=>"000000011",
  17904=>"001000000",
  17905=>"111111111",
  17906=>"100111111",
  17907=>"000100000",
  17908=>"111000000",
  17909=>"011111111",
  17910=>"000000000",
  17911=>"111101000",
  17912=>"000110110",
  17913=>"000100111",
  17914=>"000000000",
  17915=>"111101111",
  17916=>"011010000",
  17917=>"000100111",
  17918=>"100111111",
  17919=>"000000000",
  17920=>"000010011",
  17921=>"111001001",
  17922=>"111111111",
  17923=>"000000111",
  17924=>"000010001",
  17925=>"000000000",
  17926=>"000000000",
  17927=>"000000001",
  17928=>"111111111",
  17929=>"000111111",
  17930=>"111101000",
  17931=>"010101111",
  17932=>"000000100",
  17933=>"000000000",
  17934=>"000100111",
  17935=>"001001010",
  17936=>"111111101",
  17937=>"111111000",
  17938=>"000010000",
  17939=>"111100001",
  17940=>"000000000",
  17941=>"000000000",
  17942=>"000110011",
  17943=>"100110100",
  17944=>"000000000",
  17945=>"000011011",
  17946=>"000000111",
  17947=>"000110111",
  17948=>"111111111",
  17949=>"000000000",
  17950=>"010110000",
  17951=>"111111111",
  17952=>"100010011",
  17953=>"000000000",
  17954=>"100110110",
  17955=>"111001111",
  17956=>"000000000",
  17957=>"000000000",
  17958=>"111010111",
  17959=>"111111001",
  17960=>"000010111",
  17961=>"000000110",
  17962=>"111111000",
  17963=>"111111111",
  17964=>"111111111",
  17965=>"000000001",
  17966=>"111111111",
  17967=>"111111000",
  17968=>"111011000",
  17969=>"000001111",
  17970=>"110110100",
  17971=>"100100100",
  17972=>"001000000",
  17973=>"100000100",
  17974=>"111011111",
  17975=>"111111110",
  17976=>"111111110",
  17977=>"100111011",
  17978=>"111111111",
  17979=>"111111111",
  17980=>"111110111",
  17981=>"010000000",
  17982=>"111111111",
  17983=>"111110101",
  17984=>"000000100",
  17985=>"000100110",
  17986=>"111111110",
  17987=>"111110111",
  17988=>"111111100",
  17989=>"000000100",
  17990=>"000000000",
  17991=>"000001001",
  17992=>"111111110",
  17993=>"000000000",
  17994=>"111111111",
  17995=>"111000000",
  17996=>"100110000",
  17997=>"000000001",
  17998=>"100101000",
  17999=>"111111111",
  18000=>"000000011",
  18001=>"111111001",
  18002=>"000000000",
  18003=>"000001001",
  18004=>"001011000",
  18005=>"100110000",
  18006=>"111111111",
  18007=>"000010010",
  18008=>"001001000",
  18009=>"101000000",
  18010=>"111111111",
  18011=>"111111111",
  18012=>"000000000",
  18013=>"110000000",
  18014=>"000011011",
  18015=>"000000001",
  18016=>"000000000",
  18017=>"111111111",
  18018=>"011100111",
  18019=>"000000000",
  18020=>"011011111",
  18021=>"111111011",
  18022=>"011111111",
  18023=>"110110110",
  18024=>"000000000",
  18025=>"000000000",
  18026=>"110111011",
  18027=>"000000000",
  18028=>"011001000",
  18029=>"000000001",
  18030=>"000000000",
  18031=>"000000000",
  18032=>"111111010",
  18033=>"000000000",
  18034=>"000000001",
  18035=>"111111111",
  18036=>"000000000",
  18037=>"010110010",
  18038=>"111000100",
  18039=>"111111111",
  18040=>"001000000",
  18041=>"000000000",
  18042=>"000000000",
  18043=>"000000000",
  18044=>"111111110",
  18045=>"000000011",
  18046=>"011111111",
  18047=>"111111111",
  18048=>"111111000",
  18049=>"000000100",
  18050=>"111100000",
  18051=>"000000110",
  18052=>"111111111",
  18053=>"000000000",
  18054=>"111011111",
  18055=>"111111111",
  18056=>"000000000",
  18057=>"110010010",
  18058=>"000000000",
  18059=>"111111111",
  18060=>"111111111",
  18061=>"000000000",
  18062=>"100100100",
  18063=>"111111011",
  18064=>"111111000",
  18065=>"001111111",
  18066=>"000000000",
  18067=>"111111111",
  18068=>"111010000",
  18069=>"111111111",
  18070=>"000100001",
  18071=>"000000000",
  18072=>"000000001",
  18073=>"000100111",
  18074=>"110110111",
  18075=>"111111110",
  18076=>"111100100",
  18077=>"101001000",
  18078=>"001000000",
  18079=>"010010000",
  18080=>"000000111",
  18081=>"000111110",
  18082=>"111111001",
  18083=>"111111111",
  18084=>"011011100",
  18085=>"001000000",
  18086=>"111000000",
  18087=>"100100100",
  18088=>"111111111",
  18089=>"111111111",
  18090=>"000000101",
  18091=>"000000000",
  18092=>"111100111",
  18093=>"000110110",
  18094=>"101110101",
  18095=>"000001111",
  18096=>"011111000",
  18097=>"001001011",
  18098=>"010111011",
  18099=>"100100110",
  18100=>"000111111",
  18101=>"000000000",
  18102=>"111111111",
  18103=>"011100111",
  18104=>"000000000",
  18105=>"111111111",
  18106=>"000000000",
  18107=>"111011010",
  18108=>"000000000",
  18109=>"100000000",
  18110=>"000000000",
  18111=>"111101101",
  18112=>"000000000",
  18113=>"111000000",
  18114=>"111111111",
  18115=>"001000011",
  18116=>"111111111",
  18117=>"000000000",
  18118=>"011011000",
  18119=>"000000000",
  18120=>"000000000",
  18121=>"111110111",
  18122=>"111111111",
  18123=>"000000011",
  18124=>"111110100",
  18125=>"011111111",
  18126=>"100110111",
  18127=>"000000000",
  18128=>"101111111",
  18129=>"010000111",
  18130=>"011111111",
  18131=>"000000010",
  18132=>"000000000",
  18133=>"101000111",
  18134=>"000000000",
  18135=>"000000000",
  18136=>"000000011",
  18137=>"110110000",
  18138=>"000000000",
  18139=>"000000000",
  18140=>"111111111",
  18141=>"000000000",
  18142=>"111111111",
  18143=>"000000011",
  18144=>"011111111",
  18145=>"000100111",
  18146=>"000000000",
  18147=>"001011011",
  18148=>"111111111",
  18149=>"000000000",
  18150=>"111111111",
  18151=>"110110111",
  18152=>"100000000",
  18153=>"111111111",
  18154=>"001000000",
  18155=>"111111111",
  18156=>"000000000",
  18157=>"000100000",
  18158=>"011111111",
  18159=>"101111111",
  18160=>"111111111",
  18161=>"101111000",
  18162=>"111111100",
  18163=>"000000000",
  18164=>"111011111",
  18165=>"110100000",
  18166=>"100000000",
  18167=>"111111110",
  18168=>"000000000",
  18169=>"111111111",
  18170=>"000110111",
  18171=>"000000100",
  18172=>"111011011",
  18173=>"111111111",
  18174=>"100100110",
  18175=>"111111111",
  18176=>"111110010",
  18177=>"001000000",
  18178=>"000000111",
  18179=>"000000011",
  18180=>"000000000",
  18181=>"011000000",
  18182=>"000000001",
  18183=>"111111111",
  18184=>"111111111",
  18185=>"000110110",
  18186=>"011110000",
  18187=>"000000000",
  18188=>"000000000",
  18189=>"000000000",
  18190=>"111111111",
  18191=>"111111111",
  18192=>"001001001",
  18193=>"011011011",
  18194=>"000000000",
  18195=>"111011000",
  18196=>"000000111",
  18197=>"000000000",
  18198=>"000000101",
  18199=>"111001001",
  18200=>"111111100",
  18201=>"111011011",
  18202=>"100100000",
  18203=>"011000000",
  18204=>"111110000",
  18205=>"000010011",
  18206=>"000000000",
  18207=>"100110000",
  18208=>"111111111",
  18209=>"000000000",
  18210=>"000010000",
  18211=>"000000000",
  18212=>"111011001",
  18213=>"000000000",
  18214=>"100111100",
  18215=>"011011000",
  18216=>"000000000",
  18217=>"100000001",
  18218=>"101000110",
  18219=>"111111100",
  18220=>"100111110",
  18221=>"001011000",
  18222=>"111100000",
  18223=>"000111111",
  18224=>"000000001",
  18225=>"000000100",
  18226=>"111111111",
  18227=>"010010100",
  18228=>"100000000",
  18229=>"000000010",
  18230=>"000000001",
  18231=>"011000000",
  18232=>"000000000",
  18233=>"011000000",
  18234=>"000000000",
  18235=>"111000000",
  18236=>"000000000",
  18237=>"000111111",
  18238=>"000001000",
  18239=>"000000000",
  18240=>"111111111",
  18241=>"000000000",
  18242=>"001000011",
  18243=>"011011000",
  18244=>"011111111",
  18245=>"000000000",
  18246=>"000000000",
  18247=>"111111111",
  18248=>"110000000",
  18249=>"110110110",
  18250=>"101111111",
  18251=>"111111100",
  18252=>"000000111",
  18253=>"011100101",
  18254=>"111110110",
  18255=>"010000000",
  18256=>"011110000",
  18257=>"000000011",
  18258=>"000000000",
  18259=>"000000111",
  18260=>"000000000",
  18261=>"011011011",
  18262=>"111111111",
  18263=>"000111111",
  18264=>"111111111",
  18265=>"111111111",
  18266=>"110100011",
  18267=>"000000000",
  18268=>"111111111",
  18269=>"000000000",
  18270=>"000000010",
  18271=>"111111111",
  18272=>"100000000",
  18273=>"000011111",
  18274=>"001001001",
  18275=>"000001011",
  18276=>"110110100",
  18277=>"000010110",
  18278=>"000000001",
  18279=>"101000000",
  18280=>"001001101",
  18281=>"000000000",
  18282=>"000000000",
  18283=>"101111011",
  18284=>"000000000",
  18285=>"000001001",
  18286=>"000000000",
  18287=>"111111111",
  18288=>"111111111",
  18289=>"000000000",
  18290=>"111111111",
  18291=>"001001000",
  18292=>"100111111",
  18293=>"111111111",
  18294=>"100000100",
  18295=>"110011001",
  18296=>"111111111",
  18297=>"101111111",
  18298=>"000000000",
  18299=>"001000110",
  18300=>"111111111",
  18301=>"111111111",
  18302=>"000011011",
  18303=>"011010000",
  18304=>"110110110",
  18305=>"000000111",
  18306=>"000000000",
  18307=>"000000001",
  18308=>"010111111",
  18309=>"000000000",
  18310=>"110110111",
  18311=>"000000100",
  18312=>"100100110",
  18313=>"000000000",
  18314=>"101100100",
  18315=>"000000000",
  18316=>"000000000",
  18317=>"111111111",
  18318=>"011011011",
  18319=>"001111111",
  18320=>"000000000",
  18321=>"000000100",
  18322=>"011111010",
  18323=>"000000000",
  18324=>"000000000",
  18325=>"011000000",
  18326=>"001000000",
  18327=>"111111011",
  18328=>"111111011",
  18329=>"000111111",
  18330=>"000000000",
  18331=>"111111111",
  18332=>"000000111",
  18333=>"111111110",
  18334=>"000000010",
  18335=>"000000000",
  18336=>"000000000",
  18337=>"100001000",
  18338=>"111111111",
  18339=>"000000110",
  18340=>"001011111",
  18341=>"100000000",
  18342=>"101101101",
  18343=>"000000000",
  18344=>"000101111",
  18345=>"000000000",
  18346=>"111111111",
  18347=>"000000000",
  18348=>"000000000",
  18349=>"111110111",
  18350=>"110100000",
  18351=>"111111111",
  18352=>"110110111",
  18353=>"111111011",
  18354=>"000010001",
  18355=>"000000000",
  18356=>"101001001",
  18357=>"000000111",
  18358=>"000000000",
  18359=>"111101001",
  18360=>"000000111",
  18361=>"111010000",
  18362=>"000000000",
  18363=>"111111111",
  18364=>"111110000",
  18365=>"100000100",
  18366=>"000000000",
  18367=>"001101111",
  18368=>"000000000",
  18369=>"000110000",
  18370=>"111111111",
  18371=>"000111111",
  18372=>"000101111",
  18373=>"111110110",
  18374=>"000000000",
  18375=>"001000000",
  18376=>"000000000",
  18377=>"000000000",
  18378=>"000000001",
  18379=>"111111111",
  18380=>"010111010",
  18381=>"110111111",
  18382=>"000000000",
  18383=>"000000000",
  18384=>"000000000",
  18385=>"111111111",
  18386=>"111111010",
  18387=>"111111111",
  18388=>"111101111",
  18389=>"000000000",
  18390=>"111110111",
  18391=>"000000000",
  18392=>"000000000",
  18393=>"110000000",
  18394=>"000010000",
  18395=>"111111111",
  18396=>"000001111",
  18397=>"000000000",
  18398=>"111111111",
  18399=>"010000001",
  18400=>"100000000",
  18401=>"000000000",
  18402=>"111111111",
  18403=>"000000100",
  18404=>"111111110",
  18405=>"100100111",
  18406=>"001111111",
  18407=>"001000000",
  18408=>"000000000",
  18409=>"111000000",
  18410=>"100110110",
  18411=>"000000000",
  18412=>"100000000",
  18413=>"000011001",
  18414=>"011000000",
  18415=>"010011010",
  18416=>"111111010",
  18417=>"110111111",
  18418=>"000000000",
  18419=>"000000000",
  18420=>"100000110",
  18421=>"000000000",
  18422=>"111100000",
  18423=>"000000000",
  18424=>"111111111",
  18425=>"110110001",
  18426=>"111111100",
  18427=>"111000000",
  18428=>"011000000",
  18429=>"110110000",
  18430=>"000000000",
  18431=>"000100100",
  18432=>"110111111",
  18433=>"000000110",
  18434=>"111111111",
  18435=>"111111011",
  18436=>"000001111",
  18437=>"000010000",
  18438=>"111101101",
  18439=>"111111111",
  18440=>"101100010",
  18441=>"101100111",
  18442=>"000001101",
  18443=>"000000011",
  18444=>"100110111",
  18445=>"001001000",
  18446=>"111110111",
  18447=>"000000000",
  18448=>"111010000",
  18449=>"000000111",
  18450=>"110111111",
  18451=>"010010000",
  18452=>"001001000",
  18453=>"000000000",
  18454=>"001011111",
  18455=>"111111100",
  18456=>"110110110",
  18457=>"000110110",
  18458=>"110111110",
  18459=>"000011000",
  18460=>"000100100",
  18461=>"000000000",
  18462=>"000000011",
  18463=>"111100100",
  18464=>"111001001",
  18465=>"111111111",
  18466=>"000101001",
  18467=>"000000000",
  18468=>"111111111",
  18469=>"011000011",
  18470=>"000000000",
  18471=>"111000100",
  18472=>"000000010",
  18473=>"110111110",
  18474=>"000010010",
  18475=>"011011001",
  18476=>"000000011",
  18477=>"111111110",
  18478=>"000101101",
  18479=>"010000000",
  18480=>"010000000",
  18481=>"111100100",
  18482=>"100100000",
  18483=>"111100010",
  18484=>"110000000",
  18485=>"110100000",
  18486=>"000000000",
  18487=>"010000000",
  18488=>"000000000",
  18489=>"000000000",
  18490=>"100000000",
  18491=>"000000000",
  18492=>"000000000",
  18493=>"001001001",
  18494=>"111111111",
  18495=>"100110100",
  18496=>"001000101",
  18497=>"100000001",
  18498=>"111110111",
  18499=>"110110111",
  18500=>"000001001",
  18501=>"001001111",
  18502=>"111000000",
  18503=>"000000000",
  18504=>"011010000",
  18505=>"000000001",
  18506=>"111111111",
  18507=>"101111111",
  18508=>"100000000",
  18509=>"110100000",
  18510=>"111010000",
  18511=>"111100110",
  18512=>"000101111",
  18513=>"000010010",
  18514=>"000000000",
  18515=>"111111011",
  18516=>"110100000",
  18517=>"111111111",
  18518=>"111111111",
  18519=>"000100000",
  18520=>"000000110",
  18521=>"111000000",
  18522=>"101101001",
  18523=>"111011111",
  18524=>"000111000",
  18525=>"111010000",
  18526=>"000000000",
  18527=>"000100100",
  18528=>"000000000",
  18529=>"000000000",
  18530=>"111100101",
  18531=>"000000000",
  18532=>"000001001",
  18533=>"000000000",
  18534=>"000000001",
  18535=>"111111111",
  18536=>"111111011",
  18537=>"011011011",
  18538=>"101001111",
  18539=>"111111111",
  18540=>"110000001",
  18541=>"111111111",
  18542=>"000010000",
  18543=>"100000000",
  18544=>"111111111",
  18545=>"110000011",
  18546=>"011000100",
  18547=>"000000001",
  18548=>"110100011",
  18549=>"111111111",
  18550=>"100100101",
  18551=>"110100000",
  18552=>"000000000",
  18553=>"111111111",
  18554=>"111111111",
  18555=>"000000000",
  18556=>"110000111",
  18557=>"111100100",
  18558=>"111111001",
  18559=>"000111011",
  18560=>"000000000",
  18561=>"001000000",
  18562=>"111101101",
  18563=>"111011010",
  18564=>"000000000",
  18565=>"111111111",
  18566=>"000000000",
  18567=>"111111111",
  18568=>"101111111",
  18569=>"101101101",
  18570=>"000000101",
  18571=>"110110111",
  18572=>"000100000",
  18573=>"111111110",
  18574=>"111110010",
  18575=>"000000101",
  18576=>"111011000",
  18577=>"100000000",
  18578=>"000000000",
  18579=>"000000000",
  18580=>"100111111",
  18581=>"111010000",
  18582=>"111001000",
  18583=>"000000000",
  18584=>"111011011",
  18585=>"101000000",
  18586=>"000000011",
  18587=>"111111000",
  18588=>"100000000",
  18589=>"111111000",
  18590=>"011111011",
  18591=>"110011011",
  18592=>"111111111",
  18593=>"000000000",
  18594=>"000111111",
  18595=>"010010111",
  18596=>"000100101",
  18597=>"000000000",
  18598=>"100000100",
  18599=>"000000000",
  18600=>"011011000",
  18601=>"000001011",
  18602=>"111101111",
  18603=>"111110111",
  18604=>"001001010",
  18605=>"001001001",
  18606=>"000000010",
  18607=>"010000110",
  18608=>"011111111",
  18609=>"011011110",
  18610=>"111111100",
  18611=>"111111000",
  18612=>"111111111",
  18613=>"011011111",
  18614=>"110100000",
  18615=>"101000100",
  18616=>"000000000",
  18617=>"000000000",
  18618=>"011000000",
  18619=>"110100000",
  18620=>"000010110",
  18621=>"111111001",
  18622=>"000100000",
  18623=>"000101111",
  18624=>"000000000",
  18625=>"000101010",
  18626=>"111111001",
  18627=>"111111111",
  18628=>"000000101",
  18629=>"000000001",
  18630=>"110110111",
  18631=>"111011011",
  18632=>"011011010",
  18633=>"100111111",
  18634=>"110010000",
  18635=>"111111101",
  18636=>"000000000",
  18637=>"011011011",
  18638=>"101001001",
  18639=>"011001001",
  18640=>"000000101",
  18641=>"000011111",
  18642=>"111111111",
  18643=>"100000011",
  18644=>"110111111",
  18645=>"110000000",
  18646=>"000000000",
  18647=>"000000000",
  18648=>"000010000",
  18649=>"111111010",
  18650=>"000000100",
  18651=>"111111110",
  18652=>"001001001",
  18653=>"010111111",
  18654=>"111111111",
  18655=>"001001011",
  18656=>"110000000",
  18657=>"010011011",
  18658=>"111110000",
  18659=>"111101001",
  18660=>"111111111",
  18661=>"011011010",
  18662=>"011111111",
  18663=>"111000000",
  18664=>"100111111",
  18665=>"110111110",
  18666=>"111011001",
  18667=>"100100000",
  18668=>"100000111",
  18669=>"111111111",
  18670=>"111111111",
  18671=>"111011001",
  18672=>"111000000",
  18673=>"000000000",
  18674=>"111100100",
  18675=>"001111000",
  18676=>"111111111",
  18677=>"110000011",
  18678=>"100111111",
  18679=>"110110000",
  18680=>"010000001",
  18681=>"010110110",
  18682=>"110100000",
  18683=>"110000110",
  18684=>"101100100",
  18685=>"110111111",
  18686=>"111111111",
  18687=>"100110111",
  18688=>"010001001",
  18689=>"010010010",
  18690=>"111000000",
  18691=>"011001000",
  18692=>"100111111",
  18693=>"010000000",
  18694=>"010000000",
  18695=>"101001001",
  18696=>"101101111",
  18697=>"000000000",
  18698=>"111111110",
  18699=>"011001010",
  18700=>"000000000",
  18701=>"100000000",
  18702=>"011001000",
  18703=>"000000000",
  18704=>"000000000",
  18705=>"111001001",
  18706=>"111110110",
  18707=>"111111111",
  18708=>"011111101",
  18709=>"111010000",
  18710=>"000100100",
  18711=>"010000000",
  18712=>"000000000",
  18713=>"111111111",
  18714=>"111100000",
  18715=>"000001001",
  18716=>"111001011",
  18717=>"111111111",
  18718=>"111000000",
  18719=>"111111111",
  18720=>"100100000",
  18721=>"010111111",
  18722=>"111111111",
  18723=>"100000111",
  18724=>"100000001",
  18725=>"010000000",
  18726=>"111011011",
  18727=>"101111111",
  18728=>"111111111",
  18729=>"000000000",
  18730=>"010111111",
  18731=>"110111001",
  18732=>"101111100",
  18733=>"100000000",
  18734=>"111110111",
  18735=>"000000000",
  18736=>"000000000",
  18737=>"100100000",
  18738=>"111011000",
  18739=>"111101001",
  18740=>"001000100",
  18741=>"110100000",
  18742=>"000110000",
  18743=>"010000010",
  18744=>"000000111",
  18745=>"111000001",
  18746=>"111101000",
  18747=>"000000000",
  18748=>"001001000",
  18749=>"000101101",
  18750=>"110110101",
  18751=>"111111111",
  18752=>"000000011",
  18753=>"000000000",
  18754=>"000000000",
  18755=>"111111110",
  18756=>"000000000",
  18757=>"111111111",
  18758=>"111111111",
  18759=>"110111111",
  18760=>"110110110",
  18761=>"000000000",
  18762=>"001001011",
  18763=>"010000000",
  18764=>"111001000",
  18765=>"111111111",
  18766=>"111101101",
  18767=>"110110110",
  18768=>"110110000",
  18769=>"111111111",
  18770=>"000000000",
  18771=>"011011000",
  18772=>"111111111",
  18773=>"111111111",
  18774=>"101001001",
  18775=>"100100111",
  18776=>"111111111",
  18777=>"111100111",
  18778=>"111100111",
  18779=>"010000010",
  18780=>"111011111",
  18781=>"111111111",
  18782=>"000000000",
  18783=>"000000111",
  18784=>"000000001",
  18785=>"111000000",
  18786=>"011010100",
  18787=>"000000000",
  18788=>"100001001",
  18789=>"111111111",
  18790=>"110110111",
  18791=>"011001000",
  18792=>"000000000",
  18793=>"111111111",
  18794=>"000000000",
  18795=>"111111111",
  18796=>"111111111",
  18797=>"011111011",
  18798=>"111110000",
  18799=>"111111111",
  18800=>"111011011",
  18801=>"001001111",
  18802=>"111111011",
  18803=>"100100110",
  18804=>"111111111",
  18805=>"111111111",
  18806=>"110111000",
  18807=>"000100100",
  18808=>"000000001",
  18809=>"000000000",
  18810=>"000000000",
  18811=>"000000000",
  18812=>"111111001",
  18813=>"111111000",
  18814=>"100111111",
  18815=>"111110000",
  18816=>"010000001",
  18817=>"101101000",
  18818=>"000000100",
  18819=>"111111011",
  18820=>"111100110",
  18821=>"000000000",
  18822=>"000000110",
  18823=>"101111111",
  18824=>"000000000",
  18825=>"111100100",
  18826=>"000110100",
  18827=>"000000000",
  18828=>"001001111",
  18829=>"011010110",
  18830=>"000010010",
  18831=>"000001010",
  18832=>"011111011",
  18833=>"001001001",
  18834=>"100110110",
  18835=>"000101000",
  18836=>"101001000",
  18837=>"101000101",
  18838=>"000101111",
  18839=>"111111111",
  18840=>"000000000",
  18841=>"000000000",
  18842=>"111111001",
  18843=>"000000111",
  18844=>"000000000",
  18845=>"000000011",
  18846=>"010000000",
  18847=>"000000000",
  18848=>"111111111",
  18849=>"011010010",
  18850=>"010010110",
  18851=>"111001111",
  18852=>"010011111",
  18853=>"000100100",
  18854=>"001000000",
  18855=>"000101100",
  18856=>"111010000",
  18857=>"011001100",
  18858=>"000010110",
  18859=>"111011001",
  18860=>"111111100",
  18861=>"111111111",
  18862=>"110110010",
  18863=>"000101000",
  18864=>"011011111",
  18865=>"110111010",
  18866=>"111010010",
  18867=>"111101100",
  18868=>"011111111",
  18869=>"111111111",
  18870=>"000000000",
  18871=>"000110010",
  18872=>"000011011",
  18873=>"001001111",
  18874=>"111111101",
  18875=>"000010111",
  18876=>"000000100",
  18877=>"000011101",
  18878=>"000000000",
  18879=>"011011010",
  18880=>"111110111",
  18881=>"111111111",
  18882=>"111111111",
  18883=>"111111111",
  18884=>"000010111",
  18885=>"000000100",
  18886=>"111011000",
  18887=>"000000000",
  18888=>"010011010",
  18889=>"111111011",
  18890=>"000000000",
  18891=>"000000000",
  18892=>"000000000",
  18893=>"011000000",
  18894=>"000000000",
  18895=>"000000000",
  18896=>"111111111",
  18897=>"000000000",
  18898=>"111111010",
  18899=>"000000000",
  18900=>"111110100",
  18901=>"000001011",
  18902=>"001010010",
  18903=>"010000000",
  18904=>"111000000",
  18905=>"111100000",
  18906=>"000110111",
  18907=>"111111111",
  18908=>"100001000",
  18909=>"001000000",
  18910=>"000000000",
  18911=>"000000110",
  18912=>"000000000",
  18913=>"000000001",
  18914=>"010010000",
  18915=>"111100111",
  18916=>"111101000",
  18917=>"111111111",
  18918=>"000000001",
  18919=>"111111111",
  18920=>"000000010",
  18921=>"101001001",
  18922=>"000000000",
  18923=>"101101000",
  18924=>"111111111",
  18925=>"111011001",
  18926=>"000000000",
  18927=>"010000000",
  18928=>"110000100",
  18929=>"111110110",
  18930=>"000011000",
  18931=>"111111010",
  18932=>"011001001",
  18933=>"000100111",
  18934=>"000000000",
  18935=>"100101111",
  18936=>"000000000",
  18937=>"010010000",
  18938=>"001001011",
  18939=>"111111111",
  18940=>"110011000",
  18941=>"110111111",
  18942=>"111100111",
  18943=>"111111101",
  18944=>"001011100",
  18945=>"000000000",
  18946=>"001001111",
  18947=>"111011100",
  18948=>"110110110",
  18949=>"001001111",
  18950=>"000000000",
  18951=>"111011111",
  18952=>"111001000",
  18953=>"000000111",
  18954=>"111100111",
  18955=>"101111111",
  18956=>"000000100",
  18957=>"111000000",
  18958=>"000000111",
  18959=>"001000000",
  18960=>"101011000",
  18961=>"111111111",
  18962=>"111000000",
  18963=>"000011011",
  18964=>"000100100",
  18965=>"011001001",
  18966=>"000101001",
  18967=>"001100100",
  18968=>"000000110",
  18969=>"001001000",
  18970=>"101000111",
  18971=>"110011001",
  18972=>"111111111",
  18973=>"000000000",
  18974=>"000001111",
  18975=>"000110111",
  18976=>"000111100",
  18977=>"111111000",
  18978=>"111111111",
  18979=>"000000000",
  18980=>"000000111",
  18981=>"001000000",
  18982=>"000000000",
  18983=>"000001000",
  18984=>"000010000",
  18985=>"101000000",
  18986=>"111111101",
  18987=>"111111111",
  18988=>"101111000",
  18989=>"000100111",
  18990=>"100000001",
  18991=>"010000001",
  18992=>"010011111",
  18993=>"101111000",
  18994=>"000111111",
  18995=>"000111001",
  18996=>"000000111",
  18997=>"111110110",
  18998=>"110110010",
  18999=>"111111111",
  19000=>"011001001",
  19001=>"001000111",
  19002=>"000001000",
  19003=>"100001001",
  19004=>"001001111",
  19005=>"111111000",
  19006=>"111110000",
  19007=>"101111111",
  19008=>"101000111",
  19009=>"111000101",
  19010=>"000011110",
  19011=>"111111111",
  19012=>"111111000",
  19013=>"001111101",
  19014=>"111100110",
  19015=>"111001100",
  19016=>"000011011",
  19017=>"000000000",
  19018=>"111000001",
  19019=>"101000011",
  19020=>"000000000",
  19021=>"111111010",
  19022=>"111101100",
  19023=>"111111111",
  19024=>"000000000",
  19025=>"001000000",
  19026=>"111011011",
  19027=>"110110111",
  19028=>"101000000",
  19029=>"000111111",
  19030=>"111111110",
  19031=>"000111111",
  19032=>"100000000",
  19033=>"111000000",
  19034=>"111101101",
  19035=>"100101001",
  19036=>"100000000",
  19037=>"000011111",
  19038=>"111111111",
  19039=>"001000010",
  19040=>"000000100",
  19041=>"001000000",
  19042=>"000000000",
  19043=>"111010000",
  19044=>"111111000",
  19045=>"111001111",
  19046=>"011001101",
  19047=>"111111111",
  19048=>"000111111",
  19049=>"111001111",
  19050=>"111111111",
  19051=>"111001000",
  19052=>"101111111",
  19053=>"000000011",
  19054=>"111111111",
  19055=>"000011000",
  19056=>"000011010",
  19057=>"000000001",
  19058=>"000000111",
  19059=>"111111100",
  19060=>"000111111",
  19061=>"000000100",
  19062=>"000011111",
  19063=>"101111000",
  19064=>"000000111",
  19065=>"000000110",
  19066=>"111000000",
  19067=>"000001000",
  19068=>"000010010",
  19069=>"011111111",
  19070=>"010000000",
  19071=>"000000000",
  19072=>"000111001",
  19073=>"000010011",
  19074=>"001000000",
  19075=>"000000000",
  19076=>"111111111",
  19077=>"001001111",
  19078=>"110010000",
  19079=>"000001111",
  19080=>"001111011",
  19081=>"111111000",
  19082=>"000010010",
  19083=>"111000000",
  19084=>"101111111",
  19085=>"000111111",
  19086=>"000000000",
  19087=>"000111111",
  19088=>"011111111",
  19089=>"111111000",
  19090=>"111111000",
  19091=>"111111000",
  19092=>"000110111",
  19093=>"101000101",
  19094=>"000000000",
  19095=>"111000000",
  19096=>"000000110",
  19097=>"000000011",
  19098=>"110010010",
  19099=>"000000000",
  19100=>"100111111",
  19101=>"111111000",
  19102=>"000000000",
  19103=>"111100000",
  19104=>"111111000",
  19105=>"111111000",
  19106=>"101000101",
  19107=>"000000111",
  19108=>"111000000",
  19109=>"100100100",
  19110=>"111111111",
  19111=>"000100001",
  19112=>"000000011",
  19113=>"000000100",
  19114=>"000111000",
  19115=>"000010111",
  19116=>"111001000",
  19117=>"110110000",
  19118=>"000000000",
  19119=>"100000011",
  19120=>"101001000",
  19121=>"100100000",
  19122=>"111111001",
  19123=>"110111111",
  19124=>"111111000",
  19125=>"000000000",
  19126=>"000111111",
  19127=>"111111000",
  19128=>"110111111",
  19129=>"111111000",
  19130=>"000000001",
  19131=>"111111000",
  19132=>"011111111",
  19133=>"011111001",
  19134=>"101111111",
  19135=>"111000000",
  19136=>"011111011",
  19137=>"110000111",
  19138=>"111001000",
  19139=>"000000000",
  19140=>"001111111",
  19141=>"000000111",
  19142=>"111111000",
  19143=>"110111111",
  19144=>"000111111",
  19145=>"000111111",
  19146=>"000010111",
  19147=>"111111111",
  19148=>"101001001",
  19149=>"000000111",
  19150=>"111111000",
  19151=>"111101000",
  19152=>"111011000",
  19153=>"000000000",
  19154=>"101001000",
  19155=>"000000000",
  19156=>"000111111",
  19157=>"111111111",
  19158=>"001000000",
  19159=>"111111000",
  19160=>"000000111",
  19161=>"000100010",
  19162=>"111100111",
  19163=>"000000111",
  19164=>"001011111",
  19165=>"000000111",
  19166=>"101111000",
  19167=>"000000000",
  19168=>"011000000",
  19169=>"111011000",
  19170=>"100000100",
  19171=>"000100100",
  19172=>"100010111",
  19173=>"011111000",
  19174=>"111100111",
  19175=>"000000000",
  19176=>"000000000",
  19177=>"111111111",
  19178=>"010000001",
  19179=>"111000000",
  19180=>"000000001",
  19181=>"111110100",
  19182=>"111001001",
  19183=>"000110111",
  19184=>"100111111",
  19185=>"111100111",
  19186=>"000111111",
  19187=>"001001000",
  19188=>"111111011",
  19189=>"100100111",
  19190=>"101100110",
  19191=>"000000000",
  19192=>"000000010",
  19193=>"000000011",
  19194=>"000000111",
  19195=>"000000000",
  19196=>"000110011",
  19197=>"000001111",
  19198=>"101000000",
  19199=>"000000111",
  19200=>"000000111",
  19201=>"000000111",
  19202=>"000011011",
  19203=>"111111010",
  19204=>"110110111",
  19205=>"000000000",
  19206=>"111000000",
  19207=>"100111111",
  19208=>"111010000",
  19209=>"111111000",
  19210=>"000001000",
  19211=>"001000011",
  19212=>"001000011",
  19213=>"000000000",
  19214=>"111100000",
  19215=>"000000100",
  19216=>"000100111",
  19217=>"111101100",
  19218=>"000001001",
  19219=>"000111111",
  19220=>"110000010",
  19221=>"111010111",
  19222=>"000100110",
  19223=>"010010011",
  19224=>"111001001",
  19225=>"000110001",
  19226=>"000001111",
  19227=>"110111000",
  19228=>"000001101",
  19229=>"000111111",
  19230=>"000011000",
  19231=>"010111100",
  19232=>"000100111",
  19233=>"111000000",
  19234=>"000001111",
  19235=>"110111011",
  19236=>"111111001",
  19237=>"111111001",
  19238=>"101111111",
  19239=>"101101111",
  19240=>"111111111",
  19241=>"000001000",
  19242=>"010111111",
  19243=>"000000000",
  19244=>"111111011",
  19245=>"100000001",
  19246=>"101100000",
  19247=>"000000000",
  19248=>"111111111",
  19249=>"000000000",
  19250=>"111111111",
  19251=>"000000000",
  19252=>"111111111",
  19253=>"001001000",
  19254=>"000000000",
  19255=>"111001000",
  19256=>"111111000",
  19257=>"111000001",
  19258=>"111111111",
  19259=>"111111010",
  19260=>"000000000",
  19261=>"000010001",
  19262=>"000111111",
  19263=>"111000010",
  19264=>"111100000",
  19265=>"001001111",
  19266=>"000000110",
  19267=>"111111111",
  19268=>"111000000",
  19269=>"111111000",
  19270=>"000110100",
  19271=>"011000000",
  19272=>"001000000",
  19273=>"000000000",
  19274=>"011111111",
  19275=>"000000000",
  19276=>"111000000",
  19277=>"111011000",
  19278=>"111000000",
  19279=>"000000000",
  19280=>"011001000",
  19281=>"111111000",
  19282=>"100000000",
  19283=>"111100001",
  19284=>"000000111",
  19285=>"111011000",
  19286=>"000000000",
  19287=>"111111000",
  19288=>"000000000",
  19289=>"000000011",
  19290=>"000111111",
  19291=>"010111011",
  19292=>"111000001",
  19293=>"000000101",
  19294=>"000000000",
  19295=>"111111010",
  19296=>"100111101",
  19297=>"011111111",
  19298=>"000100101",
  19299=>"000011000",
  19300=>"000000111",
  19301=>"000000000",
  19302=>"111000000",
  19303=>"010010010",
  19304=>"001001011",
  19305=>"000110110",
  19306=>"111111000",
  19307=>"111000111",
  19308=>"000110110",
  19309=>"111111010",
  19310=>"111110000",
  19311=>"000000111",
  19312=>"111111011",
  19313=>"000000000",
  19314=>"111100000",
  19315=>"111111111",
  19316=>"111110000",
  19317=>"000000000",
  19318=>"000000110",
  19319=>"000000011",
  19320=>"000000000",
  19321=>"000000000",
  19322=>"111111000",
  19323=>"111111111",
  19324=>"110000110",
  19325=>"000010111",
  19326=>"000110001",
  19327=>"111111111",
  19328=>"001001001",
  19329=>"001000011",
  19330=>"110111001",
  19331=>"000111000",
  19332=>"000001111",
  19333=>"000000000",
  19334=>"001100111",
  19335=>"010111110",
  19336=>"110110000",
  19337=>"000000000",
  19338=>"000001000",
  19339=>"111110111",
  19340=>"111000111",
  19341=>"100100110",
  19342=>"010011010",
  19343=>"001111000",
  19344=>"000000000",
  19345=>"000001111",
  19346=>"000011011",
  19347=>"000000011",
  19348=>"000000111",
  19349=>"000001000",
  19350=>"000000111",
  19351=>"111110000",
  19352=>"111011000",
  19353=>"111111110",
  19354=>"111000000",
  19355=>"111111111",
  19356=>"000000111",
  19357=>"000000000",
  19358=>"000000111",
  19359=>"111111100",
  19360=>"000000000",
  19361=>"001110100",
  19362=>"000111111",
  19363=>"000000111",
  19364=>"000000110",
  19365=>"000110110",
  19366=>"111100111",
  19367=>"011011001",
  19368=>"000000001",
  19369=>"111110110",
  19370=>"111001001",
  19371=>"000000111",
  19372=>"000000000",
  19373=>"101111110",
  19374=>"000000111",
  19375=>"111111111",
  19376=>"000000111",
  19377=>"111000000",
  19378=>"000000000",
  19379=>"000101111",
  19380=>"000000000",
  19381=>"111110111",
  19382=>"000000111",
  19383=>"111001000",
  19384=>"101111000",
  19385=>"101001100",
  19386=>"110110100",
  19387=>"000001111",
  19388=>"111101100",
  19389=>"000000100",
  19390=>"000100111",
  19391=>"110111101",
  19392=>"111111101",
  19393=>"000111111",
  19394=>"000011000",
  19395=>"000000111",
  19396=>"000001111",
  19397=>"001001111",
  19398=>"111011000",
  19399=>"000011111",
  19400=>"111000000",
  19401=>"011101111",
  19402=>"000110011",
  19403=>"000000000",
  19404=>"111110000",
  19405=>"111110000",
  19406=>"011011000",
  19407=>"000111111",
  19408=>"011011000",
  19409=>"001000001",
  19410=>"001000111",
  19411=>"111000000",
  19412=>"010010110",
  19413=>"000111111",
  19414=>"000000001",
  19415=>"011000000",
  19416=>"001100100",
  19417=>"000110000",
  19418=>"010100111",
  19419=>"000000010",
  19420=>"111111111",
  19421=>"000111111",
  19422=>"000001011",
  19423=>"111100100",
  19424=>"000000010",
  19425=>"000000000",
  19426=>"110110000",
  19427=>"000100000",
  19428=>"011111100",
  19429=>"100001111",
  19430=>"011000000",
  19431=>"111000110",
  19432=>"000011111",
  19433=>"101111111",
  19434=>"011000000",
  19435=>"101011111",
  19436=>"111111110",
  19437=>"111111000",
  19438=>"000010010",
  19439=>"111111000",
  19440=>"100111111",
  19441=>"111000000",
  19442=>"111000000",
  19443=>"000000010",
  19444=>"000000111",
  19445=>"000111111",
  19446=>"110100101",
  19447=>"111000000",
  19448=>"011011011",
  19449=>"000000111",
  19450=>"000000000",
  19451=>"111111000",
  19452=>"000000000",
  19453=>"111011011",
  19454=>"000001000",
  19455=>"001000001",
  19456=>"001001011",
  19457=>"000110110",
  19458=>"001101111",
  19459=>"111110010",
  19460=>"111101111",
  19461=>"111001000",
  19462=>"110111010",
  19463=>"111100111",
  19464=>"111000000",
  19465=>"000000000",
  19466=>"111111111",
  19467=>"100100101",
  19468=>"100100100",
  19469=>"110110111",
  19470=>"110111001",
  19471=>"010111111",
  19472=>"000000001",
  19473=>"000001000",
  19474=>"101000101",
  19475=>"000011011",
  19476=>"110100000",
  19477=>"000000111",
  19478=>"111000000",
  19479=>"000000000",
  19480=>"110110000",
  19481=>"000001000",
  19482=>"000000000",
  19483=>"110000000",
  19484=>"001001111",
  19485=>"111111111",
  19486=>"000010110",
  19487=>"111111001",
  19488=>"100000000",
  19489=>"000000000",
  19490=>"101001001",
  19491=>"110110110",
  19492=>"011011010",
  19493=>"110110010",
  19494=>"111101001",
  19495=>"111011000",
  19496=>"111111100",
  19497=>"111111111",
  19498=>"000000111",
  19499=>"001001001",
  19500=>"000010000",
  19501=>"010111010",
  19502=>"001000000",
  19503=>"111011011",
  19504=>"011111111",
  19505=>"010111110",
  19506=>"100110111",
  19507=>"111111111",
  19508=>"111000000",
  19509=>"111100110",
  19510=>"101000000",
  19511=>"000000111",
  19512=>"001111111",
  19513=>"000000111",
  19514=>"100111111",
  19515=>"001111111",
  19516=>"111101111",
  19517=>"111100111",
  19518=>"110100000",
  19519=>"100100000",
  19520=>"000000101",
  19521=>"001001001",
  19522=>"000001001",
  19523=>"010000001",
  19524=>"111111100",
  19525=>"100111111",
  19526=>"111001000",
  19527=>"000001001",
  19528=>"000000000",
  19529=>"011011011",
  19530=>"100000000",
  19531=>"100111111",
  19532=>"110110001",
  19533=>"010000000",
  19534=>"000110110",
  19535=>"000000000",
  19536=>"101000000",
  19537=>"000111111",
  19538=>"000000000",
  19539=>"110110010",
  19540=>"000000000",
  19541=>"101001101",
  19542=>"111111100",
  19543=>"111110100",
  19544=>"111111111",
  19545=>"001001001",
  19546=>"111101101",
  19547=>"011011000",
  19548=>"000000000",
  19549=>"000001001",
  19550=>"000000001",
  19551=>"111111000",
  19552=>"011111111",
  19553=>"000000000",
  19554=>"110111111",
  19555=>"001010111",
  19556=>"100000000",
  19557=>"111110101",
  19558=>"100000101",
  19559=>"000011000",
  19560=>"011011011",
  19561=>"000000000",
  19562=>"010111111",
  19563=>"100110000",
  19564=>"111111000",
  19565=>"000010000",
  19566=>"000100101",
  19567=>"111111111",
  19568=>"000000000",
  19569=>"111111101",
  19570=>"000100111",
  19571=>"100000000",
  19572=>"000000110",
  19573=>"000111111",
  19574=>"000011111",
  19575=>"111111111",
  19576=>"000000000",
  19577=>"001111001",
  19578=>"000010000",
  19579=>"111111111",
  19580=>"000000000",
  19581=>"000100111",
  19582=>"110111110",
  19583=>"000000000",
  19584=>"000011111",
  19585=>"111111111",
  19586=>"101111000",
  19587=>"111111011",
  19588=>"000000000",
  19589=>"000000111",
  19590=>"111111111",
  19591=>"011001111",
  19592=>"010110010",
  19593=>"000000001",
  19594=>"000000111",
  19595=>"000000000",
  19596=>"111111111",
  19597=>"000101111",
  19598=>"111111001",
  19599=>"010111000",
  19600=>"101001111",
  19601=>"000000000",
  19602=>"111001011",
  19603=>"011000000",
  19604=>"000000111",
  19605=>"110010111",
  19606=>"000111111",
  19607=>"000011001",
  19608=>"000000111",
  19609=>"110011111",
  19610=>"111111110",
  19611=>"110001001",
  19612=>"010110110",
  19613=>"001001111",
  19614=>"110111110",
  19615=>"111111111",
  19616=>"111111111",
  19617=>"011111111",
  19618=>"000000100",
  19619=>"111100110",
  19620=>"001001000",
  19621=>"100111011",
  19622=>"000000000",
  19623=>"110111011",
  19624=>"111111110",
  19625=>"001001001",
  19626=>"111010000",
  19627=>"001000000",
  19628=>"111111111",
  19629=>"001000001",
  19630=>"000000110",
  19631=>"101100110",
  19632=>"000111111",
  19633=>"001000000",
  19634=>"011111110",
  19635=>"111110111",
  19636=>"111011000",
  19637=>"000000000",
  19638=>"000111111",
  19639=>"111110010",
  19640=>"101001001",
  19641=>"111111111",
  19642=>"001001001",
  19643=>"110100000",
  19644=>"000111111",
  19645=>"001000100",
  19646=>"111111100",
  19647=>"011111111",
  19648=>"101000000",
  19649=>"001001111",
  19650=>"001000000",
  19651=>"111111111",
  19652=>"000000110",
  19653=>"000000100",
  19654=>"010011011",
  19655=>"011011000",
  19656=>"000000000",
  19657=>"101100000",
  19658=>"001000000",
  19659=>"000000000",
  19660=>"110111000",
  19661=>"001011010",
  19662=>"111110000",
  19663=>"101101101",
  19664=>"001001111",
  19665=>"001000111",
  19666=>"001110110",
  19667=>"111000000",
  19668=>"101111111",
  19669=>"000000101",
  19670=>"001001001",
  19671=>"001000001",
  19672=>"011100101",
  19673=>"111101111",
  19674=>"000111111",
  19675=>"001001000",
  19676=>"100100000",
  19677=>"111110101",
  19678=>"100111111",
  19679=>"010000010",
  19680=>"001001001",
  19681=>"000000000",
  19682=>"001101101",
  19683=>"000000000",
  19684=>"000010100",
  19685=>"110100100",
  19686=>"000000000",
  19687=>"111010111",
  19688=>"111111010",
  19689=>"110010010",
  19690=>"110111110",
  19691=>"000011000",
  19692=>"001000010",
  19693=>"111001111",
  19694=>"001101111",
  19695=>"001000000",
  19696=>"000001001",
  19697=>"000000000",
  19698=>"110100000",
  19699=>"111000000",
  19700=>"110110110",
  19701=>"111011000",
  19702=>"000000001",
  19703=>"111111111",
  19704=>"111011000",
  19705=>"110111111",
  19706=>"111000000",
  19707=>"111011000",
  19708=>"000000000",
  19709=>"000011111",
  19710=>"111001000",
  19711=>"100111111",
  19712=>"111101111",
  19713=>"110110000",
  19714=>"000000000",
  19715=>"000000000",
  19716=>"110111110",
  19717=>"000111111",
  19718=>"111100111",
  19719=>"100000001",
  19720=>"111111111",
  19721=>"111111111",
  19722=>"001000100",
  19723=>"010000000",
  19724=>"101101101",
  19725=>"001000100",
  19726=>"110111101",
  19727=>"000000000",
  19728=>"000000101",
  19729=>"000000000",
  19730=>"111111111",
  19731=>"111111111",
  19732=>"000000100",
  19733=>"111111100",
  19734=>"100100100",
  19735=>"111101111",
  19736=>"101100010",
  19737=>"011001000",
  19738=>"111111111",
  19739=>"000000111",
  19740=>"100000000",
  19741=>"000000001",
  19742=>"000000000",
  19743=>"000110110",
  19744=>"100100001",
  19745=>"000000111",
  19746=>"010010000",
  19747=>"000000000",
  19748=>"000000110",
  19749=>"000100101",
  19750=>"011111010",
  19751=>"000000000",
  19752=>"001001111",
  19753=>"000000000",
  19754=>"110111111",
  19755=>"000000000",
  19756=>"110100110",
  19757=>"001000000",
  19758=>"111111111",
  19759=>"110000010",
  19760=>"000100100",
  19761=>"110110100",
  19762=>"111111111",
  19763=>"010110011",
  19764=>"001001001",
  19765=>"011000010",
  19766=>"000000011",
  19767=>"011111111",
  19768=>"000000000",
  19769=>"011111001",
  19770=>"111001001",
  19771=>"101001110",
  19772=>"110110111",
  19773=>"111111001",
  19774=>"001000000",
  19775=>"111101000",
  19776=>"011111111",
  19777=>"111101000",
  19778=>"101111111",
  19779=>"001001001",
  19780=>"001000101",
  19781=>"110110000",
  19782=>"111111011",
  19783=>"000000000",
  19784=>"000000001",
  19785=>"110110111",
  19786=>"110000000",
  19787=>"000000011",
  19788=>"000000001",
  19789=>"011000110",
  19790=>"101000000",
  19791=>"000000100",
  19792=>"111000000",
  19793=>"001001011",
  19794=>"111111000",
  19795=>"000000000",
  19796=>"000011000",
  19797=>"000000001",
  19798=>"111111110",
  19799=>"100000000",
  19800=>"001000000",
  19801=>"000000011",
  19802=>"101001001",
  19803=>"000000000",
  19804=>"111011000",
  19805=>"000000100",
  19806=>"111111001",
  19807=>"000001001",
  19808=>"001001001",
  19809=>"101001000",
  19810=>"001001011",
  19811=>"111111011",
  19812=>"111111111",
  19813=>"000000000",
  19814=>"000111111",
  19815=>"101001111",
  19816=>"110100101",
  19817=>"001000000",
  19818=>"000010011",
  19819=>"101111101",
  19820=>"110100100",
  19821=>"011111111",
  19822=>"111111111",
  19823=>"001000000",
  19824=>"001001000",
  19825=>"000001001",
  19826=>"000000011",
  19827=>"000011001",
  19828=>"110010010",
  19829=>"001001111",
  19830=>"101000000",
  19831=>"110111110",
  19832=>"111111000",
  19833=>"001001111",
  19834=>"010000000",
  19835=>"000001101",
  19836=>"110000000",
  19837=>"111111111",
  19838=>"111111011",
  19839=>"001001111",
  19840=>"000101101",
  19841=>"001101001",
  19842=>"110110111",
  19843=>"100000000",
  19844=>"110111111",
  19845=>"010000000",
  19846=>"000000001",
  19847=>"001000001",
  19848=>"000000011",
  19849=>"111111111",
  19850=>"000000000",
  19851=>"000000010",
  19852=>"100111111",
  19853=>"100110110",
  19854=>"111001101",
  19855=>"000010111",
  19856=>"101000000",
  19857=>"101111111",
  19858=>"100111111",
  19859=>"101100100",
  19860=>"000001011",
  19861=>"000000010",
  19862=>"110111100",
  19863=>"001001001",
  19864=>"000001101",
  19865=>"000110110",
  19866=>"000001001",
  19867=>"100101000",
  19868=>"010000000",
  19869=>"010010111",
  19870=>"000001101",
  19871=>"011111111",
  19872=>"000001001",
  19873=>"011001001",
  19874=>"111111111",
  19875=>"111011000",
  19876=>"111111111",
  19877=>"010010000",
  19878=>"100001111",
  19879=>"111000000",
  19880=>"111011001",
  19881=>"000000101",
  19882=>"111000000",
  19883=>"000100110",
  19884=>"000000000",
  19885=>"001001101",
  19886=>"111000000",
  19887=>"000100101",
  19888=>"000000100",
  19889=>"001001000",
  19890=>"110110110",
  19891=>"000000100",
  19892=>"001011111",
  19893=>"111001001",
  19894=>"000000000",
  19895=>"110110111",
  19896=>"001001111",
  19897=>"110000000",
  19898=>"000000000",
  19899=>"111111111",
  19900=>"001001000",
  19901=>"001000000",
  19902=>"000000000",
  19903=>"001000000",
  19904=>"111000001",
  19905=>"011111111",
  19906=>"011000011",
  19907=>"110111111",
  19908=>"101000101",
  19909=>"000000001",
  19910=>"000000000",
  19911=>"111111011",
  19912=>"111100000",
  19913=>"001001100",
  19914=>"101000000",
  19915=>"111111111",
  19916=>"011011011",
  19917=>"110111111",
  19918=>"001000100",
  19919=>"010010011",
  19920=>"111000000",
  19921=>"100111001",
  19922=>"000111101",
  19923=>"000001011",
  19924=>"110100000",
  19925=>"000001111",
  19926=>"001110110",
  19927=>"011011011",
  19928=>"000000001",
  19929=>"001001001",
  19930=>"110010000",
  19931=>"111111100",
  19932=>"000000101",
  19933=>"110111001",
  19934=>"101001001",
  19935=>"111111011",
  19936=>"011011011",
  19937=>"001110111",
  19938=>"111111111",
  19939=>"000000110",
  19940=>"000000111",
  19941=>"000010111",
  19942=>"110110111",
  19943=>"111000000",
  19944=>"000000000",
  19945=>"101001001",
  19946=>"000001000",
  19947=>"100100001",
  19948=>"000110111",
  19949=>"100100000",
  19950=>"001000111",
  19951=>"001001001",
  19952=>"000000001",
  19953=>"000000000",
  19954=>"101101101",
  19955=>"000000111",
  19956=>"110111111",
  19957=>"111111111",
  19958=>"001001110",
  19959=>"011111100",
  19960=>"010010000",
  19961=>"011000000",
  19962=>"101101100",
  19963=>"111010111",
  19964=>"001111011",
  19965=>"001001101",
  19966=>"111000000",
  19967=>"001111111",
  19968=>"111111000",
  19969=>"100000110",
  19970=>"000000000",
  19971=>"110111111",
  19972=>"111111000",
  19973=>"111111000",
  19974=>"111000000",
  19975=>"010000000",
  19976=>"111111111",
  19977=>"000000000",
  19978=>"111111101",
  19979=>"000000111",
  19980=>"111001011",
  19981=>"110010010",
  19982=>"000011011",
  19983=>"110100111",
  19984=>"010011000",
  19985=>"111000101",
  19986=>"011000000",
  19987=>"111111000",
  19988=>"111111111",
  19989=>"000111111",
  19990=>"010000100",
  19991=>"111000000",
  19992=>"111111111",
  19993=>"101000000",
  19994=>"000000001",
  19995=>"110000000",
  19996=>"011111111",
  19997=>"001000001",
  19998=>"111011011",
  19999=>"111111111",
  20000=>"111111110",
  20001=>"100001000",
  20002=>"011111011",
  20003=>"000111001",
  20004=>"001001000",
  20005=>"000000110",
  20006=>"111000000",
  20007=>"100100111",
  20008=>"000000111",
  20009=>"000000000",
  20010=>"111100100",
  20011=>"000111110",
  20012=>"011111000",
  20013=>"000100111",
  20014=>"000000001",
  20015=>"000110110",
  20016=>"000000100",
  20017=>"111000101",
  20018=>"001111111",
  20019=>"000001001",
  20020=>"110100101",
  20021=>"111001001",
  20022=>"010010110",
  20023=>"111011001",
  20024=>"000100111",
  20025=>"111111101",
  20026=>"000101000",
  20027=>"000000000",
  20028=>"011001111",
  20029=>"000000001",
  20030=>"000000100",
  20031=>"000111111",
  20032=>"111111111",
  20033=>"000110111",
  20034=>"001000000",
  20035=>"000101000",
  20036=>"111111011",
  20037=>"011000000",
  20038=>"000000000",
  20039=>"111111111",
  20040=>"000110110",
  20041=>"000000000",
  20042=>"111000000",
  20043=>"111111101",
  20044=>"111111111",
  20045=>"000000000",
  20046=>"001000000",
  20047=>"111111111",
  20048=>"000101111",
  20049=>"000111000",
  20050=>"111111111",
  20051=>"111111110",
  20052=>"000000000",
  20053=>"000000100",
  20054=>"000110111",
  20055=>"000000000",
  20056=>"111111111",
  20057=>"001011111",
  20058=>"000111110",
  20059=>"000110111",
  20060=>"110000000",
  20061=>"000111111",
  20062=>"111011110",
  20063=>"000111110",
  20064=>"111111001",
  20065=>"111001001",
  20066=>"000110111",
  20067=>"111110010",
  20068=>"111011011",
  20069=>"000000001",
  20070=>"000000000",
  20071=>"001000110",
  20072=>"000111001",
  20073=>"111111001",
  20074=>"100111111",
  20075=>"000011111",
  20076=>"110000001",
  20077=>"010000000",
  20078=>"000000000",
  20079=>"000000000",
  20080=>"000000110",
  20081=>"000000001",
  20082=>"101111110",
  20083=>"111101000",
  20084=>"000001000",
  20085=>"111111000",
  20086=>"000111111",
  20087=>"111111100",
  20088=>"001011010",
  20089=>"111010011",
  20090=>"111101001",
  20091=>"000000000",
  20092=>"000011001",
  20093=>"000001001",
  20094=>"111111000",
  20095=>"010110010",
  20096=>"111000000",
  20097=>"000000001",
  20098=>"111010000",
  20099=>"000110000",
  20100=>"100000101",
  20101=>"000000000",
  20102=>"110111111",
  20103=>"111001001",
  20104=>"000111111",
  20105=>"111000000",
  20106=>"000000111",
  20107=>"010010111",
  20108=>"000001001",
  20109=>"000110000",
  20110=>"111100000",
  20111=>"000000111",
  20112=>"111111111",
  20113=>"111111000",
  20114=>"111111101",
  20115=>"111111000",
  20116=>"000010010",
  20117=>"111010000",
  20118=>"110111111",
  20119=>"000101111",
  20120=>"110000000",
  20121=>"111001000",
  20122=>"000000011",
  20123=>"111111111",
  20124=>"001001000",
  20125=>"111101111",
  20126=>"000000111",
  20127=>"111101110",
  20128=>"000111110",
  20129=>"000011011",
  20130=>"111101111",
  20131=>"000000110",
  20132=>"111001011",
  20133=>"111101001",
  20134=>"111111101",
  20135=>"000100100",
  20136=>"000011011",
  20137=>"111110111",
  20138=>"011001000",
  20139=>"000000001",
  20140=>"111111111",
  20141=>"000111011",
  20142=>"000111111",
  20143=>"000000000",
  20144=>"111111111",
  20145=>"011001000",
  20146=>"101101111",
  20147=>"101000000",
  20148=>"011010110",
  20149=>"000000000",
  20150=>"110111111",
  20151=>"100000000",
  20152=>"110110110",
  20153=>"101000100",
  20154=>"111000110",
  20155=>"100000001",
  20156=>"000000000",
  20157=>"000000101",
  20158=>"000000000",
  20159=>"111111111",
  20160=>"000000100",
  20161=>"111111111",
  20162=>"111110000",
  20163=>"000000000",
  20164=>"111111111",
  20165=>"000000000",
  20166=>"010000000",
  20167=>"111111111",
  20168=>"000000000",
  20169=>"000001000",
  20170=>"011000000",
  20171=>"111111111",
  20172=>"010110000",
  20173=>"111111111",
  20174=>"100100100",
  20175=>"000000000",
  20176=>"111001000",
  20177=>"111111111",
  20178=>"111111111",
  20179=>"111111000",
  20180=>"100100101",
  20181=>"111111100",
  20182=>"000000000",
  20183=>"111111000",
  20184=>"001000000",
  20185=>"100100000",
  20186=>"000000000",
  20187=>"000011010",
  20188=>"111110000",
  20189=>"000100100",
  20190=>"001101101",
  20191=>"000000000",
  20192=>"000000111",
  20193=>"001000000",
  20194=>"000000110",
  20195=>"000111111",
  20196=>"111000001",
  20197=>"000000011",
  20198=>"000000000",
  20199=>"011111111",
  20200=>"111000000",
  20201=>"111111110",
  20202=>"110110110",
  20203=>"010000000",
  20204=>"110111110",
  20205=>"000000000",
  20206=>"111111011",
  20207=>"111111111",
  20208=>"000111111",
  20209=>"110110111",
  20210=>"000000000",
  20211=>"000000110",
  20212=>"000111111",
  20213=>"001111111",
  20214=>"001001001",
  20215=>"000111111",
  20216=>"111011000",
  20217=>"000000000",
  20218=>"000111111",
  20219=>"100111001",
  20220=>"000100100",
  20221=>"011000000",
  20222=>"100101001",
  20223=>"000111111",
  20224=>"000000000",
  20225=>"000000001",
  20226=>"111000000",
  20227=>"000110110",
  20228=>"000000011",
  20229=>"001001001",
  20230=>"011001000",
  20231=>"111111111",
  20232=>"100100000",
  20233=>"111011011",
  20234=>"111111011",
  20235=>"000101111",
  20236=>"111111001",
  20237=>"001001111",
  20238=>"111000000",
  20239=>"111111111",
  20240=>"000000000",
  20241=>"111000000",
  20242=>"000000000",
  20243=>"000000101",
  20244=>"111111000",
  20245=>"000000000",
  20246=>"001011011",
  20247=>"111000111",
  20248=>"111000111",
  20249=>"111111111",
  20250=>"000000000",
  20251=>"111011001",
  20252=>"111111111",
  20253=>"111101101",
  20254=>"110111000",
  20255=>"111000000",
  20256=>"111111101",
  20257=>"001000000",
  20258=>"101100100",
  20259=>"110110110",
  20260=>"000000000",
  20261=>"111111111",
  20262=>"100100110",
  20263=>"111001001",
  20264=>"111000100",
  20265=>"000110000",
  20266=>"000011000",
  20267=>"111000000",
  20268=>"000110110",
  20269=>"111110000",
  20270=>"111000111",
  20271=>"000000111",
  20272=>"000000000",
  20273=>"110000000",
  20274=>"111111110",
  20275=>"111000000",
  20276=>"110110111",
  20277=>"111111111",
  20278=>"000000000",
  20279=>"000000011",
  20280=>"001000100",
  20281=>"111110111",
  20282=>"111000011",
  20283=>"111111011",
  20284=>"010011000",
  20285=>"011111111",
  20286=>"000000111",
  20287=>"111110111",
  20288=>"111000000",
  20289=>"000000111",
  20290=>"000000001",
  20291=>"001001111",
  20292=>"000000111",
  20293=>"100001111",
  20294=>"110000000",
  20295=>"111000000",
  20296=>"111111111",
  20297=>"111111111",
  20298=>"000000010",
  20299=>"111001000",
  20300=>"110000001",
  20301=>"000000000",
  20302=>"000001111",
  20303=>"111100100",
  20304=>"001000000",
  20305=>"001000111",
  20306=>"111110111",
  20307=>"111111111",
  20308=>"000111111",
  20309=>"111011000",
  20310=>"100100110",
  20311=>"110111111",
  20312=>"000000000",
  20313=>"011000111",
  20314=>"000000110",
  20315=>"111111000",
  20316=>"000111111",
  20317=>"111111001",
  20318=>"111000110",
  20319=>"000110001",
  20320=>"111000000",
  20321=>"111000000",
  20322=>"110100100",
  20323=>"011011111",
  20324=>"000001111",
  20325=>"010000000",
  20326=>"000000001",
  20327=>"001000000",
  20328=>"111111001",
  20329=>"000001000",
  20330=>"111100100",
  20331=>"000011111",
  20332=>"100111110",
  20333=>"110000000",
  20334=>"011000000",
  20335=>"000000000",
  20336=>"110000000",
  20337=>"000000111",
  20338=>"000000111",
  20339=>"111111111",
  20340=>"000000100",
  20341=>"111111111",
  20342=>"111111111",
  20343=>"001000000",
  20344=>"111111111",
  20345=>"100000111",
  20346=>"000000000",
  20347=>"000111111",
  20348=>"000000000",
  20349=>"111000000",
  20350=>"000010010",
  20351=>"111000000",
  20352=>"000011111",
  20353=>"011000111",
  20354=>"110100000",
  20355=>"000000000",
  20356=>"110000111",
  20357=>"000000000",
  20358=>"000000000",
  20359=>"010011000",
  20360=>"111000000",
  20361=>"110000001",
  20362=>"111000000",
  20363=>"000000000",
  20364=>"000000000",
  20365=>"101111000",
  20366=>"100100110",
  20367=>"111000000",
  20368=>"000000000",
  20369=>"000011001",
  20370=>"111100000",
  20371=>"000000001",
  20372=>"101101111",
  20373=>"111000000",
  20374=>"000111011",
  20375=>"000011011",
  20376=>"000000000",
  20377=>"111110111",
  20378=>"110111111",
  20379=>"111100000",
  20380=>"111011000",
  20381=>"101101111",
  20382=>"001000000",
  20383=>"111111111",
  20384=>"011011000",
  20385=>"111001001",
  20386=>"000111111",
  20387=>"000000000",
  20388=>"000110110",
  20389=>"000100111",
  20390=>"100000000",
  20391=>"111001000",
  20392=>"010000110",
  20393=>"110010010",
  20394=>"000000000",
  20395=>"011001001",
  20396=>"010011011",
  20397=>"000001000",
  20398=>"000110100",
  20399=>"111111110",
  20400=>"111000100",
  20401=>"000000100",
  20402=>"111111111",
  20403=>"001000111",
  20404=>"000000000",
  20405=>"100111111",
  20406=>"000000111",
  20407=>"000000110",
  20408=>"000111100",
  20409=>"011111001",
  20410=>"010000000",
  20411=>"000010111",
  20412=>"001100001",
  20413=>"111111110",
  20414=>"000111000",
  20415=>"110100000",
  20416=>"111111111",
  20417=>"000000000",
  20418=>"000000000",
  20419=>"000000011",
  20420=>"011111101",
  20421=>"100110100",
  20422=>"101001000",
  20423=>"000011000",
  20424=>"111110000",
  20425=>"011111111",
  20426=>"110111111",
  20427=>"111001111",
  20428=>"111000000",
  20429=>"001011000",
  20430=>"111111001",
  20431=>"000000000",
  20432=>"000000000",
  20433=>"110010001",
  20434=>"111111111",
  20435=>"111001011",
  20436=>"010100110",
  20437=>"000001011",
  20438=>"001000000",
  20439=>"000100100",
  20440=>"011000000",
  20441=>"000000011",
  20442=>"011000111",
  20443=>"000011011",
  20444=>"000000101",
  20445=>"000000101",
  20446=>"111111111",
  20447=>"110111111",
  20448=>"000000000",
  20449=>"000000000",
  20450=>"111111101",
  20451=>"010000000",
  20452=>"110000000",
  20453=>"111111111",
  20454=>"111111000",
  20455=>"000000000",
  20456=>"010110111",
  20457=>"111111111",
  20458=>"000000000",
  20459=>"111110000",
  20460=>"000000000",
  20461=>"000110110",
  20462=>"001000000",
  20463=>"010000000",
  20464=>"111100111",
  20465=>"111011100",
  20466=>"011111111",
  20467=>"101101111",
  20468=>"111111011",
  20469=>"000000100",
  20470=>"100101001",
  20471=>"111111110",
  20472=>"100000000",
  20473=>"010000011",
  20474=>"000001000",
  20475=>"000000000",
  20476=>"111111111",
  20477=>"000000000",
  20478=>"000111111",
  20479=>"111011111",
  20480=>"011111111",
  20481=>"000111000",
  20482=>"000000101",
  20483=>"000000000",
  20484=>"100100110",
  20485=>"000001111",
  20486=>"001000000",
  20487=>"000000100",
  20488=>"111111111",
  20489=>"111111111",
  20490=>"000001111",
  20491=>"111000000",
  20492=>"111111111",
  20493=>"111111100",
  20494=>"111111010",
  20495=>"111101100",
  20496=>"111111111",
  20497=>"000010011",
  20498=>"000001111",
  20499=>"000000110",
  20500=>"000000000",
  20501=>"000000111",
  20502=>"000000000",
  20503=>"111110000",
  20504=>"100000111",
  20505=>"111111001",
  20506=>"111110110",
  20507=>"011000000",
  20508=>"111111111",
  20509=>"001100011",
  20510=>"000000110",
  20511=>"000000111",
  20512=>"100100101",
  20513=>"111111111",
  20514=>"111111011",
  20515=>"111111111",
  20516=>"000001111",
  20517=>"111001001",
  20518=>"100010011",
  20519=>"011011010",
  20520=>"000000101",
  20521=>"111111111",
  20522=>"000000000",
  20523=>"111000000",
  20524=>"010110110",
  20525=>"111111000",
  20526=>"110111111",
  20527=>"111111111",
  20528=>"111111110",
  20529=>"000000000",
  20530=>"100111111",
  20531=>"000000000",
  20532=>"000000111",
  20533=>"111101100",
  20534=>"001000000",
  20535=>"101000000",
  20536=>"000111111",
  20537=>"011100110",
  20538=>"111111111",
  20539=>"111111111",
  20540=>"111110111",
  20541=>"011000000",
  20542=>"000000000",
  20543=>"011000100",
  20544=>"000000000",
  20545=>"110111111",
  20546=>"010000000",
  20547=>"000000000",
  20548=>"001001111",
  20549=>"111111111",
  20550=>"000000111",
  20551=>"000000000",
  20552=>"110111111",
  20553=>"000000111",
  20554=>"000000000",
  20555=>"000000111",
  20556=>"000100111",
  20557=>"111111111",
  20558=>"111101000",
  20559=>"000001010",
  20560=>"111000011",
  20561=>"000001001",
  20562=>"000000000",
  20563=>"001000000",
  20564=>"001001011",
  20565=>"000000000",
  20566=>"101011111",
  20567=>"000111100",
  20568=>"001001001",
  20569=>"100000100",
  20570=>"111001000",
  20571=>"010010010",
  20572=>"111111110",
  20573=>"000000000",
  20574=>"001001101",
  20575=>"000000000",
  20576=>"000010110",
  20577=>"000000001",
  20578=>"000000000",
  20579=>"000000000",
  20580=>"000000000",
  20581=>"001000000",
  20582=>"111111111",
  20583=>"000000000",
  20584=>"011111111",
  20585=>"110000000",
  20586=>"000000111",
  20587=>"001000001",
  20588=>"111110110",
  20589=>"011111110",
  20590=>"000000101",
  20591=>"001000001",
  20592=>"110111010",
  20593=>"000111111",
  20594=>"100000000",
  20595=>"010011000",
  20596=>"000000000",
  20597=>"101001001",
  20598=>"000000000",
  20599=>"000000000",
  20600=>"000000000",
  20601=>"111111000",
  20602=>"000000010",
  20603=>"110100111",
  20604=>"100100100",
  20605=>"001000001",
  20606=>"000000000",
  20607=>"110100111",
  20608=>"101100001",
  20609=>"100111111",
  20610=>"000000000",
  20611=>"110100000",
  20612=>"001001000",
  20613=>"001001111",
  20614=>"001111011",
  20615=>"011111111",
  20616=>"111111111",
  20617=>"111110000",
  20618=>"000000000",
  20619=>"111111110",
  20620=>"011111111",
  20621=>"000000000",
  20622=>"101000000",
  20623=>"111111111",
  20624=>"000000000",
  20625=>"000000011",
  20626=>"101111111",
  20627=>"111111111",
  20628=>"001001100",
  20629=>"111111001",
  20630=>"111001000",
  20631=>"000000000",
  20632=>"000000001",
  20633=>"000110110",
  20634=>"101111001",
  20635=>"001001001",
  20636=>"001000001",
  20637=>"100100110",
  20638=>"110110110",
  20639=>"111111011",
  20640=>"101000000",
  20641=>"101100010",
  20642=>"111110111",
  20643=>"100000111",
  20644=>"001100110",
  20645=>"011000011",
  20646=>"000000101",
  20647=>"011111000",
  20648=>"111100100",
  20649=>"000000000",
  20650=>"001000001",
  20651=>"000010110",
  20652=>"001000111",
  20653=>"100100100",
  20654=>"110110110",
  20655=>"000000000",
  20656=>"111110000",
  20657=>"111101001",
  20658=>"110111111",
  20659=>"000000000",
  20660=>"110111010",
  20661=>"110000000",
  20662=>"100100000",
  20663=>"111011011",
  20664=>"101000000",
  20665=>"111111111",
  20666=>"000000000",
  20667=>"111001001",
  20668=>"000100000",
  20669=>"001111111",
  20670=>"111111101",
  20671=>"111011110",
  20672=>"111111111",
  20673=>"000000000",
  20674=>"101000000",
  20675=>"000000111",
  20676=>"000010111",
  20677=>"111001000",
  20678=>"111111000",
  20679=>"010010010",
  20680=>"100000000",
  20681=>"111011111",
  20682=>"000000000",
  20683=>"111111111",
  20684=>"000010111",
  20685=>"000000000",
  20686=>"001000000",
  20687=>"001000000",
  20688=>"000000000",
  20689=>"000111111",
  20690=>"000110111",
  20691=>"111111111",
  20692=>"111111010",
  20693=>"101000000",
  20694=>"001101111",
  20695=>"110110100",
  20696=>"000000110",
  20697=>"110110110",
  20698=>"111111111",
  20699=>"111111111",
  20700=>"111100110",
  20701=>"110110000",
  20702=>"000011011",
  20703=>"011000001",
  20704=>"111000000",
  20705=>"000000000",
  20706=>"111000111",
  20707=>"101000111",
  20708=>"000001000",
  20709=>"001001001",
  20710=>"001000100",
  20711=>"100000111",
  20712=>"111011000",
  20713=>"000110110",
  20714=>"111111110",
  20715=>"001000000",
  20716=>"001001101",
  20717=>"111101001",
  20718=>"000111111",
  20719=>"000111111",
  20720=>"000000100",
  20721=>"111111111",
  20722=>"000101101",
  20723=>"111000000",
  20724=>"111111111",
  20725=>"000000000",
  20726=>"000000100",
  20727=>"001000000",
  20728=>"111111111",
  20729=>"111111100",
  20730=>"000000001",
  20731=>"001000111",
  20732=>"110110110",
  20733=>"100110000",
  20734=>"001001111",
  20735=>"111111011",
  20736=>"111000011",
  20737=>"110110110",
  20738=>"000000111",
  20739=>"111111111",
  20740=>"000000000",
  20741=>"111111111",
  20742=>"100100000",
  20743=>"100100000",
  20744=>"000000000",
  20745=>"000000000",
  20746=>"111111001",
  20747=>"000000000",
  20748=>"000000001",
  20749=>"000000100",
  20750=>"000000111",
  20751=>"111111111",
  20752=>"000000000",
  20753=>"000000000",
  20754=>"110110000",
  20755=>"000000010",
  20756=>"000000000",
  20757=>"011001000",
  20758=>"110111111",
  20759=>"111111111",
  20760=>"111111000",
  20761=>"100100000",
  20762=>"000001001",
  20763=>"010110010",
  20764=>"111111111",
  20765=>"011111111",
  20766=>"001000001",
  20767=>"111010010",
  20768=>"111011001",
  20769=>"111111111",
  20770=>"011000000",
  20771=>"111111101",
  20772=>"111100000",
  20773=>"111100000",
  20774=>"110110110",
  20775=>"011010000",
  20776=>"000101111",
  20777=>"000000010",
  20778=>"111111000",
  20779=>"110110011",
  20780=>"111101101",
  20781=>"101101100",
  20782=>"110111000",
  20783=>"000000000",
  20784=>"000111011",
  20785=>"111110110",
  20786=>"111111111",
  20787=>"000111111",
  20788=>"110000000",
  20789=>"111111011",
  20790=>"011001011",
  20791=>"000000001",
  20792=>"111011001",
  20793=>"000000111",
  20794=>"111001001",
  20795=>"111000000",
  20796=>"111000110",
  20797=>"000000000",
  20798=>"011001000",
  20799=>"111111111",
  20800=>"111101100",
  20801=>"111111111",
  20802=>"000010011",
  20803=>"111111111",
  20804=>"111100100",
  20805=>"111011011",
  20806=>"001111111",
  20807=>"001001000",
  20808=>"011011001",
  20809=>"000000000",
  20810=>"111111000",
  20811=>"100000000",
  20812=>"000000001",
  20813=>"110111010",
  20814=>"111001111",
  20815=>"000110100",
  20816=>"111111101",
  20817=>"110101101",
  20818=>"111111111",
  20819=>"111111100",
  20820=>"111111111",
  20821=>"001011011",
  20822=>"111111000",
  20823=>"000000000",
  20824=>"111111101",
  20825=>"000110111",
  20826=>"100000000",
  20827=>"000000000",
  20828=>"100100000",
  20829=>"000011010",
  20830=>"100100111",
  20831=>"111110000",
  20832=>"110110000",
  20833=>"100101000",
  20834=>"100110111",
  20835=>"111111111",
  20836=>"000001111",
  20837=>"000000000",
  20838=>"111101111",
  20839=>"111110110",
  20840=>"110100000",
  20841=>"001111110",
  20842=>"000000000",
  20843=>"000110110",
  20844=>"011110111",
  20845=>"000000100",
  20846=>"001001001",
  20847=>"111111111",
  20848=>"000000111",
  20849=>"011000111",
  20850=>"100111111",
  20851=>"010000000",
  20852=>"000000010",
  20853=>"000000100",
  20854=>"000000111",
  20855=>"001000000",
  20856=>"000000000",
  20857=>"111110110",
  20858=>"000000000",
  20859=>"011001011",
  20860=>"011011011",
  20861=>"101000000",
  20862=>"000000000",
  20863=>"111101000",
  20864=>"111100111",
  20865=>"111011111",
  20866=>"111011011",
  20867=>"000000000",
  20868=>"011110000",
  20869=>"111111000",
  20870=>"000001111",
  20871=>"111011000",
  20872=>"000000000",
  20873=>"111111110",
  20874=>"000000000",
  20875=>"000000000",
  20876=>"111000000",
  20877=>"100101011",
  20878=>"111111111",
  20879=>"111111111",
  20880=>"000000000",
  20881=>"000000111",
  20882=>"000110111",
  20883=>"111001011",
  20884=>"111000111",
  20885=>"000000011",
  20886=>"000000000",
  20887=>"100000000",
  20888=>"000000000",
  20889=>"111111110",
  20890=>"001000101",
  20891=>"000000011",
  20892=>"101000001",
  20893=>"000000111",
  20894=>"000101101",
  20895=>"000000000",
  20896=>"111111111",
  20897=>"111110110",
  20898=>"110000011",
  20899=>"111011000",
  20900=>"111111111",
  20901=>"000010010",
  20902=>"000000000",
  20903=>"111111000",
  20904=>"000001001",
  20905=>"000000000",
  20906=>"001000000",
  20907=>"111101000",
  20908=>"001000000",
  20909=>"111000000",
  20910=>"111000110",
  20911=>"010000000",
  20912=>"001000100",
  20913=>"000000000",
  20914=>"000000100",
  20915=>"111011010",
  20916=>"100000100",
  20917=>"000000000",
  20918=>"100000000",
  20919=>"011111110",
  20920=>"000111111",
  20921=>"111100000",
  20922=>"000000001",
  20923=>"001000000",
  20924=>"000111111",
  20925=>"111111110",
  20926=>"111111100",
  20927=>"111101101",
  20928=>"000000000",
  20929=>"100110110",
  20930=>"101100101",
  20931=>"000001000",
  20932=>"111111100",
  20933=>"001000000",
  20934=>"111011010",
  20935=>"000000000",
  20936=>"011110000",
  20937=>"000000000",
  20938=>"000000000",
  20939=>"000000000",
  20940=>"111111111",
  20941=>"111011000",
  20942=>"000000000",
  20943=>"111111111",
  20944=>"100100100",
  20945=>"111111111",
  20946=>"011011001",
  20947=>"000000000",
  20948=>"000000100",
  20949=>"111111111",
  20950=>"000000000",
  20951=>"111111011",
  20952=>"111100111",
  20953=>"011001111",
  20954=>"000000000",
  20955=>"011000000",
  20956=>"011011111",
  20957=>"000000000",
  20958=>"110111000",
  20959=>"110100110",
  20960=>"011111111",
  20961=>"110111001",
  20962=>"111000011",
  20963=>"111111111",
  20964=>"111111000",
  20965=>"111011101",
  20966=>"111111100",
  20967=>"000000000",
  20968=>"110010000",
  20969=>"011001111",
  20970=>"101111111",
  20971=>"110111111",
  20972=>"000100111",
  20973=>"111001001",
  20974=>"100000000",
  20975=>"000000000",
  20976=>"101001100",
  20977=>"111000000",
  20978=>"100000000",
  20979=>"110000000",
  20980=>"111111111",
  20981=>"010000000",
  20982=>"100100100",
  20983=>"111111101",
  20984=>"000000000",
  20985=>"001101111",
  20986=>"110110110",
  20987=>"101000001",
  20988=>"000000110",
  20989=>"111000000",
  20990=>"001000000",
  20991=>"100000000",
  20992=>"110011011",
  20993=>"000111110",
  20994=>"000000000",
  20995=>"001111000",
  20996=>"001001101",
  20997=>"000000000",
  20998=>"000000111",
  20999=>"000000111",
  21000=>"000000000",
  21001=>"000000000",
  21002=>"101101111",
  21003=>"000011111",
  21004=>"011111110",
  21005=>"100111000",
  21006=>"001000000",
  21007=>"000010000",
  21008=>"111111110",
  21009=>"101000000",
  21010=>"111000000",
  21011=>"111111111",
  21012=>"111111111",
  21013=>"110111111",
  21014=>"110000000",
  21015=>"100000000",
  21016=>"110100100",
  21017=>"011011111",
  21018=>"010011011",
  21019=>"100111000",
  21020=>"111111111",
  21021=>"110111100",
  21022=>"111111110",
  21023=>"111111101",
  21024=>"111101001",
  21025=>"100100000",
  21026=>"000000000",
  21027=>"000011000",
  21028=>"011000000",
  21029=>"001101000",
  21030=>"000000000",
  21031=>"000111011",
  21032=>"111111110",
  21033=>"000000000",
  21034=>"000000000",
  21035=>"000110000",
  21036=>"000000000",
  21037=>"001000000",
  21038=>"111111000",
  21039=>"100100110",
  21040=>"000000001",
  21041=>"111000100",
  21042=>"100100100",
  21043=>"010111100",
  21044=>"110010111",
  21045=>"000000000",
  21046=>"000000000",
  21047=>"111111111",
  21048=>"000110110",
  21049=>"000000000",
  21050=>"000000000",
  21051=>"111111000",
  21052=>"001001111",
  21053=>"000111011",
  21054=>"000000000",
  21055=>"000010011",
  21056=>"000000000",
  21057=>"111111111",
  21058=>"000000001",
  21059=>"000000011",
  21060=>"111111000",
  21061=>"010111111",
  21062=>"000100110",
  21063=>"111111111",
  21064=>"001001011",
  21065=>"000000001",
  21066=>"000000000",
  21067=>"011001001",
  21068=>"000000000",
  21069=>"111001111",
  21070=>"100000000",
  21071=>"001000000",
  21072=>"001011011",
  21073=>"000000000",
  21074=>"010110110",
  21075=>"111111001",
  21076=>"111111111",
  21077=>"000010010",
  21078=>"000111001",
  21079=>"100111111",
  21080=>"101111110",
  21081=>"000000000",
  21082=>"000000000",
  21083=>"001111111",
  21084=>"100000101",
  21085=>"101000000",
  21086=>"111111111",
  21087=>"111111110",
  21088=>"110001000",
  21089=>"001000000",
  21090=>"111110000",
  21091=>"111111111",
  21092=>"111110010",
  21093=>"000000001",
  21094=>"001001000",
  21095=>"110000000",
  21096=>"011111111",
  21097=>"010000000",
  21098=>"000100111",
  21099=>"100100000",
  21100=>"000011001",
  21101=>"000110000",
  21102=>"100111110",
  21103=>"111111011",
  21104=>"100101001",
  21105=>"111000000",
  21106=>"111101000",
  21107=>"000001001",
  21108=>"000101111",
  21109=>"110110000",
  21110=>"111111111",
  21111=>"110010000",
  21112=>"100000000",
  21113=>"000000101",
  21114=>"111101100",
  21115=>"001000000",
  21116=>"011011000",
  21117=>"101001111",
  21118=>"111001000",
  21119=>"111111111",
  21120=>"010000001",
  21121=>"000111111",
  21122=>"000000000",
  21123=>"000100000",
  21124=>"100000000",
  21125=>"000110111",
  21126=>"000111111",
  21127=>"111101111",
  21128=>"000110000",
  21129=>"000110110",
  21130=>"111100110",
  21131=>"111111110",
  21132=>"001010111",
  21133=>"111111110",
  21134=>"111110010",
  21135=>"000001101",
  21136=>"111111011",
  21137=>"111111111",
  21138=>"111011001",
  21139=>"111111110",
  21140=>"000111111",
  21141=>"111100100",
  21142=>"000111011",
  21143=>"000100110",
  21144=>"011101101",
  21145=>"111111111",
  21146=>"001101001",
  21147=>"111011111",
  21148=>"011111001",
  21149=>"111001000",
  21150=>"100100100",
  21151=>"000111111",
  21152=>"000111111",
  21153=>"011111111",
  21154=>"000000000",
  21155=>"001001001",
  21156=>"100000000",
  21157=>"000110110",
  21158=>"000100111",
  21159=>"000000000",
  21160=>"000100110",
  21161=>"000000000",
  21162=>"001000000",
  21163=>"000000000",
  21164=>"000001000",
  21165=>"011111111",
  21166=>"001001000",
  21167=>"111111000",
  21168=>"001111111",
  21169=>"001000111",
  21170=>"111110111",
  21171=>"000000000",
  21172=>"000000100",
  21173=>"111000000",
  21174=>"111011011",
  21175=>"111011000",
  21176=>"000111011",
  21177=>"100000001",
  21178=>"101001111",
  21179=>"111001001",
  21180=>"000000000",
  21181=>"111111111",
  21182=>"110111111",
  21183=>"111011111",
  21184=>"010110010",
  21185=>"100100000",
  21186=>"001011111",
  21187=>"101000000",
  21188=>"000000000",
  21189=>"000000000",
  21190=>"111111111",
  21191=>"000111111",
  21192=>"100111111",
  21193=>"000000001",
  21194=>"001111000",
  21195=>"111000111",
  21196=>"000000000",
  21197=>"000100110",
  21198=>"001000000",
  21199=>"111111111",
  21200=>"000000000",
  21201=>"111111111",
  21202=>"000000000",
  21203=>"000001111",
  21204=>"111110000",
  21205=>"001111111",
  21206=>"111010000",
  21207=>"000000000",
  21208=>"111011010",
  21209=>"111111111",
  21210=>"000000000",
  21211=>"000111011",
  21212=>"111111011",
  21213=>"000000111",
  21214=>"000000100",
  21215=>"000100000",
  21216=>"111111111",
  21217=>"111101101",
  21218=>"000111111",
  21219=>"111111111",
  21220=>"000000110",
  21221=>"111111110",
  21222=>"001001000",
  21223=>"111111111",
  21224=>"111111011",
  21225=>"010110111",
  21226=>"000000000",
  21227=>"111101000",
  21228=>"111111010",
  21229=>"111011001",
  21230=>"111000000",
  21231=>"111101110",
  21232=>"111110110",
  21233=>"100000000",
  21234=>"110100111",
  21235=>"000001010",
  21236=>"001111111",
  21237=>"011011011",
  21238=>"000000000",
  21239=>"100000000",
  21240=>"111000000",
  21241=>"111111111",
  21242=>"001111111",
  21243=>"111000000",
  21244=>"000001011",
  21245=>"000000000",
  21246=>"111111111",
  21247=>"010111111",
  21248=>"001000000",
  21249=>"011111011",
  21250=>"111111110",
  21251=>"100110110",
  21252=>"000111111",
  21253=>"000010000",
  21254=>"111111111",
  21255=>"001111000",
  21256=>"001101101",
  21257=>"111111111",
  21258=>"000000000",
  21259=>"001111111",
  21260=>"000000110",
  21261=>"111111111",
  21262=>"111111111",
  21263=>"000110111",
  21264=>"111111111",
  21265=>"001001000",
  21266=>"010000010",
  21267=>"001001011",
  21268=>"000000000",
  21269=>"000101000",
  21270=>"011011011",
  21271=>"000000001",
  21272=>"111110110",
  21273=>"111111000",
  21274=>"000011000",
  21275=>"100100110",
  21276=>"111111111",
  21277=>"000000000",
  21278=>"000000000",
  21279=>"000000001",
  21280=>"011110010",
  21281=>"000110110",
  21282=>"000010110",
  21283=>"011011000",
  21284=>"000011001",
  21285=>"111111111",
  21286=>"100100110",
  21287=>"011000000",
  21288=>"111111110",
  21289=>"110110110",
  21290=>"001111010",
  21291=>"100111010",
  21292=>"100101101",
  21293=>"000000111",
  21294=>"000000000",
  21295=>"000000000",
  21296=>"000000000",
  21297=>"111001001",
  21298=>"000010110",
  21299=>"111111111",
  21300=>"111111111",
  21301=>"000000000",
  21302=>"000100111",
  21303=>"111000000",
  21304=>"000000001",
  21305=>"000000100",
  21306=>"000000100",
  21307=>"000000000",
  21308=>"110111111",
  21309=>"000100000",
  21310=>"110100100",
  21311=>"110011111",
  21312=>"000000000",
  21313=>"111111110",
  21314=>"001011111",
  21315=>"111100000",
  21316=>"111100111",
  21317=>"000000111",
  21318=>"110110111",
  21319=>"101000001",
  21320=>"000000001",
  21321=>"111001000",
  21322=>"000111110",
  21323=>"110110010",
  21324=>"111111000",
  21325=>"001000001",
  21326=>"000111110",
  21327=>"000000000",
  21328=>"110110100",
  21329=>"111100110",
  21330=>"001111111",
  21331=>"110110100",
  21332=>"111111111",
  21333=>"111110111",
  21334=>"111111111",
  21335=>"000000010",
  21336=>"000111111",
  21337=>"111111111",
  21338=>"000010111",
  21339=>"000000000",
  21340=>"001011111",
  21341=>"000000000",
  21342=>"011110110",
  21343=>"111001011",
  21344=>"000110100",
  21345=>"000000000",
  21346=>"110100110",
  21347=>"000000000",
  21348=>"000010110",
  21349=>"000000000",
  21350=>"011011000",
  21351=>"001011111",
  21352=>"011011001",
  21353=>"000110000",
  21354=>"010111000",
  21355=>"010011000",
  21356=>"000011001",
  21357=>"111111111",
  21358=>"000100110",
  21359=>"000000010",
  21360=>"000000000",
  21361=>"000000000",
  21362=>"111011010",
  21363=>"110111111",
  21364=>"000001001",
  21365=>"100111111",
  21366=>"111001011",
  21367=>"100100001",
  21368=>"111000000",
  21369=>"001111111",
  21370=>"000000001",
  21371=>"111101001",
  21372=>"010111111",
  21373=>"000000000",
  21374=>"000100110",
  21375=>"111110110",
  21376=>"000000000",
  21377=>"111000111",
  21378=>"000010000",
  21379=>"000000001",
  21380=>"000000000",
  21381=>"111101111",
  21382=>"011001000",
  21383=>"000100100",
  21384=>"110000000",
  21385=>"111111100",
  21386=>"111111001",
  21387=>"111111111",
  21388=>"111111111",
  21389=>"010010011",
  21390=>"001001110",
  21391=>"111110110",
  21392=>"111111111",
  21393=>"000000000",
  21394=>"001011011",
  21395=>"001011010",
  21396=>"001000000",
  21397=>"011010000",
  21398=>"000000000",
  21399=>"000000000",
  21400=>"000111011",
  21401=>"111000100",
  21402=>"000000001",
  21403=>"000000000",
  21404=>"000000000",
  21405=>"011000000",
  21406=>"111110110",
  21407=>"110111111",
  21408=>"111000001",
  21409=>"000000011",
  21410=>"011111110",
  21411=>"000000011",
  21412=>"000110000",
  21413=>"000000000",
  21414=>"100000011",
  21415=>"111011001",
  21416=>"000000000",
  21417=>"001111111",
  21418=>"111111000",
  21419=>"111111010",
  21420=>"111111111",
  21421=>"110111100",
  21422=>"000000111",
  21423=>"100111111",
  21424=>"011011111",
  21425=>"000000000",
  21426=>"101111011",
  21427=>"000000111",
  21428=>"110101001",
  21429=>"001001000",
  21430=>"111111110",
  21431=>"111111111",
  21432=>"000010110",
  21433=>"111001000",
  21434=>"000000000",
  21435=>"100111110",
  21436=>"111111111",
  21437=>"111111111",
  21438=>"000110000",
  21439=>"011111111",
  21440=>"000010000",
  21441=>"111111011",
  21442=>"111000000",
  21443=>"000011111",
  21444=>"000000010",
  21445=>"000100100",
  21446=>"000100110",
  21447=>"111111111",
  21448=>"101101111",
  21449=>"000100100",
  21450=>"000011000",
  21451=>"111011010",
  21452=>"000000111",
  21453=>"000110010",
  21454=>"000000000",
  21455=>"111101000",
  21456=>"000000010",
  21457=>"110111111",
  21458=>"000000001",
  21459=>"000100111",
  21460=>"110110000",
  21461=>"000001001",
  21462=>"100000000",
  21463=>"000000000",
  21464=>"001111001",
  21465=>"000001000",
  21466=>"100000000",
  21467=>"000010000",
  21468=>"001101111",
  21469=>"000000000",
  21470=>"111111111",
  21471=>"000001011",
  21472=>"000000100",
  21473=>"100111111",
  21474=>"000000111",
  21475=>"000000000",
  21476=>"000110110",
  21477=>"000000000",
  21478=>"001010010",
  21479=>"000000111",
  21480=>"011111110",
  21481=>"111001111",
  21482=>"111110000",
  21483=>"111011110",
  21484=>"111001000",
  21485=>"000000000",
  21486=>"100100111",
  21487=>"000000000",
  21488=>"100000111",
  21489=>"111100000",
  21490=>"000011010",
  21491=>"000011111",
  21492=>"101111010",
  21493=>"111000000",
  21494=>"000010111",
  21495=>"000000000",
  21496=>"100100110",
  21497=>"110110010",
  21498=>"111111111",
  21499=>"000000000",
  21500=>"110111110",
  21501=>"011111111",
  21502=>"000110110",
  21503=>"010000110",
  21504=>"010010000",
  21505=>"010000000",
  21506=>"100000000",
  21507=>"000000000",
  21508=>"110000100",
  21509=>"101000000",
  21510=>"000000000",
  21511=>"111111111",
  21512=>"000011111",
  21513=>"111111001",
  21514=>"111111111",
  21515=>"000000001",
  21516=>"111111111",
  21517=>"011101111",
  21518=>"011001000",
  21519=>"000000000",
  21520=>"111111111",
  21521=>"000000000",
  21522=>"001000000",
  21523=>"000011110",
  21524=>"111110110",
  21525=>"000000110",
  21526=>"000100111",
  21527=>"000000000",
  21528=>"111110110",
  21529=>"000001001",
  21530=>"101101000",
  21531=>"011011011",
  21532=>"111111111",
  21533=>"111111111",
  21534=>"111010100",
  21535=>"000000000",
  21536=>"011011000",
  21537=>"111111111",
  21538=>"110110110",
  21539=>"100100010",
  21540=>"111000001",
  21541=>"000010110",
  21542=>"000000000",
  21543=>"110111001",
  21544=>"000000000",
  21545=>"100000000",
  21546=>"110110111",
  21547=>"111111001",
  21548=>"111111111",
  21549=>"100001001",
  21550=>"111011010",
  21551=>"011111110",
  21552=>"111110000",
  21553=>"111110100",
  21554=>"010000001",
  21555=>"111111111",
  21556=>"011000000",
  21557=>"101000000",
  21558=>"000000000",
  21559=>"000000000",
  21560=>"000000001",
  21561=>"000100000",
  21562=>"000000000",
  21563=>"111000000",
  21564=>"101111111",
  21565=>"011010101",
  21566=>"110000000",
  21567=>"011011011",
  21568=>"000010001",
  21569=>"111111111",
  21570=>"000000001",
  21571=>"000010000",
  21572=>"000100000",
  21573=>"000011011",
  21574=>"110000000",
  21575=>"111111111",
  21576=>"100100000",
  21577=>"000100110",
  21578=>"000111000",
  21579=>"010011001",
  21580=>"000000001",
  21581=>"010111000",
  21582=>"111111111",
  21583=>"000111000",
  21584=>"000000000",
  21585=>"000000000",
  21586=>"000000100",
  21587=>"100100000",
  21588=>"001001011",
  21589=>"000011111",
  21590=>"000100100",
  21591=>"000000000",
  21592=>"000000000",
  21593=>"111000000",
  21594=>"000110011",
  21595=>"000011011",
  21596=>"100000000",
  21597=>"111111110",
  21598=>"000001011",
  21599=>"001111000",
  21600=>"111111111",
  21601=>"001000000",
  21602=>"000100000",
  21603=>"000000011",
  21604=>"111101111",
  21605=>"110100110",
  21606=>"100111111",
  21607=>"111100000",
  21608=>"011111111",
  21609=>"000000000",
  21610=>"000000000",
  21611=>"001011111",
  21612=>"000000010",
  21613=>"000000010",
  21614=>"011111111",
  21615=>"000000100",
  21616=>"000000100",
  21617=>"111111111",
  21618=>"111111101",
  21619=>"111111111",
  21620=>"100000011",
  21621=>"111100100",
  21622=>"000000100",
  21623=>"001000000",
  21624=>"111001000",
  21625=>"000000000",
  21626=>"111111111",
  21627=>"111111111",
  21628=>"001011111",
  21629=>"111111111",
  21630=>"111111111",
  21631=>"000000110",
  21632=>"000000000",
  21633=>"000011001",
  21634=>"111010000",
  21635=>"111111100",
  21636=>"111111010",
  21637=>"111111111",
  21638=>"110111111",
  21639=>"000110111",
  21640=>"000000000",
  21641=>"001111000",
  21642=>"011111111",
  21643=>"011011110",
  21644=>"000100111",
  21645=>"000000000",
  21646=>"011001011",
  21647=>"101110110",
  21648=>"111101000",
  21649=>"111111111",
  21650=>"000000000",
  21651=>"011001000",
  21652=>"001111000",
  21653=>"111111111",
  21654=>"000011010",
  21655=>"110111111",
  21656=>"000000010",
  21657=>"111110111",
  21658=>"000000000",
  21659=>"000000000",
  21660=>"000000000",
  21661=>"111000000",
  21662=>"000000000",
  21663=>"010000000",
  21664=>"000000000",
  21665=>"001000000",
  21666=>"000000000",
  21667=>"000000000",
  21668=>"111111110",
  21669=>"010111110",
  21670=>"111111111",
  21671=>"101100100",
  21672=>"111111011",
  21673=>"111001000",
  21674=>"000000000",
  21675=>"111001001",
  21676=>"111101111",
  21677=>"110010000",
  21678=>"000000010",
  21679=>"111111000",
  21680=>"000110000",
  21681=>"000000000",
  21682=>"001101001",
  21683=>"011000000",
  21684=>"010000111",
  21685=>"111110000",
  21686=>"111111001",
  21687=>"000000111",
  21688=>"111000010",
  21689=>"000000000",
  21690=>"000001111",
  21691=>"000111111",
  21692=>"001111111",
  21693=>"000110111",
  21694=>"111010010",
  21695=>"000000000",
  21696=>"111100000",
  21697=>"111111000",
  21698=>"000000111",
  21699=>"111111111",
  21700=>"111111000",
  21701=>"111111111",
  21702=>"111111101",
  21703=>"000001001",
  21704=>"110000000",
  21705=>"111101111",
  21706=>"001111111",
  21707=>"000111111",
  21708=>"111111000",
  21709=>"110100000",
  21710=>"110111010",
  21711=>"111111111",
  21712=>"000110100",
  21713=>"100000001",
  21714=>"011011000",
  21715=>"110000111",
  21716=>"011111111",
  21717=>"000000000",
  21718=>"111110110",
  21719=>"001000000",
  21720=>"111111111",
  21721=>"000000001",
  21722=>"111111111",
  21723=>"111111110",
  21724=>"111111111",
  21725=>"000011111",
  21726=>"000001011",
  21727=>"111110111",
  21728=>"111111111",
  21729=>"110111000",
  21730=>"000000000",
  21731=>"010110010",
  21732=>"101101111",
  21733=>"000000000",
  21734=>"011000011",
  21735=>"111110010",
  21736=>"111111111",
  21737=>"000000010",
  21738=>"110110111",
  21739=>"011010010",
  21740=>"000111111",
  21741=>"001000100",
  21742=>"111111001",
  21743=>"000000000",
  21744=>"000000000",
  21745=>"010000011",
  21746=>"111111001",
  21747=>"000110000",
  21748=>"111111111",
  21749=>"010110010",
  21750=>"111111111",
  21751=>"000001011",
  21752=>"000110111",
  21753=>"111111011",
  21754=>"110111111",
  21755=>"000100110",
  21756=>"111001001",
  21757=>"111111111",
  21758=>"110100000",
  21759=>"100100100",
  21760=>"000000010",
  21761=>"101100101",
  21762=>"000011001",
  21763=>"111111111",
  21764=>"000111111",
  21765=>"111111111",
  21766=>"011011011",
  21767=>"000111000",
  21768=>"111110000",
  21769=>"000000000",
  21770=>"000000000",
  21771=>"011111111",
  21772=>"111001111",
  21773=>"100111111",
  21774=>"010010000",
  21775=>"011011111",
  21776=>"111111000",
  21777=>"000000000",
  21778=>"101101100",
  21779=>"000011111",
  21780=>"000000000",
  21781=>"000000111",
  21782=>"111110010",
  21783=>"000000000",
  21784=>"000000000",
  21785=>"000100111",
  21786=>"000000000",
  21787=>"000111101",
  21788=>"000000100",
  21789=>"111111111",
  21790=>"010000110",
  21791=>"111111100",
  21792=>"011001100",
  21793=>"100100001",
  21794=>"111111111",
  21795=>"000000110",
  21796=>"111100110",
  21797=>"000000000",
  21798=>"011111111",
  21799=>"000000000",
  21800=>"110110000",
  21801=>"000000100",
  21802=>"000000000",
  21803=>"100111100",
  21804=>"111111000",
  21805=>"000000000",
  21806=>"000011111",
  21807=>"111111011",
  21808=>"111111011",
  21809=>"100000000",
  21810=>"011001000",
  21811=>"000000100",
  21812=>"000011011",
  21813=>"111111111",
  21814=>"010010011",
  21815=>"111111100",
  21816=>"010111000",
  21817=>"000000111",
  21818=>"101101111",
  21819=>"000011110",
  21820=>"010110111",
  21821=>"010010101",
  21822=>"000110111",
  21823=>"100100111",
  21824=>"100110000",
  21825=>"000101111",
  21826=>"000110000",
  21827=>"000000000",
  21828=>"110111011",
  21829=>"010000000",
  21830=>"000000000",
  21831=>"111111111",
  21832=>"111111111",
  21833=>"000110110",
  21834=>"011111110",
  21835=>"111110010",
  21836=>"001000000",
  21837=>"000000100",
  21838=>"000000001",
  21839=>"011011111",
  21840=>"000010011",
  21841=>"101111111",
  21842=>"100000000",
  21843=>"111111000",
  21844=>"101101111",
  21845=>"010000010",
  21846=>"010000000",
  21847=>"000000000",
  21848=>"111100000",
  21849=>"001111111",
  21850=>"000000101",
  21851=>"000000010",
  21852=>"111111000",
  21853=>"000000100",
  21854=>"111011001",
  21855=>"010110110",
  21856=>"000011111",
  21857=>"000000000",
  21858=>"111001001",
  21859=>"101100000",
  21860=>"000100000",
  21861=>"100111111",
  21862=>"100000000",
  21863=>"110111011",
  21864=>"011111110",
  21865=>"111111010",
  21866=>"111111101",
  21867=>"000001001",
  21868=>"100100100",
  21869=>"001111111",
  21870=>"110111111",
  21871=>"000000000",
  21872=>"000001111",
  21873=>"111001000",
  21874=>"000000000",
  21875=>"000111111",
  21876=>"001001101",
  21877=>"010000000",
  21878=>"000000111",
  21879=>"000000000",
  21880=>"111111111",
  21881=>"001001000",
  21882=>"110111111",
  21883=>"110110100",
  21884=>"001101100",
  21885=>"111110011",
  21886=>"111111000",
  21887=>"111111111",
  21888=>"000000000",
  21889=>"000000011",
  21890=>"000000000",
  21891=>"111011011",
  21892=>"111001001",
  21893=>"000000000",
  21894=>"000000000",
  21895=>"110110111",
  21896=>"111111111",
  21897=>"000000000",
  21898=>"000001001",
  21899=>"000111000",
  21900=>"110000000",
  21901=>"001001001",
  21902=>"100000000",
  21903=>"010111011",
  21904=>"111111000",
  21905=>"010000000",
  21906=>"111001111",
  21907=>"101001111",
  21908=>"100111111",
  21909=>"000000000",
  21910=>"111111111",
  21911=>"111111101",
  21912=>"111111111",
  21913=>"000000100",
  21914=>"111111111",
  21915=>"111111111",
  21916=>"001011111",
  21917=>"011111111",
  21918=>"000000000",
  21919=>"111111111",
  21920=>"011111111",
  21921=>"101111111",
  21922=>"000000101",
  21923=>"111111111",
  21924=>"011000000",
  21925=>"111110111",
  21926=>"110110111",
  21927=>"100111111",
  21928=>"000000000",
  21929=>"110011010",
  21930=>"000100111",
  21931=>"010110100",
  21932=>"111111000",
  21933=>"111111111",
  21934=>"000000000",
  21935=>"111111011",
  21936=>"000000000",
  21937=>"100100100",
  21938=>"000110110",
  21939=>"110111111",
  21940=>"110000000",
  21941=>"111111110",
  21942=>"001000100",
  21943=>"111000000",
  21944=>"111111100",
  21945=>"000000110",
  21946=>"111111100",
  21947=>"000000000",
  21948=>"111110110",
  21949=>"111100000",
  21950=>"000000000",
  21951=>"011011001",
  21952=>"011000000",
  21953=>"111111111",
  21954=>"000110011",
  21955=>"000000000",
  21956=>"110110111",
  21957=>"011011001",
  21958=>"100111010",
  21959=>"110100111",
  21960=>"111110111",
  21961=>"010010000",
  21962=>"011111111",
  21963=>"111011111",
  21964=>"111101111",
  21965=>"000000000",
  21966=>"110110110",
  21967=>"111111111",
  21968=>"000000000",
  21969=>"001011111",
  21970=>"100100110",
  21971=>"001000000",
  21972=>"011000000",
  21973=>"111111111",
  21974=>"001001001",
  21975=>"100100110",
  21976=>"111111111",
  21977=>"111011001",
  21978=>"000111111",
  21979=>"000000110",
  21980=>"111111111",
  21981=>"000011001",
  21982=>"000000011",
  21983=>"100110110",
  21984=>"111011110",
  21985=>"000100000",
  21986=>"100100100",
  21987=>"000000001",
  21988=>"000000100",
  21989=>"111110010",
  21990=>"100111111",
  21991=>"000000000",
  21992=>"000000111",
  21993=>"010010000",
  21994=>"001011111",
  21995=>"111111111",
  21996=>"011011000",
  21997=>"110111110",
  21998=>"000001111",
  21999=>"011111001",
  22000=>"011111111",
  22001=>"000000111",
  22002=>"111111011",
  22003=>"110011111",
  22004=>"011100000",
  22005=>"000000100",
  22006=>"100100111",
  22007=>"000000000",
  22008=>"111011011",
  22009=>"111100001",
  22010=>"010110110",
  22011=>"000000001",
  22012=>"110000101",
  22013=>"111111110",
  22014=>"111111111",
  22015=>"111111111",
  22016=>"000000011",
  22017=>"000100110",
  22018=>"000000000",
  22019=>"111110111",
  22020=>"111000000",
  22021=>"111111001",
  22022=>"111111111",
  22023=>"100110111",
  22024=>"000101101",
  22025=>"000001000",
  22026=>"000000000",
  22027=>"111111111",
  22028=>"001001111",
  22029=>"000110111",
  22030=>"111111011",
  22031=>"111000000",
  22032=>"011000001",
  22033=>"011000000",
  22034=>"000100001",
  22035=>"110111111",
  22036=>"111111001",
  22037=>"000000111",
  22038=>"000000100",
  22039=>"011011001",
  22040=>"000000111",
  22041=>"100111101",
  22042=>"000010111",
  22043=>"000111001",
  22044=>"111001000",
  22045=>"111000000",
  22046=>"000100111",
  22047=>"000111111",
  22048=>"111111111",
  22049=>"100111000",
  22050=>"000000001",
  22051=>"111111111",
  22052=>"110111111",
  22053=>"011010010",
  22054=>"000100111",
  22055=>"111000000",
  22056=>"000111111",
  22057=>"111111111",
  22058=>"110000000",
  22059=>"111000000",
  22060=>"111011000",
  22061=>"111111100",
  22062=>"110111111",
  22063=>"111000100",
  22064=>"111110111",
  22065=>"111111111",
  22066=>"111000000",
  22067=>"000000000",
  22068=>"100001000",
  22069=>"111111111",
  22070=>"001000001",
  22071=>"111010000",
  22072=>"110000100",
  22073=>"111000000",
  22074=>"000000000",
  22075=>"111110110",
  22076=>"000000000",
  22077=>"000000000",
  22078=>"000000000",
  22079=>"000100001",
  22080=>"111111000",
  22081=>"111011000",
  22082=>"111111111",
  22083=>"000000110",
  22084=>"011001000",
  22085=>"110100000",
  22086=>"110111000",
  22087=>"111010000",
  22088=>"111101111",
  22089=>"111100100",
  22090=>"100100000",
  22091=>"111011101",
  22092=>"000000000",
  22093=>"000000001",
  22094=>"101000000",
  22095=>"111111001",
  22096=>"110000000",
  22097=>"100100100",
  22098=>"110100000",
  22099=>"100101111",
  22100=>"000000000",
  22101=>"011111111",
  22102=>"111000000",
  22103=>"111111000",
  22104=>"000000001",
  22105=>"111111100",
  22106=>"111000000",
  22107=>"000000111",
  22108=>"111110000",
  22109=>"010000000",
  22110=>"011001101",
  22111=>"000000111",
  22112=>"000100000",
  22113=>"111111111",
  22114=>"111110000",
  22115=>"000000110",
  22116=>"000101111",
  22117=>"110111111",
  22118=>"011010010",
  22119=>"000111011",
  22120=>"000111000",
  22121=>"000100100",
  22122=>"110000000",
  22123=>"000000111",
  22124=>"000101100",
  22125=>"010100000",
  22126=>"111001001",
  22127=>"001001011",
  22128=>"111100100",
  22129=>"000100110",
  22130=>"100001000",
  22131=>"111111011",
  22132=>"001010000",
  22133=>"100111111",
  22134=>"111111011",
  22135=>"000000000",
  22136=>"000000011",
  22137=>"100101001",
  22138=>"000000000",
  22139=>"000011000",
  22140=>"000000110",
  22141=>"000000000",
  22142=>"000110100",
  22143=>"010000000",
  22144=>"000000111",
  22145=>"000110111",
  22146=>"110111100",
  22147=>"111011111",
  22148=>"000111101",
  22149=>"101100100",
  22150=>"000000000",
  22151=>"111010000",
  22152=>"111111111",
  22153=>"111111100",
  22154=>"110000000",
  22155=>"001111111",
  22156=>"111000001",
  22157=>"000000000",
  22158=>"000000110",
  22159=>"011111000",
  22160=>"110100000",
  22161=>"111101011",
  22162=>"010110100",
  22163=>"110110000",
  22164=>"000110111",
  22165=>"000000111",
  22166=>"011111111",
  22167=>"111000000",
  22168=>"111111111",
  22169=>"100000000",
  22170=>"000010010",
  22171=>"000111111",
  22172=>"000000001",
  22173=>"111111111",
  22174=>"100111111",
  22175=>"000000000",
  22176=>"001010100",
  22177=>"000000000",
  22178=>"000000111",
  22179=>"000000101",
  22180=>"010000000",
  22181=>"100000101",
  22182=>"110111111",
  22183=>"010111111",
  22184=>"111011000",
  22185=>"000100111",
  22186=>"011000000",
  22187=>"000000111",
  22188=>"111010110",
  22189=>"110110111",
  22190=>"111000000",
  22191=>"000100111",
  22192=>"110111001",
  22193=>"000110111",
  22194=>"110000010",
  22195=>"111111100",
  22196=>"000000011",
  22197=>"100100001",
  22198=>"111111111",
  22199=>"111100000",
  22200=>"000000010",
  22201=>"000100110",
  22202=>"010011000",
  22203=>"111101101",
  22204=>"011011000",
  22205=>"110110111",
  22206=>"101000111",
  22207=>"111010001",
  22208=>"110110100",
  22209=>"000000000",
  22210=>"111000000",
  22211=>"011111111",
  22212=>"000000000",
  22213=>"111111000",
  22214=>"000000000",
  22215=>"110100100",
  22216=>"000001000",
  22217=>"000000000",
  22218=>"001100101",
  22219=>"100000000",
  22220=>"100100111",
  22221=>"101111110",
  22222=>"111000000",
  22223=>"111000000",
  22224=>"110000011",
  22225=>"000011111",
  22226=>"111111100",
  22227=>"011100000",
  22228=>"111111010",
  22229=>"100100111",
  22230=>"011111000",
  22231=>"000000000",
  22232=>"100000000",
  22233=>"000101111",
  22234=>"000000000",
  22235=>"000000101",
  22236=>"111111011",
  22237=>"110111111",
  22238=>"111111000",
  22239=>"111110000",
  22240=>"111001000",
  22241=>"111011111",
  22242=>"011001010",
  22243=>"001000000",
  22244=>"111111111",
  22245=>"000000111",
  22246=>"100100111",
  22247=>"110110100",
  22248=>"111111111",
  22249=>"111101111",
  22250=>"000000000",
  22251=>"000111110",
  22252=>"111111101",
  22253=>"111011000",
  22254=>"000000100",
  22255=>"000000100",
  22256=>"111011110",
  22257=>"000100111",
  22258=>"000111111",
  22259=>"011011011",
  22260=>"111110101",
  22261=>"111110000",
  22262=>"100010111",
  22263=>"111111010",
  22264=>"100100111",
  22265=>"111111111",
  22266=>"101111011",
  22267=>"110110110",
  22268=>"001011011",
  22269=>"110100111",
  22270=>"111110000",
  22271=>"011110000",
  22272=>"001011011",
  22273=>"011010010",
  22274=>"111111000",
  22275=>"111111111",
  22276=>"111000000",
  22277=>"111100000",
  22278=>"000000000",
  22279=>"111000000",
  22280=>"001011110",
  22281=>"100111111",
  22282=>"001000111",
  22283=>"111000000",
  22284=>"100110110",
  22285=>"111011000",
  22286=>"110011111",
  22287=>"111111110",
  22288=>"011011011",
  22289=>"111111001",
  22290=>"000000000",
  22291=>"110100101",
  22292=>"000100111",
  22293=>"111011000",
  22294=>"000100110",
  22295=>"000101101",
  22296=>"000000000",
  22297=>"011000001",
  22298=>"111111111",
  22299=>"111000000",
  22300=>"111111111",
  22301=>"111111111",
  22302=>"111111000",
  22303=>"011000101",
  22304=>"000001111",
  22305=>"000100000",
  22306=>"000111110",
  22307=>"100100111",
  22308=>"011011011",
  22309=>"111110110",
  22310=>"100111010",
  22311=>"011000000",
  22312=>"010111011",
  22313=>"111011000",
  22314=>"110100111",
  22315=>"001000000",
  22316=>"101111111",
  22317=>"101100000",
  22318=>"111111010",
  22319=>"000000000",
  22320=>"111111111",
  22321=>"001011111",
  22322=>"000111111",
  22323=>"100110111",
  22324=>"110110100",
  22325=>"011000011",
  22326=>"000000000",
  22327=>"111100000",
  22328=>"000000111",
  22329=>"000000000",
  22330=>"000000000",
  22331=>"000000000",
  22332=>"110110000",
  22333=>"000010111",
  22334=>"011111011",
  22335=>"111000100",
  22336=>"111100100",
  22337=>"000111111",
  22338=>"101000000",
  22339=>"000100100",
  22340=>"110110110",
  22341=>"011111111",
  22342=>"011011000",
  22343=>"001000111",
  22344=>"010010000",
  22345=>"011111000",
  22346=>"111000000",
  22347=>"111001000",
  22348=>"110111111",
  22349=>"111111111",
  22350=>"000000100",
  22351=>"001001011",
  22352=>"001000000",
  22353=>"010100000",
  22354=>"111110111",
  22355=>"001111001",
  22356=>"000000000",
  22357=>"000000011",
  22358=>"111111000",
  22359=>"000000100",
  22360=>"000000000",
  22361=>"101111000",
  22362=>"110111111",
  22363=>"110000000",
  22364=>"000000101",
  22365=>"111000000",
  22366=>"011111000",
  22367=>"111111101",
  22368=>"000110111",
  22369=>"100100111",
  22370=>"000001111",
  22371=>"111111111",
  22372=>"000000000",
  22373=>"111011011",
  22374=>"111111000",
  22375=>"000000011",
  22376=>"110100000",
  22377=>"000111111",
  22378=>"111111110",
  22379=>"110110000",
  22380=>"101001111",
  22381=>"100000000",
  22382=>"001000000",
  22383=>"111111000",
  22384=>"111111000",
  22385=>"111110110",
  22386=>"100000111",
  22387=>"000110000",
  22388=>"111000000",
  22389=>"111100100",
  22390=>"000000100",
  22391=>"110111111",
  22392=>"111111111",
  22393=>"011001000",
  22394=>"001000000",
  22395=>"111000000",
  22396=>"111111001",
  22397=>"100111110",
  22398=>"001111110",
  22399=>"111111111",
  22400=>"111100111",
  22401=>"100100100",
  22402=>"111111111",
  22403=>"111111111",
  22404=>"000011011",
  22405=>"100110100",
  22406=>"000000110",
  22407=>"000000000",
  22408=>"000000000",
  22409=>"001111111",
  22410=>"000110100",
  22411=>"100100110",
  22412=>"100110110",
  22413=>"100100100",
  22414=>"000000000",
  22415=>"111110110",
  22416=>"000111111",
  22417=>"111111111",
  22418=>"000111111",
  22419=>"111011000",
  22420=>"111111111",
  22421=>"111111000",
  22422=>"111111111",
  22423=>"110000111",
  22424=>"100110001",
  22425=>"000110111",
  22426=>"110110110",
  22427=>"000011111",
  22428=>"000000000",
  22429=>"000111000",
  22430=>"011010000",
  22431=>"111111000",
  22432=>"011000000",
  22433=>"010110111",
  22434=>"000000000",
  22435=>"011000000",
  22436=>"000110110",
  22437=>"000000000",
  22438=>"111111000",
  22439=>"111011111",
  22440=>"000000000",
  22441=>"110010011",
  22442=>"000000000",
  22443=>"011011011",
  22444=>"011001000",
  22445=>"000110000",
  22446=>"111110000",
  22447=>"000000000",
  22448=>"111000000",
  22449=>"000000000",
  22450=>"000000000",
  22451=>"111000000",
  22452=>"000000000",
  22453=>"000000000",
  22454=>"100100000",
  22455=>"111000001",
  22456=>"000000000",
  22457=>"111111000",
  22458=>"011000000",
  22459=>"111000111",
  22460=>"111100111",
  22461=>"100100000",
  22462=>"100100000",
  22463=>"110110011",
  22464=>"000000011",
  22465=>"111111111",
  22466=>"000100111",
  22467=>"111000000",
  22468=>"111000000",
  22469=>"001111000",
  22470=>"111100000",
  22471=>"111111000",
  22472=>"000000001",
  22473=>"000000000",
  22474=>"110111000",
  22475=>"000000000",
  22476=>"000010111",
  22477=>"000111000",
  22478=>"100000000",
  22479=>"111110000",
  22480=>"100100100",
  22481=>"001110111",
  22482=>"111111111",
  22483=>"111011111",
  22484=>"000001000",
  22485=>"111100000",
  22486=>"000000000",
  22487=>"111010011",
  22488=>"111110111",
  22489=>"111001001",
  22490=>"111010001",
  22491=>"000000110",
  22492=>"001011011",
  22493=>"100111111",
  22494=>"000000111",
  22495=>"011010000",
  22496=>"000100110",
  22497=>"000110111",
  22498=>"110000000",
  22499=>"000000000",
  22500=>"111110110",
  22501=>"000001000",
  22502=>"100000111",
  22503=>"111111011",
  22504=>"111001000",
  22505=>"010010100",
  22506=>"000011011",
  22507=>"111000101",
  22508=>"100000011",
  22509=>"001000000",
  22510=>"101111111",
  22511=>"111111111",
  22512=>"011000000",
  22513=>"111111000",
  22514=>"011011111",
  22515=>"101100000",
  22516=>"000011001",
  22517=>"111000101",
  22518=>"000010011",
  22519=>"000111111",
  22520=>"100101000",
  22521=>"001000000",
  22522=>"010010011",
  22523=>"111111000",
  22524=>"100111111",
  22525=>"000010010",
  22526=>"111100000",
  22527=>"101001000",
  22528=>"001001001",
  22529=>"011111101",
  22530=>"000000000",
  22531=>"000111111",
  22532=>"111111100",
  22533=>"000111011",
  22534=>"100000000",
  22535=>"111101111",
  22536=>"111000000",
  22537=>"111010000",
  22538=>"111111111",
  22539=>"000011111",
  22540=>"000110110",
  22541=>"111100000",
  22542=>"100001011",
  22543=>"111111111",
  22544=>"000001101",
  22545=>"110110111",
  22546=>"000100100",
  22547=>"000010011",
  22548=>"010011011",
  22549=>"000000000",
  22550=>"111111110",
  22551=>"000001011",
  22552=>"000000000",
  22553=>"100111111",
  22554=>"000100111",
  22555=>"111111110",
  22556=>"111001000",
  22557=>"101111111",
  22558=>"111011111",
  22559=>"110000000",
  22560=>"111000000",
  22561=>"000000000",
  22562=>"000000100",
  22563=>"101000000",
  22564=>"000010111",
  22565=>"111001000",
  22566=>"111000000",
  22567=>"110010000",
  22568=>"110110111",
  22569=>"000111111",
  22570=>"000100000",
  22571=>"111111111",
  22572=>"001000000",
  22573=>"111110111",
  22574=>"111111100",
  22575=>"010111111",
  22576=>"111111111",
  22577=>"000001011",
  22578=>"100000001",
  22579=>"101100000",
  22580=>"110100000",
  22581=>"001011110",
  22582=>"100000001",
  22583=>"000000000",
  22584=>"111100100",
  22585=>"101001111",
  22586=>"001011000",
  22587=>"010111111",
  22588=>"000000000",
  22589=>"111111010",
  22590=>"100000100",
  22591=>"111101000",
  22592=>"000111101",
  22593=>"000000001",
  22594=>"000100110",
  22595=>"000000011",
  22596=>"000110110",
  22597=>"000000100",
  22598=>"010010000",
  22599=>"000000000",
  22600=>"111101111",
  22601=>"000111111",
  22602=>"010011111",
  22603=>"101111111",
  22604=>"101111001",
  22605=>"111000111",
  22606=>"000000000",
  22607=>"111111111",
  22608=>"100100000",
  22609=>"111111110",
  22610=>"111111010",
  22611=>"000000110",
  22612=>"000001000",
  22613=>"011111111",
  22614=>"000000100",
  22615=>"111101101",
  22616=>"000000000",
  22617=>"111100111",
  22618=>"101000000",
  22619=>"001000000",
  22620=>"011011000",
  22621=>"000111111",
  22622=>"000111111",
  22623=>"000100011",
  22624=>"000000000",
  22625=>"110111111",
  22626=>"000000100",
  22627=>"011001000",
  22628=>"011111110",
  22629=>"100000000",
  22630=>"110100110",
  22631=>"111100000",
  22632=>"111011111",
  22633=>"111101100",
  22634=>"000000101",
  22635=>"000000111",
  22636=>"111000000",
  22637=>"000000110",
  22638=>"101101111",
  22639=>"000000000",
  22640=>"111111100",
  22641=>"010010111",
  22642=>"011000000",
  22643=>"000000001",
  22644=>"111111000",
  22645=>"000111111",
  22646=>"111101111",
  22647=>"000000100",
  22648=>"111111111",
  22649=>"000110000",
  22650=>"000000001",
  22651=>"000000000",
  22652=>"001000110",
  22653=>"101111011",
  22654=>"000000000",
  22655=>"110111111",
  22656=>"000000000",
  22657=>"000000110",
  22658=>"000000000",
  22659=>"000000010",
  22660=>"001000100",
  22661=>"111000000",
  22662=>"110111111",
  22663=>"110111111",
  22664=>"111110111",
  22665=>"000000111",
  22666=>"111011000",
  22667=>"111011001",
  22668=>"000000000",
  22669=>"111100000",
  22670=>"110000001",
  22671=>"000111101",
  22672=>"111000000",
  22673=>"111101000",
  22674=>"111100100",
  22675=>"000011101",
  22676=>"001001000",
  22677=>"000100111",
  22678=>"000000111",
  22679=>"000000011",
  22680=>"111011010",
  22681=>"110111111",
  22682=>"001000000",
  22683=>"011000000",
  22684=>"000111110",
  22685=>"001001000",
  22686=>"001101001",
  22687=>"111001000",
  22688=>"000110001",
  22689=>"110000000",
  22690=>"000000100",
  22691=>"111111000",
  22692=>"001001011",
  22693=>"110111111",
  22694=>"010010111",
  22695=>"111101101",
  22696=>"110011000",
  22697=>"011100000",
  22698=>"000000100",
  22699=>"111001111",
  22700=>"011101111",
  22701=>"111111100",
  22702=>"000000001",
  22703=>"000111000",
  22704=>"000010000",
  22705=>"111111111",
  22706=>"110111110",
  22707=>"110000000",
  22708=>"111111110",
  22709=>"111111111",
  22710=>"000000111",
  22711=>"000000000",
  22712=>"000000000",
  22713=>"000100000",
  22714=>"101100101",
  22715=>"111110010",
  22716=>"000110110",
  22717=>"111111010",
  22718=>"000100100",
  22719=>"000001111",
  22720=>"000000001",
  22721=>"000000000",
  22722=>"100111001",
  22723=>"000111111",
  22724=>"111111111",
  22725=>"110100100",
  22726=>"000111110",
  22727=>"111101100",
  22728=>"000110111",
  22729=>"000000111",
  22730=>"000000000",
  22731=>"111100000",
  22732=>"000010011",
  22733=>"100111111",
  22734=>"110111111",
  22735=>"100100000",
  22736=>"111111100",
  22737=>"001111011",
  22738=>"100000000",
  22739=>"111000000",
  22740=>"000000111",
  22741=>"100001000",
  22742=>"111010110",
  22743=>"000000000",
  22744=>"001001000",
  22745=>"111111011",
  22746=>"000000000",
  22747=>"111111111",
  22748=>"111001000",
  22749=>"001110111",
  22750=>"011011000",
  22751=>"111101111",
  22752=>"111111011",
  22753=>"011001101",
  22754=>"000000010",
  22755=>"111010010",
  22756=>"001111111",
  22757=>"110000011",
  22758=>"100100101",
  22759=>"111000000",
  22760=>"111111111",
  22761=>"110110111",
  22762=>"001000111",
  22763=>"111111110",
  22764=>"000000101",
  22765=>"010000000",
  22766=>"111010000",
  22767=>"000000000",
  22768=>"000101111",
  22769=>"000000011",
  22770=>"000011111",
  22771=>"111010111",
  22772=>"000000000",
  22773=>"000101100",
  22774=>"000011000",
  22775=>"111010110",
  22776=>"000111111",
  22777=>"100111111",
  22778=>"000111111",
  22779=>"111111111",
  22780=>"000100110",
  22781=>"011000000",
  22782=>"110000000",
  22783=>"111111111",
  22784=>"110011011",
  22785=>"001000100",
  22786=>"111000000",
  22787=>"111111000",
  22788=>"000001000",
  22789=>"000111001",
  22790=>"000000100",
  22791=>"000110111",
  22792=>"111111000",
  22793=>"000010000",
  22794=>"111000000",
  22795=>"000000000",
  22796=>"111111111",
  22797=>"111111101",
  22798=>"000100111",
  22799=>"111111000",
  22800=>"101101111",
  22801=>"011000000",
  22802=>"000000000",
  22803=>"000110101",
  22804=>"111000000",
  22805=>"011100111",
  22806=>"111111011",
  22807=>"000001011",
  22808=>"011001001",
  22809=>"111101110",
  22810=>"111001001",
  22811=>"110100000",
  22812=>"011110110",
  22813=>"111110111",
  22814=>"111000000",
  22815=>"110111101",
  22816=>"111111000",
  22817=>"011111111",
  22818=>"110110010",
  22819=>"000000111",
  22820=>"111101101",
  22821=>"001000001",
  22822=>"111100000",
  22823=>"010000110",
  22824=>"111111111",
  22825=>"001001111",
  22826=>"010111011",
  22827=>"111111111",
  22828=>"000110111",
  22829=>"111111101",
  22830=>"010010000",
  22831=>"100100111",
  22832=>"001001100",
  22833=>"111000000",
  22834=>"000000001",
  22835=>"000000000",
  22836=>"010100110",
  22837=>"011010000",
  22838=>"111100110",
  22839=>"000000000",
  22840=>"000000000",
  22841=>"110111111",
  22842=>"111100110",
  22843=>"011000001",
  22844=>"101000000",
  22845=>"000000000",
  22846=>"101101111",
  22847=>"000101111",
  22848=>"100000001",
  22849=>"110000001",
  22850=>"000000000",
  22851=>"101000000",
  22852=>"110100000",
  22853=>"111100110",
  22854=>"000000001",
  22855=>"101001111",
  22856=>"000000001",
  22857=>"000000000",
  22858=>"000000001",
  22859=>"100101111",
  22860=>"111101111",
  22861=>"000110010",
  22862=>"100000000",
  22863=>"000101111",
  22864=>"001001111",
  22865=>"101111111",
  22866=>"000000000",
  22867=>"000101101",
  22868=>"000000100",
  22869=>"001001001",
  22870=>"111111111",
  22871=>"000011111",
  22872=>"000111111",
  22873=>"011000000",
  22874=>"001111110",
  22875=>"111111110",
  22876=>"000010000",
  22877=>"100000001",
  22878=>"111011000",
  22879=>"000101100",
  22880=>"111010000",
  22881=>"111101000",
  22882=>"111111001",
  22883=>"000100110",
  22884=>"001011110",
  22885=>"101100000",
  22886=>"110000111",
  22887=>"111001010",
  22888=>"011011000",
  22889=>"000110100",
  22890=>"000111011",
  22891=>"101111111",
  22892=>"111000000",
  22893=>"100000000",
  22894=>"000010000",
  22895=>"111001001",
  22896=>"000111111",
  22897=>"111000000",
  22898=>"111111111",
  22899=>"100111011",
  22900=>"110111100",
  22901=>"111001000",
  22902=>"111000010",
  22903=>"110111111",
  22904=>"111111111",
  22905=>"010010011",
  22906=>"000000101",
  22907=>"001000000",
  22908=>"000100001",
  22909=>"111001000",
  22910=>"111000000",
  22911=>"111111111",
  22912=>"000110110",
  22913=>"110100110",
  22914=>"000001111",
  22915=>"111000000",
  22916=>"000011111",
  22917=>"000000000",
  22918=>"001111111",
  22919=>"000011001",
  22920=>"110100000",
  22921=>"100000000",
  22922=>"001000000",
  22923=>"000111111",
  22924=>"111101101",
  22925=>"100100111",
  22926=>"111111111",
  22927=>"110111111",
  22928=>"001000000",
  22929=>"111111111",
  22930=>"000110110",
  22931=>"100100000",
  22932=>"111111111",
  22933=>"111110000",
  22934=>"000000000",
  22935=>"001000000",
  22936=>"001001001",
  22937=>"111100111",
  22938=>"111110010",
  22939=>"000100101",
  22940=>"100111111",
  22941=>"111000000",
  22942=>"111101101",
  22943=>"110110111",
  22944=>"111111111",
  22945=>"001011001",
  22946=>"110000100",
  22947=>"000000000",
  22948=>"000101111",
  22949=>"111111111",
  22950=>"110000000",
  22951=>"111111000",
  22952=>"000000000",
  22953=>"011111111",
  22954=>"011011011",
  22955=>"111000001",
  22956=>"111111111",
  22957=>"011111010",
  22958=>"111100000",
  22959=>"100001011",
  22960=>"000000100",
  22961=>"000000000",
  22962=>"011011001",
  22963=>"011001000",
  22964=>"100000000",
  22965=>"111001100",
  22966=>"000000011",
  22967=>"111000011",
  22968=>"000000000",
  22969=>"111111011",
  22970=>"110110110",
  22971=>"011011001",
  22972=>"101101001",
  22973=>"000111111",
  22974=>"111110110",
  22975=>"101100111",
  22976=>"011011011",
  22977=>"111111111",
  22978=>"111000000",
  22979=>"010000000",
  22980=>"111111111",
  22981=>"110111111",
  22982=>"111111111",
  22983=>"000000000",
  22984=>"101011011",
  22985=>"100111111",
  22986=>"100000001",
  22987=>"110110000",
  22988=>"000000100",
  22989=>"111111100",
  22990=>"111000100",
  22991=>"000000110",
  22992=>"010011000",
  22993=>"111001001",
  22994=>"001011000",
  22995=>"111111101",
  22996=>"100111111",
  22997=>"111111111",
  22998=>"000000000",
  22999=>"000011011",
  23000=>"000000111",
  23001=>"111000101",
  23002=>"101111000",
  23003=>"000000000",
  23004=>"000000001",
  23005=>"111011111",
  23006=>"111111001",
  23007=>"100001111",
  23008=>"110110110",
  23009=>"111111000",
  23010=>"000000000",
  23011=>"111111000",
  23012=>"101111000",
  23013=>"000000101",
  23014=>"010111100",
  23015=>"000000111",
  23016=>"111100100",
  23017=>"100000001",
  23018=>"011111000",
  23019=>"111111111",
  23020=>"000000000",
  23021=>"101000001",
  23022=>"001001001",
  23023=>"111111111",
  23024=>"101100101",
  23025=>"000100111",
  23026=>"000000000",
  23027=>"111010000",
  23028=>"001000100",
  23029=>"010111111",
  23030=>"000000000",
  23031=>"000111100",
  23032=>"000000001",
  23033=>"001111111",
  23034=>"111111111",
  23035=>"000000000",
  23036=>"111110100",
  23037=>"000001000",
  23038=>"000100110",
  23039=>"000000010",
  23040=>"000000000",
  23041=>"111111000",
  23042=>"110000000",
  23043=>"011111111",
  23044=>"001000000",
  23045=>"011011001",
  23046=>"000000000",
  23047=>"100100101",
  23048=>"000000000",
  23049=>"000000000",
  23050=>"011000000",
  23051=>"111111111",
  23052=>"000000000",
  23053=>"110000000",
  23054=>"000000111",
  23055=>"000000000",
  23056=>"110011111",
  23057=>"000000000",
  23058=>"001000111",
  23059=>"101111111",
  23060=>"111111000",
  23061=>"111111111",
  23062=>"111001000",
  23063=>"110111100",
  23064=>"111111011",
  23065=>"001000001",
  23066=>"011000011",
  23067=>"111110000",
  23068=>"011111111",
  23069=>"000000110",
  23070=>"111111101",
  23071=>"100101001",
  23072=>"000001001",
  23073=>"110110110",
  23074=>"000000000",
  23075=>"111101111",
  23076=>"111101011",
  23077=>"000000000",
  23078=>"111111111",
  23079=>"011001000",
  23080=>"000000000",
  23081=>"000000000",
  23082=>"000100101",
  23083=>"111111111",
  23084=>"000000000",
  23085=>"110111111",
  23086=>"001000001",
  23087=>"111111111",
  23088=>"000000000",
  23089=>"000000000",
  23090=>"000000000",
  23091=>"100111111",
  23092=>"111111011",
  23093=>"001011011",
  23094=>"000000011",
  23095=>"001001000",
  23096=>"110000000",
  23097=>"110000000",
  23098=>"001000000",
  23099=>"111111111",
  23100=>"101111111",
  23101=>"000000001",
  23102=>"111100110",
  23103=>"111000100",
  23104=>"000000000",
  23105=>"011010010",
  23106=>"111011000",
  23107=>"111101111",
  23108=>"000000000",
  23109=>"111111111",
  23110=>"111111111",
  23111=>"110110111",
  23112=>"111111110",
  23113=>"000000001",
  23114=>"011111110",
  23115=>"001000001",
  23116=>"111001000",
  23117=>"111111111",
  23118=>"111111111",
  23119=>"111110000",
  23120=>"011011000",
  23121=>"001001000",
  23122=>"111111111",
  23123=>"010000000",
  23124=>"000001000",
  23125=>"000011110",
  23126=>"011010000",
  23127=>"111110000",
  23128=>"111111111",
  23129=>"101000000",
  23130=>"001101111",
  23131=>"000000001",
  23132=>"000000000",
  23133=>"111110111",
  23134=>"000000000",
  23135=>"001000000",
  23136=>"100100000",
  23137=>"111111101",
  23138=>"101000000",
  23139=>"110000000",
  23140=>"111111100",
  23141=>"111111111",
  23142=>"111111111",
  23143=>"100100100",
  23144=>"111111111",
  23145=>"000000000",
  23146=>"000000100",
  23147=>"001011011",
  23148=>"000001111",
  23149=>"111111111",
  23150=>"000001001",
  23151=>"000000000",
  23152=>"000001101",
  23153=>"000000100",
  23154=>"000000000",
  23155=>"111111111",
  23156=>"000000011",
  23157=>"111000000",
  23158=>"000000100",
  23159=>"000000100",
  23160=>"110010000",
  23161=>"011001001",
  23162=>"110000000",
  23163=>"111111111",
  23164=>"111111001",
  23165=>"000000000",
  23166=>"111111110",
  23167=>"000000000",
  23168=>"000000000",
  23169=>"000000001",
  23170=>"100000111",
  23171=>"110000111",
  23172=>"111111101",
  23173=>"000000111",
  23174=>"000010000",
  23175=>"000000000",
  23176=>"111111111",
  23177=>"111111111",
  23178=>"111111010",
  23179=>"111111111",
  23180=>"111111111",
  23181=>"000000000",
  23182=>"101100101",
  23183=>"111111111",
  23184=>"111111111",
  23185=>"000011011",
  23186=>"011010010",
  23187=>"011001101",
  23188=>"010111111",
  23189=>"000000000",
  23190=>"111111111",
  23191=>"000000000",
  23192=>"101001011",
  23193=>"001101111",
  23194=>"000001001",
  23195=>"011011111",
  23196=>"000000111",
  23197=>"000000000",
  23198=>"111111001",
  23199=>"111111111",
  23200=>"111111111",
  23201=>"100111111",
  23202=>"000000111",
  23203=>"111111001",
  23204=>"111111111",
  23205=>"000100111",
  23206=>"010010010",
  23207=>"001100000",
  23208=>"100111111",
  23209=>"000000000",
  23210=>"000000000",
  23211=>"000000000",
  23212=>"101101111",
  23213=>"100100100",
  23214=>"001011111",
  23215=>"000000011",
  23216=>"000100000",
  23217=>"100100110",
  23218=>"010011000",
  23219=>"111001001",
  23220=>"111111011",
  23221=>"111111000",
  23222=>"111110011",
  23223=>"111011000",
  23224=>"011011111",
  23225=>"111111001",
  23226=>"000000000",
  23227=>"101101111",
  23228=>"111111111",
  23229=>"111000110",
  23230=>"000000000",
  23231=>"001000000",
  23232=>"011000000",
  23233=>"111000000",
  23234=>"000010000",
  23235=>"000000111",
  23236=>"000010111",
  23237=>"111110110",
  23238=>"000001000",
  23239=>"011111111",
  23240=>"111111111",
  23241=>"111000100",
  23242=>"111101011",
  23243=>"111111111",
  23244=>"011000000",
  23245=>"000000001",
  23246=>"000000000",
  23247=>"000100000",
  23248=>"001000000",
  23249=>"111111111",
  23250=>"000000000",
  23251=>"000101001",
  23252=>"000000111",
  23253=>"111111011",
  23254=>"000010111",
  23255=>"111111101",
  23256=>"000000100",
  23257=>"000000110",
  23258=>"000000010",
  23259=>"000000011",
  23260=>"111101001",
  23261=>"111111001",
  23262=>"110001000",
  23263=>"111101111",
  23264=>"011011100",
  23265=>"100100111",
  23266=>"000001111",
  23267=>"000001111",
  23268=>"111111111",
  23269=>"000000011",
  23270=>"000110010",
  23271=>"111111111",
  23272=>"000000000",
  23273=>"001001111",
  23274=>"011000000",
  23275=>"000000000",
  23276=>"010110111",
  23277=>"111010110",
  23278=>"111111111",
  23279=>"111111111",
  23280=>"001111111",
  23281=>"000000101",
  23282=>"111000001",
  23283=>"111111011",
  23284=>"101111111",
  23285=>"000000000",
  23286=>"000001111",
  23287=>"111111111",
  23288=>"000000000",
  23289=>"011010000",
  23290=>"000000000",
  23291=>"000010111",
  23292=>"001000111",
  23293=>"111101001",
  23294=>"111011111",
  23295=>"011111111",
  23296=>"011000001",
  23297=>"101111101",
  23298=>"110110110",
  23299=>"000000000",
  23300=>"101101111",
  23301=>"000110110",
  23302=>"000000111",
  23303=>"000000000",
  23304=>"000001011",
  23305=>"111000000",
  23306=>"100100100",
  23307=>"000001111",
  23308=>"000110111",
  23309=>"000000000",
  23310=>"111111111",
  23311=>"011000000",
  23312=>"011111111",
  23313=>"000001011",
  23314=>"111110000",
  23315=>"010110111",
  23316=>"000000000",
  23317=>"101000000",
  23318=>"100110110",
  23319=>"111111100",
  23320=>"110101101",
  23321=>"101111000",
  23322=>"111011011",
  23323=>"000000000",
  23324=>"111111101",
  23325=>"000000000",
  23326=>"111111111",
  23327=>"000000000",
  23328=>"100000000",
  23329=>"111011001",
  23330=>"000111111",
  23331=>"000000000",
  23332=>"001000000",
  23333=>"111111111",
  23334=>"111111111",
  23335=>"000000000",
  23336=>"100100000",
  23337=>"010000000",
  23338=>"110010001",
  23339=>"011001000",
  23340=>"000100000",
  23341=>"111111101",
  23342=>"000111000",
  23343=>"000001000",
  23344=>"111111111",
  23345=>"000000000",
  23346=>"001001001",
  23347=>"110110111",
  23348=>"000000000",
  23349=>"000011011",
  23350=>"111000100",
  23351=>"000111110",
  23352=>"000000000",
  23353=>"000000000",
  23354=>"000000110",
  23355=>"000000000",
  23356=>"011100111",
  23357=>"001100111",
  23358=>"001100100",
  23359=>"111111111",
  23360=>"110111111",
  23361=>"111111100",
  23362=>"000000000",
  23363=>"000000000",
  23364=>"111101110",
  23365=>"000100110",
  23366=>"001000000",
  23367=>"000001000",
  23368=>"110110111",
  23369=>"111111100",
  23370=>"101000001",
  23371=>"111111100",
  23372=>"011110101",
  23373=>"000100110",
  23374=>"100000000",
  23375=>"000110110",
  23376=>"111011011",
  23377=>"000101101",
  23378=>"111000111",
  23379=>"010000000",
  23380=>"000000000",
  23381=>"000000001",
  23382=>"000000110",
  23383=>"000110010",
  23384=>"000000000",
  23385=>"101000010",
  23386=>"111111000",
  23387=>"000000000",
  23388=>"110010111",
  23389=>"111100111",
  23390=>"000101101",
  23391=>"111111111",
  23392=>"000000000",
  23393=>"000000001",
  23394=>"000000000",
  23395=>"111111111",
  23396=>"111111111",
  23397=>"111111111",
  23398=>"000000000",
  23399=>"111111000",
  23400=>"111111101",
  23401=>"000011001",
  23402=>"010111111",
  23403=>"000000101",
  23404=>"111111111",
  23405=>"111111111",
  23406=>"100110111",
  23407=>"111111000",
  23408=>"000000000",
  23409=>"111111011",
  23410=>"001001001",
  23411=>"111111111",
  23412=>"011000000",
  23413=>"000000000",
  23414=>"111111111",
  23415=>"000000000",
  23416=>"100110111",
  23417=>"000000000",
  23418=>"000000001",
  23419=>"101100101",
  23420=>"111110110",
  23421=>"000110111",
  23422=>"010000000",
  23423=>"100100000",
  23424=>"100010111",
  23425=>"001001001",
  23426=>"111111111",
  23427=>"000000000",
  23428=>"111000000",
  23429=>"000000000",
  23430=>"111101111",
  23431=>"111111011",
  23432=>"000000111",
  23433=>"110110110",
  23434=>"111111001",
  23435=>"000000000",
  23436=>"111100111",
  23437=>"111111111",
  23438=>"000101001",
  23439=>"111111111",
  23440=>"010000000",
  23441=>"111011000",
  23442=>"010111111",
  23443=>"000000011",
  23444=>"000000001",
  23445=>"000110000",
  23446=>"111101000",
  23447=>"100000110",
  23448=>"111001111",
  23449=>"001001111",
  23450=>"000000001",
  23451=>"111111111",
  23452=>"001111111",
  23453=>"000000000",
  23454=>"010111111",
  23455=>"000101111",
  23456=>"111111111",
  23457=>"100001001",
  23458=>"111111111",
  23459=>"000010111",
  23460=>"111101101",
  23461=>"111111110",
  23462=>"000000000",
  23463=>"011010000",
  23464=>"111111111",
  23465=>"000000111",
  23466=>"001000000",
  23467=>"010111011",
  23468=>"100000000",
  23469=>"010000000",
  23470=>"001111111",
  23471=>"110110100",
  23472=>"111111111",
  23473=>"000000000",
  23474=>"000000000",
  23475=>"011001111",
  23476=>"000000000",
  23477=>"000000001",
  23478=>"111101111",
  23479=>"111001011",
  23480=>"110001101",
  23481=>"010111111",
  23482=>"000000000",
  23483=>"111111010",
  23484=>"110111111",
  23485=>"010000011",
  23486=>"111111111",
  23487=>"101101101",
  23488=>"001000000",
  23489=>"000000000",
  23490=>"000101111",
  23491=>"111111111",
  23492=>"100000100",
  23493=>"110000100",
  23494=>"111111111",
  23495=>"100111111",
  23496=>"000000011",
  23497=>"000001000",
  23498=>"110111111",
  23499=>"111110100",
  23500=>"011111000",
  23501=>"000000000",
  23502=>"010011011",
  23503=>"111010111",
  23504=>"111111111",
  23505=>"000111111",
  23506=>"010000000",
  23507=>"000000100",
  23508=>"011000000",
  23509=>"110100101",
  23510=>"000111000",
  23511=>"010000000",
  23512=>"000000111",
  23513=>"111111011",
  23514=>"010000000",
  23515=>"000000000",
  23516=>"000000000",
  23517=>"010000010",
  23518=>"100101111",
  23519=>"000100100",
  23520=>"000000000",
  23521=>"111111110",
  23522=>"000000000",
  23523=>"000000001",
  23524=>"111111111",
  23525=>"111011111",
  23526=>"000000100",
  23527=>"000000000",
  23528=>"111111111",
  23529=>"000000011",
  23530=>"011111111",
  23531=>"001001001",
  23532=>"100110110",
  23533=>"000101101",
  23534=>"111011111",
  23535=>"111111111",
  23536=>"000111111",
  23537=>"010000000",
  23538=>"000100100",
  23539=>"000000000",
  23540=>"100000000",
  23541=>"100000111",
  23542=>"111111011",
  23543=>"011011001",
  23544=>"100000000",
  23545=>"110000101",
  23546=>"000000000",
  23547=>"000001001",
  23548=>"100100000",
  23549=>"111100111",
  23550=>"010110111",
  23551=>"111111111",
  23552=>"001100100",
  23553=>"111111000",
  23554=>"000100111",
  23555=>"111111111",
  23556=>"111011010",
  23557=>"010100001",
  23558=>"000000000",
  23559=>"111111111",
  23560=>"111111000",
  23561=>"111011111",
  23562=>"000000000",
  23563=>"111001000",
  23564=>"001001000",
  23565=>"000011111",
  23566=>"000000111",
  23567=>"000000000",
  23568=>"011000000",
  23569=>"111111111",
  23570=>"000000101",
  23571=>"000000000",
  23572=>"000000000",
  23573=>"100000100",
  23574=>"000100000",
  23575=>"111111110",
  23576=>"111111111",
  23577=>"110111111",
  23578=>"011011110",
  23579=>"000000000",
  23580=>"111111111",
  23581=>"001111111",
  23582=>"001011011",
  23583=>"011001000",
  23584=>"001001101",
  23585=>"000110111",
  23586=>"101101000",
  23587=>"011111001",
  23588=>"100110111",
  23589=>"111000000",
  23590=>"000000001",
  23591=>"111111001",
  23592=>"000000100",
  23593=>"100000000",
  23594=>"000000100",
  23595=>"100000000",
  23596=>"111011001",
  23597=>"111111111",
  23598=>"000000001",
  23599=>"010011111",
  23600=>"000001011",
  23601=>"011111010",
  23602=>"111111111",
  23603=>"111011011",
  23604=>"100101111",
  23605=>"111111110",
  23606=>"001111000",
  23607=>"101101111",
  23608=>"000000000",
  23609=>"100110001",
  23610=>"000000000",
  23611=>"111110101",
  23612=>"000100111",
  23613=>"000001001",
  23614=>"000100101",
  23615=>"110100000",
  23616=>"100100111",
  23617=>"001000000",
  23618=>"111111111",
  23619=>"100110111",
  23620=>"100000000",
  23621=>"001001100",
  23622=>"011111000",
  23623=>"000000001",
  23624=>"000001001",
  23625=>"000000000",
  23626=>"000000111",
  23627=>"110011011",
  23628=>"000000011",
  23629=>"111111100",
  23630=>"111000000",
  23631=>"111111011",
  23632=>"100111010",
  23633=>"101001101",
  23634=>"000000000",
  23635=>"101000000",
  23636=>"000110111",
  23637=>"101000000",
  23638=>"000111111",
  23639=>"011111111",
  23640=>"110110000",
  23641=>"000000000",
  23642=>"111110111",
  23643=>"000001111",
  23644=>"000011000",
  23645=>"011000111",
  23646=>"110111001",
  23647=>"111111101",
  23648=>"000110111",
  23649=>"000111000",
  23650=>"111000000",
  23651=>"111111000",
  23652=>"111111111",
  23653=>"001000001",
  23654=>"111111100",
  23655=>"111111111",
  23656=>"000001001",
  23657=>"110111000",
  23658=>"010010000",
  23659=>"110000000",
  23660=>"010111111",
  23661=>"000000000",
  23662=>"001001001",
  23663=>"111101101",
  23664=>"010000000",
  23665=>"111110110",
  23666=>"000000001",
  23667=>"000010000",
  23668=>"000000000",
  23669=>"011000000",
  23670=>"111011100",
  23671=>"001111011",
  23672=>"000000000",
  23673=>"110110100",
  23674=>"001000001",
  23675=>"000100000",
  23676=>"000011110",
  23677=>"001100111",
  23678=>"001000000",
  23679=>"000000000",
  23680=>"000000000",
  23681=>"111111111",
  23682=>"000000000",
  23683=>"000010011",
  23684=>"111111111",
  23685=>"000000000",
  23686=>"111000001",
  23687=>"111101000",
  23688=>"111111111",
  23689=>"111011111",
  23690=>"001001000",
  23691=>"000000000",
  23692=>"110111111",
  23693=>"111111100",
  23694=>"000000001",
  23695=>"111111111",
  23696=>"111101111",
  23697=>"000000000",
  23698=>"110111111",
  23699=>"111110110",
  23700=>"000010010",
  23701=>"111111111",
  23702=>"000000000",
  23703=>"111110100",
  23704=>"001011001",
  23705=>"011110111",
  23706=>"001001110",
  23707=>"100000000",
  23708=>"001000000",
  23709=>"101011110",
  23710=>"000000010",
  23711=>"001001011",
  23712=>"000000111",
  23713=>"111001101",
  23714=>"100000100",
  23715=>"000101000",
  23716=>"011111111",
  23717=>"001111011",
  23718=>"000000000",
  23719=>"011011111",
  23720=>"111000000",
  23721=>"000000000",
  23722=>"000000000",
  23723=>"100100000",
  23724=>"101111111",
  23725=>"101000000",
  23726=>"001000000",
  23727=>"000000101",
  23728=>"000000100",
  23729=>"101001100",
  23730=>"011111111",
  23731=>"111111111",
  23732=>"111110000",
  23733=>"110000000",
  23734=>"001001001",
  23735=>"111001011",
  23736=>"000001100",
  23737=>"111011100",
  23738=>"001000110",
  23739=>"000100000",
  23740=>"111100000",
  23741=>"110110000",
  23742=>"001000000",
  23743=>"000001011",
  23744=>"000000000",
  23745=>"000110000",
  23746=>"000000000",
  23747=>"011111000",
  23748=>"100101111",
  23749=>"000000001",
  23750=>"000000111",
  23751=>"000000000",
  23752=>"000000111",
  23753=>"000000000",
  23754=>"111111010",
  23755=>"111111111",
  23756=>"110111111",
  23757=>"111111111",
  23758=>"111011001",
  23759=>"001011000",
  23760=>"111000000",
  23761=>"111111111",
  23762=>"011000000",
  23763=>"000010111",
  23764=>"111111111",
  23765=>"111111011",
  23766=>"000000000",
  23767=>"111111111",
  23768=>"101100000",
  23769=>"111011011",
  23770=>"000000100",
  23771=>"000000000",
  23772=>"101000000",
  23773=>"111111101",
  23774=>"111111100",
  23775=>"110000000",
  23776=>"000000000",
  23777=>"110111011",
  23778=>"100000000",
  23779=>"111111001",
  23780=>"000000111",
  23781=>"001001000",
  23782=>"000001111",
  23783=>"111111000",
  23784=>"000000000",
  23785=>"111111111",
  23786=>"001111101",
  23787=>"000000000",
  23788=>"000000001",
  23789=>"111111001",
  23790=>"011010100",
  23791=>"101011000",
  23792=>"100100110",
  23793=>"111111111",
  23794=>"100100100",
  23795=>"000100110",
  23796=>"111111111",
  23797=>"111111111",
  23798=>"111100101",
  23799=>"111101101",
  23800=>"111111111",
  23801=>"111110111",
  23802=>"000001011",
  23803=>"111011001",
  23804=>"111110110",
  23805=>"000000100",
  23806=>"110110000",
  23807=>"001111111",
  23808=>"000110111",
  23809=>"111011001",
  23810=>"000000000",
  23811=>"001001000",
  23812=>"000100000",
  23813=>"110110110",
  23814=>"000000111",
  23815=>"000110111",
  23816=>"001000000",
  23817=>"001000000",
  23818=>"000000001",
  23819=>"001001000",
  23820=>"111110100",
  23821=>"000000111",
  23822=>"000000011",
  23823=>"000000111",
  23824=>"111111111",
  23825=>"001101111",
  23826=>"010000000",
  23827=>"000000000",
  23828=>"000000100",
  23829=>"011001000",
  23830=>"111101100",
  23831=>"111111110",
  23832=>"100110011",
  23833=>"111111111",
  23834=>"110111111",
  23835=>"110100000",
  23836=>"000000111",
  23837=>"111101100",
  23838=>"000000000",
  23839=>"001111101",
  23840=>"111111100",
  23841=>"111110011",
  23842=>"111111111",
  23843=>"000000011",
  23844=>"000000000",
  23845=>"000000111",
  23846=>"111111111",
  23847=>"100101111",
  23848=>"000100100",
  23849=>"001001111",
  23850=>"100100000",
  23851=>"100110010",
  23852=>"100110110",
  23853=>"110110101",
  23854=>"000000000",
  23855=>"111111111",
  23856=>"000000000",
  23857=>"111111111",
  23858=>"110110110",
  23859=>"111000000",
  23860=>"000000000",
  23861=>"111101100",
  23862=>"100110000",
  23863=>"001101111",
  23864=>"111000000",
  23865=>"111111011",
  23866=>"111010010",
  23867=>"111111000",
  23868=>"000000100",
  23869=>"000100000",
  23870=>"000001000",
  23871=>"000000000",
  23872=>"000000000",
  23873=>"111111000",
  23874=>"110111000",
  23875=>"111111111",
  23876=>"111111000",
  23877=>"110010000",
  23878=>"011110110",
  23879=>"000000000",
  23880=>"000000000",
  23881=>"000000000",
  23882=>"000000000",
  23883=>"000010111",
  23884=>"001000100",
  23885=>"000000000",
  23886=>"000100011",
  23887=>"110110101",
  23888=>"001001001",
  23889=>"000000000",
  23890=>"000000111",
  23891=>"000000001",
  23892=>"111111111",
  23893=>"000000000",
  23894=>"110110111",
  23895=>"000001000",
  23896=>"111011111",
  23897=>"111100000",
  23898=>"111111111",
  23899=>"000100110",
  23900=>"000101111",
  23901=>"111001111",
  23902=>"111000000",
  23903=>"111011011",
  23904=>"101000000",
  23905=>"000001011",
  23906=>"011011000",
  23907=>"010111000",
  23908=>"111110110",
  23909=>"000000000",
  23910=>"000000000",
  23911=>"001000000",
  23912=>"000000100",
  23913=>"110000000",
  23914=>"011110000",
  23915=>"001001001",
  23916=>"000100000",
  23917=>"000000100",
  23918=>"000000000",
  23919=>"011111010",
  23920=>"111111000",
  23921=>"011011111",
  23922=>"111111111",
  23923=>"110110111",
  23924=>"000000000",
  23925=>"111111100",
  23926=>"111111000",
  23927=>"000010000",
  23928=>"000000000",
  23929=>"111111000",
  23930=>"000000000",
  23931=>"100110110",
  23932=>"010000000",
  23933=>"010010111",
  23934=>"111111100",
  23935=>"111111000",
  23936=>"011010010",
  23937=>"010010011",
  23938=>"111111111",
  23939=>"000000000",
  23940=>"110010000",
  23941=>"110110000",
  23942=>"000000000",
  23943=>"111111000",
  23944=>"110000000",
  23945=>"100110111",
  23946=>"110011001",
  23947=>"111111111",
  23948=>"000000000",
  23949=>"000000100",
  23950=>"110101001",
  23951=>"111111111",
  23952=>"000000000",
  23953=>"111001001",
  23954=>"100000001",
  23955=>"000000010",
  23956=>"110100111",
  23957=>"000000000",
  23958=>"011001000",
  23959=>"100101111",
  23960=>"111111111",
  23961=>"001001001",
  23962=>"100111000",
  23963=>"010100110",
  23964=>"000001011",
  23965=>"000000000",
  23966=>"111111111",
  23967=>"000000000",
  23968=>"001001000",
  23969=>"111000000",
  23970=>"001111111",
  23971=>"000000000",
  23972=>"000000001",
  23973=>"111111111",
  23974=>"011000000",
  23975=>"011111111",
  23976=>"001001001",
  23977=>"111111101",
  23978=>"001000110",
  23979=>"101100100",
  23980=>"111001000",
  23981=>"001100000",
  23982=>"000111111",
  23983=>"001011010",
  23984=>"010000111",
  23985=>"111111111",
  23986=>"000000000",
  23987=>"000000000",
  23988=>"000001101",
  23989=>"111110110",
  23990=>"100111111",
  23991=>"000110110",
  23992=>"110110000",
  23993=>"000000011",
  23994=>"001000000",
  23995=>"101101100",
  23996=>"111111110",
  23997=>"001000000",
  23998=>"111100000",
  23999=>"110100101",
  24000=>"111111011",
  24001=>"000011111",
  24002=>"000000001",
  24003=>"110001001",
  24004=>"111111011",
  24005=>"000000111",
  24006=>"000000001",
  24007=>"110111101",
  24008=>"000110111",
  24009=>"000010011",
  24010=>"000000001",
  24011=>"011001111",
  24012=>"100111000",
  24013=>"000000100",
  24014=>"000000000",
  24015=>"010011111",
  24016=>"111001000",
  24017=>"111101001",
  24018=>"111000001",
  24019=>"110000010",
  24020=>"101100111",
  24021=>"110111111",
  24022=>"000000000",
  24023=>"100001000",
  24024=>"100111001",
  24025=>"000110111",
  24026=>"111111000",
  24027=>"100100100",
  24028=>"111101101",
  24029=>"100110111",
  24030=>"111000000",
  24031=>"111110111",
  24032=>"010111010",
  24033=>"111111111",
  24034=>"011111000",
  24035=>"111101110",
  24036=>"010100110",
  24037=>"111111011",
  24038=>"110100100",
  24039=>"111100000",
  24040=>"111111011",
  24041=>"111111111",
  24042=>"100100100",
  24043=>"001001011",
  24044=>"001100100",
  24045=>"000000010",
  24046=>"100110110",
  24047=>"000000100",
  24048=>"001011111",
  24049=>"011110000",
  24050=>"001001000",
  24051=>"101000101",
  24052=>"111101111",
  24053=>"011000111",
  24054=>"000000001",
  24055=>"110000001",
  24056=>"010000000",
  24057=>"000000111",
  24058=>"000000000",
  24059=>"000000000",
  24060=>"000010111",
  24061=>"000000010",
  24062=>"000000000",
  24063=>"101001111",
  24064=>"111100111",
  24065=>"000110000",
  24066=>"000000100",
  24067=>"000000000",
  24068=>"111011011",
  24069=>"111001000",
  24070=>"111111111",
  24071=>"111000000",
  24072=>"011010111",
  24073=>"111111111",
  24074=>"010111111",
  24075=>"111111110",
  24076=>"100110110",
  24077=>"110000010",
  24078=>"000000100",
  24079=>"000000000",
  24080=>"110111111",
  24081=>"010000011",
  24082=>"111111111",
  24083=>"111000000",
  24084=>"001000000",
  24085=>"111111111",
  24086=>"111001101",
  24087=>"000100100",
  24088=>"110000000",
  24089=>"100000100",
  24090=>"000000001",
  24091=>"100110100",
  24092=>"011001001",
  24093=>"111111001",
  24094=>"010011111",
  24095=>"110010111",
  24096=>"111111111",
  24097=>"000000001",
  24098=>"111000001",
  24099=>"010011001",
  24100=>"011000000",
  24101=>"111011010",
  24102=>"101001001",
  24103=>"111111000",
  24104=>"111111010",
  24105=>"111111111",
  24106=>"001011011",
  24107=>"011000001",
  24108=>"000111111",
  24109=>"111010000",
  24110=>"110010111",
  24111=>"100100000",
  24112=>"000000000",
  24113=>"101000000",
  24114=>"111101100",
  24115=>"011011000",
  24116=>"110000001",
  24117=>"101111101",
  24118=>"111001001",
  24119=>"111000001",
  24120=>"111111111",
  24121=>"000000000",
  24122=>"111111111",
  24123=>"111110110",
  24124=>"101000000",
  24125=>"000000000",
  24126=>"000111111",
  24127=>"000000000",
  24128=>"010010000",
  24129=>"000000000",
  24130=>"000000000",
  24131=>"000000111",
  24132=>"001000001",
  24133=>"110000100",
  24134=>"111110111",
  24135=>"100000000",
  24136=>"001001101",
  24137=>"010111111",
  24138=>"111000000",
  24139=>"000000001",
  24140=>"111001111",
  24141=>"000000111",
  24142=>"000000000",
  24143=>"000000000",
  24144=>"110000100",
  24145=>"000000000",
  24146=>"001000000",
  24147=>"111110100",
  24148=>"000000000",
  24149=>"100100111",
  24150=>"111110000",
  24151=>"000000000",
  24152=>"000000000",
  24153=>"100000101",
  24154=>"111110111",
  24155=>"111111110",
  24156=>"000010000",
  24157=>"000000000",
  24158=>"010010111",
  24159=>"111000000",
  24160=>"111111111",
  24161=>"000110111",
  24162=>"000000000",
  24163=>"000000111",
  24164=>"111110000",
  24165=>"111001000",
  24166=>"111111111",
  24167=>"011000000",
  24168=>"011000011",
  24169=>"111101101",
  24170=>"000000000",
  24171=>"000000000",
  24172=>"110111000",
  24173=>"000000000",
  24174=>"001001111",
  24175=>"111111111",
  24176=>"110000111",
  24177=>"111011001",
  24178=>"110000000",
  24179=>"000000111",
  24180=>"111111111",
  24181=>"000000000",
  24182=>"111111111",
  24183=>"111111111",
  24184=>"111111000",
  24185=>"001001111",
  24186=>"111000000",
  24187=>"111110000",
  24188=>"000001000",
  24189=>"110111110",
  24190=>"111111000",
  24191=>"001000000",
  24192=>"111111111",
  24193=>"000000000",
  24194=>"100111111",
  24195=>"011111110",
  24196=>"101111111",
  24197=>"000000000",
  24198=>"001101111",
  24199=>"111001001",
  24200=>"000010111",
  24201=>"100101000",
  24202=>"001000000",
  24203=>"111111000",
  24204=>"111111000",
  24205=>"000000000",
  24206=>"111111111",
  24207=>"010000000",
  24208=>"000000101",
  24209=>"111110000",
  24210=>"000000001",
  24211=>"000000100",
  24212=>"000000110",
  24213=>"000000001",
  24214=>"010110010",
  24215=>"111001111",
  24216=>"001000100",
  24217=>"111111111",
  24218=>"000000000",
  24219=>"000001111",
  24220=>"000001001",
  24221=>"111111111",
  24222=>"111111100",
  24223=>"110111110",
  24224=>"011111111",
  24225=>"110010000",
  24226=>"111111111",
  24227=>"111111111",
  24228=>"001001000",
  24229=>"111111111",
  24230=>"000110111",
  24231=>"110111100",
  24232=>"000000110",
  24233=>"001001001",
  24234=>"000000001",
  24235=>"001000101",
  24236=>"000000000",
  24237=>"111111100",
  24238=>"111101101",
  24239=>"111000000",
  24240=>"010001111",
  24241=>"001001000",
  24242=>"110111110",
  24243=>"101000000",
  24244=>"000000000",
  24245=>"000000000",
  24246=>"111111110",
  24247=>"010111111",
  24248=>"001000101",
  24249=>"111111111",
  24250=>"111100000",
  24251=>"000000100",
  24252=>"000001001",
  24253=>"000111111",
  24254=>"110110110",
  24255=>"101111101",
  24256=>"000101000",
  24257=>"000000000",
  24258=>"010111111",
  24259=>"000000000",
  24260=>"111110001",
  24261=>"000010000",
  24262=>"000100000",
  24263=>"001001001",
  24264=>"000000000",
  24265=>"000000111",
  24266=>"000000111",
  24267=>"111101000",
  24268=>"111111000",
  24269=>"000000000",
  24270=>"000000001",
  24271=>"000000000",
  24272=>"111111111",
  24273=>"100100111",
  24274=>"100000000",
  24275=>"000100000",
  24276=>"110011111",
  24277=>"001001111",
  24278=>"101101101",
  24279=>"111000001",
  24280=>"000000111",
  24281=>"001001111",
  24282=>"010110111",
  24283=>"111111111",
  24284=>"100000111",
  24285=>"111111111",
  24286=>"000000000",
  24287=>"111111111",
  24288=>"001011111",
  24289=>"010000000",
  24290=>"000110000",
  24291=>"000000111",
  24292=>"000000000",
  24293=>"000110111",
  24294=>"111111111",
  24295=>"010000010",
  24296=>"111000000",
  24297=>"111111111",
  24298=>"000000011",
  24299=>"000000000",
  24300=>"000000000",
  24301=>"111010010",
  24302=>"010010011",
  24303=>"111000000",
  24304=>"011111011",
  24305=>"001101111",
  24306=>"111111110",
  24307=>"001001001",
  24308=>"100000000",
  24309=>"111000000",
  24310=>"000000001",
  24311=>"111111010",
  24312=>"111111010",
  24313=>"000011011",
  24314=>"001000101",
  24315=>"001111111",
  24316=>"000000000",
  24317=>"001001111",
  24318=>"101011111",
  24319=>"000000011",
  24320=>"000100000",
  24321=>"111011001",
  24322=>"111111111",
  24323=>"011111100",
  24324=>"101000101",
  24325=>"000000000",
  24326=>"100000111",
  24327=>"111011000",
  24328=>"111111111",
  24329=>"000000001",
  24330=>"111000000",
  24331=>"000001011",
  24332=>"100100111",
  24333=>"111100000",
  24334=>"111111111",
  24335=>"110111011",
  24336=>"111111000",
  24337=>"110000000",
  24338=>"000000000",
  24339=>"000000001",
  24340=>"000001111",
  24341=>"000011111",
  24342=>"111110110",
  24343=>"011011111",
  24344=>"000000001",
  24345=>"000000000",
  24346=>"111111010",
  24347=>"101000000",
  24348=>"100100000",
  24349=>"000001111",
  24350=>"000111111",
  24351=>"011001111",
  24352=>"000100111",
  24353=>"010010000",
  24354=>"111111111",
  24355=>"111111111",
  24356=>"001001001",
  24357=>"011011111",
  24358=>"111111111",
  24359=>"111100000",
  24360=>"000000111",
  24361=>"000000000",
  24362=>"010011000",
  24363=>"000000000",
  24364=>"000000000",
  24365=>"000000000",
  24366=>"000000000",
  24367=>"101001011",
  24368=>"110110100",
  24369=>"111000000",
  24370=>"111111111",
  24371=>"110100011",
  24372=>"011011010",
  24373=>"111111111",
  24374=>"001111000",
  24375=>"011111111",
  24376=>"111111011",
  24377=>"101101111",
  24378=>"000000101",
  24379=>"110010000",
  24380=>"001001100",
  24381=>"011011111",
  24382=>"000101000",
  24383=>"111101110",
  24384=>"111111111",
  24385=>"111111111",
  24386=>"010110111",
  24387=>"000000101",
  24388=>"001001111",
  24389=>"111111111",
  24390=>"100111111",
  24391=>"111111111",
  24392=>"000000111",
  24393=>"011010011",
  24394=>"000000000",
  24395=>"111000000",
  24396=>"011011111",
  24397=>"000000000",
  24398=>"111111111",
  24399=>"111111011",
  24400=>"011001011",
  24401=>"011001111",
  24402=>"111111111",
  24403=>"000111000",
  24404=>"001011011",
  24405=>"011011011",
  24406=>"000000011",
  24407=>"100110111",
  24408=>"111100111",
  24409=>"111001001",
  24410=>"101000000",
  24411=>"111000101",
  24412=>"000111111",
  24413=>"000000000",
  24414=>"111001000",
  24415=>"110000110",
  24416=>"011111001",
  24417=>"111100111",
  24418=>"101100001",
  24419=>"000000000",
  24420=>"111111111",
  24421=>"001001011",
  24422=>"010111011",
  24423=>"111111110",
  24424=>"100000000",
  24425=>"111111011",
  24426=>"000000000",
  24427=>"000000000",
  24428=>"000000000",
  24429=>"111111110",
  24430=>"000000000",
  24431=>"000000011",
  24432=>"000000101",
  24433=>"111001001",
  24434=>"000011111",
  24435=>"111111000",
  24436=>"000000000",
  24437=>"111111111",
  24438=>"001001111",
  24439=>"000000110",
  24440=>"111001000",
  24441=>"000000001",
  24442=>"101111111",
  24443=>"111101101",
  24444=>"001001001",
  24445=>"111001001",
  24446=>"000011111",
  24447=>"000000000",
  24448=>"000000000",
  24449=>"000000000",
  24450=>"000000001",
  24451=>"000000000",
  24452=>"111001000",
  24453=>"111111110",
  24454=>"000000000",
  24455=>"000000000",
  24456=>"000000000",
  24457=>"011011011",
  24458=>"000000000",
  24459=>"100110000",
  24460=>"001001001",
  24461=>"110110110",
  24462=>"111111000",
  24463=>"111000000",
  24464=>"111111111",
  24465=>"111111111",
  24466=>"000000000",
  24467=>"000000001",
  24468=>"010011000",
  24469=>"000000000",
  24470=>"000000001",
  24471=>"100000000",
  24472=>"000000111",
  24473=>"110000000",
  24474=>"000001111",
  24475=>"111111000",
  24476=>"110110000",
  24477=>"011001011",
  24478=>"101000000",
  24479=>"010010000",
  24480=>"101101111",
  24481=>"011011111",
  24482=>"111111001",
  24483=>"111100111",
  24484=>"011011111",
  24485=>"111111111",
  24486=>"100000000",
  24487=>"000001011",
  24488=>"111111111",
  24489=>"000000110",
  24490=>"110110110",
  24491=>"111000000",
  24492=>"000000000",
  24493=>"000001111",
  24494=>"110000001",
  24495=>"101101101",
  24496=>"000000000",
  24497=>"001101111",
  24498=>"111111111",
  24499=>"111101111",
  24500=>"000000000",
  24501=>"011011111",
  24502=>"011101000",
  24503=>"111110010",
  24504=>"000000000",
  24505=>"000000000",
  24506=>"111111111",
  24507=>"000000000",
  24508=>"111000000",
  24509=>"000000001",
  24510=>"000010000",
  24511=>"110111111",
  24512=>"011000000",
  24513=>"111101101",
  24514=>"111011000",
  24515=>"000000000",
  24516=>"010010001",
  24517=>"011111111",
  24518=>"000001111",
  24519=>"001101111",
  24520=>"101000000",
  24521=>"111111111",
  24522=>"000000111",
  24523=>"111111111",
  24524=>"000001111",
  24525=>"111111111",
  24526=>"000011011",
  24527=>"000000000",
  24528=>"000000000",
  24529=>"111111011",
  24530=>"110111111",
  24531=>"101101111",
  24532=>"011100000",
  24533=>"000010111",
  24534=>"000100110",
  24535=>"011111000",
  24536=>"111011000",
  24537=>"111001000",
  24538=>"000000000",
  24539=>"111000010",
  24540=>"111001100",
  24541=>"111111001",
  24542=>"001000000",
  24543=>"110111111",
  24544=>"000111111",
  24545=>"111111111",
  24546=>"110010000",
  24547=>"111110000",
  24548=>"111000000",
  24549=>"000011111",
  24550=>"011011111",
  24551=>"000000001",
  24552=>"001000000",
  24553=>"000000001",
  24554=>"000010111",
  24555=>"000000001",
  24556=>"010111111",
  24557=>"011011111",
  24558=>"000000000",
  24559=>"111000010",
  24560=>"000000111",
  24561=>"111111111",
  24562=>"111111111",
  24563=>"001101101",
  24564=>"111111011",
  24565=>"100111111",
  24566=>"101001000",
  24567=>"111111000",
  24568=>"111111111",
  24569=>"001101111",
  24570=>"101000000",
  24571=>"111110100",
  24572=>"101101111",
  24573=>"100110111",
  24574=>"000010000",
  24575=>"000000000",
  24576=>"111011001",
  24577=>"000111111",
  24578=>"111011001",
  24579=>"000000000",
  24580=>"001000000",
  24581=>"100111110",
  24582=>"000000001",
  24583=>"111101101",
  24584=>"000011111",
  24585=>"000101111",
  24586=>"001010010",
  24587=>"110111111",
  24588=>"000000000",
  24589=>"011000001",
  24590=>"011000001",
  24591=>"000100111",
  24592=>"001011111",
  24593=>"000000000",
  24594=>"111110100",
  24595=>"000000000",
  24596=>"000000111",
  24597=>"000000101",
  24598=>"110111111",
  24599=>"110111100",
  24600=>"001000000",
  24601=>"100110011",
  24602=>"000001001",
  24603=>"111000000",
  24604=>"000000000",
  24605=>"100000000",
  24606=>"111011101",
  24607=>"011001111",
  24608=>"000111111",
  24609=>"000000000",
  24610=>"101100100",
  24611=>"111111110",
  24612=>"111111000",
  24613=>"100000000",
  24614=>"000000000",
  24615=>"001001001",
  24616=>"000000000",
  24617=>"000111111",
  24618=>"111111000",
  24619=>"111111111",
  24620=>"001111111",
  24621=>"111111111",
  24622=>"111111110",
  24623=>"000001000",
  24624=>"111111111",
  24625=>"000000111",
  24626=>"000001000",
  24627=>"111111111",
  24628=>"111111000",
  24629=>"100000111",
  24630=>"000000100",
  24631=>"101101100",
  24632=>"111011111",
  24633=>"111011100",
  24634=>"000010010",
  24635=>"100000000",
  24636=>"111100101",
  24637=>"111111000",
  24638=>"000000010",
  24639=>"001111011",
  24640=>"011100110",
  24641=>"010010000",
  24642=>"000111011",
  24643=>"100000000",
  24644=>"000100000",
  24645=>"011011011",
  24646=>"001001111",
  24647=>"000000000",
  24648=>"000011011",
  24649=>"111101001",
  24650=>"011011010",
  24651=>"010000000",
  24652=>"101111101",
  24653=>"101111111",
  24654=>"000000000",
  24655=>"000111111",
  24656=>"000000000",
  24657=>"110000000",
  24658=>"111110111",
  24659=>"111110000",
  24660=>"010111000",
  24661=>"000000001",
  24662=>"000010111",
  24663=>"111111111",
  24664=>"100000000",
  24665=>"111001001",
  24666=>"000000001",
  24667=>"000001001",
  24668=>"000111111",
  24669=>"111111001",
  24670=>"000010000",
  24671=>"111111111",
  24672=>"110110111",
  24673=>"111111111",
  24674=>"111111111",
  24675=>"000000000",
  24676=>"111111011",
  24677=>"100000100",
  24678=>"111000000",
  24679=>"111000000",
  24680=>"110111111",
  24681=>"000000000",
  24682=>"111000110",
  24683=>"100000011",
  24684=>"100011001",
  24685=>"010011111",
  24686=>"000000000",
  24687=>"001000000",
  24688=>"111111111",
  24689=>"110000000",
  24690=>"100100110",
  24691=>"000110111",
  24692=>"110100000",
  24693=>"000000000",
  24694=>"000111111",
  24695=>"111111111",
  24696=>"101101111",
  24697=>"100000000",
  24698=>"001000000",
  24699=>"000100101",
  24700=>"000000010",
  24701=>"000000000",
  24702=>"000000000",
  24703=>"000010110",
  24704=>"000000000",
  24705=>"100110110",
  24706=>"111111111",
  24707=>"000000000",
  24708=>"110001111",
  24709=>"110000111",
  24710=>"000000000",
  24711=>"111001101",
  24712=>"010010110",
  24713=>"000000110",
  24714=>"000111011",
  24715=>"000000000",
  24716=>"011011000",
  24717=>"101100000",
  24718=>"100000000",
  24719=>"000010000",
  24720=>"101111111",
  24721=>"111110100",
  24722=>"111000100",
  24723=>"111000010",
  24724=>"111111000",
  24725=>"001111111",
  24726=>"000000100",
  24727=>"000001011",
  24728=>"000000110",
  24729=>"001001000",
  24730=>"111111111",
  24731=>"000000100",
  24732=>"100000000",
  24733=>"101110110",
  24734=>"111111000",
  24735=>"010111011",
  24736=>"101111111",
  24737=>"001111100",
  24738=>"001100111",
  24739=>"000000000",
  24740=>"100000000",
  24741=>"011011111",
  24742=>"111111000",
  24743=>"100110100",
  24744=>"001001000",
  24745=>"111111100",
  24746=>"000000001",
  24747=>"000100000",
  24748=>"111011001",
  24749=>"111101100",
  24750=>"001010000",
  24751=>"110100110",
  24752=>"000111111",
  24753=>"111111100",
  24754=>"111111111",
  24755=>"000111111",
  24756=>"000011011",
  24757=>"011001011",
  24758=>"000100100",
  24759=>"000000000",
  24760=>"000001011",
  24761=>"000000000",
  24762=>"111001000",
  24763=>"101001000",
  24764=>"000001001",
  24765=>"001101111",
  24766=>"000000000",
  24767=>"111111111",
  24768=>"000000000",
  24769=>"000000010",
  24770=>"111111111",
  24771=>"111111011",
  24772=>"000101111",
  24773=>"000000000",
  24774=>"011000000",
  24775=>"000001000",
  24776=>"000011011",
  24777=>"100110111",
  24778=>"000000001",
  24779=>"000000000",
  24780=>"000000000",
  24781=>"000000000",
  24782=>"001000011",
  24783=>"111111111",
  24784=>"011000100",
  24785=>"000010111",
  24786=>"000000000",
  24787=>"000000000",
  24788=>"001001000",
  24789=>"111111111",
  24790=>"001001011",
  24791=>"011001000",
  24792=>"000000111",
  24793=>"000010000",
  24794=>"100111111",
  24795=>"001001011",
  24796=>"111010000",
  24797=>"110100000",
  24798=>"000000000",
  24799=>"111001101",
  24800=>"000000000",
  24801=>"111111011",
  24802=>"111100000",
  24803=>"000000000",
  24804=>"000000000",
  24805=>"001100100",
  24806=>"110001001",
  24807=>"001010010",
  24808=>"000000000",
  24809=>"111111111",
  24810=>"111011111",
  24811=>"110011000",
  24812=>"110000000",
  24813=>"000000000",
  24814=>"111010001",
  24815=>"111110111",
  24816=>"011111011",
  24817=>"111100100",
  24818=>"111100100",
  24819=>"000111011",
  24820=>"011011111",
  24821=>"111111100",
  24822=>"000100100",
  24823=>"111111111",
  24824=>"101100100",
  24825=>"000000000",
  24826=>"011001000",
  24827=>"001011000",
  24828=>"000100010",
  24829=>"111100100",
  24830=>"000101100",
  24831=>"000001000",
  24832=>"001001011",
  24833=>"111111000",
  24834=>"110110111",
  24835=>"111100000",
  24836=>"111111100",
  24837=>"110001000",
  24838=>"011000001",
  24839=>"110110001",
  24840=>"111111011",
  24841=>"000000000",
  24842=>"111000111",
  24843=>"000000000",
  24844=>"111111101",
  24845=>"100100000",
  24846=>"010000000",
  24847=>"000110110",
  24848=>"111111011",
  24849=>"110000000",
  24850=>"000000000",
  24851=>"111111000",
  24852=>"100000000",
  24853=>"001000011",
  24854=>"111111000",
  24855=>"111111100",
  24856=>"111111001",
  24857=>"000001111",
  24858=>"000000000",
  24859=>"011000000",
  24860=>"100100101",
  24861=>"011111111",
  24862=>"010110010",
  24863=>"001111111",
  24864=>"111111000",
  24865=>"000000101",
  24866=>"000000111",
  24867=>"111111110",
  24868=>"111111111",
  24869=>"011111111",
  24870=>"111011011",
  24871=>"111111011",
  24872=>"111100000",
  24873=>"000000000",
  24874=>"001001000",
  24875=>"000011001",
  24876=>"000011111",
  24877=>"001111111",
  24878=>"111111111",
  24879=>"001001111",
  24880=>"000000000",
  24881=>"110010011",
  24882=>"100111110",
  24883=>"111011000",
  24884=>"000000000",
  24885=>"100000000",
  24886=>"111101101",
  24887=>"011111111",
  24888=>"000000000",
  24889=>"000111001",
  24890=>"111111000",
  24891=>"111001001",
  24892=>"001001000",
  24893=>"001101001",
  24894=>"111111111",
  24895=>"011111111",
  24896=>"111111111",
  24897=>"100110111",
  24898=>"000100101",
  24899=>"111110000",
  24900=>"000000101",
  24901=>"011111000",
  24902=>"111111111",
  24903=>"111111101",
  24904=>"000000000",
  24905=>"000000111",
  24906=>"011111000",
  24907=>"111111100",
  24908=>"100000000",
  24909=>"101100110",
  24910=>"001111001",
  24911=>"101001001",
  24912=>"111111101",
  24913=>"001011111",
  24914=>"111111111",
  24915=>"000001000",
  24916=>"000110110",
  24917=>"011001001",
  24918=>"110000000",
  24919=>"110100111",
  24920=>"000011111",
  24921=>"111111111",
  24922=>"001101100",
  24923=>"011000110",
  24924=>"000111111",
  24925=>"000111010",
  24926=>"000000110",
  24927=>"101111011",
  24928=>"000001111",
  24929=>"001111111",
  24930=>"100100110",
  24931=>"111001111",
  24932=>"001011111",
  24933=>"110111111",
  24934=>"111111011",
  24935=>"111011001",
  24936=>"110111111",
  24937=>"100111111",
  24938=>"100111111",
  24939=>"111111110",
  24940=>"000100001",
  24941=>"000000000",
  24942=>"000000000",
  24943=>"111111111",
  24944=>"000000100",
  24945=>"111011010",
  24946=>"110110111",
  24947=>"100100111",
  24948=>"000000000",
  24949=>"011011111",
  24950=>"000000111",
  24951=>"000100111",
  24952=>"000000000",
  24953=>"000001111",
  24954=>"110111111",
  24955=>"010000000",
  24956=>"001111110",
  24957=>"000000011",
  24958=>"101101001",
  24959=>"000001111",
  24960=>"010110000",
  24961=>"111011000",
  24962=>"100100100",
  24963=>"111111111",
  24964=>"000011001",
  24965=>"000000010",
  24966=>"000111110",
  24967=>"111111011",
  24968=>"001001101",
  24969=>"111000001",
  24970=>"000000001",
  24971=>"000000000",
  24972=>"101001001",
  24973=>"110100110",
  24974=>"000000000",
  24975=>"011111011",
  24976=>"111111111",
  24977=>"000000100",
  24978=>"000011001",
  24979=>"000000000",
  24980=>"111111011",
  24981=>"011110010",
  24982=>"100000010",
  24983=>"111111011",
  24984=>"100000000",
  24985=>"111111111",
  24986=>"000000000",
  24987=>"111111111",
  24988=>"111111111",
  24989=>"000110110",
  24990=>"100000000",
  24991=>"000011111",
  24992=>"011110011",
  24993=>"110100101",
  24994=>"001000000",
  24995=>"101100111",
  24996=>"011000111",
  24997=>"111111100",
  24998=>"111001011",
  24999=>"011110000",
  25000=>"000000001",
  25001=>"111111110",
  25002=>"000001000",
  25003=>"111111000",
  25004=>"000001111",
  25005=>"111111110",
  25006=>"111111111",
  25007=>"111111011",
  25008=>"000000111",
  25009=>"000000000",
  25010=>"000000001",
  25011=>"110111000",
  25012=>"000000100",
  25013=>"110111111",
  25014=>"000000000",
  25015=>"000000001",
  25016=>"011001000",
  25017=>"111101111",
  25018=>"000001000",
  25019=>"111110111",
  25020=>"000100111",
  25021=>"111111011",
  25022=>"000000000",
  25023=>"111111111",
  25024=>"111111001",
  25025=>"000100111",
  25026=>"001110111",
  25027=>"111111100",
  25028=>"100111111",
  25029=>"011001100",
  25030=>"111101111",
  25031=>"001000000",
  25032=>"000001100",
  25033=>"000101111",
  25034=>"111111111",
  25035=>"000001000",
  25036=>"101000000",
  25037=>"111111111",
  25038=>"111000100",
  25039=>"111011000",
  25040=>"111100100",
  25041=>"111011000",
  25042=>"000000000",
  25043=>"111111111",
  25044=>"000000000",
  25045=>"110110000",
  25046=>"001111111",
  25047=>"000010000",
  25048=>"000110111",
  25049=>"000110000",
  25050=>"000111111",
  25051=>"111110100",
  25052=>"000100100",
  25053=>"100000010",
  25054=>"000000111",
  25055=>"111111111",
  25056=>"111001111",
  25057=>"110110010",
  25058=>"100111011",
  25059=>"100100000",
  25060=>"111101111",
  25061=>"011011001",
  25062=>"000110000",
  25063=>"000000111",
  25064=>"001000111",
  25065=>"111111111",
  25066=>"100111111",
  25067=>"100111111",
  25068=>"111100000",
  25069=>"111110100",
  25070=>"100100111",
  25071=>"111111100",
  25072=>"110100001",
  25073=>"000000000",
  25074=>"111111111",
  25075=>"000111111",
  25076=>"001000000",
  25077=>"011001001",
  25078=>"111111101",
  25079=>"101001001",
  25080=>"111000010",
  25081=>"001001100",
  25082=>"000000100",
  25083=>"000000101",
  25084=>"111111011",
  25085=>"110111111",
  25086=>"110011011",
  25087=>"000111110",
  25088=>"000001111",
  25089=>"000111000",
  25090=>"111111111",
  25091=>"111111111",
  25092=>"111100110",
  25093=>"101100110",
  25094=>"000011011",
  25095=>"101000101",
  25096=>"000110000",
  25097=>"000000100",
  25098=>"111111000",
  25099=>"111001000",
  25100=>"000010000",
  25101=>"000000000",
  25102=>"000000011",
  25103=>"000111111",
  25104=>"000000100",
  25105=>"110111111",
  25106=>"100100111",
  25107=>"000000101",
  25108=>"111111111",
  25109=>"010000000",
  25110=>"010111101",
  25111=>"000100111",
  25112=>"111111011",
  25113=>"100100101",
  25114=>"111111111",
  25115=>"001010000",
  25116=>"100000000",
  25117=>"011111111",
  25118=>"000000010",
  25119=>"100110000",
  25120=>"111111110",
  25121=>"111100000",
  25122=>"001001111",
  25123=>"111011001",
  25124=>"000000000",
  25125=>"000000000",
  25126=>"000100100",
  25127=>"101111111",
  25128=>"011100100",
  25129=>"111011111",
  25130=>"111111111",
  25131=>"000000000",
  25132=>"000000000",
  25133=>"000000000",
  25134=>"011100001",
  25135=>"000100111",
  25136=>"000000100",
  25137=>"011101000",
  25138=>"011011011",
  25139=>"111111001",
  25140=>"011001011",
  25141=>"110110000",
  25142=>"110111011",
  25143=>"000100111",
  25144=>"000000100",
  25145=>"010110001",
  25146=>"011110101",
  25147=>"111111111",
  25148=>"111001111",
  25149=>"000000000",
  25150=>"000000000",
  25151=>"000000000",
  25152=>"000000111",
  25153=>"011000010",
  25154=>"000000111",
  25155=>"000011011",
  25156=>"110111100",
  25157=>"111000000",
  25158=>"000010111",
  25159=>"000000000",
  25160=>"011011011",
  25161=>"111001011",
  25162=>"111111111",
  25163=>"111000100",
  25164=>"000000000",
  25165=>"111110100",
  25166=>"000000000",
  25167=>"111000000",
  25168=>"000100000",
  25169=>"011000000",
  25170=>"111111010",
  25171=>"100100110",
  25172=>"100000000",
  25173=>"000000010",
  25174=>"011010111",
  25175=>"111101111",
  25176=>"111111001",
  25177=>"001000001",
  25178=>"001001001",
  25179=>"100100000",
  25180=>"111001000",
  25181=>"000000100",
  25182=>"111111110",
  25183=>"001111110",
  25184=>"110000000",
  25185=>"001000001",
  25186=>"110100000",
  25187=>"000001001",
  25188=>"101111101",
  25189=>"110111111",
  25190=>"111110001",
  25191=>"111011111",
  25192=>"000000000",
  25193=>"000000111",
  25194=>"000000010",
  25195=>"000010010",
  25196=>"000000000",
  25197=>"000000100",
  25198=>"111001011",
  25199=>"111001011",
  25200=>"110110111",
  25201=>"011011010",
  25202=>"011111111",
  25203=>"011101000",
  25204=>"000010111",
  25205=>"000100000",
  25206=>"000000000",
  25207=>"110000001",
  25208=>"100100101",
  25209=>"000000000",
  25210=>"100100000",
  25211=>"111000000",
  25212=>"110110100",
  25213=>"111111111",
  25214=>"000000000",
  25215=>"000000000",
  25216=>"000000001",
  25217=>"111000111",
  25218=>"010111001",
  25219=>"111111011",
  25220=>"000000001",
  25221=>"001111111",
  25222=>"100111000",
  25223=>"000100000",
  25224=>"000000100",
  25225=>"000000111",
  25226=>"111011000",
  25227=>"000001111",
  25228=>"000001111",
  25229=>"111110110",
  25230=>"000000111",
  25231=>"000000001",
  25232=>"111001000",
  25233=>"010000000",
  25234=>"000001111",
  25235=>"111111111",
  25236=>"010000000",
  25237=>"100111111",
  25238=>"000000100",
  25239=>"000000000",
  25240=>"000000000",
  25241=>"101110000",
  25242=>"100111111",
  25243=>"101001001",
  25244=>"000111111",
  25245=>"000000000",
  25246=>"001101111",
  25247=>"000000111",
  25248=>"000010000",
  25249=>"000000000",
  25250=>"001010000",
  25251=>"000111111",
  25252=>"000101101",
  25253=>"000000011",
  25254=>"000101111",
  25255=>"111111111",
  25256=>"111111111",
  25257=>"001110100",
  25258=>"000000111",
  25259=>"111111111",
  25260=>"000000010",
  25261=>"001111111",
  25262=>"111111001",
  25263=>"111111001",
  25264=>"000101001",
  25265=>"100101001",
  25266=>"000111000",
  25267=>"100000000",
  25268=>"011111111",
  25269=>"111111110",
  25270=>"000110000",
  25271=>"001001111",
  25272=>"011100000",
  25273=>"111111100",
  25274=>"111111011",
  25275=>"100111111",
  25276=>"111001000",
  25277=>"111111111",
  25278=>"000111111",
  25279=>"111111111",
  25280=>"000000001",
  25281=>"000000110",
  25282=>"000000000",
  25283=>"111111111",
  25284=>"111111111",
  25285=>"000000000",
  25286=>"000000101",
  25287=>"100100110",
  25288=>"110110110",
  25289=>"000000000",
  25290=>"001001001",
  25291=>"000000000",
  25292=>"000000111",
  25293=>"000110111",
  25294=>"111110110",
  25295=>"110111111",
  25296=>"000110000",
  25297=>"000000000",
  25298=>"111111111",
  25299=>"000000111",
  25300=>"001101111",
  25301=>"000000000",
  25302=>"000000000",
  25303=>"111111010",
  25304=>"000110000",
  25305=>"000000001",
  25306=>"111001111",
  25307=>"111001111",
  25308=>"110111111",
  25309=>"011011111",
  25310=>"000000000",
  25311=>"110100101",
  25312=>"011011111",
  25313=>"000011111",
  25314=>"110110000",
  25315=>"001000000",
  25316=>"000110111",
  25317=>"111111111",
  25318=>"000000000",
  25319=>"100000000",
  25320=>"111000000",
  25321=>"000000000",
  25322=>"110000000",
  25323=>"111111000",
  25324=>"011011001",
  25325=>"000110001",
  25326=>"110111100",
  25327=>"000000000",
  25328=>"100000000",
  25329=>"000000000",
  25330=>"111111101",
  25331=>"001000001",
  25332=>"110000000",
  25333=>"100110000",
  25334=>"011111111",
  25335=>"111011111",
  25336=>"100100000",
  25337=>"000000000",
  25338=>"111100100",
  25339=>"111110100",
  25340=>"110110111",
  25341=>"000010000",
  25342=>"110101111",
  25343=>"000100110",
  25344=>"100000000",
  25345=>"001000000",
  25346=>"111111111",
  25347=>"110111111",
  25348=>"000100000",
  25349=>"000000000",
  25350=>"000000000",
  25351=>"001000011",
  25352=>"000000000",
  25353=>"001001111",
  25354=>"110000000",
  25355=>"011111010",
  25356=>"000000100",
  25357=>"011000000",
  25358=>"000000000",
  25359=>"000000000",
  25360=>"110000001",
  25361=>"110111111",
  25362=>"000000111",
  25363=>"011000000",
  25364=>"111111111",
  25365=>"000111000",
  25366=>"001101001",
  25367=>"111111001",
  25368=>"110110110",
  25369=>"000110111",
  25370=>"110110111",
  25371=>"110110111",
  25372=>"110111111",
  25373=>"110111111",
  25374=>"010000000",
  25375=>"111111111",
  25376=>"000111011",
  25377=>"111001000",
  25378=>"111001001",
  25379=>"000000000",
  25380=>"000111000",
  25381=>"111110000",
  25382=>"001001001",
  25383=>"000000000",
  25384=>"101100101",
  25385=>"000000100",
  25386=>"011000100",
  25387=>"111111001",
  25388=>"111010011",
  25389=>"110111111",
  25390=>"000000000",
  25391=>"111000000",
  25392=>"000000000",
  25393=>"101111111",
  25394=>"000000000",
  25395=>"000000111",
  25396=>"111111000",
  25397=>"101111111",
  25398=>"110110110",
  25399=>"111111001",
  25400=>"000110110",
  25401=>"100110111",
  25402=>"110001000",
  25403=>"000101111",
  25404=>"000000000",
  25405=>"001000101",
  25406=>"011011000",
  25407=>"000000000",
  25408=>"000000000",
  25409=>"111111111",
  25410=>"101100111",
  25411=>"111011001",
  25412=>"000000000",
  25413=>"001111001",
  25414=>"000000000",
  25415=>"100001011",
  25416=>"000110100",
  25417=>"000100000",
  25418=>"111111101",
  25419=>"111011111",
  25420=>"000110110",
  25421=>"010000000",
  25422=>"000000000",
  25423=>"000010111",
  25424=>"110110110",
  25425=>"010000000",
  25426=>"111000011",
  25427=>"000110110",
  25428=>"111111111",
  25429=>"011001011",
  25430=>"111111111",
  25431=>"000000100",
  25432=>"110000011",
  25433=>"001001000",
  25434=>"111111000",
  25435=>"111111001",
  25436=>"000000000",
  25437=>"111111111",
  25438=>"111010001",
  25439=>"000000000",
  25440=>"110110000",
  25441=>"001000111",
  25442=>"000001000",
  25443=>"000000101",
  25444=>"000001001",
  25445=>"110000000",
  25446=>"000011111",
  25447=>"000000000",
  25448=>"110110011",
  25449=>"100110110",
  25450=>"000101100",
  25451=>"010000000",
  25452=>"000110100",
  25453=>"011111011",
  25454=>"000000111",
  25455=>"000000000",
  25456=>"110111000",
  25457=>"000000000",
  25458=>"110111111",
  25459=>"000000000",
  25460=>"100100111",
  25461=>"000000000",
  25462=>"000010001",
  25463=>"000111111",
  25464=>"100111111",
  25465=>"000000000",
  25466=>"000000000",
  25467=>"110110110",
  25468=>"111111000",
  25469=>"000000111",
  25470=>"111100110",
  25471=>"000001111",
  25472=>"111111111",
  25473=>"000000110",
  25474=>"111100100",
  25475=>"001111111",
  25476=>"001000101",
  25477=>"111111111",
  25478=>"110110110",
  25479=>"001001001",
  25480=>"001000000",
  25481=>"000000111",
  25482=>"000000100",
  25483=>"111011000",
  25484=>"101001111",
  25485=>"000000000",
  25486=>"111011001",
  25487=>"111011000",
  25488=>"000000000",
  25489=>"111111000",
  25490=>"111110001",
  25491=>"111110100",
  25492=>"010010010",
  25493=>"000000110",
  25494=>"111100110",
  25495=>"000001000",
  25496=>"010011000",
  25497=>"000000000",
  25498=>"000000000",
  25499=>"111111111",
  25500=>"101101111",
  25501=>"001011000",
  25502=>"000000001",
  25503=>"110111111",
  25504=>"100100100",
  25505=>"000001001",
  25506=>"111001011",
  25507=>"111101111",
  25508=>"001000000",
  25509=>"000000111",
  25510=>"011000000",
  25511=>"111111111",
  25512=>"110010111",
  25513=>"100110111",
  25514=>"111111000",
  25515=>"001000011",
  25516=>"100001111",
  25517=>"111110000",
  25518=>"000000011",
  25519=>"111111000",
  25520=>"000000000",
  25521=>"010011001",
  25522=>"000000000",
  25523=>"110000000",
  25524=>"111111010",
  25525=>"111010001",
  25526=>"000000011",
  25527=>"000000000",
  25528=>"111111101",
  25529=>"101101100",
  25530=>"111100100",
  25531=>"101111111",
  25532=>"110110111",
  25533=>"111110110",
  25534=>"000111110",
  25535=>"000001001",
  25536=>"000000101",
  25537=>"000000000",
  25538=>"000000000",
  25539=>"000000000",
  25540=>"011111111",
  25541=>"111101101",
  25542=>"000000110",
  25543=>"000000000",
  25544=>"100000000",
  25545=>"000000000",
  25546=>"100000000",
  25547=>"111001111",
  25548=>"011000000",
  25549=>"111111001",
  25550=>"001110111",
  25551=>"111111111",
  25552=>"010110011",
  25553=>"111101101",
  25554=>"000000000",
  25555=>"001001111",
  25556=>"111111001",
  25557=>"100111111",
  25558=>"000000000",
  25559=>"011001011",
  25560=>"001011001",
  25561=>"110100100",
  25562=>"111011001",
  25563=>"000000111",
  25564=>"111111011",
  25565=>"011111011",
  25566=>"110110100",
  25567=>"000000100",
  25568=>"000000000",
  25569=>"000000110",
  25570=>"111111010",
  25571=>"111111111",
  25572=>"001001111",
  25573=>"111000000",
  25574=>"111111000",
  25575=>"000000000",
  25576=>"000110111",
  25577=>"100111111",
  25578=>"110111111",
  25579=>"000000110",
  25580=>"111011000",
  25581=>"000000100",
  25582=>"001001000",
  25583=>"100110110",
  25584=>"010011100",
  25585=>"011111011",
  25586=>"111111111",
  25587=>"011011011",
  25588=>"111000000",
  25589=>"000000110",
  25590=>"000110111",
  25591=>"000111111",
  25592=>"111000111",
  25593=>"100000110",
  25594=>"000110110",
  25595=>"101111111",
  25596=>"000000010",
  25597=>"000100101",
  25598=>"101100110",
  25599=>"001111111",
  25600=>"000000000",
  25601=>"000000000",
  25602=>"000000000",
  25603=>"111111111",
  25604=>"100110111",
  25605=>"011011001",
  25606=>"000000100",
  25607=>"000000000",
  25608=>"000000001",
  25609=>"101100000",
  25610=>"111111111",
  25611=>"111111111",
  25612=>"001011111",
  25613=>"001111110",
  25614=>"111100000",
  25615=>"111111110",
  25616=>"000001111",
  25617=>"001000000",
  25618=>"000001000",
  25619=>"111101111",
  25620=>"011011011",
  25621=>"000010111",
  25622=>"110111111",
  25623=>"111111110",
  25624=>"011011100",
  25625=>"000001011",
  25626=>"111111001",
  25627=>"000000000",
  25628=>"000000111",
  25629=>"000000000",
  25630=>"110110111",
  25631=>"111101111",
  25632=>"111111000",
  25633=>"111111110",
  25634=>"111111011",
  25635=>"111011001",
  25636=>"111111001",
  25637=>"100000000",
  25638=>"111111111",
  25639=>"111000111",
  25640=>"111111111",
  25641=>"000000000",
  25642=>"111100101",
  25643=>"110100100",
  25644=>"111100000",
  25645=>"100100110",
  25646=>"000011011",
  25647=>"100110000",
  25648=>"111111111",
  25649=>"111001011",
  25650=>"000000000",
  25651=>"100100111",
  25652=>"000110100",
  25653=>"000011111",
  25654=>"111001001",
  25655=>"011010000",
  25656=>"111000000",
  25657=>"111100000",
  25658=>"100000000",
  25659=>"111011011",
  25660=>"000100111",
  25661=>"111111111",
  25662=>"100100000",
  25663=>"000000000",
  25664=>"000100100",
  25665=>"100100000",
  25666=>"111100100",
  25667=>"000000001",
  25668=>"000001000",
  25669=>"111011011",
  25670=>"111000000",
  25671=>"111111111",
  25672=>"011010000",
  25673=>"111111111",
  25674=>"000111111",
  25675=>"111000000",
  25676=>"111111111",
  25677=>"000000000",
  25678=>"000010111",
  25679=>"011111111",
  25680=>"111111111",
  25681=>"001001011",
  25682=>"111011011",
  25683=>"001001000",
  25684=>"000000111",
  25685=>"000100100",
  25686=>"111110110",
  25687=>"111111111",
  25688=>"111011111",
  25689=>"001000011",
  25690=>"111111101",
  25691=>"000111111",
  25692=>"000000010",
  25693=>"000000000",
  25694=>"111111000",
  25695=>"100010000",
  25696=>"000000111",
  25697=>"111111010",
  25698=>"111000001",
  25699=>"111111111",
  25700=>"001110111",
  25701=>"000111111",
  25702=>"011011010",
  25703=>"000000000",
  25704=>"111111111",
  25705=>"111111111",
  25706=>"011000000",
  25707=>"001001101",
  25708=>"011000011",
  25709=>"111001101",
  25710=>"011000000",
  25711=>"111111100",
  25712=>"000000000",
  25713=>"101010011",
  25714=>"111111000",
  25715=>"001000000",
  25716=>"111111111",
  25717=>"001001001",
  25718=>"000000000",
  25719=>"000000000",
  25720=>"111111111",
  25721=>"000000100",
  25722=>"000001001",
  25723=>"111000000",
  25724=>"000001001",
  25725=>"011111111",
  25726=>"001000001",
  25727=>"111111000",
  25728=>"111111111",
  25729=>"111111100",
  25730=>"000000000",
  25731=>"001010010",
  25732=>"001000100",
  25733=>"101101111",
  25734=>"000000000",
  25735=>"011111011",
  25736=>"111111111",
  25737=>"000000000",
  25738=>"111111111",
  25739=>"111111110",
  25740=>"011000000",
  25741=>"111111111",
  25742=>"000000111",
  25743=>"001000000",
  25744=>"111111111",
  25745=>"111111111",
  25746=>"111111111",
  25747=>"011000000",
  25748=>"001001000",
  25749=>"111101100",
  25750=>"011010011",
  25751=>"111111111",
  25752=>"101101110",
  25753=>"000000100",
  25754=>"001000000",
  25755=>"000000000",
  25756=>"111110110",
  25757=>"000000000",
  25758=>"000000000",
  25759=>"101100101",
  25760=>"000000001",
  25761=>"111111111",
  25762=>"111110111",
  25763=>"111111100",
  25764=>"000001001",
  25765=>"110111111",
  25766=>"111111111",
  25767=>"100100100",
  25768=>"111111010",
  25769=>"000100111",
  25770=>"111000000",
  25771=>"000111111",
  25772=>"111111111",
  25773=>"011010011",
  25774=>"100100111",
  25775=>"111111111",
  25776=>"111000000",
  25777=>"000000111",
  25778=>"000000000",
  25779=>"000000000",
  25780=>"100100101",
  25781=>"111101111",
  25782=>"111011001",
  25783=>"111111111",
  25784=>"100100101",
  25785=>"111111111",
  25786=>"000000000",
  25787=>"111111111",
  25788=>"010011011",
  25789=>"000000000",
  25790=>"111111111",
  25791=>"000110010",
  25792=>"000000000",
  25793=>"111110110",
  25794=>"000000000",
  25795=>"010000000",
  25796=>"111011000",
  25797=>"111000000",
  25798=>"000111111",
  25799=>"111111111",
  25800=>"100100111",
  25801=>"111001001",
  25802=>"111011111",
  25803=>"111111001",
  25804=>"111110111",
  25805=>"000110100",
  25806=>"000000000",
  25807=>"000100000",
  25808=>"111111111",
  25809=>"000000000",
  25810=>"000110000",
  25811=>"111111111",
  25812=>"101100111",
  25813=>"111011001",
  25814=>"111000010",
  25815=>"100100000",
  25816=>"111111001",
  25817=>"101111111",
  25818=>"000000000",
  25819=>"000000011",
  25820=>"001000011",
  25821=>"010010111",
  25822=>"111011011",
  25823=>"000000110",
  25824=>"000000000",
  25825=>"000000000",
  25826=>"001000000",
  25827=>"111111000",
  25828=>"111111100",
  25829=>"110100000",
  25830=>"111111111",
  25831=>"111111111",
  25832=>"001111111",
  25833=>"001000110",
  25834=>"000000000",
  25835=>"111000000",
  25836=>"000111111",
  25837=>"111111111",
  25838=>"111110111",
  25839=>"000111111",
  25840=>"111111111",
  25841=>"000000000",
  25842=>"001111111",
  25843=>"111001111",
  25844=>"110100000",
  25845=>"001001000",
  25846=>"000000000",
  25847=>"111011011",
  25848=>"000000000",
  25849=>"000000000",
  25850=>"111000110",
  25851=>"111111000",
  25852=>"111101001",
  25853=>"000000001",
  25854=>"110111011",
  25855=>"111111000",
  25856=>"000000000",
  25857=>"000000000",
  25858=>"111111111",
  25859=>"110110100",
  25860=>"100101111",
  25861=>"000000000",
  25862=>"101101101",
  25863=>"000000000",
  25864=>"000110100",
  25865=>"000000000",
  25866=>"000100111",
  25867=>"101111111",
  25868=>"011011111",
  25869=>"111111111",
  25870=>"111001000",
  25871=>"111100110",
  25872=>"000000100",
  25873=>"000000110",
  25874=>"111111111",
  25875=>"010000011",
  25876=>"000001001",
  25877=>"000000001",
  25878=>"011011011",
  25879=>"000000000",
  25880=>"100110011",
  25881=>"000000000",
  25882=>"000100100",
  25883=>"001000000",
  25884=>"100000000",
  25885=>"111111111",
  25886=>"000110110",
  25887=>"000000000",
  25888=>"111111001",
  25889=>"011111111",
  25890=>"010010011",
  25891=>"101111111",
  25892=>"001000001",
  25893=>"100111111",
  25894=>"000110110",
  25895=>"111111011",
  25896=>"111111111",
  25897=>"000000000",
  25898=>"000000000",
  25899=>"111111111",
  25900=>"111111111",
  25901=>"111111111",
  25902=>"000111000",
  25903=>"000000001",
  25904=>"001011111",
  25905=>"000000000",
  25906=>"110010011",
  25907=>"000000010",
  25908=>"000000000",
  25909=>"000000000",
  25910=>"000010000",
  25911=>"111000000",
  25912=>"000001000",
  25913=>"000000010",
  25914=>"000110111",
  25915=>"001101111",
  25916=>"110100011",
  25917=>"111010010",
  25918=>"110110110",
  25919=>"100111111",
  25920=>"111111111",
  25921=>"111110111",
  25922=>"000000000",
  25923=>"111111111",
  25924=>"000000000",
  25925=>"000000000",
  25926=>"000000111",
  25927=>"111111111",
  25928=>"111000000",
  25929=>"011111111",
  25930=>"101111011",
  25931=>"111011000",
  25932=>"010000111",
  25933=>"111111111",
  25934=>"111011000",
  25935=>"000000000",
  25936=>"000000000",
  25937=>"000110100",
  25938=>"100000111",
  25939=>"110010000",
  25940=>"000000000",
  25941=>"101110110",
  25942=>"110000000",
  25943=>"111111111",
  25944=>"111001111",
  25945=>"000000000",
  25946=>"000000001",
  25947=>"011111111",
  25948=>"111111011",
  25949=>"111111111",
  25950=>"111011000",
  25951=>"111011000",
  25952=>"111111000",
  25953=>"111010111",
  25954=>"000001001",
  25955=>"000001111",
  25956=>"111111111",
  25957=>"000000000",
  25958=>"000000111",
  25959=>"111011111",
  25960=>"111000001",
  25961=>"000000001",
  25962=>"110111111",
  25963=>"010011011",
  25964=>"001000011",
  25965=>"011000011",
  25966=>"000000111",
  25967=>"110110110",
  25968=>"010110000",
  25969=>"000000000",
  25970=>"000000000",
  25971=>"110110110",
  25972=>"111111011",
  25973=>"101111111",
  25974=>"111111111",
  25975=>"000000000",
  25976=>"000000110",
  25977=>"000000010",
  25978=>"110110110",
  25979=>"000000000",
  25980=>"010000000",
  25981=>"111111000",
  25982=>"000000000",
  25983=>"100111111",
  25984=>"000001111",
  25985=>"110010000",
  25986=>"111111111",
  25987=>"111111000",
  25988=>"000000001",
  25989=>"100101101",
  25990=>"011010000",
  25991=>"000000011",
  25992=>"010000000",
  25993=>"000000110",
  25994=>"111001001",
  25995=>"111101001",
  25996=>"001000111",
  25997=>"000001001",
  25998=>"000111001",
  25999=>"111111111",
  26000=>"000000100",
  26001=>"000011111",
  26002=>"000000111",
  26003=>"011011110",
  26004=>"111111111",
  26005=>"000000000",
  26006=>"111111111",
  26007=>"111101011",
  26008=>"000001101",
  26009=>"111001000",
  26010=>"111111111",
  26011=>"000000001",
  26012=>"111111111",
  26013=>"010000000",
  26014=>"011111001",
  26015=>"110111000",
  26016=>"000001111",
  26017=>"111110010",
  26018=>"111100100",
  26019=>"001001011",
  26020=>"110100000",
  26021=>"110111111",
  26022=>"110110000",
  26023=>"110110110",
  26024=>"000000100",
  26025=>"011000000",
  26026=>"111111111",
  26027=>"111111111",
  26028=>"111111111",
  26029=>"001001000",
  26030=>"100000111",
  26031=>"111111111",
  26032=>"000000110",
  26033=>"011011011",
  26034=>"001000000",
  26035=>"111000001",
  26036=>"000000100",
  26037=>"000000100",
  26038=>"111111111",
  26039=>"111111010",
  26040=>"110110011",
  26041=>"111111011",
  26042=>"000000000",
  26043=>"111101111",
  26044=>"000000000",
  26045=>"100000001",
  26046=>"000111111",
  26047=>"111111111",
  26048=>"111000010",
  26049=>"000000000",
  26050=>"111001111",
  26051=>"000011010",
  26052=>"111110111",
  26053=>"100010101",
  26054=>"111000000",
  26055=>"001001000",
  26056=>"000000000",
  26057=>"100000000",
  26058=>"000000000",
  26059=>"111111111",
  26060=>"000001000",
  26061=>"111011111",
  26062=>"110110000",
  26063=>"110110011",
  26064=>"111111111",
  26065=>"111111100",
  26066=>"000100100",
  26067=>"111011001",
  26068=>"110110110",
  26069=>"000000100",
  26070=>"000000000",
  26071=>"110110111",
  26072=>"111000000",
  26073=>"100000000",
  26074=>"000000000",
  26075=>"000000000",
  26076=>"001011001",
  26077=>"111001001",
  26078=>"000111111",
  26079=>"000000111",
  26080=>"001000000",
  26081=>"000110111",
  26082=>"000000000",
  26083=>"111110100",
  26084=>"111110111",
  26085=>"100000000",
  26086=>"111111011",
  26087=>"000111111",
  26088=>"000000000",
  26089=>"000001001",
  26090=>"001111111",
  26091=>"000000101",
  26092=>"111000000",
  26093=>"100100100",
  26094=>"111111111",
  26095=>"111110110",
  26096=>"000000000",
  26097=>"111111100",
  26098=>"011000000",
  26099=>"001001000",
  26100=>"001000000",
  26101=>"111111111",
  26102=>"010000000",
  26103=>"000000000",
  26104=>"111111111",
  26105=>"000000000",
  26106=>"111001001",
  26107=>"110110010",
  26108=>"000000000",
  26109=>"000011111",
  26110=>"000000000",
  26111=>"000000000",
  26112=>"001111110",
  26113=>"001111100",
  26114=>"000000111",
  26115=>"111101111",
  26116=>"000111111",
  26117=>"000000000",
  26118=>"001000000",
  26119=>"111011000",
  26120=>"111111000",
  26121=>"111001001",
  26122=>"111111111",
  26123=>"011111111",
  26124=>"100000000",
  26125=>"111000010",
  26126=>"000000000",
  26127=>"000000000",
  26128=>"111001001",
  26129=>"001101000",
  26130=>"110111111",
  26131=>"001000000",
  26132=>"111101101",
  26133=>"000111111",
  26134=>"000010011",
  26135=>"101100100",
  26136=>"111111011",
  26137=>"000100001",
  26138=>"000000000",
  26139=>"110000001",
  26140=>"111110100",
  26141=>"000010111",
  26142=>"111011011",
  26143=>"001001111",
  26144=>"011011111",
  26145=>"000000000",
  26146=>"100000000",
  26147=>"000000000",
  26148=>"111111111",
  26149=>"111111111",
  26150=>"111011011",
  26151=>"111111001",
  26152=>"111001000",
  26153=>"001001111",
  26154=>"111110110",
  26155=>"111111100",
  26156=>"000000000",
  26157=>"000000000",
  26158=>"010111111",
  26159=>"000011011",
  26160=>"000000000",
  26161=>"000000000",
  26162=>"000001011",
  26163=>"100100111",
  26164=>"010000000",
  26165=>"100110110",
  26166=>"000111111",
  26167=>"000110000",
  26168=>"111111111",
  26169=>"000010000",
  26170=>"000000000",
  26171=>"000000000",
  26172=>"010011111",
  26173=>"110010000",
  26174=>"110111111",
  26175=>"000000000",
  26176=>"000000000",
  26177=>"111111111",
  26178=>"111111111",
  26179=>"000000000",
  26180=>"111001001",
  26181=>"000000000",
  26182=>"110000000",
  26183=>"111111111",
  26184=>"000000000",
  26185=>"000000000",
  26186=>"000111000",
  26187=>"011000000",
  26188=>"000000000",
  26189=>"000011001",
  26190=>"100010010",
  26191=>"111111111",
  26192=>"111011111",
  26193=>"100110000",
  26194=>"000000010",
  26195=>"111111111",
  26196=>"000000110",
  26197=>"111111111",
  26198=>"111101100",
  26199=>"000000010",
  26200=>"000011000",
  26201=>"000000000",
  26202=>"000000110",
  26203=>"111110100",
  26204=>"011111111",
  26205=>"110000000",
  26206=>"110111011",
  26207=>"001001111",
  26208=>"000000000",
  26209=>"000000001",
  26210=>"111111110",
  26211=>"000000000",
  26212=>"111111000",
  26213=>"011111111",
  26214=>"111110000",
  26215=>"000001101",
  26216=>"101001000",
  26217=>"000000010",
  26218=>"000000111",
  26219=>"111011000",
  26220=>"011111111",
  26221=>"000110111",
  26222=>"111111000",
  26223=>"000000000",
  26224=>"001111110",
  26225=>"010000000",
  26226=>"111111011",
  26227=>"111111111",
  26228=>"000000000",
  26229=>"011111111",
  26230=>"000000111",
  26231=>"000000000",
  26232=>"000000000",
  26233=>"111111111",
  26234=>"000100101",
  26235=>"000010000",
  26236=>"011011011",
  26237=>"000000000",
  26238=>"000111111",
  26239=>"001110111",
  26240=>"000011000",
  26241=>"000001011",
  26242=>"001101111",
  26243=>"000111111",
  26244=>"111111001",
  26245=>"011111011",
  26246=>"110111111",
  26247=>"101001000",
  26248=>"111111111",
  26249=>"100000111",
  26250=>"111111000",
  26251=>"111111111",
  26252=>"111110100",
  26253=>"110111111",
  26254=>"000000000",
  26255=>"001011001",
  26256=>"111111111",
  26257=>"001101100",
  26258=>"000101101",
  26259=>"000000111",
  26260=>"011001000",
  26261=>"110111111",
  26262=>"111011001",
  26263=>"111100100",
  26264=>"010111110",
  26265=>"000000000",
  26266=>"000100111",
  26267=>"111001100",
  26268=>"111111111",
  26269=>"011001000",
  26270=>"111111111",
  26271=>"011011111",
  26272=>"111111111",
  26273=>"000000110",
  26274=>"111111111",
  26275=>"001001111",
  26276=>"011001000",
  26277=>"101101111",
  26278=>"111000000",
  26279=>"101111111",
  26280=>"111010000",
  26281=>"000000000",
  26282=>"111000000",
  26283=>"000111111",
  26284=>"000011111",
  26285=>"011011001",
  26286=>"000010000",
  26287=>"111010000",
  26288=>"111111111",
  26289=>"000001101",
  26290=>"000000000",
  26291=>"111000111",
  26292=>"100000000",
  26293=>"111111111",
  26294=>"111101101",
  26295=>"111000000",
  26296=>"000000000",
  26297=>"000000000",
  26298=>"000000000",
  26299=>"011011111",
  26300=>"000000000",
  26301=>"000100000",
  26302=>"000000001",
  26303=>"000101111",
  26304=>"000100100",
  26305=>"111111111",
  26306=>"101111111",
  26307=>"111001000",
  26308=>"000000000",
  26309=>"000000000",
  26310=>"000010010",
  26311=>"111110110",
  26312=>"110100010",
  26313=>"011010000",
  26314=>"011111111",
  26315=>"101010011",
  26316=>"000000000",
  26317=>"110100000",
  26318=>"111010000",
  26319=>"101110110",
  26320=>"100000100",
  26321=>"110000000",
  26322=>"111111111",
  26323=>"111000000",
  26324=>"000000100",
  26325=>"111001000",
  26326=>"111110110",
  26327=>"000000000",
  26328=>"111111111",
  26329=>"111011000",
  26330=>"000000000",
  26331=>"111001011",
  26332=>"111111111",
  26333=>"000000111",
  26334=>"011111111",
  26335=>"000000011",
  26336=>"111111111",
  26337=>"111111111",
  26338=>"100000000",
  26339=>"111111101",
  26340=>"000101111",
  26341=>"000010010",
  26342=>"000011001",
  26343=>"111111011",
  26344=>"010000000",
  26345=>"001011000",
  26346=>"111111111",
  26347=>"000000000",
  26348=>"000000000",
  26349=>"001011011",
  26350=>"000000000",
  26351=>"001010000",
  26352=>"111000000",
  26353=>"000000000",
  26354=>"011001001",
  26355=>"111110000",
  26356=>"111111111",
  26357=>"000010111",
  26358=>"001101111",
  26359=>"000000000",
  26360=>"000000000",
  26361=>"111100100",
  26362=>"111111100",
  26363=>"100100111",
  26364=>"101111111",
  26365=>"000000000",
  26366=>"111000000",
  26367=>"100100000",
  26368=>"000000000",
  26369=>"000000000",
  26370=>"111111011",
  26371=>"000000001",
  26372=>"000011000",
  26373=>"011000000",
  26374=>"000000000",
  26375=>"000010000",
  26376=>"111001111",
  26377=>"111101001",
  26378=>"101000000",
  26379=>"111111111",
  26380=>"000000000",
  26381=>"111111111",
  26382=>"111111111",
  26383=>"100100100",
  26384=>"111111111",
  26385=>"001111111",
  26386=>"000000000",
  26387=>"111111111",
  26388=>"111111111",
  26389=>"000000111",
  26390=>"011011011",
  26391=>"000000001",
  26392=>"111110110",
  26393=>"111111111",
  26394=>"111111111",
  26395=>"100000000",
  26396=>"011111110",
  26397=>"111111101",
  26398=>"000000011",
  26399=>"000111000",
  26400=>"110111100",
  26401=>"000000000",
  26402=>"110110111",
  26403=>"111001011",
  26404=>"000001011",
  26405=>"000000000",
  26406=>"111111111",
  26407=>"011100100",
  26408=>"001100100",
  26409=>"000100111",
  26410=>"110111111",
  26411=>"110011011",
  26412=>"111111111",
  26413=>"011011001",
  26414=>"111111110",
  26415=>"010010010",
  26416=>"111011100",
  26417=>"101100000",
  26418=>"111000000",
  26419=>"111111111",
  26420=>"100110100",
  26421=>"000111111",
  26422=>"100100111",
  26423=>"001111100",
  26424=>"000000000",
  26425=>"000000111",
  26426=>"001000000",
  26427=>"110111111",
  26428=>"000000000",
  26429=>"000000000",
  26430=>"011111111",
  26431=>"000100110",
  26432=>"000000000",
  26433=>"111111111",
  26434=>"111011000",
  26435=>"000001000",
  26436=>"000000000",
  26437=>"111111111",
  26438=>"000000110",
  26439=>"110110111",
  26440=>"110111111",
  26441=>"000000000",
  26442=>"101110110",
  26443=>"100100000",
  26444=>"111011001",
  26445=>"000001011",
  26446=>"000000000",
  26447=>"100110110",
  26448=>"000000011",
  26449=>"000000111",
  26450=>"000000111",
  26451=>"111111111",
  26452=>"000000000",
  26453=>"110111111",
  26454=>"111111111",
  26455=>"111111111",
  26456=>"111111111",
  26457=>"100000000",
  26458=>"000101100",
  26459=>"010010010",
  26460=>"000011011",
  26461=>"111111111",
  26462=>"000010010",
  26463=>"000101001",
  26464=>"111111111",
  26465=>"111000000",
  26466=>"111111111",
  26467=>"111101011",
  26468=>"110100100",
  26469=>"111110010",
  26470=>"111111001",
  26471=>"000000000",
  26472=>"001000000",
  26473=>"000000000",
  26474=>"011111000",
  26475=>"111111111",
  26476=>"111001000",
  26477=>"000000000",
  26478=>"000000000",
  26479=>"001001011",
  26480=>"111111101",
  26481=>"111101111",
  26482=>"111111000",
  26483=>"011001000",
  26484=>"111100101",
  26485=>"010111111",
  26486=>"111111000",
  26487=>"111111111",
  26488=>"000000010",
  26489=>"000101111",
  26490=>"011000000",
  26491=>"111000001",
  26492=>"000101101",
  26493=>"111111111",
  26494=>"000000000",
  26495=>"000000000",
  26496=>"000000101",
  26497=>"111000000",
  26498=>"101101100",
  26499=>"000000000",
  26500=>"011011111",
  26501=>"000000000",
  26502=>"000011010",
  26503=>"100111111",
  26504=>"000000000",
  26505=>"001000001",
  26506=>"100000001",
  26507=>"111101111",
  26508=>"001001001",
  26509=>"011000000",
  26510=>"100110100",
  26511=>"000000000",
  26512=>"111111110",
  26513=>"101111111",
  26514=>"111111111",
  26515=>"001000000",
  26516=>"000000101",
  26517=>"111110100",
  26518=>"000100100",
  26519=>"000000000",
  26520=>"000111111",
  26521=>"100000000",
  26522=>"000000000",
  26523=>"000111111",
  26524=>"111011001",
  26525=>"111011011",
  26526=>"000000111",
  26527=>"000000000",
  26528=>"111100110",
  26529=>"111111111",
  26530=>"010000000",
  26531=>"111001111",
  26532=>"000000000",
  26533=>"111111101",
  26534=>"000000000",
  26535=>"111101101",
  26536=>"111100000",
  26537=>"111100100",
  26538=>"000111111",
  26539=>"001010010",
  26540=>"111000111",
  26541=>"111101010",
  26542=>"111111111",
  26543=>"111111111",
  26544=>"000000000",
  26545=>"111100000",
  26546=>"001000000",
  26547=>"111111111",
  26548=>"111111110",
  26549=>"111111011",
  26550=>"000000000",
  26551=>"111111111",
  26552=>"000010010",
  26553=>"100000000",
  26554=>"101100100",
  26555=>"100110110",
  26556=>"000000000",
  26557=>"111111111",
  26558=>"111111111",
  26559=>"001011010",
  26560=>"100110110",
  26561=>"011111110",
  26562=>"000000000",
  26563=>"000000000",
  26564=>"111111000",
  26565=>"001000010",
  26566=>"011011001",
  26567=>"110100100",
  26568=>"000000000",
  26569=>"000000111",
  26570=>"111111111",
  26571=>"110111010",
  26572=>"000000001",
  26573=>"000001001",
  26574=>"010000110",
  26575=>"011111111",
  26576=>"111111111",
  26577=>"110111111",
  26578=>"011011001",
  26579=>"111111111",
  26580=>"100110110",
  26581=>"100100000",
  26582=>"100000000",
  26583=>"001001000",
  26584=>"011110110",
  26585=>"111110000",
  26586=>"111100101",
  26587=>"011010010",
  26588=>"010000000",
  26589=>"111111111",
  26590=>"000000000",
  26591=>"011000010",
  26592=>"000000010",
  26593=>"000010000",
  26594=>"110111111",
  26595=>"000000000",
  26596=>"000000000",
  26597=>"000000101",
  26598=>"000110011",
  26599=>"101001111",
  26600=>"111111111",
  26601=>"000001001",
  26602=>"011000011",
  26603=>"110110111",
  26604=>"011011000",
  26605=>"000000111",
  26606=>"111111111",
  26607=>"000000000",
  26608=>"011000000",
  26609=>"000000110",
  26610=>"000000000",
  26611=>"111000000",
  26612=>"000000000",
  26613=>"100100111",
  26614=>"000000000",
  26615=>"000000010",
  26616=>"001000000",
  26617=>"000100110",
  26618=>"111111011",
  26619=>"110111000",
  26620=>"000000111",
  26621=>"001111111",
  26622=>"000000011",
  26623=>"000000000",
  26624=>"010110110",
  26625=>"111111111",
  26626=>"111111111",
  26627=>"001011000",
  26628=>"000000000",
  26629=>"011011110",
  26630=>"100001001",
  26631=>"000000000",
  26632=>"101111011",
  26633=>"011011001",
  26634=>"111111111",
  26635=>"100000000",
  26636=>"000011011",
  26637=>"000001001",
  26638=>"110100000",
  26639=>"111111111",
  26640=>"111001000",
  26641=>"000000000",
  26642=>"011111111",
  26643=>"111011101",
  26644=>"111101000",
  26645=>"011111111",
  26646=>"111101111",
  26647=>"000000000",
  26648=>"000000000",
  26649=>"000000011",
  26650=>"000111001",
  26651=>"000111001",
  26652=>"001001000",
  26653=>"110110110",
  26654=>"000000011",
  26655=>"000001011",
  26656=>"101101111",
  26657=>"000000000",
  26658=>"110010110",
  26659=>"111110111",
  26660=>"111111111",
  26661=>"111001000",
  26662=>"000000000",
  26663=>"000111111",
  26664=>"111111101",
  26665=>"011011011",
  26666=>"000000000",
  26667=>"111000000",
  26668=>"000000000",
  26669=>"111100000",
  26670=>"110111111",
  26671=>"000000000",
  26672=>"111001001",
  26673=>"000000000",
  26674=>"000100001",
  26675=>"000001000",
  26676=>"001001000",
  26677=>"000011000",
  26678=>"000101111",
  26679=>"110111101",
  26680=>"111111111",
  26681=>"111111111",
  26682=>"100000111",
  26683=>"000000000",
  26684=>"101101100",
  26685=>"000011011",
  26686=>"001001101",
  26687=>"111111111",
  26688=>"001111111",
  26689=>"101111111",
  26690=>"111000000",
  26691=>"000001000",
  26692=>"010011011",
  26693=>"111011001",
  26694=>"011000000",
  26695=>"000000000",
  26696=>"001011010",
  26697=>"001110111",
  26698=>"111111111",
  26699=>"110111111",
  26700=>"101100111",
  26701=>"001101000",
  26702=>"111011111",
  26703=>"111011011",
  26704=>"111001011",
  26705=>"000000000",
  26706=>"111111111",
  26707=>"111110000",
  26708=>"000000000",
  26709=>"000000000",
  26710=>"011000001",
  26711=>"111111110",
  26712=>"111111001",
  26713=>"111111000",
  26714=>"101100000",
  26715=>"001100111",
  26716=>"000011000",
  26717=>"111111111",
  26718=>"111111111",
  26719=>"000000111",
  26720=>"100000000",
  26721=>"011011001",
  26722=>"111111111",
  26723=>"000000000",
  26724=>"111101001",
  26725=>"100111111",
  26726=>"111111111",
  26727=>"111111110",
  26728=>"000001010",
  26729=>"000100100",
  26730=>"100000000",
  26731=>"111111111",
  26732=>"000000000",
  26733=>"000000011",
  26734=>"000000000",
  26735=>"111111111",
  26736=>"001111000",
  26737=>"111111111",
  26738=>"001111111",
  26739=>"000000000",
  26740=>"111111111",
  26741=>"000000101",
  26742=>"000111111",
  26743=>"111001000",
  26744=>"110000000",
  26745=>"000011011",
  26746=>"000000000",
  26747=>"011111110",
  26748=>"000000000",
  26749=>"101111111",
  26750=>"000000000",
  26751=>"011111100",
  26752=>"111111111",
  26753=>"111111101",
  26754=>"000000000",
  26755=>"111110000",
  26756=>"111111111",
  26757=>"000000111",
  26758=>"000000000",
  26759=>"000011111",
  26760=>"000000101",
  26761=>"111000001",
  26762=>"111110000",
  26763=>"000000000",
  26764=>"000000000",
  26765=>"111111111",
  26766=>"000001111",
  26767=>"010111110",
  26768=>"001000000",
  26769=>"111111000",
  26770=>"111111111",
  26771=>"010011000",
  26772=>"111111001",
  26773=>"001001011",
  26774=>"100000111",
  26775=>"000000000",
  26776=>"011111101",
  26777=>"111111011",
  26778=>"000000000",
  26779=>"111111111",
  26780=>"000000111",
  26781=>"000000000",
  26782=>"001101100",
  26783=>"111111111",
  26784=>"111100101",
  26785=>"000000100",
  26786=>"010110000",
  26787=>"000000000",
  26788=>"110110111",
  26789=>"000001001",
  26790=>"111111111",
  26791=>"000111001",
  26792=>"110110011",
  26793=>"000000000",
  26794=>"000000111",
  26795=>"100101101",
  26796=>"101001100",
  26797=>"000000000",
  26798=>"111111111",
  26799=>"100100001",
  26800=>"111111111",
  26801=>"100100100",
  26802=>"111111001",
  26803=>"000000000",
  26804=>"000001111",
  26805=>"111100000",
  26806=>"011111111",
  26807=>"101110111",
  26808=>"000000001",
  26809=>"000000101",
  26810=>"111100001",
  26811=>"000000111",
  26812=>"111111000",
  26813=>"101111111",
  26814=>"101000100",
  26815=>"010000001",
  26816=>"000000100",
  26817=>"000000000",
  26818=>"011000101",
  26819=>"111111111",
  26820=>"000000000",
  26821=>"111111111",
  26822=>"111111111",
  26823=>"110010000",
  26824=>"111111001",
  26825=>"001000101",
  26826=>"111011011",
  26827=>"111000000",
  26828=>"001001101",
  26829=>"111110111",
  26830=>"000000001",
  26831=>"000100111",
  26832=>"000000000",
  26833=>"111111111",
  26834=>"010000111",
  26835=>"000000100",
  26836=>"111111000",
  26837=>"011011110",
  26838=>"000000000",
  26839=>"000000001",
  26840=>"000000000",
  26841=>"111111101",
  26842=>"111100111",
  26843=>"000000111",
  26844=>"000000101",
  26845=>"000000101",
  26846=>"111111011",
  26847=>"111111111",
  26848=>"111111111",
  26849=>"100100110",
  26850=>"010110000",
  26851=>"000111111",
  26852=>"000000000",
  26853=>"000000111",
  26854=>"000111011",
  26855=>"111001000",
  26856=>"111010110",
  26857=>"000000000",
  26858=>"100000100",
  26859=>"111111111",
  26860=>"000000111",
  26861=>"111111111",
  26862=>"111111111",
  26863=>"001001101",
  26864=>"110100100",
  26865=>"000000000",
  26866=>"111000100",
  26867=>"111101111",
  26868=>"000100111",
  26869=>"000000100",
  26870=>"000010000",
  26871=>"111111111",
  26872=>"000000111",
  26873=>"001001011",
  26874=>"111111111",
  26875=>"100110110",
  26876=>"111111111",
  26877=>"111000000",
  26878=>"001001000",
  26879=>"000100000",
  26880=>"111111001",
  26881=>"011111111",
  26882=>"000011111",
  26883=>"000000010",
  26884=>"111111111",
  26885=>"111111111",
  26886=>"111101111",
  26887=>"000000111",
  26888=>"000000000",
  26889=>"100000000",
  26890=>"111111111",
  26891=>"000101011",
  26892=>"000011111",
  26893=>"011110111",
  26894=>"111111111",
  26895=>"100100000",
  26896=>"110000000",
  26897=>"111000000",
  26898=>"111111111",
  26899=>"001000000",
  26900=>"000100100",
  26901=>"111111010",
  26902=>"011111101",
  26903=>"000000000",
  26904=>"000000000",
  26905=>"101000000",
  26906=>"111111001",
  26907=>"111111111",
  26908=>"011011011",
  26909=>"011011111",
  26910=>"111111111",
  26911=>"001011011",
  26912=>"000000000",
  26913=>"100100000",
  26914=>"111111111",
  26915=>"011011001",
  26916=>"100010000",
  26917=>"111111111",
  26918=>"000111111",
  26919=>"011111011",
  26920=>"011001011",
  26921=>"100100110",
  26922=>"111001001",
  26923=>"000100010",
  26924=>"000000000",
  26925=>"010000000",
  26926=>"101000111",
  26927=>"101101111",
  26928=>"111111111",
  26929=>"000000000",
  26930=>"111111110",
  26931=>"000000010",
  26932=>"000000111",
  26933=>"001111111",
  26934=>"000000000",
  26935=>"001011001",
  26936=>"111111111",
  26937=>"111101000",
  26938=>"000000000",
  26939=>"000000110",
  26940=>"111111111",
  26941=>"000000000",
  26942=>"101001101",
  26943=>"000000000",
  26944=>"111111111",
  26945=>"000000101",
  26946=>"000000000",
  26947=>"111111111",
  26948=>"110100000",
  26949=>"111111111",
  26950=>"000000000",
  26951=>"110111110",
  26952=>"111111111",
  26953=>"111111101",
  26954=>"111111001",
  26955=>"111001111",
  26956=>"101100111",
  26957=>"011001011",
  26958=>"000000001",
  26959=>"000000111",
  26960=>"000110000",
  26961=>"000000000",
  26962=>"001000000",
  26963=>"111111111",
  26964=>"000000000",
  26965=>"011010011",
  26966=>"000000011",
  26967=>"111111111",
  26968=>"000000000",
  26969=>"111111111",
  26970=>"111111011",
  26971=>"111111101",
  26972=>"001001000",
  26973=>"000000000",
  26974=>"011111111",
  26975=>"010000000",
  26976=>"110000000",
  26977=>"111111001",
  26978=>"010000010",
  26979=>"000000000",
  26980=>"000000000",
  26981=>"001001001",
  26982=>"011111111",
  26983=>"000000000",
  26984=>"111111111",
  26985=>"000000000",
  26986=>"000100100",
  26987=>"000000111",
  26988=>"000011010",
  26989=>"111111111",
  26990=>"000000000",
  26991=>"101000100",
  26992=>"000000011",
  26993=>"111111111",
  26994=>"111111111",
  26995=>"111000000",
  26996=>"111111111",
  26997=>"000000101",
  26998=>"111111011",
  26999=>"000000000",
  27000=>"100100111",
  27001=>"000000000",
  27002=>"111111111",
  27003=>"101111001",
  27004=>"000000110",
  27005=>"000000000",
  27006=>"111111110",
  27007=>"111111111",
  27008=>"111111111",
  27009=>"100111111",
  27010=>"111010000",
  27011=>"111111111",
  27012=>"000010010",
  27013=>"000100111",
  27014=>"111100111",
  27015=>"111111111",
  27016=>"000000111",
  27017=>"000000000",
  27018=>"000000000",
  27019=>"000000000",
  27020=>"111111111",
  27021=>"000000000",
  27022=>"111100000",
  27023=>"000011111",
  27024=>"000011000",
  27025=>"000000100",
  27026=>"000000000",
  27027=>"111111111",
  27028=>"000000000",
  27029=>"111111111",
  27030=>"111111111",
  27031=>"011010011",
  27032=>"000000000",
  27033=>"100111101",
  27034=>"000000010",
  27035=>"011001111",
  27036=>"111111100",
  27037=>"111111000",
  27038=>"111111111",
  27039=>"010111000",
  27040=>"111111111",
  27041=>"000000000",
  27042=>"100100000",
  27043=>"010010000",
  27044=>"111100000",
  27045=>"000000000",
  27046=>"001111110",
  27047=>"111111111",
  27048=>"111111111",
  27049=>"000000000",
  27050=>"000000000",
  27051=>"111111111",
  27052=>"100110010",
  27053=>"010000101",
  27054=>"000000000",
  27055=>"000000000",
  27056=>"001000100",
  27057=>"000000010",
  27058=>"000000001",
  27059=>"000000000",
  27060=>"100000011",
  27061=>"111101001",
  27062=>"111101000",
  27063=>"101001000",
  27064=>"111111000",
  27065=>"111011011",
  27066=>"010000000",
  27067=>"000000000",
  27068=>"111111111",
  27069=>"000000000",
  27070=>"111011001",
  27071=>"000111011",
  27072=>"111111111",
  27073=>"110111111",
  27074=>"000000000",
  27075=>"111111111",
  27076=>"001100100",
  27077=>"111110111",
  27078=>"000000011",
  27079=>"000000000",
  27080=>"011001000",
  27081=>"001100100",
  27082=>"001011011",
  27083=>"100100111",
  27084=>"000000000",
  27085=>"110000000",
  27086=>"100110101",
  27087=>"000000000",
  27088=>"000000111",
  27089=>"000010111",
  27090=>"001000000",
  27091=>"111111011",
  27092=>"110100001",
  27093=>"110100000",
  27094=>"110100001",
  27095=>"011110100",
  27096=>"111111011",
  27097=>"000000000",
  27098=>"111111111",
  27099=>"111111111",
  27100=>"100000000",
  27101=>"101000111",
  27102=>"100001111",
  27103=>"000111111",
  27104=>"001100101",
  27105=>"000011111",
  27106=>"111111000",
  27107=>"001000001",
  27108=>"111001111",
  27109=>"001111010",
  27110=>"111000000",
  27111=>"000000000",
  27112=>"000000000",
  27113=>"111011001",
  27114=>"111111101",
  27115=>"000111101",
  27116=>"100000100",
  27117=>"000010010",
  27118=>"001111001",
  27119=>"111111101",
  27120=>"111011001",
  27121=>"000000000",
  27122=>"000001001",
  27123=>"001100100",
  27124=>"110110100",
  27125=>"000000000",
  27126=>"001000001",
  27127=>"111111011",
  27128=>"000100111",
  27129=>"000000000",
  27130=>"000000000",
  27131=>"000000000",
  27132=>"111101000",
  27133=>"000001000",
  27134=>"000111001",
  27135=>"101000000",
  27136=>"110100110",
  27137=>"111111001",
  27138=>"000000000",
  27139=>"111111111",
  27140=>"100000000",
  27141=>"111000000",
  27142=>"000000001",
  27143=>"111111111",
  27144=>"001001011",
  27145=>"000000000",
  27146=>"000000000",
  27147=>"111110111",
  27148=>"001111111",
  27149=>"111111111",
  27150=>"111111000",
  27151=>"111111100",
  27152=>"000000001",
  27153=>"000000011",
  27154=>"110100110",
  27155=>"000000101",
  27156=>"111011001",
  27157=>"001001001",
  27158=>"000000001",
  27159=>"001001011",
  27160=>"110110100",
  27161=>"101110111",
  27162=>"101101111",
  27163=>"111010000",
  27164=>"000000011",
  27165=>"100001111",
  27166=>"110111111",
  27167=>"011011011",
  27168=>"110110000",
  27169=>"110110110",
  27170=>"111111111",
  27171=>"001001111",
  27172=>"101100111",
  27173=>"111111011",
  27174=>"000000000",
  27175=>"110111111",
  27176=>"000000000",
  27177=>"000000000",
  27178=>"010010111",
  27179=>"100000111",
  27180=>"111001111",
  27181=>"000101111",
  27182=>"111111011",
  27183=>"110111111",
  27184=>"100000000",
  27185=>"111111110",
  27186=>"111011011",
  27187=>"010010000",
  27188=>"000011000",
  27189=>"111111100",
  27190=>"000000000",
  27191=>"111100000",
  27192=>"010110000",
  27193=>"111111111",
  27194=>"000000000",
  27195=>"000000000",
  27196=>"000111111",
  27197=>"100100100",
  27198=>"000000000",
  27199=>"111111111",
  27200=>"101000001",
  27201=>"010010001",
  27202=>"111111111",
  27203=>"100100000",
  27204=>"111011000",
  27205=>"000100110",
  27206=>"111111110",
  27207=>"111111111",
  27208=>"100100011",
  27209=>"000000000",
  27210=>"111111111",
  27211=>"111111111",
  27212=>"000000001",
  27213=>"111111010",
  27214=>"100000000",
  27215=>"000000000",
  27216=>"011111111",
  27217=>"011111111",
  27218=>"100000000",
  27219=>"100111011",
  27220=>"000000000",
  27221=>"011001001",
  27222=>"111110110",
  27223=>"110111111",
  27224=>"010000111",
  27225=>"111111111",
  27226=>"111111101",
  27227=>"100110000",
  27228=>"111011000",
  27229=>"100111111",
  27230=>"000000000",
  27231=>"001001011",
  27232=>"000000000",
  27233=>"000000001",
  27234=>"000000000",
  27235=>"010000000",
  27236=>"111000000",
  27237=>"000000110",
  27238=>"001101111",
  27239=>"111010000",
  27240=>"001011111",
  27241=>"001000000",
  27242=>"010011011",
  27243=>"000000000",
  27244=>"000000100",
  27245=>"111111111",
  27246=>"100101111",
  27247=>"000000000",
  27248=>"111111011",
  27249=>"000001111",
  27250=>"000001001",
  27251=>"111111111",
  27252=>"000000000",
  27253=>"111111111",
  27254=>"000001111",
  27255=>"000000000",
  27256=>"000000100",
  27257=>"111011111",
  27258=>"011001001",
  27259=>"000000000",
  27260=>"111111111",
  27261=>"111100110",
  27262=>"111111110",
  27263=>"010010011",
  27264=>"000000100",
  27265=>"110000000",
  27266=>"000000000",
  27267=>"111111111",
  27268=>"111111011",
  27269=>"110000111",
  27270=>"111111011",
  27271=>"111111111",
  27272=>"000000000",
  27273=>"111001000",
  27274=>"001111111",
  27275=>"011011011",
  27276=>"000000011",
  27277=>"001000111",
  27278=>"000000111",
  27279=>"000000011",
  27280=>"000001101",
  27281=>"000000000",
  27282=>"000000000",
  27283=>"111111100",
  27284=>"000010000",
  27285=>"111111111",
  27286=>"000000111",
  27287=>"000000000",
  27288=>"000000010",
  27289=>"111111111",
  27290=>"000000000",
  27291=>"000000000",
  27292=>"111111111",
  27293=>"100100000",
  27294=>"111111111",
  27295=>"000000000",
  27296=>"000000011",
  27297=>"010000000",
  27298=>"000110111",
  27299=>"000000000",
  27300=>"110111111",
  27301=>"101001000",
  27302=>"111111111",
  27303=>"111111111",
  27304=>"000000000",
  27305=>"111100100",
  27306=>"000010000",
  27307=>"111100111",
  27308=>"000000001",
  27309=>"000010110",
  27310=>"111111111",
  27311=>"001001000",
  27312=>"000011111",
  27313=>"111110100",
  27314=>"010111010",
  27315=>"011110000",
  27316=>"111110010",
  27317=>"111111111",
  27318=>"111111111",
  27319=>"000000100",
  27320=>"000000100",
  27321=>"000000100",
  27322=>"000000000",
  27323=>"110010000",
  27324=>"111111000",
  27325=>"111111111",
  27326=>"111000110",
  27327=>"000100111",
  27328=>"000000000",
  27329=>"100110111",
  27330=>"000100100",
  27331=>"111111011",
  27332=>"011001000",
  27333=>"000000000",
  27334=>"000001001",
  27335=>"111100000",
  27336=>"100101101",
  27337=>"000000001",
  27338=>"011110100",
  27339=>"111111111",
  27340=>"110110110",
  27341=>"000000000",
  27342=>"000000000",
  27343=>"000000000",
  27344=>"011000000",
  27345=>"001000000",
  27346=>"000110111",
  27347=>"000000000",
  27348=>"000000100",
  27349=>"000000010",
  27350=>"110000000",
  27351=>"010100000",
  27352=>"111111111",
  27353=>"011011111",
  27354=>"000000000",
  27355=>"111111111",
  27356=>"001011011",
  27357=>"110110111",
  27358=>"010011000",
  27359=>"000000000",
  27360=>"001011111",
  27361=>"000000000",
  27362=>"111111111",
  27363=>"111111111",
  27364=>"011111101",
  27365=>"000000000",
  27366=>"111111111",
  27367=>"111111111",
  27368=>"111111111",
  27369=>"111111111",
  27370=>"000010111",
  27371=>"111111001",
  27372=>"000111101",
  27373=>"000000111",
  27374=>"000000000",
  27375=>"000000000",
  27376=>"000000001",
  27377=>"000000000",
  27378=>"111100000",
  27379=>"110111111",
  27380=>"111111011",
  27381=>"111100100",
  27382=>"111100001",
  27383=>"000000000",
  27384=>"111111111",
  27385=>"000000000",
  27386=>"111111001",
  27387=>"000000000",
  27388=>"110100100",
  27389=>"000100110",
  27390=>"110000000",
  27391=>"101111111",
  27392=>"000010011",
  27393=>"101001000",
  27394=>"111111111",
  27395=>"000000000",
  27396=>"111000000",
  27397=>"000000000",
  27398=>"111000111",
  27399=>"111111111",
  27400=>"000100111",
  27401=>"110000000",
  27402=>"000000000",
  27403=>"000000001",
  27404=>"000000000",
  27405=>"001001001",
  27406=>"000010010",
  27407=>"000000000",
  27408=>"111001000",
  27409=>"000010000",
  27410=>"000000111",
  27411=>"000000000",
  27412=>"011010000",
  27413=>"111101111",
  27414=>"111111111",
  27415=>"100010000",
  27416=>"000000001",
  27417=>"011111111",
  27418=>"011001000",
  27419=>"000110100",
  27420=>"111111100",
  27421=>"000111111",
  27422=>"011111110",
  27423=>"010000100",
  27424=>"101011111",
  27425=>"000000000",
  27426=>"111111111",
  27427=>"000000000",
  27428=>"111111111",
  27429=>"000000000",
  27430=>"000111000",
  27431=>"011011111",
  27432=>"111000000",
  27433=>"000110111",
  27434=>"001000000",
  27435=>"111011111",
  27436=>"101110100",
  27437=>"000000000",
  27438=>"010000111",
  27439=>"000000000",
  27440=>"111111111",
  27441=>"000111111",
  27442=>"000001001",
  27443=>"011000000",
  27444=>"010000010",
  27445=>"101110111",
  27446=>"000011001",
  27447=>"111111011",
  27448=>"111111111",
  27449=>"000000011",
  27450=>"111111111",
  27451=>"111111111",
  27452=>"000000000",
  27453=>"000100101",
  27454=>"000000000",
  27455=>"000000000",
  27456=>"000000000",
  27457=>"111111111",
  27458=>"010000110",
  27459=>"000000000",
  27460=>"000000000",
  27461=>"011000000",
  27462=>"111101111",
  27463=>"111101111",
  27464=>"111111111",
  27465=>"000000010",
  27466=>"111111111",
  27467=>"011011111",
  27468=>"100100100",
  27469=>"000000000",
  27470=>"000000000",
  27471=>"000000100",
  27472=>"000011111",
  27473=>"111111111",
  27474=>"100111111",
  27475=>"111111011",
  27476=>"000001111",
  27477=>"011011011",
  27478=>"110110111",
  27479=>"111111111",
  27480=>"111111111",
  27481=>"011111111",
  27482=>"111000111",
  27483=>"001100000",
  27484=>"000000000",
  27485=>"111111100",
  27486=>"000011111",
  27487=>"111111111",
  27488=>"000100111",
  27489=>"111111001",
  27490=>"111111111",
  27491=>"001000000",
  27492=>"110011000",
  27493=>"000000000",
  27494=>"000000100",
  27495=>"100110010",
  27496=>"110110110",
  27497=>"111111111",
  27498=>"000000111",
  27499=>"000000000",
  27500=>"011101101",
  27501=>"010111111",
  27502=>"010111111",
  27503=>"000000000",
  27504=>"000000000",
  27505=>"000101111",
  27506=>"010111110",
  27507=>"000100100",
  27508=>"110111111",
  27509=>"000000000",
  27510=>"000011001",
  27511=>"101010000",
  27512=>"111101111",
  27513=>"111111110",
  27514=>"111001001",
  27515=>"100111111",
  27516=>"001111111",
  27517=>"000000000",
  27518=>"000000000",
  27519=>"000111111",
  27520=>"000000010",
  27521=>"000000000",
  27522=>"101100111",
  27523=>"001111111",
  27524=>"111111001",
  27525=>"111111011",
  27526=>"101110111",
  27527=>"111111111",
  27528=>"001000101",
  27529=>"000000011",
  27530=>"000000000",
  27531=>"110111000",
  27532=>"000000001",
  27533=>"000000100",
  27534=>"110111111",
  27535=>"010000000",
  27536=>"111111111",
  27537=>"111011111",
  27538=>"111111111",
  27539=>"000100111",
  27540=>"000000000",
  27541=>"010010000",
  27542=>"010110111",
  27543=>"100100000",
  27544=>"111110000",
  27545=>"000000000",
  27546=>"100110111",
  27547=>"110111111",
  27548=>"000000000",
  27549=>"000000100",
  27550=>"000000100",
  27551=>"100111111",
  27552=>"000000000",
  27553=>"000001001",
  27554=>"000000000",
  27555=>"001011011",
  27556=>"111111111",
  27557=>"111111111",
  27558=>"111111111",
  27559=>"101111111",
  27560=>"010010000",
  27561=>"111000000",
  27562=>"000001000",
  27563=>"110110000",
  27564=>"000000000",
  27565=>"111110111",
  27566=>"000001101",
  27567=>"111111011",
  27568=>"111001111",
  27569=>"000010010",
  27570=>"000010011",
  27571=>"000000001",
  27572=>"001001101",
  27573=>"110100001",
  27574=>"000000001",
  27575=>"000000000",
  27576=>"011000000",
  27577=>"101110111",
  27578=>"000000101",
  27579=>"000000000",
  27580=>"111111111",
  27581=>"111000000",
  27582=>"011011000",
  27583=>"100000001",
  27584=>"111111100",
  27585=>"111111111",
  27586=>"111111111",
  27587=>"011111111",
  27588=>"111111001",
  27589=>"111111011",
  27590=>"000010001",
  27591=>"000000000",
  27592=>"000111111",
  27593=>"000000000",
  27594=>"000000000",
  27595=>"100000010",
  27596=>"111111110",
  27597=>"110100000",
  27598=>"101100000",
  27599=>"111111101",
  27600=>"110111011",
  27601=>"001101100",
  27602=>"000001000",
  27603=>"000000001",
  27604=>"000000000",
  27605=>"000000000",
  27606=>"110110000",
  27607=>"000111111",
  27608=>"011111000",
  27609=>"111111111",
  27610=>"100100111",
  27611=>"110111111",
  27612=>"011011111",
  27613=>"000100001",
  27614=>"100110000",
  27615=>"110100100",
  27616=>"101101100",
  27617=>"110100000",
  27618=>"111111011",
  27619=>"111111111",
  27620=>"011000000",
  27621=>"000111111",
  27622=>"001011011",
  27623=>"000000000",
  27624=>"000000000",
  27625=>"101001000",
  27626=>"000000000",
  27627=>"000000000",
  27628=>"110111110",
  27629=>"010011001",
  27630=>"111111111",
  27631=>"111111100",
  27632=>"010000000",
  27633=>"000000000",
  27634=>"111111011",
  27635=>"111111011",
  27636=>"011011111",
  27637=>"000101111",
  27638=>"000000000",
  27639=>"000000110",
  27640=>"000110111",
  27641=>"110110110",
  27642=>"111010110",
  27643=>"001001000",
  27644=>"011001001",
  27645=>"001001001",
  27646=>"001000110",
  27647=>"000000000",
  27648=>"000000000",
  27649=>"111011111",
  27650=>"001101111",
  27651=>"110111111",
  27652=>"110111000",
  27653=>"000000001",
  27654=>"111111111",
  27655=>"101000000",
  27656=>"111111111",
  27657=>"000100000",
  27658=>"111100101",
  27659=>"111111111",
  27660=>"100100100",
  27661=>"000000000",
  27662=>"100000011",
  27663=>"111000111",
  27664=>"000000000",
  27665=>"111110000",
  27666=>"110000000",
  27667=>"111111111",
  27668=>"000111111",
  27669=>"000000011",
  27670=>"111111111",
  27671=>"000000111",
  27672=>"111111111",
  27673=>"011011111",
  27674=>"000000000",
  27675=>"001101110",
  27676=>"100000110",
  27677=>"000100111",
  27678=>"010000000",
  27679=>"111111111",
  27680=>"111100101",
  27681=>"111111000",
  27682=>"111011101",
  27683=>"111111111",
  27684=>"000000010",
  27685=>"110111111",
  27686=>"111100100",
  27687=>"011001000",
  27688=>"000000110",
  27689=>"000000000",
  27690=>"001101111",
  27691=>"111100101",
  27692=>"000000110",
  27693=>"011111100",
  27694=>"001111001",
  27695=>"111111111",
  27696=>"111111011",
  27697=>"000000000",
  27698=>"100100100",
  27699=>"011111111",
  27700=>"000001000",
  27701=>"110100000",
  27702=>"111100001",
  27703=>"111111110",
  27704=>"000001111",
  27705=>"001001111",
  27706=>"000000000",
  27707=>"000010111",
  27708=>"111000000",
  27709=>"111000000",
  27710=>"001011100",
  27711=>"111111111",
  27712=>"111000000",
  27713=>"111111111",
  27714=>"000000000",
  27715=>"001000000",
  27716=>"000010000",
  27717=>"001001001",
  27718=>"110110110",
  27719=>"111111111",
  27720=>"011111011",
  27721=>"001001000",
  27722=>"111001000",
  27723=>"101001101",
  27724=>"001001000",
  27725=>"100111111",
  27726=>"000001000",
  27727=>"000000000",
  27728=>"111001111",
  27729=>"111111010",
  27730=>"111110111",
  27731=>"110000000",
  27732=>"001111111",
  27733=>"000000000",
  27734=>"111000000",
  27735=>"111111111",
  27736=>"000000000",
  27737=>"001000000",
  27738=>"001010100",
  27739=>"110111111",
  27740=>"111001111",
  27741=>"111111111",
  27742=>"110111111",
  27743=>"010110110",
  27744=>"000000000",
  27745=>"000000000",
  27746=>"000000001",
  27747=>"110111010",
  27748=>"000000000",
  27749=>"000000000",
  27750=>"000111111",
  27751=>"010011000",
  27752=>"000100100",
  27753=>"001001001",
  27754=>"000000000",
  27755=>"011111111",
  27756=>"000010011",
  27757=>"111111111",
  27758=>"000000000",
  27759=>"000000010",
  27760=>"011011111",
  27761=>"000001110",
  27762=>"011010000",
  27763=>"000000000",
  27764=>"000111111",
  27765=>"110010000",
  27766=>"111111111",
  27767=>"111111000",
  27768=>"111011001",
  27769=>"101111111",
  27770=>"000000000",
  27771=>"000000000",
  27772=>"010110110",
  27773=>"011000001",
  27774=>"000000000",
  27775=>"000000000",
  27776=>"111111111",
  27777=>"001111111",
  27778=>"000000000",
  27779=>"010001011",
  27780=>"001001111",
  27781=>"000000000",
  27782=>"111111110",
  27783=>"000010011",
  27784=>"000100000",
  27785=>"111000001",
  27786=>"111111000",
  27787=>"100100010",
  27788=>"000000110",
  27789=>"111011111",
  27790=>"100001000",
  27791=>"101111111",
  27792=>"000001011",
  27793=>"111111111",
  27794=>"000000110",
  27795=>"111111001",
  27796=>"000000000",
  27797=>"111111111",
  27798=>"000000000",
  27799=>"001101100",
  27800=>"111100110",
  27801=>"000001001",
  27802=>"111111111",
  27803=>"111111111",
  27804=>"000000000",
  27805=>"111001001",
  27806=>"111111101",
  27807=>"100000000",
  27808=>"100100111",
  27809=>"111100000",
  27810=>"111110110",
  27811=>"111111111",
  27812=>"000000000",
  27813=>"100000000",
  27814=>"011001101",
  27815=>"010011000",
  27816=>"111111111",
  27817=>"000000000",
  27818=>"000000000",
  27819=>"000000000",
  27820=>"000011010",
  27821=>"110110110",
  27822=>"000111111",
  27823=>"000011111",
  27824=>"111110110",
  27825=>"011111001",
  27826=>"111111110",
  27827=>"000000000",
  27828=>"111111111",
  27829=>"000110100",
  27830=>"111111111",
  27831=>"111111010",
  27832=>"010011100",
  27833=>"100000111",
  27834=>"000000000",
  27835=>"000000100",
  27836=>"011111111",
  27837=>"111111110",
  27838=>"100000100",
  27839=>"001001111",
  27840=>"000000000",
  27841=>"001001001",
  27842=>"111000000",
  27843=>"000100000",
  27844=>"001111011",
  27845=>"011011000",
  27846=>"101101000",
  27847=>"001111100",
  27848=>"111111011",
  27849=>"110111111",
  27850=>"010111011",
  27851=>"010010000",
  27852=>"110110110",
  27853=>"001011000",
  27854=>"111111111",
  27855=>"000010111",
  27856=>"011000000",
  27857=>"111010010",
  27858=>"111111111",
  27859=>"100001101",
  27860=>"000000000",
  27861=>"111011000",
  27862=>"111110000",
  27863=>"000000000",
  27864=>"100100100",
  27865=>"000001001",
  27866=>"000010110",
  27867=>"000000111",
  27868=>"111001000",
  27869=>"000100111",
  27870=>"000000100",
  27871=>"011001000",
  27872=>"001111111",
  27873=>"111001111",
  27874=>"000000100",
  27875=>"000000101",
  27876=>"101110111",
  27877=>"111001100",
  27878=>"111111111",
  27879=>"000001100",
  27880=>"000000000",
  27881=>"000000101",
  27882=>"000000111",
  27883=>"101001100",
  27884=>"111111000",
  27885=>"000000000",
  27886=>"111101000",
  27887=>"110000000",
  27888=>"111111000",
  27889=>"110000110",
  27890=>"000000000",
  27891=>"101101101",
  27892=>"110000000",
  27893=>"010111111",
  27894=>"000000010",
  27895=>"111011111",
  27896=>"100110111",
  27897=>"000000000",
  27898=>"000100111",
  27899=>"011000000",
  27900=>"000110111",
  27901=>"000000100",
  27902=>"111010111",
  27903=>"000000000",
  27904=>"000100101",
  27905=>"001011110",
  27906=>"000000000",
  27907=>"100000110",
  27908=>"111111111",
  27909=>"010000000",
  27910=>"001000000",
  27911=>"111001111",
  27912=>"111111101",
  27913=>"111111000",
  27914=>"000000000",
  27915=>"001111111",
  27916=>"111110000",
  27917=>"110111111",
  27918=>"000000000",
  27919=>"101001000",
  27920=>"111111111",
  27921=>"000000000",
  27922=>"000000000",
  27923=>"011000001",
  27924=>"000001001",
  27925=>"111000000",
  27926=>"100110100",
  27927=>"000000111",
  27928=>"110110100",
  27929=>"111111111",
  27930=>"000000000",
  27931=>"000000000",
  27932=>"111111111",
  27933=>"001001011",
  27934=>"000000001",
  27935=>"000011111",
  27936=>"000000011",
  27937=>"011011000",
  27938=>"000000000",
  27939=>"111011011",
  27940=>"010111111",
  27941=>"111111110",
  27942=>"000000000",
  27943=>"101001111",
  27944=>"000000000",
  27945=>"000000000",
  27946=>"000001111",
  27947=>"111001111",
  27948=>"010011111",
  27949=>"000000110",
  27950=>"000000000",
  27951=>"111111000",
  27952=>"000000000",
  27953=>"011001111",
  27954=>"110110001",
  27955=>"000000000",
  27956=>"111111111",
  27957=>"011111111",
  27958=>"000001111",
  27959=>"000000000",
  27960=>"000000110",
  27961=>"001000111",
  27962=>"000000100",
  27963=>"001111011",
  27964=>"111110111",
  27965=>"110110111",
  27966=>"000000000",
  27967=>"100100101",
  27968=>"000000000",
  27969=>"100100110",
  27970=>"111101111",
  27971=>"111000000",
  27972=>"100100111",
  27973=>"111111111",
  27974=>"000000011",
  27975=>"100000000",
  27976=>"000000000",
  27977=>"111111100",
  27978=>"111011111",
  27979=>"000000000",
  27980=>"010011011",
  27981=>"000000000",
  27982=>"010000111",
  27983=>"110110100",
  27984=>"000110110",
  27985=>"111111111",
  27986=>"011001000",
  27987=>"111111001",
  27988=>"111111111",
  27989=>"011011011",
  27990=>"000000111",
  27991=>"111000000",
  27992=>"000000100",
  27993=>"110111111",
  27994=>"010110111",
  27995=>"111111000",
  27996=>"111111000",
  27997=>"111100000",
  27998=>"111011000",
  27999=>"100111111",
  28000=>"111001111",
  28001=>"000000000",
  28002=>"000000000",
  28003=>"111111111",
  28004=>"111111111",
  28005=>"000000001",
  28006=>"000011111",
  28007=>"001001111",
  28008=>"000000000",
  28009=>"000110110",
  28010=>"111111111",
  28011=>"111111111",
  28012=>"010000000",
  28013=>"111111111",
  28014=>"000000000",
  28015=>"110110000",
  28016=>"001000000",
  28017=>"011000000",
  28018=>"011011011",
  28019=>"110111111",
  28020=>"000000000",
  28021=>"000001111",
  28022=>"100100110",
  28023=>"000000001",
  28024=>"111111111",
  28025=>"000000110",
  28026=>"000000000",
  28027=>"111111111",
  28028=>"000000000",
  28029=>"000000001",
  28030=>"000000110",
  28031=>"001000100",
  28032=>"011010000",
  28033=>"000000111",
  28034=>"000110111",
  28035=>"111001111",
  28036=>"001111000",
  28037=>"000000000",
  28038=>"000000000",
  28039=>"011111111",
  28040=>"000000000",
  28041=>"011011010",
  28042=>"101101111",
  28043=>"111111111",
  28044=>"111111111",
  28045=>"111111001",
  28046=>"000100100",
  28047=>"000000000",
  28048=>"111111100",
  28049=>"111111111",
  28050=>"111111110",
  28051=>"111111111",
  28052=>"000000000",
  28053=>"000000000",
  28054=>"000001011",
  28055=>"000000000",
  28056=>"000111111",
  28057=>"111100100",
  28058=>"000000111",
  28059=>"000000110",
  28060=>"111101111",
  28061=>"000110000",
  28062=>"000000000",
  28063=>"111111111",
  28064=>"110100100",
  28065=>"001000000",
  28066=>"110100100",
  28067=>"101000000",
  28068=>"100100111",
  28069=>"111111111",
  28070=>"000000000",
  28071=>"001001110",
  28072=>"000010000",
  28073=>"011001011",
  28074=>"111111111",
  28075=>"010000000",
  28076=>"000000000",
  28077=>"110111001",
  28078=>"000000000",
  28079=>"000000000",
  28080=>"001000000",
  28081=>"000001111",
  28082=>"000111111",
  28083=>"111111111",
  28084=>"111111111",
  28085=>"000000100",
  28086=>"111111111",
  28087=>"110100000",
  28088=>"100111111",
  28089=>"001000000",
  28090=>"110110111",
  28091=>"000000000",
  28092=>"111111111",
  28093=>"100000101",
  28094=>"000001111",
  28095=>"011011010",
  28096=>"110110100",
  28097=>"000000000",
  28098=>"000000000",
  28099=>"000000000",
  28100=>"111001001",
  28101=>"111111010",
  28102=>"000000000",
  28103=>"000000000",
  28104=>"111111111",
  28105=>"000000000",
  28106=>"001001000",
  28107=>"011111110",
  28108=>"111011000",
  28109=>"111111111",
  28110=>"000000000",
  28111=>"000000111",
  28112=>"000000000",
  28113=>"000000000",
  28114=>"111111011",
  28115=>"000000000",
  28116=>"000100100",
  28117=>"000100111",
  28118=>"000000111",
  28119=>"000000000",
  28120=>"000000000",
  28121=>"000100100",
  28122=>"110000010",
  28123=>"111111111",
  28124=>"111111111",
  28125=>"111111011",
  28126=>"100000000",
  28127=>"000000110",
  28128=>"110111111",
  28129=>"111110000",
  28130=>"000001011",
  28131=>"111011001",
  28132=>"000011011",
  28133=>"000000000",
  28134=>"000000000",
  28135=>"000011111",
  28136=>"001001011",
  28137=>"111111000",
  28138=>"000000000",
  28139=>"000001001",
  28140=>"111000110",
  28141=>"001001001",
  28142=>"111111111",
  28143=>"111111011",
  28144=>"000000000",
  28145=>"011000000",
  28146=>"111111111",
  28147=>"111000000",
  28148=>"000000110",
  28149=>"000000110",
  28150=>"000011011",
  28151=>"100110100",
  28152=>"111111111",
  28153=>"010010010",
  28154=>"111111111",
  28155=>"111111111",
  28156=>"111111111",
  28157=>"000000000",
  28158=>"111111011",
  28159=>"000000000",
  28160=>"110000000",
  28161=>"001000100",
  28162=>"111110000",
  28163=>"010011000",
  28164=>"000001011",
  28165=>"001000100",
  28166=>"100100111",
  28167=>"111111111",
  28168=>"000011111",
  28169=>"000000000",
  28170=>"101100101",
  28171=>"100000010",
  28172=>"100110010",
  28173=>"011000000",
  28174=>"111110111",
  28175=>"110111111",
  28176=>"101100111",
  28177=>"000000000",
  28178=>"100000100",
  28179=>"000000111",
  28180=>"000000000",
  28181=>"001001001",
  28182=>"111111111",
  28183=>"110110110",
  28184=>"111111111",
  28185=>"110100110",
  28186=>"111101001",
  28187=>"110100100",
  28188=>"101001000",
  28189=>"010111111",
  28190=>"111111000",
  28191=>"110110100",
  28192=>"001000001",
  28193=>"011011111",
  28194=>"111110111",
  28195=>"111111111",
  28196=>"110111111",
  28197=>"111111111",
  28198=>"000000000",
  28199=>"000000000",
  28200=>"000000001",
  28201=>"010000000",
  28202=>"000000000",
  28203=>"000010100",
  28204=>"100000000",
  28205=>"000000000",
  28206=>"111111100",
  28207=>"001001001",
  28208=>"001111000",
  28209=>"011000001",
  28210=>"111111001",
  28211=>"100111111",
  28212=>"000000001",
  28213=>"110100000",
  28214=>"110111101",
  28215=>"110110010",
  28216=>"011111111",
  28217=>"111000111",
  28218=>"100101111",
  28219=>"000100110",
  28220=>"111111111",
  28221=>"000000000",
  28222=>"000000100",
  28223=>"101101111",
  28224=>"101111111",
  28225=>"011000111",
  28226=>"000000001",
  28227=>"111111001",
  28228=>"111111111",
  28229=>"001001000",
  28230=>"111111000",
  28231=>"001111111",
  28232=>"100000000",
  28233=>"000000000",
  28234=>"001111010",
  28235=>"000010011",
  28236=>"101111100",
  28237=>"000001001",
  28238=>"111100100",
  28239=>"000000000",
  28240=>"000000001",
  28241=>"011011011",
  28242=>"000000000",
  28243=>"111011111",
  28244=>"110110000",
  28245=>"000000000",
  28246=>"111111101",
  28247=>"100111111",
  28248=>"111101001",
  28249=>"000011000",
  28250=>"111111000",
  28251=>"110001011",
  28252=>"110001001",
  28253=>"111111011",
  28254=>"010000000",
  28255=>"111111011",
  28256=>"000000100",
  28257=>"101111111",
  28258=>"101001100",
  28259=>"111111111",
  28260=>"011000000",
  28261=>"101100111",
  28262=>"000000110",
  28263=>"101101111",
  28264=>"100000001",
  28265=>"000000101",
  28266=>"111111000",
  28267=>"111111111",
  28268=>"111111100",
  28269=>"000100110",
  28270=>"000000110",
  28271=>"111011000",
  28272=>"000110111",
  28273=>"011011011",
  28274=>"100000000",
  28275=>"100000011",
  28276=>"100110100",
  28277=>"100000100",
  28278=>"000010111",
  28279=>"111111111",
  28280=>"000100001",
  28281=>"001000000",
  28282=>"111111111",
  28283=>"000000000",
  28284=>"111111111",
  28285=>"110000000",
  28286=>"111111111",
  28287=>"000110000",
  28288=>"110110110",
  28289=>"000100000",
  28290=>"001000010",
  28291=>"110110000",
  28292=>"111101111",
  28293=>"001000000",
  28294=>"000000000",
  28295=>"011000000",
  28296=>"000000000",
  28297=>"011001000",
  28298=>"010110110",
  28299=>"000000000",
  28300=>"110100000",
  28301=>"100010011",
  28302=>"000000001",
  28303=>"000000000",
  28304=>"011011011",
  28305=>"000000000",
  28306=>"111111111",
  28307=>"011011100",
  28308=>"011011111",
  28309=>"111100100",
  28310=>"011111111",
  28311=>"000010000",
  28312=>"000110111",
  28313=>"111111111",
  28314=>"000111111",
  28315=>"000000000",
  28316=>"000010000",
  28317=>"000000000",
  28318=>"100000000",
  28319=>"000000011",
  28320=>"000000000",
  28321=>"101001001",
  28322=>"110100000",
  28323=>"000110000",
  28324=>"111111111",
  28325=>"000000000",
  28326=>"000000000",
  28327=>"011111000",
  28328=>"111011011",
  28329=>"111110000",
  28330=>"000000010",
  28331=>"111001111",
  28332=>"011111111",
  28333=>"000000000",
  28334=>"111111110",
  28335=>"011010100",
  28336=>"000000000",
  28337=>"100001000",
  28338=>"011001001",
  28339=>"011000010",
  28340=>"111110111",
  28341=>"111111111",
  28342=>"111111011",
  28343=>"000000100",
  28344=>"100000000",
  28345=>"111111111",
  28346=>"100000000",
  28347=>"010000011",
  28348=>"111111111",
  28349=>"000000000",
  28350=>"010000000",
  28351=>"111111111",
  28352=>"000100100",
  28353=>"011111111",
  28354=>"111111111",
  28355=>"111111111",
  28356=>"111000000",
  28357=>"000000010",
  28358=>"111111111",
  28359=>"111111011",
  28360=>"001000000",
  28361=>"111111111",
  28362=>"001001000",
  28363=>"011011001",
  28364=>"101001000",
  28365=>"111111000",
  28366=>"011001001",
  28367=>"000000000",
  28368=>"111100000",
  28369=>"111111110",
  28370=>"111111100",
  28371=>"000000000",
  28372=>"001100000",
  28373=>"001110110",
  28374=>"000000000",
  28375=>"111111111",
  28376=>"000000000",
  28377=>"000000000",
  28378=>"000000000",
  28379=>"111111111",
  28380=>"000000010",
  28381=>"111111111",
  28382=>"001000000",
  28383=>"111111000",
  28384=>"000111011",
  28385=>"011010111",
  28386=>"111111011",
  28387=>"010000000",
  28388=>"000111111",
  28389=>"011011011",
  28390=>"000000000",
  28391=>"000000000",
  28392=>"001111111",
  28393=>"111111111",
  28394=>"001000111",
  28395=>"111101101",
  28396=>"111111110",
  28397=>"000000001",
  28398=>"000000000",
  28399=>"111111111",
  28400=>"000000000",
  28401=>"000000000",
  28402=>"111111111",
  28403=>"000011011",
  28404=>"111111011",
  28405=>"111111111",
  28406=>"111111111",
  28407=>"001111001",
  28408=>"000000000",
  28409=>"000000000",
  28410=>"000000000",
  28411=>"000000000",
  28412=>"001011001",
  28413=>"111111111",
  28414=>"011111011",
  28415=>"000110110",
  28416=>"000000011",
  28417=>"100100000",
  28418=>"000000111",
  28419=>"001110110",
  28420=>"111111111",
  28421=>"011010000",
  28422=>"111111100",
  28423=>"111010111",
  28424=>"110111111",
  28425=>"000000000",
  28426=>"111010000",
  28427=>"000000011",
  28428=>"111111111",
  28429=>"111111111",
  28430=>"000000000",
  28431=>"011111110",
  28432=>"110110100",
  28433=>"101001111",
  28434=>"000000001",
  28435=>"111111111",
  28436=>"111111111",
  28437=>"000000000",
  28438=>"111111111",
  28439=>"100000000",
  28440=>"000000000",
  28441=>"111101000",
  28442=>"000000001",
  28443=>"111001000",
  28444=>"111111111",
  28445=>"111111111",
  28446=>"010010000",
  28447=>"111111111",
  28448=>"001000111",
  28449=>"001111111",
  28450=>"111111111",
  28451=>"111111000",
  28452=>"111011010",
  28453=>"111101111",
  28454=>"001011001",
  28455=>"011011011",
  28456=>"111100100",
  28457=>"000000000",
  28458=>"001000000",
  28459=>"111000000",
  28460=>"000000000",
  28461=>"110100110",
  28462=>"110010000",
  28463=>"000000000",
  28464=>"000000000",
  28465=>"010111011",
  28466=>"000000000",
  28467=>"001000000",
  28468=>"111111111",
  28469=>"000000000",
  28470=>"010110111",
  28471=>"000111110",
  28472=>"000000000",
  28473=>"000100100",
  28474=>"111011111",
  28475=>"010000011",
  28476=>"000000000",
  28477=>"111000000",
  28478=>"000111111",
  28479=>"011011010",
  28480=>"111111100",
  28481=>"000000000",
  28482=>"111111001",
  28483=>"000000000",
  28484=>"000000000",
  28485=>"000110110",
  28486=>"110111111",
  28487=>"111000011",
  28488=>"011011011",
  28489=>"000010110",
  28490=>"110001000",
  28491=>"001000001",
  28492=>"111101101",
  28493=>"100001000",
  28494=>"111111111",
  28495=>"011001000",
  28496=>"000000000",
  28497=>"111111111",
  28498=>"000000111",
  28499=>"000000110",
  28500=>"000000000",
  28501=>"000000000",
  28502=>"000000000",
  28503=>"000000000",
  28504=>"000000000",
  28505=>"111111111",
  28506=>"101101111",
  28507=>"111111111",
  28508=>"001011000",
  28509=>"000000000",
  28510=>"100000000",
  28511=>"110110000",
  28512=>"000000000",
  28513=>"111111111",
  28514=>"111111111",
  28515=>"100111000",
  28516=>"111111001",
  28517=>"101100000",
  28518=>"111000000",
  28519=>"000100001",
  28520=>"100110110",
  28521=>"111011011",
  28522=>"111111100",
  28523=>"000000000",
  28524=>"000110110",
  28525=>"000000000",
  28526=>"000110110",
  28527=>"010010010",
  28528=>"000000000",
  28529=>"000000110",
  28530=>"001111111",
  28531=>"111100110",
  28532=>"011011000",
  28533=>"000000001",
  28534=>"100111011",
  28535=>"100000000",
  28536=>"110110110",
  28537=>"000001000",
  28538=>"000000000",
  28539=>"000001000",
  28540=>"110000110",
  28541=>"111011010",
  28542=>"111101000",
  28543=>"000000000",
  28544=>"111111001",
  28545=>"000001001",
  28546=>"100100000",
  28547=>"000000100",
  28548=>"000000110",
  28549=>"000000111",
  28550=>"000000010",
  28551=>"110111010",
  28552=>"111110010",
  28553=>"000000110",
  28554=>"100111000",
  28555=>"000000000",
  28556=>"111111111",
  28557=>"111111110",
  28558=>"000000000",
  28559=>"000001001",
  28560=>"000000000",
  28561=>"010000110",
  28562=>"111011010",
  28563=>"100110000",
  28564=>"000001001",
  28565=>"000010000",
  28566=>"101101000",
  28567=>"111001000",
  28568=>"000000000",
  28569=>"111101100",
  28570=>"111111100",
  28571=>"001101111",
  28572=>"000000001",
  28573=>"111100000",
  28574=>"011000000",
  28575=>"000000000",
  28576=>"111111111",
  28577=>"100100000",
  28578=>"100000000",
  28579=>"000011111",
  28580=>"101000001",
  28581=>"010111010",
  28582=>"111111011",
  28583=>"000000000",
  28584=>"000000000",
  28585=>"001000111",
  28586=>"000000000",
  28587=>"000100100",
  28588=>"110000000",
  28589=>"111111100",
  28590=>"001111111",
  28591=>"101000111",
  28592=>"011000000",
  28593=>"111111111",
  28594=>"000000000",
  28595=>"100101001",
  28596=>"101111111",
  28597=>"000000000",
  28598=>"011111011",
  28599=>"011010110",
  28600=>"011000000",
  28601=>"000101111",
  28602=>"011111110",
  28603=>"110110110",
  28604=>"111111111",
  28605=>"011010100",
  28606=>"111001000",
  28607=>"110000000",
  28608=>"111101101",
  28609=>"111110000",
  28610=>"111011000",
  28611=>"111111010",
  28612=>"111011001",
  28613=>"011000100",
  28614=>"000111111",
  28615=>"110111111",
  28616=>"000000000",
  28617=>"111110000",
  28618=>"000000001",
  28619=>"000000000",
  28620=>"000000000",
  28621=>"000000000",
  28622=>"001000000",
  28623=>"010011011",
  28624=>"000000000",
  28625=>"001001001",
  28626=>"000000000",
  28627=>"011011011",
  28628=>"100100100",
  28629=>"000000000",
  28630=>"100010111",
  28631=>"111110000",
  28632=>"101100000",
  28633=>"000000010",
  28634=>"000000100",
  28635=>"111111111",
  28636=>"000000001",
  28637=>"001001011",
  28638=>"001001000",
  28639=>"100100100",
  28640=>"001000000",
  28641=>"000000000",
  28642=>"000000000",
  28643=>"111000000",
  28644=>"111001111",
  28645=>"000000001",
  28646=>"110011111",
  28647=>"010010110",
  28648=>"111111101",
  28649=>"000000000",
  28650=>"111000000",
  28651=>"111111111",
  28652=>"111011000",
  28653=>"000100000",
  28654=>"111111001",
  28655=>"000001000",
  28656=>"011111101",
  28657=>"000000011",
  28658=>"111111111",
  28659=>"001001000",
  28660=>"100000000",
  28661=>"111110010",
  28662=>"111111111",
  28663=>"111000000",
  28664=>"111111111",
  28665=>"111111111",
  28666=>"111111111",
  28667=>"000000000",
  28668=>"001001000",
  28669=>"110100000",
  28670=>"001001111",
  28671=>"000000101",
  28672=>"010100100",
  28673=>"111111111",
  28674=>"111111111",
  28675=>"000000000",
  28676=>"000000000",
  28677=>"011111111",
  28678=>"111111011",
  28679=>"111111111",
  28680=>"000110111",
  28681=>"111111111",
  28682=>"111000111",
  28683=>"111111111",
  28684=>"100100110",
  28685=>"000000110",
  28686=>"000000111",
  28687=>"000000000",
  28688=>"000000000",
  28689=>"000000100",
  28690=>"111010000",
  28691=>"111001000",
  28692=>"111111111",
  28693=>"000000010",
  28694=>"000000000",
  28695=>"010011111",
  28696=>"000000000",
  28697=>"000100100",
  28698=>"000000000",
  28699=>"110110111",
  28700=>"111111111",
  28701=>"100100100",
  28702=>"000000000",
  28703=>"000000110",
  28704=>"111111111",
  28705=>"111111111",
  28706=>"111111111",
  28707=>"111111111",
  28708=>"000000000",
  28709=>"111111110",
  28710=>"000000000",
  28711=>"010011000",
  28712=>"111000000",
  28713=>"000000000",
  28714=>"100111000",
  28715=>"000111111",
  28716=>"000000000",
  28717=>"111000000",
  28718=>"111111111",
  28719=>"000000001",
  28720=>"111110111",
  28721=>"000111000",
  28722=>"000000000",
  28723=>"000000000",
  28724=>"000000100",
  28725=>"111101000",
  28726=>"000110000",
  28727=>"111111111",
  28728=>"000000000",
  28729=>"000000000",
  28730=>"100000000",
  28731=>"111111110",
  28732=>"111111000",
  28733=>"111110111",
  28734=>"000011001",
  28735=>"000110000",
  28736=>"111111000",
  28737=>"000000000",
  28738=>"000000100",
  28739=>"110111000",
  28740=>"000000000",
  28741=>"111111111",
  28742=>"001111111",
  28743=>"000000001",
  28744=>"000000000",
  28745=>"111111111",
  28746=>"111111111",
  28747=>"000000000",
  28748=>"111111111",
  28749=>"111011101",
  28750=>"000011100",
  28751=>"000110110",
  28752=>"111000000",
  28753=>"000000000",
  28754=>"101101100",
  28755=>"111110110",
  28756=>"111111110",
  28757=>"000000100",
  28758=>"111100000",
  28759=>"111111111",
  28760=>"110101111",
  28761=>"111111111",
  28762=>"000101101",
  28763=>"000000000",
  28764=>"000000000",
  28765=>"000000000",
  28766=>"011011111",
  28767=>"000000000",
  28768=>"111100000",
  28769=>"000110001",
  28770=>"100110111",
  28771=>"000110111",
  28772=>"111111111",
  28773=>"000010000",
  28774=>"100101111",
  28775=>"000000000",
  28776=>"111100111",
  28777=>"000000000",
  28778=>"000000000",
  28779=>"000000000",
  28780=>"100110100",
  28781=>"000000000",
  28782=>"110100111",
  28783=>"111000000",
  28784=>"111111111",
  28785=>"000000000",
  28786=>"010110011",
  28787=>"000000000",
  28788=>"100000000",
  28789=>"110111111",
  28790=>"001001001",
  28791=>"101111111",
  28792=>"111111111",
  28793=>"000111111",
  28794=>"010111010",
  28795=>"000000000",
  28796=>"111110111",
  28797=>"111111111",
  28798=>"111001000",
  28799=>"000100000",
  28800=>"101000000",
  28801=>"000000101",
  28802=>"000000000",
  28803=>"111111111",
  28804=>"001000000",
  28805=>"111111111",
  28806=>"100111110",
  28807=>"111000000",
  28808=>"000000000",
  28809=>"111111111",
  28810=>"110000000",
  28811=>"000111111",
  28812=>"000000000",
  28813=>"000000000",
  28814=>"110111001",
  28815=>"111000000",
  28816=>"000111010",
  28817=>"100100001",
  28818=>"000000000",
  28819=>"000000000",
  28820=>"111110000",
  28821=>"100100100",
  28822=>"000000011",
  28823=>"111000000",
  28824=>"010110010",
  28825=>"100111111",
  28826=>"101101111",
  28827=>"111111011",
  28828=>"111111001",
  28829=>"011110110",
  28830=>"110010000",
  28831=>"111101101",
  28832=>"000000001",
  28833=>"000000000",
  28834=>"000000000",
  28835=>"111111111",
  28836=>"110110110",
  28837=>"111111111",
  28838=>"000010000",
  28839=>"011011111",
  28840=>"000000000",
  28841=>"010100000",
  28842=>"000001111",
  28843=>"000000000",
  28844=>"000000000",
  28845=>"110110110",
  28846=>"111001001",
  28847=>"000000000",
  28848=>"000010000",
  28849=>"110111000",
  28850=>"010111010",
  28851=>"000111010",
  28852=>"000100110",
  28853=>"111111111",
  28854=>"000011000",
  28855=>"000000000",
  28856=>"111100111",
  28857=>"000000000",
  28858=>"001000000",
  28859=>"100000000",
  28860=>"010011101",
  28861=>"000000000",
  28862=>"111111111",
  28863=>"000000000",
  28864=>"101101000",
  28865=>"000000000",
  28866=>"111111111",
  28867=>"101111111",
  28868=>"000010000",
  28869=>"111111111",
  28870=>"111101100",
  28871=>"110110001",
  28872=>"011111010",
  28873=>"000000000",
  28874=>"110110111",
  28875=>"001001111",
  28876=>"000000000",
  28877=>"000000000",
  28878=>"111111000",
  28879=>"000000111",
  28880=>"000000111",
  28881=>"000000101",
  28882=>"111111110",
  28883=>"110110111",
  28884=>"000001101",
  28885=>"111111001",
  28886=>"000000100",
  28887=>"111111111",
  28888=>"000000000",
  28889=>"000000000",
  28890=>"000000000",
  28891=>"111111111",
  28892=>"111111111",
  28893=>"111111111",
  28894=>"000000000",
  28895=>"110110000",
  28896=>"000100101",
  28897=>"000000000",
  28898=>"000111111",
  28899=>"101001111",
  28900=>"101000000",
  28901=>"000000000",
  28902=>"111111111",
  28903=>"111000110",
  28904=>"000000100",
  28905=>"000010110",
  28906=>"101111111",
  28907=>"111111111",
  28908=>"000010010",
  28909=>"111100111",
  28910=>"100101001",
  28911=>"010100100",
  28912=>"111111111",
  28913=>"111000000",
  28914=>"001001011",
  28915=>"000000000",
  28916=>"011001000",
  28917=>"000000000",
  28918=>"111111110",
  28919=>"000000000",
  28920=>"000100111",
  28921=>"001000111",
  28922=>"110110111",
  28923=>"000000001",
  28924=>"000000000",
  28925=>"111101100",
  28926=>"000000000",
  28927=>"100100111",
  28928=>"000000000",
  28929=>"010011001",
  28930=>"000111111",
  28931=>"100111000",
  28932=>"100100111",
  28933=>"111111111",
  28934=>"101001101",
  28935=>"000010110",
  28936=>"110000110",
  28937=>"000000111",
  28938=>"111111101",
  28939=>"011011110",
  28940=>"011011000",
  28941=>"100001111",
  28942=>"000000110",
  28943=>"100001111",
  28944=>"110100000",
  28945=>"000000000",
  28946=>"000000111",
  28947=>"000000000",
  28948=>"111111000",
  28949=>"111111111",
  28950=>"000000000",
  28951=>"100000000",
  28952=>"100000000",
  28953=>"000000000",
  28954=>"000000000",
  28955=>"111011111",
  28956=>"000100100",
  28957=>"111111111",
  28958=>"111011001",
  28959=>"000000000",
  28960=>"111111111",
  28961=>"111111111",
  28962=>"011111001",
  28963=>"111111111",
  28964=>"000111111",
  28965=>"111100111",
  28966=>"000000000",
  28967=>"111111111",
  28968=>"000000011",
  28969=>"111100000",
  28970=>"111111000",
  28971=>"111111111",
  28972=>"000000000",
  28973=>"100100100",
  28974=>"111111111",
  28975=>"111111111",
  28976=>"111111111",
  28977=>"110100100",
  28978=>"000100111",
  28979=>"111100100",
  28980=>"111111111",
  28981=>"001000111",
  28982=>"000000000",
  28983=>"111000000",
  28984=>"000000000",
  28985=>"000000000",
  28986=>"010010000",
  28987=>"111111111",
  28988=>"111111111",
  28989=>"110100000",
  28990=>"111100111",
  28991=>"111111001",
  28992=>"111111011",
  28993=>"000000111",
  28994=>"111111111",
  28995=>"111110111",
  28996=>"010000000",
  28997=>"111011000",
  28998=>"111110100",
  28999=>"000000000",
  29000=>"000000000",
  29001=>"111111001",
  29002=>"111110100",
  29003=>"000000000",
  29004=>"111011011",
  29005=>"111111111",
  29006=>"000010100",
  29007=>"011011011",
  29008=>"000000110",
  29009=>"010110111",
  29010=>"000000000",
  29011=>"000000000",
  29012=>"000000000",
  29013=>"011001011",
  29014=>"111111111",
  29015=>"111011111",
  29016=>"100111110",
  29017=>"000000000",
  29018=>"111111111",
  29019=>"111110110",
  29020=>"111111111",
  29021=>"110111111",
  29022=>"111111101",
  29023=>"001011111",
  29024=>"111111111",
  29025=>"000011001",
  29026=>"000000110",
  29027=>"111111111",
  29028=>"110100100",
  29029=>"110110110",
  29030=>"111111111",
  29031=>"000000100",
  29032=>"001011001",
  29033=>"000000000",
  29034=>"000100111",
  29035=>"000110111",
  29036=>"111100000",
  29037=>"111011111",
  29038=>"111111111",
  29039=>"000000000",
  29040=>"111000111",
  29041=>"111111111",
  29042=>"111000000",
  29043=>"000000000",
  29044=>"000000000",
  29045=>"111111101",
  29046=>"000000000",
  29047=>"000000000",
  29048=>"111111111",
  29049=>"010111111",
  29050=>"100100111",
  29051=>"000000000",
  29052=>"111111111",
  29053=>"111111111",
  29054=>"111111111",
  29055=>"000000001",
  29056=>"110111111",
  29057=>"111111100",
  29058=>"111111111",
  29059=>"001011000",
  29060=>"110010000",
  29061=>"000000000",
  29062=>"111111101",
  29063=>"001011000",
  29064=>"000000000",
  29065=>"100100000",
  29066=>"101111111",
  29067=>"010000010",
  29068=>"111111111",
  29069=>"111111111",
  29070=>"110000000",
  29071=>"000000000",
  29072=>"000000000",
  29073=>"110110110",
  29074=>"110111111",
  29075=>"111111111",
  29076=>"111111011",
  29077=>"000001111",
  29078=>"110000100",
  29079=>"011001001",
  29080=>"000000000",
  29081=>"101101111",
  29082=>"111101001",
  29083=>"001000000",
  29084=>"000000000",
  29085=>"111110000",
  29086=>"000000000",
  29087=>"000000000",
  29088=>"111000000",
  29089=>"001011011",
  29090=>"000000000",
  29091=>"000000000",
  29092=>"111111111",
  29093=>"000100111",
  29094=>"000000000",
  29095=>"000000101",
  29096=>"111111111",
  29097=>"000000000",
  29098=>"000000000",
  29099=>"000000010",
  29100=>"000000000",
  29101=>"000000000",
  29102=>"000000000",
  29103=>"010000000",
  29104=>"111111111",
  29105=>"110111111",
  29106=>"111100000",
  29107=>"110111111",
  29108=>"111101111",
  29109=>"000000000",
  29110=>"111111011",
  29111=>"110100000",
  29112=>"111111111",
  29113=>"011000000",
  29114=>"100100111",
  29115=>"111111111",
  29116=>"000000000",
  29117=>"111110000",
  29118=>"000111111",
  29119=>"000000000",
  29120=>"111111000",
  29121=>"000111011",
  29122=>"111111111",
  29123=>"111111111",
  29124=>"000000010",
  29125=>"100100001",
  29126=>"110100000",
  29127=>"100100100",
  29128=>"000000000",
  29129=>"000000000",
  29130=>"111110111",
  29131=>"000000011",
  29132=>"000000000",
  29133=>"000110000",
  29134=>"000000000",
  29135=>"000000000",
  29136=>"001111111",
  29137=>"100101000",
  29138=>"111111111",
  29139=>"111111111",
  29140=>"111101000",
  29141=>"111111111",
  29142=>"100000000",
  29143=>"000100111",
  29144=>"000000000",
  29145=>"110110111",
  29146=>"110000000",
  29147=>"111111111",
  29148=>"111000000",
  29149=>"110110100",
  29150=>"111111111",
  29151=>"000000101",
  29152=>"000010000",
  29153=>"000000000",
  29154=>"111111010",
  29155=>"111111101",
  29156=>"111110010",
  29157=>"001000000",
  29158=>"000000000",
  29159=>"111111111",
  29160=>"110110100",
  29161=>"001001101",
  29162=>"000000000",
  29163=>"010110111",
  29164=>"111111010",
  29165=>"001000000",
  29166=>"111111110",
  29167=>"000000010",
  29168=>"000000000",
  29169=>"000000111",
  29170=>"001111111",
  29171=>"000000000",
  29172=>"000000000",
  29173=>"111100100",
  29174=>"000000000",
  29175=>"101111111",
  29176=>"000000000",
  29177=>"000010010",
  29178=>"110010000",
  29179=>"011110111",
  29180=>"111000000",
  29181=>"111111001",
  29182=>"111111111",
  29183=>"000110000",
  29184=>"001111111",
  29185=>"110111000",
  29186=>"010100100",
  29187=>"000000010",
  29188=>"110110111",
  29189=>"000000001",
  29190=>"111111111",
  29191=>"111111100",
  29192=>"011001011",
  29193=>"000000001",
  29194=>"001001001",
  29195=>"101100000",
  29196=>"101001111",
  29197=>"111110110",
  29198=>"111111110",
  29199=>"111111111",
  29200=>"111111111",
  29201=>"010000000",
  29202=>"111100000",
  29203=>"101100000",
  29204=>"000000000",
  29205=>"111111010",
  29206=>"100000000",
  29207=>"001001001",
  29208=>"110110110",
  29209=>"111111000",
  29210=>"001001001",
  29211=>"000000100",
  29212=>"111111111",
  29213=>"111110111",
  29214=>"000100111",
  29215=>"110000000",
  29216=>"001000100",
  29217=>"110010000",
  29218=>"011011111",
  29219=>"000000001",
  29220=>"000000011",
  29221=>"111111111",
  29222=>"010010000",
  29223=>"100100100",
  29224=>"101101111",
  29225=>"010000000",
  29226=>"000000000",
  29227=>"100011000",
  29228=>"010110111",
  29229=>"000100111",
  29230=>"000111001",
  29231=>"000000000",
  29232=>"000000101",
  29233=>"001101111",
  29234=>"001001001",
  29235=>"111111111",
  29236=>"000000000",
  29237=>"000001101",
  29238=>"000101111",
  29239=>"010010110",
  29240=>"001101000",
  29241=>"001001000",
  29242=>"000000000",
  29243=>"111111111",
  29244=>"111111111",
  29245=>"011010000",
  29246=>"011011011",
  29247=>"001001001",
  29248=>"000000001",
  29249=>"100100111",
  29250=>"110000011",
  29251=>"111010000",
  29252=>"000000000",
  29253=>"001010011",
  29254=>"011000010",
  29255=>"000011011",
  29256=>"011111111",
  29257=>"000001001",
  29258=>"100000111",
  29259=>"000000001",
  29260=>"010111000",
  29261=>"101101111",
  29262=>"111111111",
  29263=>"000001101",
  29264=>"111111101",
  29265=>"011111111",
  29266=>"000100111",
  29267=>"101000000",
  29268=>"111000000",
  29269=>"000000011",
  29270=>"111111111",
  29271=>"111111111",
  29272=>"000000000",
  29273=>"000000000",
  29274=>"010111111",
  29275=>"110100000",
  29276=>"110000000",
  29277=>"111000000",
  29278=>"010110110",
  29279=>"011011011",
  29280=>"000001010",
  29281=>"110111111",
  29282=>"111111111",
  29283=>"111110111",
  29284=>"110110010",
  29285=>"100100101",
  29286=>"111111111",
  29287=>"111111111",
  29288=>"111101101",
  29289=>"000001111",
  29290=>"111110110",
  29291=>"111111010",
  29292=>"100110111",
  29293=>"111111101",
  29294=>"111111110",
  29295=>"000000101",
  29296=>"000000000",
  29297=>"000001001",
  29298=>"000000000",
  29299=>"001000000",
  29300=>"000000000",
  29301=>"000000000",
  29302=>"000000001",
  29303=>"100100000",
  29304=>"000000000",
  29305=>"110111010",
  29306=>"001000000",
  29307=>"000000101",
  29308=>"000100100",
  29309=>"000100100",
  29310=>"000000001",
  29311=>"110111010",
  29312=>"000000000",
  29313=>"110110110",
  29314=>"000100110",
  29315=>"111011010",
  29316=>"111111111",
  29317=>"000001101",
  29318=>"100110000",
  29319=>"111011000",
  29320=>"110010111",
  29321=>"111111000",
  29322=>"110000000",
  29323=>"110100100",
  29324=>"011001000",
  29325=>"111111111",
  29326=>"000001111",
  29327=>"111111110",
  29328=>"000000001",
  29329=>"000000000",
  29330=>"001001011",
  29331=>"110110110",
  29332=>"111110110",
  29333=>"111111011",
  29334=>"010010000",
  29335=>"000000100",
  29336=>"010111111",
  29337=>"101000101",
  29338=>"000100100",
  29339=>"111000000",
  29340=>"011111111",
  29341=>"111000000",
  29342=>"001010000",
  29343=>"100111011",
  29344=>"000000000",
  29345=>"001011010",
  29346=>"001000001",
  29347=>"111111001",
  29348=>"000010100",
  29349=>"001111110",
  29350=>"110110010",
  29351=>"000000110",
  29352=>"111111111",
  29353=>"111001001",
  29354=>"000100100",
  29355=>"000000011",
  29356=>"001001111",
  29357=>"000100111",
  29358=>"111111111",
  29359=>"001001101",
  29360=>"010000000",
  29361=>"001001011",
  29362=>"111111111",
  29363=>"110010111",
  29364=>"000000000",
  29365=>"000000111",
  29366=>"000000000",
  29367=>"111111011",
  29368=>"010000000",
  29369=>"000000000",
  29370=>"000000000",
  29371=>"111110110",
  29372=>"010010010",
  29373=>"110111111",
  29374=>"111001000",
  29375=>"110110111",
  29376=>"111111111",
  29377=>"000000001",
  29378=>"110000110",
  29379=>"111111000",
  29380=>"100000000",
  29381=>"101001000",
  29382=>"111111111",
  29383=>"101111101",
  29384=>"111111111",
  29385=>"001001001",
  29386=>"100110111",
  29387=>"111111111",
  29388=>"111011001",
  29389=>"111110000",
  29390=>"111111111",
  29391=>"011110110",
  29392=>"000100101",
  29393=>"111111011",
  29394=>"011001001",
  29395=>"111111011",
  29396=>"111111001",
  29397=>"110110100",
  29398=>"000110111",
  29399=>"111110000",
  29400=>"000000011",
  29401=>"000000001",
  29402=>"000000001",
  29403=>"111111111",
  29404=>"111110000",
  29405=>"110111110",
  29406=>"011011000",
  29407=>"001111100",
  29408=>"111000000",
  29409=>"000010010",
  29410=>"111111011",
  29411=>"011011010",
  29412=>"100111111",
  29413=>"011011011",
  29414=>"010010001",
  29415=>"111111111",
  29416=>"110010111",
  29417=>"000001001",
  29418=>"100000000",
  29419=>"011111111",
  29420=>"111111111",
  29421=>"000000000",
  29422=>"000100100",
  29423=>"001111111",
  29424=>"110111111",
  29425=>"111111011",
  29426=>"110010110",
  29427=>"000000000",
  29428=>"000111111",
  29429=>"100000100",
  29430=>"111111111",
  29431=>"000000010",
  29432=>"000000001",
  29433=>"111001011",
  29434=>"111001111",
  29435=>"111111111",
  29436=>"000000000",
  29437=>"000000110",
  29438=>"111110110",
  29439=>"111111011",
  29440=>"000000000",
  29441=>"000000000",
  29442=>"001001000",
  29443=>"000000000",
  29444=>"001000000",
  29445=>"111111101",
  29446=>"100000100",
  29447=>"111111111",
  29448=>"001001000",
  29449=>"000000000",
  29450=>"111001000",
  29451=>"100101100",
  29452=>"000000111",
  29453=>"110111110",
  29454=>"001001001",
  29455=>"111111111",
  29456=>"101101001",
  29457=>"011011001",
  29458=>"100000000",
  29459=>"001001001",
  29460=>"101100000",
  29461=>"111000010",
  29462=>"001001111",
  29463=>"001001001",
  29464=>"100111111",
  29465=>"000000001",
  29466=>"000101110",
  29467=>"111111000",
  29468=>"100101111",
  29469=>"000000000",
  29470=>"100110000",
  29471=>"000000000",
  29472=>"100111011",
  29473=>"111111111",
  29474=>"000000000",
  29475=>"000000000",
  29476=>"000000001",
  29477=>"111000000",
  29478=>"111111111",
  29479=>"001000111",
  29480=>"000000000",
  29481=>"101001000",
  29482=>"001000001",
  29483=>"000000111",
  29484=>"111111110",
  29485=>"110111110",
  29486=>"111111111",
  29487=>"111001001",
  29488=>"100001000",
  29489=>"110001001",
  29490=>"110110110",
  29491=>"000000000",
  29492=>"111110000",
  29493=>"000011011",
  29494=>"000001001",
  29495=>"010110000",
  29496=>"000110111",
  29497=>"001001101",
  29498=>"000000000",
  29499=>"111111111",
  29500=>"000010011",
  29501=>"111111011",
  29502=>"100111101",
  29503=>"010110110",
  29504=>"000000000",
  29505=>"000000001",
  29506=>"001011011",
  29507=>"110111111",
  29508=>"011101111",
  29509=>"110111111",
  29510=>"000100100",
  29511=>"011001000",
  29512=>"111111111",
  29513=>"111110110",
  29514=>"000000000",
  29515=>"001001001",
  29516=>"001000000",
  29517=>"000000100",
  29518=>"000000000",
  29519=>"110011101",
  29520=>"001001111",
  29521=>"011011011",
  29522=>"111111111",
  29523=>"010011010",
  29524=>"000000000",
  29525=>"011011011",
  29526=>"110111111",
  29527=>"001001101",
  29528=>"111111111",
  29529=>"111111111",
  29530=>"000000000",
  29531=>"000000111",
  29532=>"111111111",
  29533=>"000000000",
  29534=>"001000000",
  29535=>"000000000",
  29536=>"000001001",
  29537=>"111011011",
  29538=>"101111111",
  29539=>"111101111",
  29540=>"001011100",
  29541=>"111011001",
  29542=>"110111111",
  29543=>"001001000",
  29544=>"000110110",
  29545=>"000000000",
  29546=>"100001101",
  29547=>"001000010",
  29548=>"000001001",
  29549=>"000011111",
  29550=>"000000000",
  29551=>"000000001",
  29552=>"001001001",
  29553=>"000010011",
  29554=>"010111111",
  29555=>"111111110",
  29556=>"001001001",
  29557=>"111111111",
  29558=>"000000011",
  29559=>"001111100",
  29560=>"101001101",
  29561=>"001100100",
  29562=>"111111111",
  29563=>"000000000",
  29564=>"000000000",
  29565=>"111111111",
  29566=>"111111111",
  29567=>"101011111",
  29568=>"111111100",
  29569=>"011111111",
  29570=>"000000000",
  29571=>"110110000",
  29572=>"111001101",
  29573=>"111111111",
  29574=>"011111111",
  29575=>"000100001",
  29576=>"000001011",
  29577=>"111111111",
  29578=>"111111111",
  29579=>"001000000",
  29580=>"101001001",
  29581=>"111011000",
  29582=>"000000000",
  29583=>"000000001",
  29584=>"111110110",
  29585=>"111111000",
  29586=>"111111111",
  29587=>"010010010",
  29588=>"111000000",
  29589=>"000000000",
  29590=>"000111111",
  29591=>"111111111",
  29592=>"111111111",
  29593=>"001000000",
  29594=>"001110111",
  29595=>"111111110",
  29596=>"000000000",
  29597=>"110111111",
  29598=>"000100110",
  29599=>"000000000",
  29600=>"111111111",
  29601=>"111110110",
  29602=>"000000111",
  29603=>"000110111",
  29604=>"000000000",
  29605=>"111111111",
  29606=>"111111111",
  29607=>"110110111",
  29608=>"111100000",
  29609=>"001001111",
  29610=>"000000110",
  29611=>"000000000",
  29612=>"111111110",
  29613=>"111111111",
  29614=>"001001000",
  29615=>"100000101",
  29616=>"111111111",
  29617=>"000000000",
  29618=>"111111100",
  29619=>"111001001",
  29620=>"011011001",
  29621=>"001001000",
  29622=>"011000111",
  29623=>"000000000",
  29624=>"000111111",
  29625=>"010010011",
  29626=>"111110111",
  29627=>"110110111",
  29628=>"000000000",
  29629=>"111111111",
  29630=>"111011101",
  29631=>"000011011",
  29632=>"111001000",
  29633=>"111100000",
  29634=>"001011101",
  29635=>"000011011",
  29636=>"000000001",
  29637=>"001000100",
  29638=>"000110110",
  29639=>"000111011",
  29640=>"000000000",
  29641=>"000000000",
  29642=>"000000001",
  29643=>"111111011",
  29644=>"110010000",
  29645=>"000000000",
  29646=>"001001001",
  29647=>"000010000",
  29648=>"111111111",
  29649=>"011111011",
  29650=>"110110110",
  29651=>"111111010",
  29652=>"011101001",
  29653=>"101001010",
  29654=>"000000000",
  29655=>"100000000",
  29656=>"000000000",
  29657=>"001000001",
  29658=>"110111011",
  29659=>"001101111",
  29660=>"111101110",
  29661=>"000000101",
  29662=>"110111111",
  29663=>"000000000",
  29664=>"001000000",
  29665=>"000000000",
  29666=>"000000000",
  29667=>"011010011",
  29668=>"000000001",
  29669=>"000100100",
  29670=>"011011011",
  29671=>"011111111",
  29672=>"001101101",
  29673=>"111111111",
  29674=>"101111111",
  29675=>"110110000",
  29676=>"000001000",
  29677=>"111111011",
  29678=>"111100100",
  29679=>"111101000",
  29680=>"001000101",
  29681=>"000111111",
  29682=>"001001001",
  29683=>"000000000",
  29684=>"111001000",
  29685=>"000000110",
  29686=>"101101001",
  29687=>"110110111",
  29688=>"111101000",
  29689=>"001001001",
  29690=>"100110111",
  29691=>"000011001",
  29692=>"111111110",
  29693=>"011001001",
  29694=>"000000111",
  29695=>"111111111",
  29696=>"000000110",
  29697=>"110110000",
  29698=>"101000000",
  29699=>"011110110",
  29700=>"111111111",
  29701=>"000001111",
  29702=>"010000000",
  29703=>"000000010",
  29704=>"011000111",
  29705=>"000110000",
  29706=>"111111111",
  29707=>"100111111",
  29708=>"001011111",
  29709=>"001011010",
  29710=>"000010001",
  29711=>"111111111",
  29712=>"011011011",
  29713=>"100111111",
  29714=>"000000000",
  29715=>"111111111",
  29716=>"111110000",
  29717=>"101001111",
  29718=>"111011111",
  29719=>"001111111",
  29720=>"010100110",
  29721=>"111111111",
  29722=>"000000000",
  29723=>"111111100",
  29724=>"000000000",
  29725=>"000001001",
  29726=>"000001000",
  29727=>"000000110",
  29728=>"111111111",
  29729=>"110000000",
  29730=>"000000000",
  29731=>"100111111",
  29732=>"110000000",
  29733=>"110100110",
  29734=>"111100100",
  29735=>"001011000",
  29736=>"010110100",
  29737=>"011001111",
  29738=>"110111111",
  29739=>"000000000",
  29740=>"111001111",
  29741=>"101000000",
  29742=>"000000010",
  29743=>"111011000",
  29744=>"000000111",
  29745=>"000001000",
  29746=>"000010000",
  29747=>"000011011",
  29748=>"111001101",
  29749=>"000000000",
  29750=>"110000111",
  29751=>"000000000",
  29752=>"000000000",
  29753=>"011111011",
  29754=>"111111110",
  29755=>"000000101",
  29756=>"011000000",
  29757=>"111111000",
  29758=>"011011001",
  29759=>"000000000",
  29760=>"001001000",
  29761=>"101101000",
  29762=>"111010000",
  29763=>"111011000",
  29764=>"001001001",
  29765=>"011001000",
  29766=>"111111111",
  29767=>"111100111",
  29768=>"000010111",
  29769=>"000000000",
  29770=>"011011000",
  29771=>"000000000",
  29772=>"001111011",
  29773=>"111111111",
  29774=>"000000000",
  29775=>"111000000",
  29776=>"110111111",
  29777=>"110111111",
  29778=>"110000000",
  29779=>"000000001",
  29780=>"011001011",
  29781=>"001100000",
  29782=>"010100000",
  29783=>"000000000",
  29784=>"001111100",
  29785=>"000000000",
  29786=>"111111111",
  29787=>"000000000",
  29788=>"000111111",
  29789=>"000000111",
  29790=>"000111111",
  29791=>"111000000",
  29792=>"000000000",
  29793=>"000001101",
  29794=>"000000000",
  29795=>"000000001",
  29796=>"001011111",
  29797=>"110111111",
  29798=>"011001000",
  29799=>"000000000",
  29800=>"000000001",
  29801=>"111111111",
  29802=>"000000000",
  29803=>"100110110",
  29804=>"001001101",
  29805=>"111111001",
  29806=>"000010000",
  29807=>"000110111",
  29808=>"000110111",
  29809=>"111111111",
  29810=>"000000000",
  29811=>"100100111",
  29812=>"110100000",
  29813=>"111001000",
  29814=>"000000000",
  29815=>"111111111",
  29816=>"000000000",
  29817=>"100111111",
  29818=>"111110000",
  29819=>"000000111",
  29820=>"110111111",
  29821=>"111000000",
  29822=>"000000001",
  29823=>"001001001",
  29824=>"111111111",
  29825=>"111111110",
  29826=>"000000000",
  29827=>"000000110",
  29828=>"000000100",
  29829=>"111111111",
  29830=>"111111111",
  29831=>"000000000",
  29832=>"111101100",
  29833=>"001000000",
  29834=>"000000000",
  29835=>"000000000",
  29836=>"100111111",
  29837=>"111111110",
  29838=>"011011000",
  29839=>"000000000",
  29840=>"000110110",
  29841=>"101100111",
  29842=>"000000000",
  29843=>"000111111",
  29844=>"011001001",
  29845=>"110011111",
  29846=>"000001111",
  29847=>"001000000",
  29848=>"000000000",
  29849=>"111111001",
  29850=>"000000000",
  29851=>"000000000",
  29852=>"000100100",
  29853=>"100000110",
  29854=>"111111111",
  29855=>"000000010",
  29856=>"000101101",
  29857=>"111001001",
  29858=>"111111111",
  29859=>"000001110",
  29860=>"001001001",
  29861=>"010011000",
  29862=>"001001101",
  29863=>"111000000",
  29864=>"000000000",
  29865=>"000000001",
  29866=>"000000100",
  29867=>"000101000",
  29868=>"010010000",
  29869=>"000000111",
  29870=>"111111011",
  29871=>"100111011",
  29872=>"000000000",
  29873=>"110110111",
  29874=>"111111111",
  29875=>"100000111",
  29876=>"111110000",
  29877=>"111000101",
  29878=>"110110111",
  29879=>"000000000",
  29880=>"000001011",
  29881=>"000000000",
  29882=>"000110011",
  29883=>"110000000",
  29884=>"000000000",
  29885=>"110111110",
  29886=>"111111111",
  29887=>"100001000",
  29888=>"100000000",
  29889=>"110011011",
  29890=>"111111111",
  29891=>"010010011",
  29892=>"000000000",
  29893=>"000011000",
  29894=>"000100010",
  29895=>"000001001",
  29896=>"000010011",
  29897=>"100001001",
  29898=>"100000000",
  29899=>"000100100",
  29900=>"001001001",
  29901=>"000100100",
  29902=>"000000000",
  29903=>"111111000",
  29904=>"001000100",
  29905=>"111000000",
  29906=>"111011011",
  29907=>"000000000",
  29908=>"000000000",
  29909=>"110111110",
  29910=>"000000001",
  29911=>"101001001",
  29912=>"101101000",
  29913=>"001000000",
  29914=>"100110111",
  29915=>"000000000",
  29916=>"110110110",
  29917=>"111111010",
  29918=>"111111111",
  29919=>"000000100",
  29920=>"111111111",
  29921=>"001000100",
  29922=>"000000000",
  29923=>"000000000",
  29924=>"111110000",
  29925=>"000000001",
  29926=>"010111001",
  29927=>"111111111",
  29928=>"111111111",
  29929=>"000100010",
  29930=>"000000001",
  29931=>"100100000",
  29932=>"000000001",
  29933=>"000011111",
  29934=>"000000111",
  29935=>"000000000",
  29936=>"011000010",
  29937=>"110111111",
  29938=>"000000001",
  29939=>"000001111",
  29940=>"010000000",
  29941=>"111000000",
  29942=>"101101111",
  29943=>"111110101",
  29944=>"000000000",
  29945=>"000100111",
  29946=>"111111111",
  29947=>"000000101",
  29948=>"000000000",
  29949=>"111111101",
  29950=>"000100110",
  29951=>"111111110",
  29952=>"000000000",
  29953=>"001000000",
  29954=>"110110000",
  29955=>"111111111",
  29956=>"000001001",
  29957=>"011011010",
  29958=>"111011111",
  29959=>"111111111",
  29960=>"000000000",
  29961=>"000000000",
  29962=>"010010111",
  29963=>"111111111",
  29964=>"111101001",
  29965=>"111110101",
  29966=>"000000000",
  29967=>"111110111",
  29968=>"000100100",
  29969=>"000000000",
  29970=>"000000100",
  29971=>"000000001",
  29972=>"000000000",
  29973=>"111010011",
  29974=>"011001011",
  29975=>"110111001",
  29976=>"001111111",
  29977=>"000111111",
  29978=>"000000000",
  29979=>"111000111",
  29980=>"011011111",
  29981=>"010000111",
  29982=>"000000000",
  29983=>"100101111",
  29984=>"110111011",
  29985=>"000110111",
  29986=>"111111011",
  29987=>"000101111",
  29988=>"111110110",
  29989=>"000010011",
  29990=>"000110111",
  29991=>"110110000",
  29992=>"000000000",
  29993=>"000110111",
  29994=>"101111111",
  29995=>"100100000",
  29996=>"111111111",
  29997=>"001000101",
  29998=>"000001001",
  29999=>"000000001",
  30000=>"000011110",
  30001=>"111000000",
  30002=>"000010010",
  30003=>"000000100",
  30004=>"000000000",
  30005=>"000000111",
  30006=>"110110111",
  30007=>"001000000",
  30008=>"101000000",
  30009=>"100000100",
  30010=>"110110110",
  30011=>"000000000",
  30012=>"000000000",
  30013=>"111111111",
  30014=>"111111111",
  30015=>"111111111",
  30016=>"001000000",
  30017=>"110000000",
  30018=>"111111111",
  30019=>"110100000",
  30020=>"000000000",
  30021=>"000000000",
  30022=>"111111111",
  30023=>"000000000",
  30024=>"000000000",
  30025=>"000000001",
  30026=>"000000000",
  30027=>"010010000",
  30028=>"111000111",
  30029=>"000001011",
  30030=>"111111111",
  30031=>"000000000",
  30032=>"000010111",
  30033=>"000000000",
  30034=>"110110111",
  30035=>"111111101",
  30036=>"000000000",
  30037=>"001000001",
  30038=>"000000000",
  30039=>"110111110",
  30040=>"111111111",
  30041=>"000011111",
  30042=>"111101010",
  30043=>"000000000",
  30044=>"000000000",
  30045=>"100000000",
  30046=>"000000000",
  30047=>"110111111",
  30048=>"000000000",
  30049=>"000000000",
  30050=>"000000000",
  30051=>"000000000",
  30052=>"011011000",
  30053=>"000000000",
  30054=>"000000010",
  30055=>"111111111",
  30056=>"001011111",
  30057=>"000000000",
  30058=>"001001001",
  30059=>"111111001",
  30060=>"001001111",
  30061=>"010000000",
  30062=>"111110110",
  30063=>"000000000",
  30064=>"111011111",
  30065=>"000000000",
  30066=>"010001111",
  30067=>"111001001",
  30068=>"000110111",
  30069=>"000000000",
  30070=>"000000000",
  30071=>"000000111",
  30072=>"000000000",
  30073=>"111000000",
  30074=>"111110000",
  30075=>"000000000",
  30076=>"000001000",
  30077=>"111111111",
  30078=>"100100100",
  30079=>"000000001",
  30080=>"100000000",
  30081=>"100001111",
  30082=>"100000000",
  30083=>"111100110",
  30084=>"000000000",
  30085=>"111111111",
  30086=>"100100100",
  30087=>"110100110",
  30088=>"000000000",
  30089=>"011000000",
  30090=>"110100000",
  30091=>"000000000",
  30092=>"000000001",
  30093=>"000000000",
  30094=>"000001011",
  30095=>"111111111",
  30096=>"000000000",
  30097=>"111111111",
  30098=>"101000000",
  30099=>"000000000",
  30100=>"111111000",
  30101=>"000000000",
  30102=>"111011010",
  30103=>"000011011",
  30104=>"111111111",
  30105=>"111110110",
  30106=>"000000000",
  30107=>"000010111",
  30108=>"111100100",
  30109=>"111111101",
  30110=>"000000000",
  30111=>"000011100",
  30112=>"100101111",
  30113=>"000011011",
  30114=>"111000101",
  30115=>"001001111",
  30116=>"001001000",
  30117=>"000000001",
  30118=>"111111111",
  30119=>"001111101",
  30120=>"000000000",
  30121=>"000000100",
  30122=>"110111111",
  30123=>"001000011",
  30124=>"000000000",
  30125=>"000000000",
  30126=>"000000000",
  30127=>"010101000",
  30128=>"111111000",
  30129=>"000000001",
  30130=>"000000000",
  30131=>"111100000",
  30132=>"111011001",
  30133=>"000000000",
  30134=>"000000000",
  30135=>"110111111",
  30136=>"000000000",
  30137=>"111111001",
  30138=>"000100100",
  30139=>"111111111",
  30140=>"111111111",
  30141=>"000000111",
  30142=>"000000101",
  30143=>"000000000",
  30144=>"000000000",
  30145=>"000000001",
  30146=>"111111111",
  30147=>"110111001",
  30148=>"001001001",
  30149=>"100011001",
  30150=>"001001001",
  30151=>"111101001",
  30152=>"000111111",
  30153=>"110110100",
  30154=>"000000000",
  30155=>"000100000",
  30156=>"111000000",
  30157=>"000000000",
  30158=>"111000001",
  30159=>"000001001",
  30160=>"000111000",
  30161=>"001011111",
  30162=>"110100000",
  30163=>"000010111",
  30164=>"111111111",
  30165=>"100111000",
  30166=>"100100101",
  30167=>"111100100",
  30168=>"000000000",
  30169=>"100000001",
  30170=>"000000111",
  30171=>"111111011",
  30172=>"111111111",
  30173=>"111111111",
  30174=>"000000010",
  30175=>"000000000",
  30176=>"000000000",
  30177=>"111110100",
  30178=>"111111111",
  30179=>"000111100",
  30180=>"111111011",
  30181=>"110010000",
  30182=>"111111111",
  30183=>"000000100",
  30184=>"000000111",
  30185=>"011111000",
  30186=>"000100101",
  30187=>"111111011",
  30188=>"000000001",
  30189=>"001001111",
  30190=>"001000000",
  30191=>"000000010",
  30192=>"000010011",
  30193=>"010011111",
  30194=>"000111111",
  30195=>"001001001",
  30196=>"000001010",
  30197=>"000000010",
  30198=>"000000011",
  30199=>"100100110",
  30200=>"000000000",
  30201=>"010000001",
  30202=>"111101111",
  30203=>"111100111",
  30204=>"000000000",
  30205=>"000011111",
  30206=>"011111111",
  30207=>"000000000",
  30208=>"001000000",
  30209=>"000000000",
  30210=>"111111111",
  30211=>"001000000",
  30212=>"000000000",
  30213=>"110111010",
  30214=>"011001101",
  30215=>"111001001",
  30216=>"111101001",
  30217=>"100100000",
  30218=>"110110000",
  30219=>"000100111",
  30220=>"001000010",
  30221=>"111100000",
  30222=>"110100111",
  30223=>"011010000",
  30224=>"000001111",
  30225=>"011111110",
  30226=>"111010110",
  30227=>"000000011",
  30228=>"101000000",
  30229=>"000000100",
  30230=>"110000000",
  30231=>"110010111",
  30232=>"000000110",
  30233=>"100110110",
  30234=>"000000000",
  30235=>"000000000",
  30236=>"111111111",
  30237=>"111111111",
  30238=>"010110001",
  30239=>"010000000",
  30240=>"001101111",
  30241=>"011001001",
  30242=>"110000000",
  30243=>"001101111",
  30244=>"000000000",
  30245=>"111000001",
  30246=>"010001111",
  30247=>"110000000",
  30248=>"111111111",
  30249=>"100000000",
  30250=>"001000000",
  30251=>"000000000",
  30252=>"111111111",
  30253=>"111111111",
  30254=>"111001111",
  30255=>"100000000",
  30256=>"111111011",
  30257=>"000000100",
  30258=>"011011011",
  30259=>"111111011",
  30260=>"111111111",
  30261=>"001000000",
  30262=>"111000000",
  30263=>"100111001",
  30264=>"100101111",
  30265=>"000000001",
  30266=>"000000000",
  30267=>"000111111",
  30268=>"000000000",
  30269=>"000000000",
  30270=>"000000000",
  30271=>"111110111",
  30272=>"111010010",
  30273=>"011011011",
  30274=>"000000001",
  30275=>"000000100",
  30276=>"011000000",
  30277=>"000110110",
  30278=>"011001011",
  30279=>"001001001",
  30280=>"111111111",
  30281=>"100000000",
  30282=>"101111110",
  30283=>"001000000",
  30284=>"110110000",
  30285=>"000000111",
  30286=>"101100110",
  30287=>"010000000",
  30288=>"111011000",
  30289=>"100100000",
  30290=>"111111111",
  30291=>"100111111",
  30292=>"011111111",
  30293=>"100000111",
  30294=>"110000000",
  30295=>"000100000",
  30296=>"111011010",
  30297=>"111100000",
  30298=>"000000100",
  30299=>"111111000",
  30300=>"001000000",
  30301=>"101001111",
  30302=>"010010110",
  30303=>"011011111",
  30304=>"111000000",
  30305=>"111111000",
  30306=>"100011111",
  30307=>"000000000",
  30308=>"111011111",
  30309=>"111111111",
  30310=>"000000000",
  30311=>"001001001",
  30312=>"000000111",
  30313=>"111111001",
  30314=>"110110110",
  30315=>"000111111",
  30316=>"010011001",
  30317=>"011000001",
  30318=>"111111111",
  30319=>"000000110",
  30320=>"110110111",
  30321=>"000001011",
  30322=>"111111001",
  30323=>"111101101",
  30324=>"111111111",
  30325=>"111111111",
  30326=>"101111011",
  30327=>"000000000",
  30328=>"111101111",
  30329=>"111110111",
  30330=>"011101101",
  30331=>"000000000",
  30332=>"111111111",
  30333=>"111111111",
  30334=>"101001111",
  30335=>"000000000",
  30336=>"011001111",
  30337=>"111111011",
  30338=>"000000000",
  30339=>"111011001",
  30340=>"111111110",
  30341=>"000000000",
  30342=>"110000010",
  30343=>"011011010",
  30344=>"000000000",
  30345=>"111111111",
  30346=>"111111100",
  30347=>"011000000",
  30348=>"111111111",
  30349=>"000000000",
  30350=>"010000100",
  30351=>"110111101",
  30352=>"111111111",
  30353=>"100000001",
  30354=>"101100110",
  30355=>"000000001",
  30356=>"001001001",
  30357=>"100100000",
  30358=>"111111111",
  30359=>"000000100",
  30360=>"000000000",
  30361=>"111111100",
  30362=>"000000000",
  30363=>"001000000",
  30364=>"000000000",
  30365=>"111111110",
  30366=>"010110111",
  30367=>"010111111",
  30368=>"001111111",
  30369=>"000000100",
  30370=>"111111111",
  30371=>"111111110",
  30372=>"111001001",
  30373=>"011001011",
  30374=>"001001111",
  30375=>"111111110",
  30376=>"000000000",
  30377=>"101111111",
  30378=>"111100000",
  30379=>"000000000",
  30380=>"101001111",
  30381=>"111001000",
  30382=>"101001011",
  30383=>"100111111",
  30384=>"000010000",
  30385=>"111001101",
  30386=>"001001000",
  30387=>"000000111",
  30388=>"001111000",
  30389=>"000000100",
  30390=>"000000000",
  30391=>"000000011",
  30392=>"101100000",
  30393=>"111100000",
  30394=>"001001000",
  30395=>"100001001",
  30396=>"100000000",
  30397=>"000100100",
  30398=>"111011000",
  30399=>"000001000",
  30400=>"010010010",
  30401=>"100100011",
  30402=>"001001000",
  30403=>"001011111",
  30404=>"111111111",
  30405=>"111111001",
  30406=>"001111011",
  30407=>"010000010",
  30408=>"111010111",
  30409=>"110110111",
  30410=>"000000110",
  30411=>"000000000",
  30412=>"000000000",
  30413=>"000000011",
  30414=>"000100110",
  30415=>"000000001",
  30416=>"000111111",
  30417=>"001101111",
  30418=>"010111100",
  30419=>"011000000",
  30420=>"111111111",
  30421=>"110001111",
  30422=>"111011000",
  30423=>"101000100",
  30424=>"101000101",
  30425=>"000110111",
  30426=>"111111111",
  30427=>"111000110",
  30428=>"110100111",
  30429=>"100000000",
  30430=>"000000001",
  30431=>"000000000",
  30432=>"010000000",
  30433=>"111000000",
  30434=>"111111110",
  30435=>"000000000",
  30436=>"001111110",
  30437=>"000001111",
  30438=>"111111001",
  30439=>"111001001",
  30440=>"001011000",
  30441=>"101101000",
  30442=>"111111001",
  30443=>"000000000",
  30444=>"111111111",
  30445=>"000000000",
  30446=>"111001000",
  30447=>"111111111",
  30448=>"000001011",
  30449=>"100000000",
  30450=>"000111111",
  30451=>"111100000",
  30452=>"001001101",
  30453=>"010111111",
  30454=>"101111111",
  30455=>"000000000",
  30456=>"000000000",
  30457=>"111111111",
  30458=>"110110111",
  30459=>"111111111",
  30460=>"000111111",
  30461=>"100100110",
  30462=>"111111111",
  30463=>"000000000",
  30464=>"111111111",
  30465=>"000001011",
  30466=>"011111000",
  30467=>"101000000",
  30468=>"000000000",
  30469=>"111110110",
  30470=>"011000110",
  30471=>"110000000",
  30472=>"100100010",
  30473=>"000000000",
  30474=>"000000000",
  30475=>"100100000",
  30476=>"000000000",
  30477=>"000000000",
  30478=>"111101111",
  30479=>"000000111",
  30480=>"000001111",
  30481=>"110111111",
  30482=>"111111110",
  30483=>"111111111",
  30484=>"000000000",
  30485=>"000111111",
  30486=>"110000010",
  30487=>"000001001",
  30488=>"110110011",
  30489=>"000111111",
  30490=>"000000000",
  30491=>"000000000",
  30492=>"110110011",
  30493=>"111111111",
  30494=>"111111000",
  30495=>"000000000",
  30496=>"111111111",
  30497=>"001001000",
  30498=>"100000111",
  30499=>"001011110",
  30500=>"100100101",
  30501=>"000000001",
  30502=>"110000000",
  30503=>"011111001",
  30504=>"111011111",
  30505=>"110000000",
  30506=>"111111111",
  30507=>"111111100",
  30508=>"100000110",
  30509=>"100100101",
  30510=>"111000000",
  30511=>"111111111",
  30512=>"100000000",
  30513=>"000000000",
  30514=>"111010000",
  30515=>"001000110",
  30516=>"111011001",
  30517=>"111101000",
  30518=>"100100111",
  30519=>"111111110",
  30520=>"000000111",
  30521=>"000001111",
  30522=>"111111101",
  30523=>"111000000",
  30524=>"010000000",
  30525=>"100100111",
  30526=>"000000100",
  30527=>"010110000",
  30528=>"001001111",
  30529=>"111111011",
  30530=>"000000000",
  30531=>"000000000",
  30532=>"101000000",
  30533=>"000000000",
  30534=>"000000101",
  30535=>"111111110",
  30536=>"000010000",
  30537=>"000000010",
  30538=>"110100100",
  30539=>"010000010",
  30540=>"000001001",
  30541=>"000000100",
  30542=>"110110111",
  30543=>"001001000",
  30544=>"000000000",
  30545=>"111000010",
  30546=>"111011011",
  30547=>"111111111",
  30548=>"000000000",
  30549=>"001111111",
  30550=>"111111000",
  30551=>"111111111",
  30552=>"000000000",
  30553=>"001001001",
  30554=>"000000100",
  30555=>"000000000",
  30556=>"111101000",
  30557=>"001000001",
  30558=>"011100000",
  30559=>"000000000",
  30560=>"111000000",
  30561=>"111111111",
  30562=>"000011011",
  30563=>"111111111",
  30564=>"100110111",
  30565=>"111111111",
  30566=>"111100000",
  30567=>"111101100",
  30568=>"110000011",
  30569=>"000001000",
  30570=>"011111001",
  30571=>"000111110",
  30572=>"100100100",
  30573=>"001001000",
  30574=>"111111001",
  30575=>"000000000",
  30576=>"111111110",
  30577=>"100100110",
  30578=>"111101000",
  30579=>"000110110",
  30580=>"111111001",
  30581=>"000000100",
  30582=>"111110000",
  30583=>"000000000",
  30584=>"001000000",
  30585=>"111111111",
  30586=>"111111000",
  30587=>"101111111",
  30588=>"000000011",
  30589=>"111000000",
  30590=>"111111111",
  30591=>"000000111",
  30592=>"111111110",
  30593=>"111101110",
  30594=>"001001111",
  30595=>"000000000",
  30596=>"100100000",
  30597=>"111111111",
  30598=>"000000000",
  30599=>"111111111",
  30600=>"111110000",
  30601=>"111111101",
  30602=>"000000000",
  30603=>"000000111",
  30604=>"100111111",
  30605=>"111110111",
  30606=>"000000000",
  30607=>"001000000",
  30608=>"000010010",
  30609=>"111111011",
  30610=>"011111110",
  30611=>"011001101",
  30612=>"111111111",
  30613=>"000000000",
  30614=>"000100111",
  30615=>"111111111",
  30616=>"000000010",
  30617=>"111111111",
  30618=>"000000000",
  30619=>"111111111",
  30620=>"001111111",
  30621=>"000000000",
  30622=>"000101111",
  30623=>"111111000",
  30624=>"001001101",
  30625=>"101011001",
  30626=>"111100100",
  30627=>"000111111",
  30628=>"111111111",
  30629=>"000000000",
  30630=>"011001000",
  30631=>"000010110",
  30632=>"011011011",
  30633=>"000000000",
  30634=>"000000000",
  30635=>"111001101",
  30636=>"000000000",
  30637=>"001111111",
  30638=>"111111001",
  30639=>"000111111",
  30640=>"111111111",
  30641=>"001000000",
  30642=>"100111101",
  30643=>"000000001",
  30644=>"100111111",
  30645=>"110111011",
  30646=>"100111111",
  30647=>"000000000",
  30648=>"000000011",
  30649=>"111111101",
  30650=>"000000000",
  30651=>"110000100",
  30652=>"000000000",
  30653=>"110000100",
  30654=>"001111111",
  30655=>"100000000",
  30656=>"111111000",
  30657=>"000010011",
  30658=>"111111111",
  30659=>"000000000",
  30660=>"011011110",
  30661=>"101101101",
  30662=>"101000001",
  30663=>"111111111",
  30664=>"111000111",
  30665=>"111110111",
  30666=>"100100000",
  30667=>"000000111",
  30668=>"000111111",
  30669=>"011001111",
  30670=>"001000000",
  30671=>"111111111",
  30672=>"000110110",
  30673=>"000000101",
  30674=>"001001001",
  30675=>"111111000",
  30676=>"100100110",
  30677=>"100000000",
  30678=>"101000100",
  30679=>"110110110",
  30680=>"111111000",
  30681=>"110110110",
  30682=>"000000000",
  30683=>"111011000",
  30684=>"000000000",
  30685=>"111100000",
  30686=>"000000000",
  30687=>"000000000",
  30688=>"011110110",
  30689=>"000000001",
  30690=>"000110111",
  30691=>"111110110",
  30692=>"010000101",
  30693=>"111111111",
  30694=>"011000011",
  30695=>"111101100",
  30696=>"111111111",
  30697=>"000000000",
  30698=>"111111101",
  30699=>"000010111",
  30700=>"000000011",
  30701=>"111111111",
  30702=>"011010000",
  30703=>"110000000",
  30704=>"111111111",
  30705=>"110111110",
  30706=>"010010011",
  30707=>"011001001",
  30708=>"111111111",
  30709=>"111111111",
  30710=>"111111111",
  30711=>"111001110",
  30712=>"010111111",
  30713=>"010001001",
  30714=>"110110111",
  30715=>"000110000",
  30716=>"011011111",
  30717=>"111111111",
  30718=>"111111100",
  30719=>"000001111",
  30720=>"000000000",
  30721=>"111000000",
  30722=>"000100000",
  30723=>"111101111",
  30724=>"001000000",
  30725=>"000101111",
  30726=>"000000000",
  30727=>"000000110",
  30728=>"111111011",
  30729=>"111000000",
  30730=>"011000000",
  30731=>"111111101",
  30732=>"111110000",
  30733=>"111111000",
  30734=>"111101000",
  30735=>"111100100",
  30736=>"011011001",
  30737=>"111000000",
  30738=>"000000111",
  30739=>"111111111",
  30740=>"000110000",
  30741=>"000000000",
  30742=>"000000000",
  30743=>"001011111",
  30744=>"000111111",
  30745=>"111011000",
  30746=>"001101001",
  30747=>"111111000",
  30748=>"011111111",
  30749=>"111111111",
  30750=>"000100010",
  30751=>"111011011",
  30752=>"111101101",
  30753=>"111111110",
  30754=>"000000101",
  30755=>"000000000",
  30756=>"111000001",
  30757=>"111000000",
  30758=>"001101100",
  30759=>"000011010",
  30760=>"000001001",
  30761=>"000000000",
  30762=>"101111111",
  30763=>"000001001",
  30764=>"111111111",
  30765=>"100111111",
  30766=>"110000001",
  30767=>"111111111",
  30768=>"111111101",
  30769=>"111000010",
  30770=>"010000100",
  30771=>"000111100",
  30772=>"111111111",
  30773=>"110111111",
  30774=>"010100011",
  30775=>"000001011",
  30776=>"101111000",
  30777=>"000111111",
  30778=>"000000000",
  30779=>"011000011",
  30780=>"001001111",
  30781=>"000010011",
  30782=>"110000000",
  30783=>"000100110",
  30784=>"111101000",
  30785=>"000000000",
  30786=>"100000000",
  30787=>"000000000",
  30788=>"011001001",
  30789=>"000000000",
  30790=>"001011000",
  30791=>"111111111",
  30792=>"111111110",
  30793=>"000000000",
  30794=>"011000000",
  30795=>"000000001",
  30796=>"000000000",
  30797=>"111010000",
  30798=>"000001001",
  30799=>"111011011",
  30800=>"000111111",
  30801=>"011011011",
  30802=>"000000000",
  30803=>"000010010",
  30804=>"111110110",
  30805=>"100000100",
  30806=>"000111111",
  30807=>"000000100",
  30808=>"111111111",
  30809=>"001000111",
  30810=>"000100111",
  30811=>"111001001",
  30812=>"000000000",
  30813=>"111111111",
  30814=>"011111000",
  30815=>"111010111",
  30816=>"000000001",
  30817=>"000000000",
  30818=>"000000000",
  30819=>"100111111",
  30820=>"011011000",
  30821=>"000000001",
  30822=>"101100000",
  30823=>"111111111",
  30824=>"000000011",
  30825=>"000000000",
  30826=>"000000000",
  30827=>"101100110",
  30828=>"000000000",
  30829=>"000000000",
  30830=>"000000000",
  30831=>"111011000",
  30832=>"111100000",
  30833=>"000001000",
  30834=>"111111111",
  30835=>"111111111",
  30836=>"000000000",
  30837=>"000000110",
  30838=>"100100000",
  30839=>"111111111",
  30840=>"111111111",
  30841=>"000111100",
  30842=>"010000000",
  30843=>"000000100",
  30844=>"100100110",
  30845=>"110111111",
  30846=>"010000000",
  30847=>"000000000",
  30848=>"000000000",
  30849=>"000100100",
  30850=>"000000111",
  30851=>"000111100",
  30852=>"111100100",
  30853=>"111111000",
  30854=>"000000000",
  30855=>"110001000",
  30856=>"011011111",
  30857=>"000000000",
  30858=>"000000000",
  30859=>"111011011",
  30860=>"100111111",
  30861=>"111011010",
  30862=>"000110001",
  30863=>"111111111",
  30864=>"100111111",
  30865=>"111111111",
  30866=>"000000000",
  30867=>"010000010",
  30868=>"001111000",
  30869=>"111011000",
  30870=>"000101001",
  30871=>"000000000",
  30872=>"111111100",
  30873=>"000110111",
  30874=>"111111111",
  30875=>"000000000",
  30876=>"100111111",
  30877=>"000000000",
  30878=>"000100110",
  30879=>"111111111",
  30880=>"100000000",
  30881=>"011001000",
  30882=>"000000000",
  30883=>"000000111",
  30884=>"110110000",
  30885=>"000011000",
  30886=>"000000000",
  30887=>"011000111",
  30888=>"000111100",
  30889=>"000000000",
  30890=>"111111111",
  30891=>"100000000",
  30892=>"110110111",
  30893=>"101100000",
  30894=>"111111111",
  30895=>"111011001",
  30896=>"000000000",
  30897=>"111111000",
  30898=>"111111111",
  30899=>"010011111",
  30900=>"111111000",
  30901=>"111111100",
  30902=>"000000000",
  30903=>"111111010",
  30904=>"111111111",
  30905=>"000110100",
  30906=>"110000100",
  30907=>"011110000",
  30908=>"111111011",
  30909=>"000111001",
  30910=>"010000000",
  30911=>"001001000",
  30912=>"000011111",
  30913=>"111111111",
  30914=>"111101000",
  30915=>"011000000",
  30916=>"000000000",
  30917=>"000000101",
  30918=>"010011111",
  30919=>"111111000",
  30920=>"010111000",
  30921=>"011111110",
  30922=>"111111111",
  30923=>"011010111",
  30924=>"001111101",
  30925=>"111111111",
  30926=>"111111110",
  30927=>"010011110",
  30928=>"111111001",
  30929=>"000000000",
  30930=>"111111000",
  30931=>"000000000",
  30932=>"110000101",
  30933=>"110100111",
  30934=>"000000000",
  30935=>"000000000",
  30936=>"000000100",
  30937=>"000111111",
  30938=>"000000111",
  30939=>"110111111",
  30940=>"000000100",
  30941=>"000000000",
  30942=>"111111101",
  30943=>"001101101",
  30944=>"000000000",
  30945=>"111110110",
  30946=>"110111110",
  30947=>"110111111",
  30948=>"010000000",
  30949=>"111110100",
  30950=>"000000000",
  30951=>"000000000",
  30952=>"000000000",
  30953=>"111111100",
  30954=>"111011001",
  30955=>"101111111",
  30956=>"111111001",
  30957=>"111111111",
  30958=>"111111111",
  30959=>"000001000",
  30960=>"100000111",
  30961=>"000100001",
  30962=>"011111000",
  30963=>"000000000",
  30964=>"111111111",
  30965=>"111111111",
  30966=>"101010000",
  30967=>"000000000",
  30968=>"111111111",
  30969=>"000101101",
  30970=>"000000000",
  30971=>"010011001",
  30972=>"111100110",
  30973=>"110011011",
  30974=>"000100100",
  30975=>"000000111",
  30976=>"000011111",
  30977=>"100110100",
  30978=>"111111111",
  30979=>"111111000",
  30980=>"000000000",
  30981=>"000000000",
  30982=>"000000000",
  30983=>"001111000",
  30984=>"110111110",
  30985=>"110000000",
  30986=>"111111111",
  30987=>"000111111",
  30988=>"111111111",
  30989=>"010111111",
  30990=>"000111000",
  30991=>"100000111",
  30992=>"110111111",
  30993=>"111000000",
  30994=>"000000010",
  30995=>"000011111",
  30996=>"010001111",
  30997=>"111111111",
  30998=>"100100111",
  30999=>"111111111",
  31000=>"110010001",
  31001=>"000000000",
  31002=>"111111000",
  31003=>"000000100",
  31004=>"110010110",
  31005=>"000000000",
  31006=>"000000000",
  31007=>"111100000",
  31008=>"111111100",
  31009=>"111001100",
  31010=>"000100100",
  31011=>"000000000",
  31012=>"110110110",
  31013=>"111111111",
  31014=>"000000000",
  31015=>"011010011",
  31016=>"111000100",
  31017=>"111111111",
  31018=>"000000000",
  31019=>"101100101",
  31020=>"111101111",
  31021=>"010000111",
  31022=>"100000000",
  31023=>"011010000",
  31024=>"000000000",
  31025=>"000000000",
  31026=>"011110000",
  31027=>"100101111",
  31028=>"000000000",
  31029=>"101000000",
  31030=>"000000111",
  31031=>"111111111",
  31032=>"111001001",
  31033=>"000101111",
  31034=>"000100110",
  31035=>"100101111",
  31036=>"000000000",
  31037=>"000000100",
  31038=>"111000000",
  31039=>"000000000",
  31040=>"000000000",
  31041=>"111111111",
  31042=>"000111000",
  31043=>"111111111",
  31044=>"000000000",
  31045=>"000100111",
  31046=>"111111111",
  31047=>"111100100",
  31048=>"000000000",
  31049=>"000000000",
  31050=>"111101000",
  31051=>"011111011",
  31052=>"000000101",
  31053=>"111011110",
  31054=>"000100110",
  31055=>"001001000",
  31056=>"001001001",
  31057=>"000001011",
  31058=>"001001111",
  31059=>"011110110",
  31060=>"000010010",
  31061=>"111011001",
  31062=>"110000000",
  31063=>"001111110",
  31064=>"000001010",
  31065=>"111100000",
  31066=>"110110110",
  31067=>"001111010",
  31068=>"001001001",
  31069=>"111111111",
  31070=>"000000000",
  31071=>"010110000",
  31072=>"000010000",
  31073=>"100110111",
  31074=>"111011000",
  31075=>"111111111",
  31076=>"110111111",
  31077=>"000110100",
  31078=>"111100100",
  31079=>"000000100",
  31080=>"100001101",
  31081=>"110000001",
  31082=>"000000001",
  31083=>"000010110",
  31084=>"110111111",
  31085=>"111111111",
  31086=>"011000000",
  31087=>"000000000",
  31088=>"000000000",
  31089=>"000000110",
  31090=>"111111000",
  31091=>"001000010",
  31092=>"001000101",
  31093=>"111111111",
  31094=>"000111111",
  31095=>"000110110",
  31096=>"000000111",
  31097=>"000000000",
  31098=>"010000000",
  31099=>"111101100",
  31100=>"000111010",
  31101=>"000011111",
  31102=>"100000000",
  31103=>"000000010",
  31104=>"111111011",
  31105=>"001001011",
  31106=>"110100100",
  31107=>"110111100",
  31108=>"011111111",
  31109=>"111111111",
  31110=>"101100111",
  31111=>"111110000",
  31112=>"111110111",
  31113=>"000011011",
  31114=>"000000111",
  31115=>"010000000",
  31116=>"111111101",
  31117=>"000000000",
  31118=>"001000000",
  31119=>"111001001",
  31120=>"110110000",
  31121=>"011011011",
  31122=>"011111011",
  31123=>"000000010",
  31124=>"100101111",
  31125=>"010010011",
  31126=>"000000000",
  31127=>"110110110",
  31128=>"111111000",
  31129=>"110111110",
  31130=>"000100111",
  31131=>"000000000",
  31132=>"000000000",
  31133=>"111111111",
  31134=>"111000111",
  31135=>"000000000",
  31136=>"111111111",
  31137=>"011111111",
  31138=>"000000100",
  31139=>"000110111",
  31140=>"000111111",
  31141=>"111111111",
  31142=>"000000000",
  31143=>"101111000",
  31144=>"111011000",
  31145=>"111111100",
  31146=>"000000000",
  31147=>"000000001",
  31148=>"110000000",
  31149=>"000000000",
  31150=>"000110111",
  31151=>"000011000",
  31152=>"110100000",
  31153=>"111111111",
  31154=>"011001000",
  31155=>"101000000",
  31156=>"000001000",
  31157=>"010000010",
  31158=>"000000011",
  31159=>"011000000",
  31160=>"000000000",
  31161=>"111000000",
  31162=>"111011000",
  31163=>"000000100",
  31164=>"011001111",
  31165=>"100110010",
  31166=>"000000001",
  31167=>"111111110",
  31168=>"111110100",
  31169=>"110011111",
  31170=>"111111111",
  31171=>"000000000",
  31172=>"000111111",
  31173=>"000101000",
  31174=>"101101000",
  31175=>"000001001",
  31176=>"000000000",
  31177=>"111001000",
  31178=>"000000000",
  31179=>"111111111",
  31180=>"000000000",
  31181=>"011111111",
  31182=>"001000000",
  31183=>"100100000",
  31184=>"100111011",
  31185=>"010110111",
  31186=>"100000111",
  31187=>"000111111",
  31188=>"000100001",
  31189=>"000000000",
  31190=>"100100101",
  31191=>"000000000",
  31192=>"000000110",
  31193=>"000110110",
  31194=>"011110000",
  31195=>"111111111",
  31196=>"000000000",
  31197=>"001111111",
  31198=>"111111000",
  31199=>"111100110",
  31200=>"100000001",
  31201=>"111111111",
  31202=>"111000100",
  31203=>"111111111",
  31204=>"111100101",
  31205=>"111111111",
  31206=>"000000000",
  31207=>"000000011",
  31208=>"111110111",
  31209=>"000000000",
  31210=>"000000000",
  31211=>"010111110",
  31212=>"111011001",
  31213=>"000000011",
  31214=>"111111111",
  31215=>"001000111",
  31216=>"000000010",
  31217=>"111111111",
  31218=>"001011000",
  31219=>"101101101",
  31220=>"000000100",
  31221=>"111001001",
  31222=>"000000000",
  31223=>"110100100",
  31224=>"010000111",
  31225=>"111101111",
  31226=>"000000111",
  31227=>"000000000",
  31228=>"000000111",
  31229=>"111111111",
  31230=>"000110000",
  31231=>"100111111",
  31232=>"100010110",
  31233=>"111111110",
  31234=>"010010000",
  31235=>"000000000",
  31236=>"000010000",
  31237=>"111111111",
  31238=>"111101001",
  31239=>"000000000",
  31240=>"110111000",
  31241=>"111001101",
  31242=>"100000000",
  31243=>"000000101",
  31244=>"001001111",
  31245=>"100000110",
  31246=>"000010100",
  31247=>"001000100",
  31248=>"100111111",
  31249=>"111111111",
  31250=>"100111111",
  31251=>"100001011",
  31252=>"000000000",
  31253=>"111100111",
  31254=>"000000000",
  31255=>"101000100",
  31256=>"001001001",
  31257=>"111111111",
  31258=>"000000000",
  31259=>"110111111",
  31260=>"011010111",
  31261=>"000000000",
  31262=>"010011011",
  31263=>"000000000",
  31264=>"000000000",
  31265=>"111111111",
  31266=>"101001001",
  31267=>"111010000",
  31268=>"111111100",
  31269=>"111011010",
  31270=>"000000010",
  31271=>"000100100",
  31272=>"100110010",
  31273=>"000000011",
  31274=>"111101111",
  31275=>"011111100",
  31276=>"100000000",
  31277=>"000100000",
  31278=>"000011111",
  31279=>"111111111",
  31280=>"000000001",
  31281=>"111111111",
  31282=>"011001000",
  31283=>"111010000",
  31284=>"000000000",
  31285=>"000100111",
  31286=>"000100100",
  31287=>"110110110",
  31288=>"011011011",
  31289=>"110110111",
  31290=>"111101111",
  31291=>"110110000",
  31292=>"110110110",
  31293=>"101000000",
  31294=>"111111111",
  31295=>"111100000",
  31296=>"011111110",
  31297=>"000000000",
  31298=>"111111111",
  31299=>"100000000",
  31300=>"001001001",
  31301=>"111101111",
  31302=>"011111000",
  31303=>"111000000",
  31304=>"001100100",
  31305=>"111100010",
  31306=>"000001111",
  31307=>"100010001",
  31308=>"001111010",
  31309=>"011001001",
  31310=>"111001000",
  31311=>"001001101",
  31312=>"000000111",
  31313=>"100110110",
  31314=>"101111000",
  31315=>"110111111",
  31316=>"111101101",
  31317=>"011011001",
  31318=>"000000000",
  31319=>"000010000",
  31320=>"011111110",
  31321=>"000000000",
  31322=>"110110000",
  31323=>"100100100",
  31324=>"010001000",
  31325=>"100111111",
  31326=>"001001000",
  31327=>"001001000",
  31328=>"000000011",
  31329=>"011000000",
  31330=>"111111111",
  31331=>"110110100",
  31332=>"000001101",
  31333=>"011011000",
  31334=>"111110110",
  31335=>"110110110",
  31336=>"111011111",
  31337=>"000000000",
  31338=>"011111110",
  31339=>"000010001",
  31340=>"111111111",
  31341=>"111111111",
  31342=>"111111000",
  31343=>"011011001",
  31344=>"001001010",
  31345=>"000010000",
  31346=>"000000010",
  31347=>"000000000",
  31348=>"111111111",
  31349=>"101111101",
  31350=>"000000000",
  31351=>"111111111",
  31352=>"111111110",
  31353=>"000000000",
  31354=>"110110111",
  31355=>"111001010",
  31356=>"111101111",
  31357=>"001001111",
  31358=>"000000000",
  31359=>"111111000",
  31360=>"011111011",
  31361=>"101101101",
  31362=>"000001111",
  31363=>"011001111",
  31364=>"111100101",
  31365=>"100100111",
  31366=>"110000000",
  31367=>"101000000",
  31368=>"000000000",
  31369=>"001111111",
  31370=>"111101101",
  31371=>"111000000",
  31372=>"001010110",
  31373=>"101111111",
  31374=>"110000011",
  31375=>"101111111",
  31376=>"001011111",
  31377=>"011110000",
  31378=>"110111001",
  31379=>"011011011",
  31380=>"111111111",
  31381=>"101011000",
  31382=>"011011001",
  31383=>"111001001",
  31384=>"010000000",
  31385=>"100100100",
  31386=>"111111111",
  31387=>"000000000",
  31388=>"111010000",
  31389=>"000111111",
  31390=>"100000111",
  31391=>"111111111",
  31392=>"111111111",
  31393=>"010110000",
  31394=>"001001000",
  31395=>"100100110",
  31396=>"000100100",
  31397=>"111111111",
  31398=>"000000000",
  31399=>"011001011",
  31400=>"001100000",
  31401=>"111111111",
  31402=>"111111111",
  31403=>"000000000",
  31404=>"111110111",
  31405=>"111101100",
  31406=>"000010110",
  31407=>"011000000",
  31408=>"111111111",
  31409=>"011011111",
  31410=>"000000000",
  31411=>"000000000",
  31412=>"000000000",
  31413=>"011010001",
  31414=>"001000000",
  31415=>"111100000",
  31416=>"000010110",
  31417=>"000000000",
  31418=>"100101100",
  31419=>"101101100",
  31420=>"111111101",
  31421=>"011111001",
  31422=>"011111111",
  31423=>"111111110",
  31424=>"111110100",
  31425=>"001011010",
  31426=>"000000000",
  31427=>"001001111",
  31428=>"110111000",
  31429=>"000000000",
  31430=>"100110111",
  31431=>"100000000",
  31432=>"000000011",
  31433=>"100100000",
  31434=>"000011111",
  31435=>"111001000",
  31436=>"111111110",
  31437=>"111001111",
  31438=>"111101111",
  31439=>"011001111",
  31440=>"111111111",
  31441=>"010010000",
  31442=>"111111111",
  31443=>"111111111",
  31444=>"111111100",
  31445=>"111111111",
  31446=>"000000110",
  31447=>"111111111",
  31448=>"000001000",
  31449=>"101100100",
  31450=>"010010000",
  31451=>"111001000",
  31452=>"000000100",
  31453=>"000000001",
  31454=>"000100100",
  31455=>"111000000",
  31456=>"110100100",
  31457=>"000000000",
  31458=>"000000000",
  31459=>"111000000",
  31460=>"000001111",
  31461=>"000000000",
  31462=>"000000000",
  31463=>"100000000",
  31464=>"100110100",
  31465=>"110100000",
  31466=>"111111000",
  31467=>"101101111",
  31468=>"000000000",
  31469=>"111111111",
  31470=>"000000111",
  31471=>"100100000",
  31472=>"000000100",
  31473=>"011010111",
  31474=>"111111101",
  31475=>"111011011",
  31476=>"111100000",
  31477=>"110010010",
  31478=>"001001011",
  31479=>"000000000",
  31480=>"100000100",
  31481=>"111110100",
  31482=>"111011111",
  31483=>"110110110",
  31484=>"110111101",
  31485=>"000100100",
  31486=>"001000111",
  31487=>"111101100",
  31488=>"100000000",
  31489=>"001001011",
  31490=>"100111101",
  31491=>"111000000",
  31492=>"111111111",
  31493=>"011000011",
  31494=>"111111111",
  31495=>"000000100",
  31496=>"101000100",
  31497=>"111111000",
  31498=>"111111111",
  31499=>"100100100",
  31500=>"000000000",
  31501=>"100100000",
  31502=>"100111110",
  31503=>"000110111",
  31504=>"100111101",
  31505=>"011000001",
  31506=>"110010000",
  31507=>"111101001",
  31508=>"111111111",
  31509=>"000110000",
  31510=>"100110101",
  31511=>"111111000",
  31512=>"110110111",
  31513=>"111000000",
  31514=>"110110110",
  31515=>"110111111",
  31516=>"011001001",
  31517=>"001001111",
  31518=>"001001001",
  31519=>"000010000",
  31520=>"000110100",
  31521=>"100100000",
  31522=>"110100100",
  31523=>"011000000",
  31524=>"110111111",
  31525=>"101111101",
  31526=>"100000000",
  31527=>"000100111",
  31528=>"100111111",
  31529=>"000100111",
  31530=>"000000000",
  31531=>"000001001",
  31532=>"000000000",
  31533=>"000010000",
  31534=>"000010000",
  31535=>"000110100",
  31536=>"111111111",
  31537=>"100100000",
  31538=>"000000000",
  31539=>"011111111",
  31540=>"000000010",
  31541=>"001001001",
  31542=>"110111011",
  31543=>"111100000",
  31544=>"110110111",
  31545=>"111011010",
  31546=>"111111111",
  31547=>"000000001",
  31548=>"111111111",
  31549=>"111001110",
  31550=>"000000000",
  31551=>"101100000",
  31552=>"001001111",
  31553=>"100000000",
  31554=>"111000000",
  31555=>"010000010",
  31556=>"000110110",
  31557=>"111111111",
  31558=>"111111111",
  31559=>"000000000",
  31560=>"000000000",
  31561=>"011011000",
  31562=>"010011011",
  31563=>"000000000",
  31564=>"110111111",
  31565=>"011111110",
  31566=>"111111111",
  31567=>"000110110",
  31568=>"001101111",
  31569=>"111111100",
  31570=>"011010110",
  31571=>"111100000",
  31572=>"100000000",
  31573=>"011101101",
  31574=>"100011111",
  31575=>"000000001",
  31576=>"010010000",
  31577=>"100100000",
  31578=>"111111110",
  31579=>"000000000",
  31580=>"111111111",
  31581=>"111111111",
  31582=>"111111111",
  31583=>"000100000",
  31584=>"010001011",
  31585=>"011001001",
  31586=>"000010011",
  31587=>"000000000",
  31588=>"000000001",
  31589=>"100110100",
  31590=>"110110000",
  31591=>"101100100",
  31592=>"010100111",
  31593=>"001000000",
  31594=>"001001011",
  31595=>"000000000",
  31596=>"011000101",
  31597=>"010000100",
  31598=>"111101100",
  31599=>"001001000",
  31600=>"111011111",
  31601=>"001001101",
  31602=>"000111110",
  31603=>"100100110",
  31604=>"111111111",
  31605=>"111111111",
  31606=>"111111111",
  31607=>"111110100",
  31608=>"000000110",
  31609=>"101100000",
  31610=>"011011011",
  31611=>"110101111",
  31612=>"000110110",
  31613=>"111111111",
  31614=>"111111111",
  31615=>"111111111",
  31616=>"101001001",
  31617=>"100000101",
  31618=>"111101111",
  31619=>"011010000",
  31620=>"001011111",
  31621=>"000000100",
  31622=>"110110111",
  31623=>"111111111",
  31624=>"000000000",
  31625=>"111111111",
  31626=>"000010011",
  31627=>"000000000",
  31628=>"111111111",
  31629=>"110100111",
  31630=>"100100100",
  31631=>"000011111",
  31632=>"001111000",
  31633=>"111001001",
  31634=>"100111110",
  31635=>"111111111",
  31636=>"010111100",
  31637=>"101101111",
  31638=>"100111111",
  31639=>"111111101",
  31640=>"001000101",
  31641=>"000100100",
  31642=>"001000000",
  31643=>"111100111",
  31644=>"101001111",
  31645=>"100100011",
  31646=>"011011000",
  31647=>"111111111",
  31648=>"111011001",
  31649=>"011011011",
  31650=>"000000011",
  31651=>"111111011",
  31652=>"110011011",
  31653=>"011111111",
  31654=>"000000000",
  31655=>"000000000",
  31656=>"110110100",
  31657=>"111111111",
  31658=>"111111111",
  31659=>"111111111",
  31660=>"111111111",
  31661=>"001000011",
  31662=>"000000111",
  31663=>"001001001",
  31664=>"000010010",
  31665=>"000000000",
  31666=>"111111111",
  31667=>"101001000",
  31668=>"000000010",
  31669=>"010011011",
  31670=>"001011111",
  31671=>"111111111",
  31672=>"011111110",
  31673=>"101111111",
  31674=>"111110100",
  31675=>"000000000",
  31676=>"000100110",
  31677=>"110111110",
  31678=>"101000000",
  31679=>"110110110",
  31680=>"000000001",
  31681=>"000000000",
  31682=>"000000000",
  31683=>"000000000",
  31684=>"000010010",
  31685=>"110011111",
  31686=>"111101111",
  31687=>"000000000",
  31688=>"100000100",
  31689=>"100000000",
  31690=>"011111111",
  31691=>"000010111",
  31692=>"000000010",
  31693=>"000000000",
  31694=>"000000100",
  31695=>"000011011",
  31696=>"000000011",
  31697=>"000010010",
  31698=>"001111111",
  31699=>"000001001",
  31700=>"111111111",
  31701=>"110110000",
  31702=>"101001000",
  31703=>"110100100",
  31704=>"101000001",
  31705=>"111010000",
  31706=>"100000100",
  31707=>"000000100",
  31708=>"100100100",
  31709=>"110000000",
  31710=>"011111110",
  31711=>"101001000",
  31712=>"001011000",
  31713=>"100100000",
  31714=>"000000100",
  31715=>"100000001",
  31716=>"000011111",
  31717=>"100101101",
  31718=>"100000000",
  31719=>"011111111",
  31720=>"111011011",
  31721=>"000000001",
  31722=>"011011010",
  31723=>"110011001",
  31724=>"011010110",
  31725=>"011000000",
  31726=>"000011000",
  31727=>"110010010",
  31728=>"111011011",
  31729=>"011111111",
  31730=>"111001001",
  31731=>"000000100",
  31732=>"111111001",
  31733=>"011011011",
  31734=>"011001000",
  31735=>"110000000",
  31736=>"000100100",
  31737=>"000000000",
  31738=>"111001000",
  31739=>"000000000",
  31740=>"111111111",
  31741=>"111011011",
  31742=>"111011011",
  31743=>"001111101",
  31744=>"000001001",
  31745=>"000000001",
  31746=>"000000000",
  31747=>"111000000",
  31748=>"111100100",
  31749=>"110111111",
  31750=>"111001001",
  31751=>"111111111",
  31752=>"111101101",
  31753=>"110111110",
  31754=>"101101111",
  31755=>"000000110",
  31756=>"101001001",
  31757=>"001011001",
  31758=>"000100100",
  31759=>"000000001",
  31760=>"111010010",
  31761=>"000000000",
  31762=>"111101011",
  31763=>"000000000",
  31764=>"000000000",
  31765=>"001001000",
  31766=>"010000000",
  31767=>"000001011",
  31768=>"100001111",
  31769=>"110011001",
  31770=>"000000000",
  31771=>"000100100",
  31772=>"000000000",
  31773=>"111110110",
  31774=>"000000000",
  31775=>"000001101",
  31776=>"110110110",
  31777=>"000110110",
  31778=>"001101101",
  31779=>"000000000",
  31780=>"110110110",
  31781=>"001001000",
  31782=>"000000001",
  31783=>"111111001",
  31784=>"001001000",
  31785=>"000000000",
  31786=>"001001001",
  31787=>"001001000",
  31788=>"000100101",
  31789=>"111111010",
  31790=>"100101101",
  31791=>"111111111",
  31792=>"110110000",
  31793=>"000000100",
  31794=>"110100100",
  31795=>"101011000",
  31796=>"101101101",
  31797=>"110110000",
  31798=>"111001001",
  31799=>"001111110",
  31800=>"100001101",
  31801=>"000000000",
  31802=>"001001101",
  31803=>"100000001",
  31804=>"101111111",
  31805=>"011000011",
  31806=>"100100101",
  31807=>"111011000",
  31808=>"001101000",
  31809=>"000100000",
  31810=>"000100000",
  31811=>"000000000",
  31812=>"001001000",
  31813=>"001001000",
  31814=>"000001000",
  31815=>"000000000",
  31816=>"110100000",
  31817=>"111111111",
  31818=>"001001101",
  31819=>"110110010",
  31820=>"000000001",
  31821=>"010111111",
  31822=>"000010111",
  31823=>"000101111",
  31824=>"111000000",
  31825=>"111101111",
  31826=>"001000000",
  31827=>"111110110",
  31828=>"111110110",
  31829=>"110110010",
  31830=>"110110111",
  31831=>"110100000",
  31832=>"111100111",
  31833=>"111110111",
  31834=>"000000000",
  31835=>"000000001",
  31836=>"010110110",
  31837=>"001010001",
  31838=>"111111111",
  31839=>"110000000",
  31840=>"000000000",
  31841=>"000000000",
  31842=>"000001111",
  31843=>"001001001",
  31844=>"011010011",
  31845=>"110110010",
  31846=>"110010110",
  31847=>"001001000",
  31848=>"001100111",
  31849=>"011111111",
  31850=>"010000010",
  31851=>"000000000",
  31852=>"111111101",
  31853=>"000110100",
  31854=>"111101101",
  31855=>"001001001",
  31856=>"111000000",
  31857=>"111000000",
  31858=>"000001001",
  31859=>"000000110",
  31860=>"000000000",
  31861=>"000000011",
  31862=>"101111111",
  31863=>"111111111",
  31864=>"110110110",
  31865=>"010110011",
  31866=>"000000001",
  31867=>"000001000",
  31868=>"101101100",
  31869=>"100000000",
  31870=>"000001111",
  31871=>"000000100",
  31872=>"101111111",
  31873=>"110111111",
  31874=>"000011111",
  31875=>"011111111",
  31876=>"111111111",
  31877=>"111111111",
  31878=>"000000000",
  31879=>"111001101",
  31880=>"001000000",
  31881=>"000001101",
  31882=>"000001101",
  31883=>"000000001",
  31884=>"001001000",
  31885=>"000101001",
  31886=>"000111111",
  31887=>"110111011",
  31888=>"000000000",
  31889=>"110110000",
  31890=>"000000000",
  31891=>"001110110",
  31892=>"110100100",
  31893=>"100110110",
  31894=>"101001111",
  31895=>"111111101",
  31896=>"111111101",
  31897=>"000000000",
  31898=>"000000100",
  31899=>"000000000",
  31900=>"111110000",
  31901=>"000111110",
  31902=>"110110110",
  31903=>"000001000",
  31904=>"000000000",
  31905=>"001111111",
  31906=>"111111000",
  31907=>"111110111",
  31908=>"110011011",
  31909=>"110110110",
  31910=>"010110010",
  31911=>"001001001",
  31912=>"001011111",
  31913=>"010010010",
  31914=>"001111111",
  31915=>"111000000",
  31916=>"000000001",
  31917=>"000000000",
  31918=>"111000000",
  31919=>"110010111",
  31920=>"000111111",
  31921=>"111100000",
  31922=>"011111111",
  31923=>"000000000",
  31924=>"110110110",
  31925=>"000000011",
  31926=>"011001000",
  31927=>"011011011",
  31928=>"111111111",
  31929=>"101001111",
  31930=>"110000000",
  31931=>"110010110",
  31932=>"101101101",
  31933=>"011011111",
  31934=>"010011001",
  31935=>"010010000",
  31936=>"111111111",
  31937=>"111010111",
  31938=>"111110110",
  31939=>"110111010",
  31940=>"011011111",
  31941=>"000000000",
  31942=>"100000000",
  31943=>"010010000",
  31944=>"000000001",
  31945=>"101111011",
  31946=>"000001011",
  31947=>"111111111",
  31948=>"101101000",
  31949=>"001111111",
  31950=>"000110110",
  31951=>"110110011",
  31952=>"000111100",
  31953=>"000000001",
  31954=>"111111111",
  31955=>"000000000",
  31956=>"111110000",
  31957=>"010000000",
  31958=>"111111111",
  31959=>"111010010",
  31960=>"100101101",
  31961=>"111111111",
  31962=>"011001000",
  31963=>"111111111",
  31964=>"000000000",
  31965=>"100111111",
  31966=>"010010100",
  31967=>"110110010",
  31968=>"001110110",
  31969=>"111111110",
  31970=>"101000000",
  31971=>"101111101",
  31972=>"110110110",
  31973=>"001000000",
  31974=>"111010111",
  31975=>"101100111",
  31976=>"000000000",
  31977=>"111111001",
  31978=>"010111111",
  31979=>"000010010",
  31980=>"000000001",
  31981=>"000000101",
  31982=>"011000111",
  31983=>"000000111",
  31984=>"011011010",
  31985=>"111011000",
  31986=>"000001000",
  31987=>"110000001",
  31988=>"011010111",
  31989=>"001001001",
  31990=>"000110111",
  31991=>"101101111",
  31992=>"000000000",
  31993=>"000000000",
  31994=>"000111011",
  31995=>"110111101",
  31996=>"000000101",
  31997=>"000000000",
  31998=>"100000101",
  31999=>"110100110",
  32000=>"000011111",
  32001=>"001001011",
  32002=>"111111000",
  32003=>"000000000",
  32004=>"100001001",
  32005=>"111001000",
  32006=>"000111111",
  32007=>"110010010",
  32008=>"001001111",
  32009=>"111000000",
  32010=>"111101111",
  32011=>"111111111",
  32012=>"000000000",
  32013=>"110010010",
  32014=>"111111000",
  32015=>"000110110",
  32016=>"000010010",
  32017=>"000000100",
  32018=>"000000000",
  32019=>"001000000",
  32020=>"000000000",
  32021=>"100100000",
  32022=>"000101001",
  32023=>"111101111",
  32024=>"111110110",
  32025=>"110000000",
  32026=>"010010010",
  32027=>"100100111",
  32028=>"011011011",
  32029=>"111101101",
  32030=>"000001111",
  32031=>"000011111",
  32032=>"000000001",
  32033=>"011111111",
  32034=>"000111111",
  32035=>"000010010",
  32036=>"010011000",
  32037=>"111111101",
  32038=>"111011011",
  32039=>"110010110",
  32040=>"111011011",
  32041=>"101001000",
  32042=>"001000100",
  32043=>"001001001",
  32044=>"111000000",
  32045=>"100110100",
  32046=>"000111111",
  32047=>"111100100",
  32048=>"110110110",
  32049=>"000000000",
  32050=>"110000000",
  32051=>"000000111",
  32052=>"011111111",
  32053=>"111101001",
  32054=>"000000001",
  32055=>"000001101",
  32056=>"001111111",
  32057=>"101111001",
  32058=>"000000101",
  32059=>"000100000",
  32060=>"100000000",
  32061=>"000111111",
  32062=>"000000110",
  32063=>"110110110",
  32064=>"000000100",
  32065=>"010010010",
  32066=>"000000111",
  32067=>"101101101",
  32068=>"101111111",
  32069=>"110111000",
  32070=>"000110010",
  32071=>"111111001",
  32072=>"001001000",
  32073=>"010000111",
  32074=>"000100111",
  32075=>"100100100",
  32076=>"000000110",
  32077=>"001101001",
  32078=>"111111111",
  32079=>"001001111",
  32080=>"000000000",
  32081=>"110110110",
  32082=>"100010010",
  32083=>"111000100",
  32084=>"111111111",
  32085=>"001111001",
  32086=>"010110111",
  32087=>"000111111",
  32088=>"111111110",
  32089=>"000100000",
  32090=>"000000111",
  32091=>"001001000",
  32092=>"000000000",
  32093=>"001000000",
  32094=>"001111111",
  32095=>"110100000",
  32096=>"111100101",
  32097=>"010010000",
  32098=>"011000000",
  32099=>"111111101",
  32100=>"110111110",
  32101=>"110010110",
  32102=>"001000111",
  32103=>"000000000",
  32104=>"101001001",
  32105=>"110110110",
  32106=>"000100100",
  32107=>"001001001",
  32108=>"111111111",
  32109=>"000001000",
  32110=>"101101101",
  32111=>"000000011",
  32112=>"001011111",
  32113=>"100101111",
  32114=>"111101000",
  32115=>"001001101",
  32116=>"100100000",
  32117=>"110000100",
  32118=>"010000000",
  32119=>"101001001",
  32120=>"101101101",
  32121=>"000000111",
  32122=>"110100000",
  32123=>"011011011",
  32124=>"110110110",
  32125=>"110110010",
  32126=>"110111110",
  32127=>"111100101",
  32128=>"100111000",
  32129=>"110011000",
  32130=>"100100110",
  32131=>"010011011",
  32132=>"111111111",
  32133=>"000100111",
  32134=>"000000011",
  32135=>"101100111",
  32136=>"000000000",
  32137=>"011111111",
  32138=>"101111111",
  32139=>"110011110",
  32140=>"111111011",
  32141=>"111100000",
  32142=>"111101111",
  32143=>"111010111",
  32144=>"000000000",
  32145=>"101101111",
  32146=>"111100000",
  32147=>"001001001",
  32148=>"111111111",
  32149=>"000010000",
  32150=>"000000110",
  32151=>"111111110",
  32152=>"100001101",
  32153=>"000110111",
  32154=>"111111110",
  32155=>"111111100",
  32156=>"111101101",
  32157=>"000000001",
  32158=>"111110110",
  32159=>"000000100",
  32160=>"111000110",
  32161=>"011011011",
  32162=>"110100000",
  32163=>"100000000",
  32164=>"000000101",
  32165=>"111111101",
  32166=>"000000000",
  32167=>"000111111",
  32168=>"111111111",
  32169=>"000000000",
  32170=>"000000101",
  32171=>"111111111",
  32172=>"010111111",
  32173=>"001111111",
  32174=>"111101001",
  32175=>"110110111",
  32176=>"000000000",
  32177=>"111111111",
  32178=>"111111111",
  32179=>"000000000",
  32180=>"110110110",
  32181=>"111110011",
  32182=>"111110111",
  32183=>"001011000",
  32184=>"000000000",
  32185=>"000110100",
  32186=>"111011010",
  32187=>"111111111",
  32188=>"001001011",
  32189=>"111111010",
  32190=>"100001011",
  32191=>"110110010",
  32192=>"000000000",
  32193=>"101111111",
  32194=>"000010111",
  32195=>"000000000",
  32196=>"100000011",
  32197=>"000000000",
  32198=>"000000010",
  32199=>"101101101",
  32200=>"111010011",
  32201=>"000000000",
  32202=>"000000000",
  32203=>"011111111",
  32204=>"000000111",
  32205=>"111111111",
  32206=>"000111001",
  32207=>"000100100",
  32208=>"000000001",
  32209=>"111111011",
  32210=>"110110111",
  32211=>"111111011",
  32212=>"001000011",
  32213=>"000000111",
  32214=>"101111111",
  32215=>"011011001",
  32216=>"111101000",
  32217=>"110110110",
  32218=>"111111110",
  32219=>"111110111",
  32220=>"101101000",
  32221=>"110011010",
  32222=>"111111111",
  32223=>"110100000",
  32224=>"111111100",
  32225=>"111111011",
  32226=>"111111000",
  32227=>"000000011",
  32228=>"110000010",
  32229=>"000101011",
  32230=>"000000000",
  32231=>"000000000",
  32232=>"111010011",
  32233=>"000100110",
  32234=>"000000101",
  32235=>"101000000",
  32236=>"001001111",
  32237=>"011011011",
  32238=>"101101001",
  32239=>"111011011",
  32240=>"110000111",
  32241=>"000111110",
  32242=>"101100001",
  32243=>"110111111",
  32244=>"110110010",
  32245=>"000110010",
  32246=>"111111111",
  32247=>"110110110",
  32248=>"001111001",
  32249=>"011001001",
  32250=>"100101110",
  32251=>"001111111",
  32252=>"001001111",
  32253=>"010000011",
  32254=>"000000000",
  32255=>"001000001",
  32256=>"100100100",
  32257=>"000000100",
  32258=>"111000000",
  32259=>"000000000",
  32260=>"000000000",
  32261=>"000000000",
  32262=>"011111111",
  32263=>"111111111",
  32264=>"111110000",
  32265=>"110110000",
  32266=>"001000000",
  32267=>"111111111",
  32268=>"000000110",
  32269=>"100000000",
  32270=>"011000101",
  32271=>"000111011",
  32272=>"001001000",
  32273=>"000000111",
  32274=>"111111111",
  32275=>"000000000",
  32276=>"000011000",
  32277=>"000000010",
  32278=>"000101101",
  32279=>"101001011",
  32280=>"100100100",
  32281=>"001000000",
  32282=>"100000111",
  32283=>"110111101",
  32284=>"100111111",
  32285=>"000110001",
  32286=>"100000000",
  32287=>"111111100",
  32288=>"100000100",
  32289=>"111000000",
  32290=>"111111111",
  32291=>"111111111",
  32292=>"000000001",
  32293=>"111111111",
  32294=>"111011011",
  32295=>"110111111",
  32296=>"100111101",
  32297=>"110000000",
  32298=>"000000000",
  32299=>"111111111",
  32300=>"001001000",
  32301=>"111110110",
  32302=>"000000000",
  32303=>"111111111",
  32304=>"110100000",
  32305=>"000000100",
  32306=>"111001001",
  32307=>"000000011",
  32308=>"000001000",
  32309=>"000000000",
  32310=>"011111011",
  32311=>"110111011",
  32312=>"100111000",
  32313=>"100001000",
  32314=>"000011011",
  32315=>"000000111",
  32316=>"111101111",
  32317=>"001111000",
  32318=>"110110111",
  32319=>"110100111",
  32320=>"111111011",
  32321=>"010010010",
  32322=>"111111111",
  32323=>"111100111",
  32324=>"111111111",
  32325=>"000001000",
  32326=>"000000111",
  32327=>"110100000",
  32328=>"011111111",
  32329=>"000000111",
  32330=>"000000000",
  32331=>"101100100",
  32332=>"111111111",
  32333=>"000000000",
  32334=>"000000000",
  32335=>"001001000",
  32336=>"000000000",
  32337=>"011111110",
  32338=>"011010000",
  32339=>"000000000",
  32340=>"000000000",
  32341=>"111100110",
  32342=>"100100110",
  32343=>"000000000",
  32344=>"111111111",
  32345=>"000000111",
  32346=>"010110001",
  32347=>"001011111",
  32348=>"111111111",
  32349=>"000000000",
  32350=>"001001000",
  32351=>"011011011",
  32352=>"000011111",
  32353=>"111101101",
  32354=>"000000000",
  32355=>"111111101",
  32356=>"110110110",
  32357=>"111111111",
  32358=>"011111111",
  32359=>"000110111",
  32360=>"111111111",
  32361=>"000000111",
  32362=>"001011010",
  32363=>"000000011",
  32364=>"011111101",
  32365=>"111111111",
  32366=>"000000000",
  32367=>"000000010",
  32368=>"111111111",
  32369=>"111111111",
  32370=>"000000000",
  32371=>"000001000",
  32372=>"010111000",
  32373=>"001000011",
  32374=>"111111000",
  32375=>"001011111",
  32376=>"100100111",
  32377=>"111111111",
  32378=>"101000000",
  32379=>"111111111",
  32380=>"001011111",
  32381=>"111111011",
  32382=>"111101111",
  32383=>"000010010",
  32384=>"111111111",
  32385=>"111010000",
  32386=>"111111110",
  32387=>"000000000",
  32388=>"000000000",
  32389=>"000000000",
  32390=>"111111110",
  32391=>"101101111",
  32392=>"000000000",
  32393=>"001100100",
  32394=>"111111111",
  32395=>"000010011",
  32396=>"111110000",
  32397=>"000000000",
  32398=>"111111111",
  32399=>"000000000",
  32400=>"111111111",
  32401=>"000110111",
  32402=>"111101100",
  32403=>"111101001",
  32404=>"100000000",
  32405=>"110100101",
  32406=>"000000001",
  32407=>"000000000",
  32408=>"000000000",
  32409=>"100110110",
  32410=>"101110011",
  32411=>"111111000",
  32412=>"000000011",
  32413=>"101100001",
  32414=>"011111110",
  32415=>"000001000",
  32416=>"000000000",
  32417=>"111111111",
  32418=>"110110111",
  32419=>"100100011",
  32420=>"001001001",
  32421=>"000111111",
  32422=>"110100111",
  32423=>"000111111",
  32424=>"011111101",
  32425=>"010111111",
  32426=>"000000000",
  32427=>"000000000",
  32428=>"111111111",
  32429=>"000000110",
  32430=>"111001111",
  32431=>"000000000",
  32432=>"000110000",
  32433=>"101101101",
  32434=>"111111111",
  32435=>"010110110",
  32436=>"000001111",
  32437=>"000101101",
  32438=>"000000000",
  32439=>"000000000",
  32440=>"111111111",
  32441=>"111111111",
  32442=>"100100101",
  32443=>"100111111",
  32444=>"000000001",
  32445=>"111111111",
  32446=>"011110110",
  32447=>"111111111",
  32448=>"111100000",
  32449=>"000000001",
  32450=>"111111111",
  32451=>"000000000",
  32452=>"000000000",
  32453=>"000000000",
  32454=>"001000100",
  32455=>"101111010",
  32456=>"000010111",
  32457=>"101001000",
  32458=>"100000001",
  32459=>"111111011",
  32460=>"000111111",
  32461=>"000000100",
  32462=>"001001011",
  32463=>"100011001",
  32464=>"111100000",
  32465=>"111111011",
  32466=>"110100111",
  32467=>"111111000",
  32468=>"000000100",
  32469=>"111011011",
  32470=>"000000000",
  32471=>"000000000",
  32472=>"000000100",
  32473=>"111111111",
  32474=>"011111111",
  32475=>"011111111",
  32476=>"011111111",
  32477=>"000000110",
  32478=>"001001000",
  32479=>"000000000",
  32480=>"000000000",
  32481=>"010010010",
  32482=>"011001000",
  32483=>"111111111",
  32484=>"111111111",
  32485=>"010111011",
  32486=>"000000100",
  32487=>"110000100",
  32488=>"000000000",
  32489=>"100100100",
  32490=>"000000000",
  32491=>"100000001",
  32492=>"111111111",
  32493=>"000000000",
  32494=>"101000111",
  32495=>"110111111",
  32496=>"011100000",
  32497=>"110000000",
  32498=>"000000111",
  32499=>"000000000",
  32500=>"100001000",
  32501=>"110011000",
  32502=>"011011001",
  32503=>"000000000",
  32504=>"111111111",
  32505=>"111011011",
  32506=>"111111111",
  32507=>"001000111",
  32508=>"110100000",
  32509=>"011000000",
  32510=>"011111011",
  32511=>"111111111",
  32512=>"100000110",
  32513=>"100100011",
  32514=>"000000000",
  32515=>"100111111",
  32516=>"000001001",
  32517=>"000000001",
  32518=>"001000000",
  32519=>"101111111",
  32520=>"000000000",
  32521=>"111111011",
  32522=>"111111111",
  32523=>"000000000",
  32524=>"110100110",
  32525=>"101101000",
  32526=>"000000000",
  32527=>"111000000",
  32528=>"110110000",
  32529=>"000100111",
  32530=>"000000111",
  32531=>"000100100",
  32532=>"111000000",
  32533=>"000000000",
  32534=>"011011111",
  32535=>"000100000",
  32536=>"100000101",
  32537=>"111001000",
  32538=>"111111111",
  32539=>"011111111",
  32540=>"111111111",
  32541=>"110111011",
  32542=>"000000000",
  32543=>"000110110",
  32544=>"011011000",
  32545=>"000000000",
  32546=>"111111010",
  32547=>"111111111",
  32548=>"111110000",
  32549=>"000000000",
  32550=>"000011001",
  32551=>"001000000",
  32552=>"111000000",
  32553=>"000000000",
  32554=>"001111111",
  32555=>"111011010",
  32556=>"000000000",
  32557=>"000000000",
  32558=>"111110110",
  32559=>"000001011",
  32560=>"111111111",
  32561=>"000100110",
  32562=>"001001001",
  32563=>"011110000",
  32564=>"000000000",
  32565=>"101100110",
  32566=>"011010100",
  32567=>"111111000",
  32568=>"111011011",
  32569=>"100000000",
  32570=>"010111111",
  32571=>"111111111",
  32572=>"000001001",
  32573=>"000001111",
  32574=>"100100101",
  32575=>"000000110",
  32576=>"111111000",
  32577=>"000000000",
  32578=>"001101011",
  32579=>"000000000",
  32580=>"111111111",
  32581=>"111011001",
  32582=>"000000011",
  32583=>"000001111",
  32584=>"000000001",
  32585=>"000000000",
  32586=>"000100000",
  32587=>"001101111",
  32588=>"100100110",
  32589=>"111111110",
  32590=>"111111111",
  32591=>"111110110",
  32592=>"001111111",
  32593=>"001001111",
  32594=>"111000000",
  32595=>"111101000",
  32596=>"001000000",
  32597=>"011011011",
  32598=>"000000000",
  32599=>"111111111",
  32600=>"100000001",
  32601=>"110100111",
  32602=>"111001001",
  32603=>"011001001",
  32604=>"110110111",
  32605=>"000000000",
  32606=>"000000000",
  32607=>"001001001",
  32608=>"000000111",
  32609=>"111100101",
  32610=>"111111101",
  32611=>"101101111",
  32612=>"010110000",
  32613=>"000000000",
  32614=>"010000000",
  32615=>"001101110",
  32616=>"011011010",
  32617=>"010000000",
  32618=>"100000000",
  32619=>"111100111",
  32620=>"000100100",
  32621=>"000000000",
  32622=>"000000000",
  32623=>"000000000",
  32624=>"000101111",
  32625=>"010010011",
  32626=>"000101111",
  32627=>"111110111",
  32628=>"110110111",
  32629=>"110000001",
  32630=>"111111111",
  32631=>"100000000",
  32632=>"000000001",
  32633=>"111110000",
  32634=>"111101011",
  32635=>"110111110",
  32636=>"110100000",
  32637=>"101110111",
  32638=>"111110000",
  32639=>"000000000",
  32640=>"000000000",
  32641=>"001000001",
  32642=>"000000000",
  32643=>"000000000",
  32644=>"111111111",
  32645=>"011001111",
  32646=>"011101101",
  32647=>"000001001",
  32648=>"111111111",
  32649=>"111011011",
  32650=>"001001000",
  32651=>"000000000",
  32652=>"111111111",
  32653=>"100110111",
  32654=>"111111100",
  32655=>"000000000",
  32656=>"000000000",
  32657=>"011001000",
  32658=>"000100100",
  32659=>"000000000",
  32660=>"000000010",
  32661=>"000000000",
  32662=>"000000000",
  32663=>"000000000",
  32664=>"111111111",
  32665=>"111111111",
  32666=>"000000000",
  32667=>"000100100",
  32668=>"101000000",
  32669=>"000111110",
  32670=>"000000000",
  32671=>"000110111",
  32672=>"111111100",
  32673=>"111011011",
  32674=>"111111111",
  32675=>"111111111",
  32676=>"100111111",
  32677=>"111111010",
  32678=>"000000110",
  32679=>"111111101",
  32680=>"011111000",
  32681=>"111111110",
  32682=>"000000110",
  32683=>"000000000",
  32684=>"000000000",
  32685=>"000000000",
  32686=>"001001011",
  32687=>"111111110",
  32688=>"011011011",
  32689=>"001111111",
  32690=>"000000000",
  32691=>"000000000",
  32692=>"101111111",
  32693=>"011100110",
  32694=>"111000111",
  32695=>"000000000",
  32696=>"110111111",
  32697=>"101100000",
  32698=>"110111001",
  32699=>"000000001",
  32700=>"000011111",
  32701=>"111110111",
  32702=>"111110100",
  32703=>"001001001",
  32704=>"000000000",
  32705=>"000000000",
  32706=>"111110110",
  32707=>"111111000",
  32708=>"000000000",
  32709=>"000001111",
  32710=>"101100100",
  32711=>"011000000",
  32712=>"000000000",
  32713=>"100100110",
  32714=>"101111110",
  32715=>"110110000",
  32716=>"000000000",
  32717=>"001001001",
  32718=>"110100000",
  32719=>"111011011",
  32720=>"111111001",
  32721=>"100111111",
  32722=>"111110110",
  32723=>"000000110",
  32724=>"101111111",
  32725=>"000111100",
  32726=>"111100000",
  32727=>"001111111",
  32728=>"100000010",
  32729=>"111100000",
  32730=>"111000000",
  32731=>"111101000",
  32732=>"111000000",
  32733=>"100100011",
  32734=>"001100111",
  32735=>"000000011",
  32736=>"011000000",
  32737=>"101111011",
  32738=>"001111111",
  32739=>"011010111",
  32740=>"000000111",
  32741=>"011111110",
  32742=>"000001000",
  32743=>"111111111",
  32744=>"000000000",
  32745=>"000000011",
  32746=>"111111111",
  32747=>"000000000",
  32748=>"000100000",
  32749=>"000000000",
  32750=>"111111111",
  32751=>"000000100",
  32752=>"100000100",
  32753=>"011011011",
  32754=>"111111111",
  32755=>"000000000",
  32756=>"101100000",
  32757=>"000000100",
  32758=>"001101001",
  32759=>"111111001",
  32760=>"111111011",
  32761=>"000000000",
  32762=>"000000000",
  32763=>"111110000",
  32764=>"011010011",
  32765=>"011111010",
  32766=>"000000000",
  32767=>"001001100",
  32768=>"101101000",
  32769=>"110000000",
  32770=>"101111111",
  32771=>"000000000",
  32772=>"111111111",
  32773=>"000000000",
  32774=>"000000000",
  32775=>"111111011",
  32776=>"000001001",
  32777=>"000000000",
  32778=>"000000000",
  32779=>"101100000",
  32780=>"111111110",
  32781=>"000000000",
  32782=>"000000001",
  32783=>"111111111",
  32784=>"111111111",
  32785=>"111111111",
  32786=>"111111111",
  32787=>"111111111",
  32788=>"000000000",
  32789=>"000100110",
  32790=>"001111111",
  32791=>"111111111",
  32792=>"111111000",
  32793=>"100101011",
  32794=>"111111110",
  32795=>"111111001",
  32796=>"111111111",
  32797=>"000000000",
  32798=>"001100100",
  32799=>"001000000",
  32800=>"011100111",
  32801=>"001001111",
  32802=>"111111111",
  32803=>"000000000",
  32804=>"111111111",
  32805=>"111111111",
  32806=>"000111111",
  32807=>"111111100",
  32808=>"000000000",
  32809=>"000000000",
  32810=>"100100111",
  32811=>"001000000",
  32812=>"111001101",
  32813=>"000111110",
  32814=>"111111011",
  32815=>"001001000",
  32816=>"110111000",
  32817=>"001000000",
  32818=>"000101011",
  32819=>"110000000",
  32820=>"000000101",
  32821=>"011011111",
  32822=>"000111111",
  32823=>"001000000",
  32824=>"000000010",
  32825=>"111111111",
  32826=>"111111111",
  32827=>"111100000",
  32828=>"000001011",
  32829=>"000000000",
  32830=>"000000000",
  32831=>"000000000",
  32832=>"001011111",
  32833=>"110000000",
  32834=>"001001000",
  32835=>"001101111",
  32836=>"111001001",
  32837=>"001011111",
  32838=>"111111111",
  32839=>"000000000",
  32840=>"100100000",
  32841=>"110010000",
  32842=>"111111001",
  32843=>"111111110",
  32844=>"111000010",
  32845=>"000111111",
  32846=>"111000001",
  32847=>"100111111",
  32848=>"111111111",
  32849=>"011010000",
  32850=>"011000000",
  32851=>"100100111",
  32852=>"000100111",
  32853=>"000000000",
  32854=>"000111111",
  32855=>"000000100",
  32856=>"110100000",
  32857=>"100000000",
  32858=>"011010000",
  32859=>"100000000",
  32860=>"000000000",
  32861=>"000000000",
  32862=>"000000000",
  32863=>"001001011",
  32864=>"111001001",
  32865=>"000000000",
  32866=>"000000000",
  32867=>"111100000",
  32868=>"111111000",
  32869=>"001000000",
  32870=>"001111111",
  32871=>"111100111",
  32872=>"000000000",
  32873=>"100000000",
  32874=>"000000011",
  32875=>"110100000",
  32876=>"000000000",
  32877=>"111111111",
  32878=>"000101111",
  32879=>"011011110",
  32880=>"100110111",
  32881=>"000000000",
  32882=>"010000000",
  32883=>"110111110",
  32884=>"011111011",
  32885=>"111111111",
  32886=>"001000000",
  32887=>"000001000",
  32888=>"111111011",
  32889=>"001001111",
  32890=>"001000000",
  32891=>"111111111",
  32892=>"001111111",
  32893=>"101100000",
  32894=>"000000000",
  32895=>"000111000",
  32896=>"011001011",
  32897=>"111111000",
  32898=>"000010111",
  32899=>"100111110",
  32900=>"000010000",
  32901=>"000111111",
  32902=>"111111001",
  32903=>"111111000",
  32904=>"111110100",
  32905=>"111111111",
  32906=>"000000000",
  32907=>"111111010",
  32908=>"111110010",
  32909=>"111111111",
  32910=>"110111111",
  32911=>"111111110",
  32912=>"100100000",
  32913=>"000000000",
  32914=>"000111111",
  32915=>"000000000",
  32916=>"111111111",
  32917=>"111001001",
  32918=>"110111111",
  32919=>"000110000",
  32920=>"000000000",
  32921=>"101111010",
  32922=>"000000110",
  32923=>"000000000",
  32924=>"011001011",
  32925=>"100100001",
  32926=>"000001111",
  32927=>"001001000",
  32928=>"111111011",
  32929=>"000000000",
  32930=>"000000000",
  32931=>"111111111",
  32932=>"000000110",
  32933=>"011001000",
  32934=>"011000000",
  32935=>"110100100",
  32936=>"001111000",
  32937=>"000000000",
  32938=>"111111111",
  32939=>"111111000",
  32940=>"101111111",
  32941=>"000110010",
  32942=>"000100111",
  32943=>"000111111",
  32944=>"001111001",
  32945=>"011000100",
  32946=>"111111010",
  32947=>"000000000",
  32948=>"111111110",
  32949=>"001000000",
  32950=>"100000000",
  32951=>"111111111",
  32952=>"100100110",
  32953=>"111111111",
  32954=>"111100100",
  32955=>"011111100",
  32956=>"001000000",
  32957=>"001001000",
  32958=>"011000000",
  32959=>"001111111",
  32960=>"110100001",
  32961=>"111111011",
  32962=>"000000000",
  32963=>"111111011",
  32964=>"111111111",
  32965=>"000000000",
  32966=>"000100100",
  32967=>"100110110",
  32968=>"101111111",
  32969=>"011001000",
  32970=>"100011011",
  32971=>"111111111",
  32972=>"100100111",
  32973=>"101101111",
  32974=>"000111110",
  32975=>"000000000",
  32976=>"000110100",
  32977=>"111111111",
  32978=>"000110000",
  32979=>"001111111",
  32980=>"000000000",
  32981=>"000100000",
  32982=>"111001000",
  32983=>"001000000",
  32984=>"000001010",
  32985=>"000000000",
  32986=>"111111000",
  32987=>"000001001",
  32988=>"100100000",
  32989=>"000000000",
  32990=>"010010011",
  32991=>"011000000",
  32992=>"001111100",
  32993=>"011111111",
  32994=>"000000100",
  32995=>"000100000",
  32996=>"000000000",
  32997=>"001000011",
  32998=>"001000000",
  32999=>"111111111",
  33000=>"000110001",
  33001=>"000110000",
  33002=>"111111111",
  33003=>"000010010",
  33004=>"111111111",
  33005=>"000001111",
  33006=>"101111100",
  33007=>"000111010",
  33008=>"011101111",
  33009=>"001000000",
  33010=>"111000111",
  33011=>"100000001",
  33012=>"011000000",
  33013=>"111110110",
  33014=>"100000111",
  33015=>"111010111",
  33016=>"111111011",
  33017=>"000000011",
  33018=>"000111000",
  33019=>"010110111",
  33020=>"111111111",
  33021=>"000100110",
  33022=>"000010111",
  33023=>"111101000",
  33024=>"000000000",
  33025=>"110110110",
  33026=>"000000001",
  33027=>"000000110",
  33028=>"111111000",
  33029=>"110000000",
  33030=>"111111111",
  33031=>"011111000",
  33032=>"011111111",
  33033=>"000000011",
  33034=>"111110000",
  33035=>"111110000",
  33036=>"000000000",
  33037=>"100101111",
  33038=>"000000000",
  33039=>"001011000",
  33040=>"111011111",
  33041=>"111001000",
  33042=>"111100100",
  33043=>"000000000",
  33044=>"000001110",
  33045=>"111111111",
  33046=>"100100000",
  33047=>"011001011",
  33048=>"000011111",
  33049=>"000000000",
  33050=>"000110111",
  33051=>"111111111",
  33052=>"011011100",
  33053=>"111111110",
  33054=>"000000111",
  33055=>"110000000",
  33056=>"110010000",
  33057=>"111110000",
  33058=>"111111111",
  33059=>"111111111",
  33060=>"000001001",
  33061=>"000000001",
  33062=>"110111111",
  33063=>"000001011",
  33064=>"010111110",
  33065=>"101111111",
  33066=>"000000000",
  33067=>"111001000",
  33068=>"001001001",
  33069=>"101011111",
  33070=>"000000000",
  33071=>"001000000",
  33072=>"111111111",
  33073=>"000000000",
  33074=>"100000001",
  33075=>"111111100",
  33076=>"110110000",
  33077=>"111111111",
  33078=>"011111011",
  33079=>"011011001",
  33080=>"000000000",
  33081=>"000011001",
  33082=>"000000000",
  33083=>"000110100",
  33084=>"111111111",
  33085=>"011111001",
  33086=>"001001000",
  33087=>"011111000",
  33088=>"000000100",
  33089=>"000000010",
  33090=>"000000000",
  33091=>"111011011",
  33092=>"000000000",
  33093=>"000000000",
  33094=>"000000101",
  33095=>"001111001",
  33096=>"000001000",
  33097=>"111011000",
  33098=>"110111110",
  33099=>"111011011",
  33100=>"111111100",
  33101=>"111110111",
  33102=>"000000000",
  33103=>"001111111",
  33104=>"000000111",
  33105=>"111111111",
  33106=>"000000111",
  33107=>"000000000",
  33108=>"000000000",
  33109=>"010010111",
  33110=>"010010111",
  33111=>"000110110",
  33112=>"100000000",
  33113=>"000000000",
  33114=>"000001000",
  33115=>"000000000",
  33116=>"000000000",
  33117=>"111000000",
  33118=>"110111001",
  33119=>"111111001",
  33120=>"000111110",
  33121=>"000000001",
  33122=>"010010111",
  33123=>"011110000",
  33124=>"000001001",
  33125=>"000000000",
  33126=>"000001101",
  33127=>"000000000",
  33128=>"111111011",
  33129=>"001000000",
  33130=>"111111111",
  33131=>"000110111",
  33132=>"111111011",
  33133=>"000000000",
  33134=>"111111011",
  33135=>"000011000",
  33136=>"000000000",
  33137=>"000000000",
  33138=>"000100100",
  33139=>"000000000",
  33140=>"000000000",
  33141=>"000000000",
  33142=>"000111111",
  33143=>"000010100",
  33144=>"100000000",
  33145=>"000111100",
  33146=>"111001011",
  33147=>"001011101",
  33148=>"101000000",
  33149=>"000000111",
  33150=>"001001011",
  33151=>"111111111",
  33152=>"110100000",
  33153=>"111111110",
  33154=>"110010000",
  33155=>"110111000",
  33156=>"000000101",
  33157=>"110111110",
  33158=>"000000110",
  33159=>"111111001",
  33160=>"111001000",
  33161=>"000000000",
  33162=>"000000000",
  33163=>"010110110",
  33164=>"111111111",
  33165=>"110110110",
  33166=>"111111000",
  33167=>"000000000",
  33168=>"010010000",
  33169=>"000000111",
  33170=>"100111111",
  33171=>"100111111",
  33172=>"001001000",
  33173=>"100000111",
  33174=>"000100000",
  33175=>"111100111",
  33176=>"111111000",
  33177=>"000000110",
  33178=>"111111110",
  33179=>"111111111",
  33180=>"000110111",
  33181=>"100110110",
  33182=>"101000111",
  33183=>"000000000",
  33184=>"111011111",
  33185=>"111111111",
  33186=>"100100100",
  33187=>"111111000",
  33188=>"111111101",
  33189=>"000000000",
  33190=>"111111000",
  33191=>"111101111",
  33192=>"111111111",
  33193=>"000000011",
  33194=>"000000000",
  33195=>"111111000",
  33196=>"010010000",
  33197=>"000000000",
  33198=>"110111110",
  33199=>"111111111",
  33200=>"111111111",
  33201=>"000000100",
  33202=>"000000000",
  33203=>"011111111",
  33204=>"000000000",
  33205=>"100111001",
  33206=>"111111111",
  33207=>"000001111",
  33208=>"000100010",
  33209=>"111111111",
  33210=>"111011000",
  33211=>"111111110",
  33212=>"111101000",
  33213=>"001000000",
  33214=>"000000000",
  33215=>"000000000",
  33216=>"000000011",
  33217=>"000000000",
  33218=>"000000000",
  33219=>"010011000",
  33220=>"000111111",
  33221=>"000001001",
  33222=>"000111111",
  33223=>"000000000",
  33224=>"000000000",
  33225=>"000000000",
  33226=>"001111000",
  33227=>"000010000",
  33228=>"001000000",
  33229=>"000000000",
  33230=>"111100000",
  33231=>"000000100",
  33232=>"110101000",
  33233=>"010111111",
  33234=>"111111111",
  33235=>"111011000",
  33236=>"000010010",
  33237=>"111111011",
  33238=>"000000111",
  33239=>"010111111",
  33240=>"111111111",
  33241=>"111111111",
  33242=>"001000000",
  33243=>"111111011",
  33244=>"111101111",
  33245=>"000000000",
  33246=>"000000000",
  33247=>"100100100",
  33248=>"111111111",
  33249=>"001000000",
  33250=>"111111111",
  33251=>"111111110",
  33252=>"011011011",
  33253=>"111111111",
  33254=>"110111000",
  33255=>"011000000",
  33256=>"111111101",
  33257=>"111111111",
  33258=>"000000101",
  33259=>"000000000",
  33260=>"000000000",
  33261=>"111101111",
  33262=>"100000111",
  33263=>"000000101",
  33264=>"000000000",
  33265=>"000000000",
  33266=>"000011001",
  33267=>"000000000",
  33268=>"001000000",
  33269=>"100001000",
  33270=>"000000000",
  33271=>"001001000",
  33272=>"000000000",
  33273=>"001001001",
  33274=>"000000000",
  33275=>"111011011",
  33276=>"001000010",
  33277=>"110111111",
  33278=>"011011011",
  33279=>"111111111",
  33280=>"111110100",
  33281=>"100000000",
  33282=>"000000000",
  33283=>"111111111",
  33284=>"000000000",
  33285=>"111110000",
  33286=>"000000000",
  33287=>"111111111",
  33288=>"100100111",
  33289=>"111111111",
  33290=>"000110110",
  33291=>"000001001",
  33292=>"000000011",
  33293=>"111101001",
  33294=>"000000000",
  33295=>"100000111",
  33296=>"111111111",
  33297=>"001001111",
  33298=>"011001000",
  33299=>"100111111",
  33300=>"000000011",
  33301=>"000000000",
  33302=>"111111111",
  33303=>"111111111",
  33304=>"001000011",
  33305=>"000110000",
  33306=>"000000100",
  33307=>"110100011",
  33308=>"111111111",
  33309=>"111111110",
  33310=>"001001000",
  33311=>"000000000",
  33312=>"001000000",
  33313=>"000000001",
  33314=>"110000000",
  33315=>"100000111",
  33316=>"000000000",
  33317=>"110000000",
  33318=>"111000000",
  33319=>"000000001",
  33320=>"001000000",
  33321=>"111111111",
  33322=>"110110000",
  33323=>"000000000",
  33324=>"111111111",
  33325=>"110110110",
  33326=>"110110110",
  33327=>"000110100",
  33328=>"101111111",
  33329=>"000111000",
  33330=>"110001001",
  33331=>"000000000",
  33332=>"110000001",
  33333=>"000001011",
  33334=>"000000000",
  33335=>"011111111",
  33336=>"100000000",
  33337=>"000100111",
  33338=>"111111111",
  33339=>"000000000",
  33340=>"000000001",
  33341=>"011111110",
  33342=>"000000000",
  33343=>"000000110",
  33344=>"111000011",
  33345=>"100111111",
  33346=>"111000001",
  33347=>"011110000",
  33348=>"000000000",
  33349=>"010100000",
  33350=>"000000111",
  33351=>"111111101",
  33352=>"110010000",
  33353=>"111111111",
  33354=>"111111110",
  33355=>"011110110",
  33356=>"000000000",
  33357=>"101000000",
  33358=>"001000000",
  33359=>"111100000",
  33360=>"111111101",
  33361=>"111111111",
  33362=>"100100110",
  33363=>"000000011",
  33364=>"000000000",
  33365=>"111111111",
  33366=>"101101101",
  33367=>"111110000",
  33368=>"111111111",
  33369=>"000000000",
  33370=>"100100000",
  33371=>"001001001",
  33372=>"101000000",
  33373=>"101111111",
  33374=>"000010111",
  33375=>"100000111",
  33376=>"000000000",
  33377=>"001001100",
  33378=>"000000000",
  33379=>"100000000",
  33380=>"000000111",
  33381=>"100011011",
  33382=>"111111111",
  33383=>"111111010",
  33384=>"111001000",
  33385=>"000000000",
  33386=>"000100110",
  33387=>"000000100",
  33388=>"000000000",
  33389=>"101100101",
  33390=>"011000000",
  33391=>"000011011",
  33392=>"000110110",
  33393=>"001000100",
  33394=>"100100011",
  33395=>"000001111",
  33396=>"010000000",
  33397=>"001011001",
  33398=>"111111111",
  33399=>"110100000",
  33400=>"111101111",
  33401=>"000000000",
  33402=>"001101000",
  33403=>"000000100",
  33404=>"000001000",
  33405=>"111111111",
  33406=>"111011011",
  33407=>"000000000",
  33408=>"000000101",
  33409=>"111111111",
  33410=>"111010000",
  33411=>"111111111",
  33412=>"101011001",
  33413=>"000000111",
  33414=>"011111111",
  33415=>"111111111",
  33416=>"111111111",
  33417=>"000111011",
  33418=>"111111110",
  33419=>"111111111",
  33420=>"111111111",
  33421=>"000000000",
  33422=>"000100110",
  33423=>"011011000",
  33424=>"111111111",
  33425=>"111100100",
  33426=>"011001011",
  33427=>"100100000",
  33428=>"000100100",
  33429=>"111011000",
  33430=>"111111000",
  33431=>"111110111",
  33432=>"000000000",
  33433=>"000011111",
  33434=>"001001001",
  33435=>"111111111",
  33436=>"011111001",
  33437=>"000000010",
  33438=>"111111111",
  33439=>"001000000",
  33440=>"000000000",
  33441=>"000000000",
  33442=>"011111111",
  33443=>"000000000",
  33444=>"001011111",
  33445=>"010000000",
  33446=>"111100100",
  33447=>"001001000",
  33448=>"000000000",
  33449=>"000000000",
  33450=>"000000000",
  33451=>"111111111",
  33452=>"001101111",
  33453=>"000000000",
  33454=>"111110100",
  33455=>"100000000",
  33456=>"011111000",
  33457=>"001001101",
  33458=>"111111111",
  33459=>"111110000",
  33460=>"110111100",
  33461=>"111011000",
  33462=>"111111111",
  33463=>"100000001",
  33464=>"111000000",
  33465=>"111111001",
  33466=>"111000000",
  33467=>"011000001",
  33468=>"000000000",
  33469=>"111101111",
  33470=>"000000000",
  33471=>"010000000",
  33472=>"000000000",
  33473=>"111111011",
  33474=>"111101111",
  33475=>"111000100",
  33476=>"000111111",
  33477=>"000000000",
  33478=>"000111011",
  33479=>"110100000",
  33480=>"111111111",
  33481=>"011111111",
  33482=>"000001111",
  33483=>"111001001",
  33484=>"000000000",
  33485=>"000000000",
  33486=>"100111000",
  33487=>"011111000",
  33488=>"000000000",
  33489=>"101101111",
  33490=>"001001000",
  33491=>"111111111",
  33492=>"001001111",
  33493=>"111100110",
  33494=>"000000000",
  33495=>"000000100",
  33496=>"000000010",
  33497=>"000000001",
  33498=>"000000000",
  33499=>"011000000",
  33500=>"000000000",
  33501=>"011000000",
  33502=>"011011111",
  33503=>"011000000",
  33504=>"110000000",
  33505=>"000000111",
  33506=>"010111111",
  33507=>"000000000",
  33508=>"001000000",
  33509=>"001100110",
  33510=>"000011000",
  33511=>"010001000",
  33512=>"111011001",
  33513=>"000000100",
  33514=>"010110111",
  33515=>"000000110",
  33516=>"001001000",
  33517=>"100000100",
  33518=>"111111011",
  33519=>"111111111",
  33520=>"010100000",
  33521=>"000000000",
  33522=>"000000000",
  33523=>"000000100",
  33524=>"101100111",
  33525=>"011010001",
  33526=>"111111110",
  33527=>"000000111",
  33528=>"000000000",
  33529=>"110000000",
  33530=>"011000000",
  33531=>"000000000",
  33532=>"111110110",
  33533=>"100000011",
  33534=>"001001001",
  33535=>"000000000",
  33536=>"110100100",
  33537=>"000000000",
  33538=>"111111111",
  33539=>"111001111",
  33540=>"000000100",
  33541=>"000000110",
  33542=>"000011110",
  33543=>"111001001",
  33544=>"000100100",
  33545=>"000000000",
  33546=>"011111111",
  33547=>"011001110",
  33548=>"000000000",
  33549=>"111111000",
  33550=>"011111111",
  33551=>"001000000",
  33552=>"111111101",
  33553=>"001001111",
  33554=>"001000001",
  33555=>"000000000",
  33556=>"110111111",
  33557=>"000000000",
  33558=>"011011011",
  33559=>"100000000",
  33560=>"001111011",
  33561=>"111111111",
  33562=>"000000000",
  33563=>"000111111",
  33564=>"011001111",
  33565=>"111000100",
  33566=>"011111111",
  33567=>"001111111",
  33568=>"110010010",
  33569=>"111111001",
  33570=>"100100111",
  33571=>"111110111",
  33572=>"001001111",
  33573=>"111111111",
  33574=>"001011111",
  33575=>"100100110",
  33576=>"111111011",
  33577=>"100000000",
  33578=>"111111111",
  33579=>"000000000",
  33580=>"000000000",
  33581=>"011011011",
  33582=>"000000000",
  33583=>"111111000",
  33584=>"110101011",
  33585=>"111111000",
  33586=>"011111111",
  33587=>"000000111",
  33588=>"100000000",
  33589=>"000000001",
  33590=>"001011111",
  33591=>"111100101",
  33592=>"000000000",
  33593=>"001001111",
  33594=>"101000000",
  33595=>"000000000",
  33596=>"011111000",
  33597=>"001000000",
  33598=>"111111111",
  33599=>"000100111",
  33600=>"001111111",
  33601=>"111011111",
  33602=>"001100101",
  33603=>"011011000",
  33604=>"000000100",
  33605=>"000010111",
  33606=>"111111110",
  33607=>"000001111",
  33608=>"100100000",
  33609=>"111111111",
  33610=>"100110111",
  33611=>"100100000",
  33612=>"001001001",
  33613=>"101100110",
  33614=>"000100111",
  33615=>"001011000",
  33616=>"100100000",
  33617=>"000000000",
  33618=>"000000011",
  33619=>"101001011",
  33620=>"111000111",
  33621=>"000111111",
  33622=>"111000000",
  33623=>"000110111",
  33624=>"000000000",
  33625=>"110111111",
  33626=>"001001011",
  33627=>"001111111",
  33628=>"000101111",
  33629=>"000000000",
  33630=>"000000000",
  33631=>"001011111",
  33632=>"000100000",
  33633=>"000000100",
  33634=>"100100101",
  33635=>"000000000",
  33636=>"111001001",
  33637=>"000010000",
  33638=>"100110111",
  33639=>"111001001",
  33640=>"100111111",
  33641=>"111111011",
  33642=>"111110000",
  33643=>"011000110",
  33644=>"000010011",
  33645=>"101111110",
  33646=>"111111111",
  33647=>"000000001",
  33648=>"100100101",
  33649=>"100000000",
  33650=>"111101001",
  33651=>"001001000",
  33652=>"000000000",
  33653=>"100000000",
  33654=>"000001011",
  33655=>"110001111",
  33656=>"000000000",
  33657=>"001000010",
  33658=>"111111100",
  33659=>"000000000",
  33660=>"100001011",
  33661=>"111111111",
  33662=>"000000000",
  33663=>"000000000",
  33664=>"111011011",
  33665=>"001001101",
  33666=>"000000000",
  33667=>"000000000",
  33668=>"000000000",
  33669=>"111110000",
  33670=>"000000101",
  33671=>"001000110",
  33672=>"100111111",
  33673=>"111011011",
  33674=>"111000000",
  33675=>"100100000",
  33676=>"000000000",
  33677=>"000100110",
  33678=>"000100111",
  33679=>"111111111",
  33680=>"000000000",
  33681=>"111010010",
  33682=>"110111000",
  33683=>"001000000",
  33684=>"000000000",
  33685=>"111011111",
  33686=>"000000111",
  33687=>"010000011",
  33688=>"000000111",
  33689=>"111100000",
  33690=>"000000100",
  33691=>"111000000",
  33692=>"001011010",
  33693=>"001001010",
  33694=>"111111101",
  33695=>"110110110",
  33696=>"001000100",
  33697=>"110110110",
  33698=>"001001001",
  33699=>"100111111",
  33700=>"000000000",
  33701=>"000000000",
  33702=>"111111111",
  33703=>"011000001",
  33704=>"111111111",
  33705=>"110110111",
  33706=>"000000000",
  33707=>"011011010",
  33708=>"100010110",
  33709=>"000000000",
  33710=>"101101111",
  33711=>"111100000",
  33712=>"101111111",
  33713=>"000000000",
  33714=>"000001001",
  33715=>"010111111",
  33716=>"111111111",
  33717=>"111111111",
  33718=>"101100000",
  33719=>"110010011",
  33720=>"111001011",
  33721=>"011000000",
  33722=>"111111011",
  33723=>"111100100",
  33724=>"000100111",
  33725=>"111001010",
  33726=>"100100100",
  33727=>"001011011",
  33728=>"000011011",
  33729=>"000000000",
  33730=>"000010000",
  33731=>"111111111",
  33732=>"100100111",
  33733=>"000000000",
  33734=>"000000111",
  33735=>"111100100",
  33736=>"000010000",
  33737=>"111111111",
  33738=>"000110000",
  33739=>"001011001",
  33740=>"000000101",
  33741=>"000000000",
  33742=>"000000000",
  33743=>"110111111",
  33744=>"000000000",
  33745=>"001000000",
  33746=>"000000000",
  33747=>"111111111",
  33748=>"000001000",
  33749=>"100111111",
  33750=>"000100100",
  33751=>"000110110",
  33752=>"000110111",
  33753=>"011011110",
  33754=>"000001001",
  33755=>"000000001",
  33756=>"000000000",
  33757=>"000000000",
  33758=>"000000000",
  33759=>"001001111",
  33760=>"000100111",
  33761=>"100000000",
  33762=>"101000000",
  33763=>"011111110",
  33764=>"101111111",
  33765=>"111111101",
  33766=>"000011111",
  33767=>"000000000",
  33768=>"111000000",
  33769=>"111111111",
  33770=>"111111100",
  33771=>"011000000",
  33772=>"100000111",
  33773=>"001000000",
  33774=>"110111110",
  33775=>"011111111",
  33776=>"001001000",
  33777=>"010000000",
  33778=>"001000000",
  33779=>"000000001",
  33780=>"001011111",
  33781=>"111101100",
  33782=>"100000000",
  33783=>"010010010",
  33784=>"000000111",
  33785=>"111111100",
  33786=>"000110100",
  33787=>"111111111",
  33788=>"000010111",
  33789=>"111111111",
  33790=>"000110100",
  33791=>"000000000",
  33792=>"111110111",
  33793=>"000000000",
  33794=>"111000100",
  33795=>"001111111",
  33796=>"000000000",
  33797=>"011000111",
  33798=>"000000000",
  33799=>"111111111",
  33800=>"000000000",
  33801=>"111101111",
  33802=>"000000000",
  33803=>"111111000",
  33804=>"000011110",
  33805=>"010111111",
  33806=>"111111111",
  33807=>"000000000",
  33808=>"001001110",
  33809=>"001000000",
  33810=>"000000111",
  33811=>"000000011",
  33812=>"000000000",
  33813=>"000000000",
  33814=>"100000000",
  33815=>"100100000",
  33816=>"001000100",
  33817=>"000000000",
  33818=>"111111111",
  33819=>"000000011",
  33820=>"011111001",
  33821=>"111111000",
  33822=>"000001001",
  33823=>"111111000",
  33824=>"010111000",
  33825=>"110111110",
  33826=>"000000000",
  33827=>"000000000",
  33828=>"100010011",
  33829=>"011000011",
  33830=>"111100000",
  33831=>"010000000",
  33832=>"111110110",
  33833=>"000000000",
  33834=>"111111111",
  33835=>"000000000",
  33836=>"001000111",
  33837=>"000000000",
  33838=>"000000100",
  33839=>"000000000",
  33840=>"111110111",
  33841=>"000000000",
  33842=>"000000011",
  33843=>"000100110",
  33844=>"000000000",
  33845=>"000000001",
  33846=>"111001001",
  33847=>"111100100",
  33848=>"111111011",
  33849=>"111111010",
  33850=>"000000111",
  33851=>"000000111",
  33852=>"000000000",
  33853=>"000111011",
  33854=>"000000000",
  33855=>"001000111",
  33856=>"111111111",
  33857=>"100000000",
  33858=>"101000000",
  33859=>"000000000",
  33860=>"011111111",
  33861=>"000000110",
  33862=>"111000000",
  33863=>"000110000",
  33864=>"011000000",
  33865=>"111000111",
  33866=>"110111111",
  33867=>"111000000",
  33868=>"111111111",
  33869=>"000000000",
  33870=>"001111111",
  33871=>"111100111",
  33872=>"000000010",
  33873=>"000000000",
  33874=>"001000101",
  33875=>"110110111",
  33876=>"000000000",
  33877=>"101111111",
  33878=>"100100100",
  33879=>"111111111",
  33880=>"100101101",
  33881=>"111011111",
  33882=>"111001001",
  33883=>"000000000",
  33884=>"001111111",
  33885=>"000111111",
  33886=>"011111111",
  33887=>"001111111",
  33888=>"000110110",
  33889=>"000111110",
  33890=>"000000100",
  33891=>"000000000",
  33892=>"000000101",
  33893=>"000000000",
  33894=>"111111000",
  33895=>"000000100",
  33896=>"111001000",
  33897=>"111111111",
  33898=>"111111111",
  33899=>"000000001",
  33900=>"100100111",
  33901=>"111111111",
  33902=>"100101101",
  33903=>"001001000",
  33904=>"000000000",
  33905=>"000000000",
  33906=>"001000101",
  33907=>"011111001",
  33908=>"000000000",
  33909=>"000111111",
  33910=>"000000000",
  33911=>"000100110",
  33912=>"000000000",
  33913=>"101000111",
  33914=>"000000000",
  33915=>"111010000",
  33916=>"100111111",
  33917=>"000000111",
  33918=>"101000010",
  33919=>"000011111",
  33920=>"001001000",
  33921=>"000111111",
  33922=>"000111111",
  33923=>"000011001",
  33924=>"110011000",
  33925=>"101100111",
  33926=>"000011011",
  33927=>"000100111",
  33928=>"111111100",
  33929=>"001000000",
  33930=>"000100000",
  33931=>"000001111",
  33932=>"000000111",
  33933=>"000000000",
  33934=>"101000011",
  33935=>"000000000",
  33936=>"100111111",
  33937=>"000000000",
  33938=>"111111111",
  33939=>"100000000",
  33940=>"001011000",
  33941=>"000000000",
  33942=>"111101000",
  33943=>"111011000",
  33944=>"111011000",
  33945=>"111000111",
  33946=>"000000000",
  33947=>"110111000",
  33948=>"111000000",
  33949=>"000000111",
  33950=>"000000111",
  33951=>"111111111",
  33952=>"101000000",
  33953=>"011110000",
  33954=>"111111011",
  33955=>"000000110",
  33956=>"100100000",
  33957=>"101111111",
  33958=>"100110100",
  33959=>"001011111",
  33960=>"010011110",
  33961=>"000000100",
  33962=>"111111101",
  33963=>"000000000",
  33964=>"111111010",
  33965=>"110110000",
  33966=>"100000000",
  33967=>"000101111",
  33968=>"000000111",
  33969=>"000000000",
  33970=>"111111111",
  33971=>"110101000",
  33972=>"000101111",
  33973=>"111011001",
  33974=>"000111111",
  33975=>"000010000",
  33976=>"011111111",
  33977=>"000001000",
  33978=>"000000000",
  33979=>"001011111",
  33980=>"000000000",
  33981=>"000011011",
  33982=>"000000111",
  33983=>"111111111",
  33984=>"000110111",
  33985=>"000001000",
  33986=>"000011111",
  33987=>"000011000",
  33988=>"000000111",
  33989=>"001000000",
  33990=>"111111000",
  33991=>"100011110",
  33992=>"000000110",
  33993=>"000000111",
  33994=>"011110110",
  33995=>"000000000",
  33996=>"111111111",
  33997=>"111111111",
  33998=>"100111111",
  33999=>"100100000",
  34000=>"000000110",
  34001=>"000000101",
  34002=>"000111111",
  34003=>"110111111",
  34004=>"111111101",
  34005=>"111100111",
  34006=>"011001000",
  34007=>"111111111",
  34008=>"101101000",
  34009=>"010110111",
  34010=>"000000000",
  34011=>"000000000",
  34012=>"111111111",
  34013=>"000110110",
  34014=>"111111011",
  34015=>"111011011",
  34016=>"000000001",
  34017=>"000011000",
  34018=>"111111000",
  34019=>"111100000",
  34020=>"111111111",
  34021=>"000000000",
  34022=>"000000111",
  34023=>"000000000",
  34024=>"111101000",
  34025=>"000100111",
  34026=>"111111111",
  34027=>"111111001",
  34028=>"000111111",
  34029=>"111101000",
  34030=>"111111111",
  34031=>"111111000",
  34032=>"001000000",
  34033=>"111110110",
  34034=>"111111111",
  34035=>"011111001",
  34036=>"000111111",
  34037=>"111111011",
  34038=>"110100001",
  34039=>"111000000",
  34040=>"001000101",
  34041=>"010000000",
  34042=>"000000011",
  34043=>"010011000",
  34044=>"000100110",
  34045=>"000100110",
  34046=>"111111111",
  34047=>"100100110",
  34048=>"000000010",
  34049=>"011011001",
  34050=>"111111000",
  34051=>"000000010",
  34052=>"011111111",
  34053=>"110111111",
  34054=>"111000000",
  34055=>"101111001",
  34056=>"000000000",
  34057=>"011011111",
  34058=>"111111111",
  34059=>"000000111",
  34060=>"000000100",
  34061=>"001111111",
  34062=>"000000110",
  34063=>"111001111",
  34064=>"000000000",
  34065=>"000000000",
  34066=>"111111010",
  34067=>"000000000",
  34068=>"000000100",
  34069=>"000000000",
  34070=>"110110110",
  34071=>"000000000",
  34072=>"001101111",
  34073=>"111000000",
  34074=>"111111111",
  34075=>"000111111",
  34076=>"010011000",
  34077=>"111111000",
  34078=>"111111111",
  34079=>"111011000",
  34080=>"000100100",
  34081=>"000000111",
  34082=>"100000001",
  34083=>"111111111",
  34084=>"000000000",
  34085=>"000000111",
  34086=>"011111000",
  34087=>"111110100",
  34088=>"000000000",
  34089=>"111001001",
  34090=>"001111000",
  34091=>"000000000",
  34092=>"000000000",
  34093=>"001111100",
  34094=>"000100000",
  34095=>"000000111",
  34096=>"000110111",
  34097=>"000001111",
  34098=>"011000000",
  34099=>"111111111",
  34100=>"100100000",
  34101=>"011011010",
  34102=>"000000001",
  34103=>"111111000",
  34104=>"111100000",
  34105=>"111111000",
  34106=>"000111101",
  34107=>"111111000",
  34108=>"000000110",
  34109=>"000001111",
  34110=>"111111111",
  34111=>"000000000",
  34112=>"010110111",
  34113=>"000000001",
  34114=>"000001010",
  34115=>"000000010",
  34116=>"011010000",
  34117=>"000000001",
  34118=>"001000000",
  34119=>"111101001",
  34120=>"110111111",
  34121=>"000000101",
  34122=>"111110111",
  34123=>"000011010",
  34124=>"111111111",
  34125=>"111111111",
  34126=>"001000000",
  34127=>"100110100",
  34128=>"100110110",
  34129=>"111100000",
  34130=>"010000000",
  34131=>"111111111",
  34132=>"000000110",
  34133=>"011011011",
  34134=>"111111111",
  34135=>"100111111",
  34136=>"111111111",
  34137=>"111111111",
  34138=>"000000000",
  34139=>"111111111",
  34140=>"101000000",
  34141=>"000000000",
  34142=>"000000000",
  34143=>"000000000",
  34144=>"100100111",
  34145=>"000111111",
  34146=>"100110110",
  34147=>"101000000",
  34148=>"000000111",
  34149=>"000000111",
  34150=>"000001000",
  34151=>"000111111",
  34152=>"110111111",
  34153=>"000011111",
  34154=>"000001001",
  34155=>"111010110",
  34156=>"110111111",
  34157=>"111110111",
  34158=>"000010001",
  34159=>"111111111",
  34160=>"000010111",
  34161=>"111111111",
  34162=>"000001000",
  34163=>"111111110",
  34164=>"111111000",
  34165=>"111110110",
  34166=>"000000000",
  34167=>"000000111",
  34168=>"111000001",
  34169=>"000110110",
  34170=>"111111111",
  34171=>"010110110",
  34172=>"111111111",
  34173=>"011000111",
  34174=>"000111000",
  34175=>"000000000",
  34176=>"000000111",
  34177=>"111000000",
  34178=>"000010001",
  34179=>"000000000",
  34180=>"000000110",
  34181=>"111010010",
  34182=>"111111111",
  34183=>"111000001",
  34184=>"000000000",
  34185=>"111111111",
  34186=>"001001101",
  34187=>"000000111",
  34188=>"000111111",
  34189=>"001001000",
  34190=>"000000111",
  34191=>"111111111",
  34192=>"000000000",
  34193=>"111000111",
  34194=>"000000000",
  34195=>"000000111",
  34196=>"000111111",
  34197=>"000000000",
  34198=>"111110110",
  34199=>"100100100",
  34200=>"111000000",
  34201=>"000011111",
  34202=>"000000000",
  34203=>"011100110",
  34204=>"100000001",
  34205=>"000110111",
  34206=>"011000000",
  34207=>"000000000",
  34208=>"100000000",
  34209=>"000001000",
  34210=>"010011000",
  34211=>"111111101",
  34212=>"111111111",
  34213=>"001111001",
  34214=>"000000000",
  34215=>"000000100",
  34216=>"100110111",
  34217=>"000111111",
  34218=>"111111111",
  34219=>"111000000",
  34220=>"010111000",
  34221=>"001001100",
  34222=>"110000000",
  34223=>"001000010",
  34224=>"101000000",
  34225=>"000000000",
  34226=>"000100000",
  34227=>"111111101",
  34228=>"111110111",
  34229=>"110111111",
  34230=>"111111111",
  34231=>"111100000",
  34232=>"111111111",
  34233=>"011000000",
  34234=>"000000101",
  34235=>"011000000",
  34236=>"111111111",
  34237=>"111111001",
  34238=>"000000000",
  34239=>"000010010",
  34240=>"001000000",
  34241=>"010000000",
  34242=>"111111000",
  34243=>"000111111",
  34244=>"111111001",
  34245=>"000111111",
  34246=>"000000001",
  34247=>"000000010",
  34248=>"001011000",
  34249=>"011000000",
  34250=>"000110111",
  34251=>"000000000",
  34252=>"111111000",
  34253=>"011101001",
  34254=>"001100000",
  34255=>"001000000",
  34256=>"000000111",
  34257=>"001000000",
  34258=>"001001001",
  34259=>"000000001",
  34260=>"001010010",
  34261=>"000000000",
  34262=>"000000000",
  34263=>"000000011",
  34264=>"000000000",
  34265=>"011111110",
  34266=>"111111000",
  34267=>"000111111",
  34268=>"000110110",
  34269=>"101111111",
  34270=>"000000000",
  34271=>"000001001",
  34272=>"001000000",
  34273=>"000000000",
  34274=>"000001000",
  34275=>"111111011",
  34276=>"111111011",
  34277=>"111000000",
  34278=>"100000111",
  34279=>"111111111",
  34280=>"011000110",
  34281=>"001011111",
  34282=>"000010011",
  34283=>"001111111",
  34284=>"000110111",
  34285=>"001011001",
  34286=>"000000001",
  34287=>"111111111",
  34288=>"111100000",
  34289=>"000000000",
  34290=>"111110110",
  34291=>"101001000",
  34292=>"000001000",
  34293=>"111111111",
  34294=>"001001000",
  34295=>"110111000",
  34296=>"111111000",
  34297=>"110111111",
  34298=>"011000000",
  34299=>"111111111",
  34300=>"010000000",
  34301=>"001011111",
  34302=>"111000000",
  34303=>"000000000",
  34304=>"111010000",
  34305=>"000000000",
  34306=>"111111111",
  34307=>"011011011",
  34308=>"111100111",
  34309=>"001001000",
  34310=>"001000011",
  34311=>"111111101",
  34312=>"100000000",
  34313=>"111111111",
  34314=>"001111001",
  34315=>"000100100",
  34316=>"000100110",
  34317=>"000100111",
  34318=>"101000000",
  34319=>"000110110",
  34320=>"111001001",
  34321=>"001000000",
  34322=>"011011000",
  34323=>"110110111",
  34324=>"111111111",
  34325=>"111111111",
  34326=>"000000011",
  34327=>"000100100",
  34328=>"001001111",
  34329=>"000000000",
  34330=>"000000110",
  34331=>"000100001",
  34332=>"111000000",
  34333=>"110111111",
  34334=>"111011101",
  34335=>"000000000",
  34336=>"111111101",
  34337=>"011100000",
  34338=>"111100100",
  34339=>"010110111",
  34340=>"000010000",
  34341=>"111110110",
  34342=>"111111011",
  34343=>"111001000",
  34344=>"001001011",
  34345=>"111111111",
  34346=>"111111111",
  34347=>"000000111",
  34348=>"000100100",
  34349=>"111111011",
  34350=>"001011100",
  34351=>"111111010",
  34352=>"000100110",
  34353=>"000111111",
  34354=>"111110111",
  34355=>"000000000",
  34356=>"000000101",
  34357=>"110110100",
  34358=>"111001001",
  34359=>"111000000",
  34360=>"100000000",
  34361=>"000000000",
  34362=>"100000000",
  34363=>"111111111",
  34364=>"111101111",
  34365=>"111111111",
  34366=>"101110110",
  34367=>"000000000",
  34368=>"100100100",
  34369=>"111111111",
  34370=>"111001000",
  34371=>"111111111",
  34372=>"000000101",
  34373=>"001001011",
  34374=>"111111110",
  34375=>"000000000",
  34376=>"111110110",
  34377=>"111111111",
  34378=>"000000000",
  34379=>"111100101",
  34380=>"000000111",
  34381=>"001010000",
  34382=>"000011000",
  34383=>"001000111",
  34384=>"111111111",
  34385=>"111111111",
  34386=>"001000000",
  34387=>"001010000",
  34388=>"111101000",
  34389=>"000000000",
  34390=>"111110111",
  34391=>"111111111",
  34392=>"100000000",
  34393=>"000000000",
  34394=>"111010000",
  34395=>"000000111",
  34396=>"111111000",
  34397=>"010111111",
  34398=>"111110110",
  34399=>"110000000",
  34400=>"000000000",
  34401=>"111111000",
  34402=>"000000100",
  34403=>"000000100",
  34404=>"100111111",
  34405=>"111100000",
  34406=>"111111111",
  34407=>"000101000",
  34408=>"111111111",
  34409=>"000000000",
  34410=>"100110110",
  34411=>"111110111",
  34412=>"111111111",
  34413=>"010011001",
  34414=>"111111111",
  34415=>"000000011",
  34416=>"100100111",
  34417=>"011011000",
  34418=>"000001111",
  34419=>"000000000",
  34420=>"000000010",
  34421=>"110000000",
  34422=>"000000111",
  34423=>"000011000",
  34424=>"111111001",
  34425=>"111111111",
  34426=>"011000000",
  34427=>"000000100",
  34428=>"111111001",
  34429=>"000000000",
  34430=>"001001000",
  34431=>"000000000",
  34432=>"011011000",
  34433=>"001001101",
  34434=>"000000000",
  34435=>"000011011",
  34436=>"110000001",
  34437=>"000111111",
  34438=>"111111111",
  34439=>"000000000",
  34440=>"111111111",
  34441=>"011000001",
  34442=>"000000000",
  34443=>"111111111",
  34444=>"000000000",
  34445=>"000000111",
  34446=>"101101001",
  34447=>"010111111",
  34448=>"101111111",
  34449=>"111001000",
  34450=>"000100000",
  34451=>"000001000",
  34452=>"000011101",
  34453=>"001001011",
  34454=>"111111110",
  34455=>"100000100",
  34456=>"000011111",
  34457=>"111111111",
  34458=>"001011111",
  34459=>"111110100",
  34460=>"111111111",
  34461=>"000111111",
  34462=>"111111101",
  34463=>"000001011",
  34464=>"110111111",
  34465=>"001000000",
  34466=>"111111111",
  34467=>"000000000",
  34468=>"011011000",
  34469=>"000000000",
  34470=>"000001101",
  34471=>"100100000",
  34472=>"111111111",
  34473=>"100100000",
  34474=>"000110111",
  34475=>"111111111",
  34476=>"000000111",
  34477=>"111111111",
  34478=>"110000011",
  34479=>"000100111",
  34480=>"000111010",
  34481=>"000000001",
  34482=>"111110010",
  34483=>"000000000",
  34484=>"111001001",
  34485=>"111010010",
  34486=>"111111111",
  34487=>"111000000",
  34488=>"111111111",
  34489=>"001000000",
  34490=>"001001111",
  34491=>"001111111",
  34492=>"011000000",
  34493=>"000000010",
  34494=>"000111111",
  34495=>"000000000",
  34496=>"111111111",
  34497=>"111111111",
  34498=>"010011111",
  34499=>"010001111",
  34500=>"001111111",
  34501=>"111111000",
  34502=>"011000000",
  34503=>"111001001",
  34504=>"000000000",
  34505=>"111100000",
  34506=>"111001110",
  34507=>"001011111",
  34508=>"000001000",
  34509=>"111111100",
  34510=>"111111100",
  34511=>"101100110",
  34512=>"000110110",
  34513=>"001001000",
  34514=>"111111111",
  34515=>"011111011",
  34516=>"001001111",
  34517=>"111111111",
  34518=>"000000111",
  34519=>"011011011",
  34520=>"000101111",
  34521=>"110111111",
  34522=>"000110110",
  34523=>"000000111",
  34524=>"111000000",
  34525=>"100000000",
  34526=>"111111111",
  34527=>"111000000",
  34528=>"111010110",
  34529=>"000000000",
  34530=>"000000000",
  34531=>"111111111",
  34532=>"001111011",
  34533=>"000000000",
  34534=>"000001001",
  34535=>"000001101",
  34536=>"110110111",
  34537=>"000000000",
  34538=>"000000111",
  34539=>"000000000",
  34540=>"000000000",
  34541=>"000000010",
  34542=>"000000110",
  34543=>"001000000",
  34544=>"110100000",
  34545=>"000010010",
  34546=>"111111111",
  34547=>"000000000",
  34548=>"111111111",
  34549=>"111111111",
  34550=>"000001001",
  34551=>"111111110",
  34552=>"000000000",
  34553=>"011111111",
  34554=>"000010111",
  34555=>"000000000",
  34556=>"011110111",
  34557=>"000010000",
  34558=>"011111111",
  34559=>"111111111",
  34560=>"111111111",
  34561=>"111111110",
  34562=>"010000000",
  34563=>"000101111",
  34564=>"100100001",
  34565=>"111011000",
  34566=>"100101101",
  34567=>"110000000",
  34568=>"000000111",
  34569=>"000000000",
  34570=>"001101111",
  34571=>"000111111",
  34572=>"000000110",
  34573=>"111101000",
  34574=>"110111000",
  34575=>"111111110",
  34576=>"000011111",
  34577=>"000000011",
  34578=>"000000000",
  34579=>"111100001",
  34580=>"001011001",
  34581=>"111111000",
  34582=>"001111111",
  34583=>"100111111",
  34584=>"000000100",
  34585=>"111111111",
  34586=>"000000000",
  34587=>"000100000",
  34588=>"000000000",
  34589=>"110000000",
  34590=>"000000000",
  34591=>"001100000",
  34592=>"111111100",
  34593=>"000000000",
  34594=>"111111000",
  34595=>"100100110",
  34596=>"101111111",
  34597=>"000111111",
  34598=>"000000110",
  34599=>"000000000",
  34600=>"111111111",
  34601=>"111111100",
  34602=>"101000000",
  34603=>"111101000",
  34604=>"000000111",
  34605=>"010001000",
  34606=>"000000000",
  34607=>"111111111",
  34608=>"110110110",
  34609=>"101100010",
  34610=>"111100100",
  34611=>"000000000",
  34612=>"111011000",
  34613=>"000000000",
  34614=>"000000001",
  34615=>"000110100",
  34616=>"011111000",
  34617=>"000100110",
  34618=>"000111111",
  34619=>"111111110",
  34620=>"011101001",
  34621=>"000000111",
  34622=>"011111011",
  34623=>"000100000",
  34624=>"000000000",
  34625=>"111111111",
  34626=>"111111110",
  34627=>"010111011",
  34628=>"000000000",
  34629=>"000111011",
  34630=>"101111011",
  34631=>"000000000",
  34632=>"000001011",
  34633=>"000000000",
  34634=>"000000000",
  34635=>"000111111",
  34636=>"000100111",
  34637=>"111111010",
  34638=>"111111111",
  34639=>"100111001",
  34640=>"000000001",
  34641=>"111110010",
  34642=>"000111111",
  34643=>"000111111",
  34644=>"000000000",
  34645=>"111110011",
  34646=>"000110111",
  34647=>"010100101",
  34648=>"000000011",
  34649=>"000000000",
  34650=>"111111011",
  34651=>"000001000",
  34652=>"000000110",
  34653=>"000111111",
  34654=>"111111000",
  34655=>"000000100",
  34656=>"111111111",
  34657=>"111111111",
  34658=>"000100110",
  34659=>"111011000",
  34660=>"000000000",
  34661=>"111001000",
  34662=>"000111101",
  34663=>"111111111",
  34664=>"011001110",
  34665=>"000111111",
  34666=>"111100000",
  34667=>"111001001",
  34668=>"000000110",
  34669=>"011111111",
  34670=>"011000000",
  34671=>"001111111",
  34672=>"001000000",
  34673=>"000000000",
  34674=>"110110101",
  34675=>"010010010",
  34676=>"000010110",
  34677=>"110111001",
  34678=>"011000000",
  34679=>"000011000",
  34680=>"000000000",
  34681=>"000000100",
  34682=>"000000000",
  34683=>"010110111",
  34684=>"111010000",
  34685=>"111111011",
  34686=>"011011011",
  34687=>"111101101",
  34688=>"000000000",
  34689=>"100100110",
  34690=>"011111010",
  34691=>"000000000",
  34692=>"000010111",
  34693=>"000000000",
  34694=>"110110100",
  34695=>"000000000",
  34696=>"000101111",
  34697=>"000000000",
  34698=>"000000000",
  34699=>"000000110",
  34700=>"111100111",
  34701=>"000000011",
  34702=>"000001011",
  34703=>"011001000",
  34704=>"000000000",
  34705=>"001000111",
  34706=>"000111111",
  34707=>"110110110",
  34708=>"111000000",
  34709=>"000000000",
  34710=>"111001111",
  34711=>"110011000",
  34712=>"000100000",
  34713=>"011101101",
  34714=>"000000100",
  34715=>"111111010",
  34716=>"001101111",
  34717=>"000000000",
  34718=>"000000000",
  34719=>"000000001",
  34720=>"000000000",
  34721=>"011111111",
  34722=>"001000011",
  34723=>"111111011",
  34724=>"100100110",
  34725=>"000000000",
  34726=>"000000000",
  34727=>"110111111",
  34728=>"000010111",
  34729=>"000010000",
  34730=>"001000000",
  34731=>"000000000",
  34732=>"000000000",
  34733=>"000000000",
  34734=>"011111110",
  34735=>"000000001",
  34736=>"111111111",
  34737=>"111111011",
  34738=>"000111111",
  34739=>"111101111",
  34740=>"110111011",
  34741=>"000111111",
  34742=>"110111111",
  34743=>"111111110",
  34744=>"000110111",
  34745=>"111111000",
  34746=>"001000000",
  34747=>"111110111",
  34748=>"111111000",
  34749=>"111111111",
  34750=>"000000000",
  34751=>"101101111",
  34752=>"001100000",
  34753=>"110101101",
  34754=>"000100111",
  34755=>"111111101",
  34756=>"111100000",
  34757=>"000000100",
  34758=>"100000000",
  34759=>"000000000",
  34760=>"000011111",
  34761=>"011111111",
  34762=>"001001111",
  34763=>"000000111",
  34764=>"011001011",
  34765=>"111111111",
  34766=>"110111111",
  34767=>"111111111",
  34768=>"000111100",
  34769=>"000001111",
  34770=>"000001011",
  34771=>"000000000",
  34772=>"100110110",
  34773=>"001111111",
  34774=>"001101111",
  34775=>"010111111",
  34776=>"000000011",
  34777=>"111111111",
  34778=>"111111000",
  34779=>"111111110",
  34780=>"000010000",
  34781=>"000000000",
  34782=>"110100000",
  34783=>"100000000",
  34784=>"000000000",
  34785=>"000000011",
  34786=>"011000000",
  34787=>"011010001",
  34788=>"111011111",
  34789=>"011010010",
  34790=>"000000001",
  34791=>"010011111",
  34792=>"000000000",
  34793=>"011011111",
  34794=>"000100100",
  34795=>"000100100",
  34796=>"100100110",
  34797=>"111110110",
  34798=>"111000000",
  34799=>"000000101",
  34800=>"111101001",
  34801=>"011001000",
  34802=>"111110111",
  34803=>"110000000",
  34804=>"000000110",
  34805=>"010010000",
  34806=>"100001111",
  34807=>"111101111",
  34808=>"000100111",
  34809=>"100100000",
  34810=>"000000110",
  34811=>"010000000",
  34812=>"000001111",
  34813=>"110100100",
  34814=>"000000001",
  34815=>"111111000",
  34816=>"000000000",
  34817=>"000000000",
  34818=>"000000000",
  34819=>"011001001",
  34820=>"001011011",
  34821=>"011111111",
  34822=>"000011111",
  34823=>"111000000",
  34824=>"010111111",
  34825=>"111111111",
  34826=>"001000000",
  34827=>"000000000",
  34828=>"000000101",
  34829=>"100100111",
  34830=>"111110100",
  34831=>"111111111",
  34832=>"010110111",
  34833=>"000000100",
  34834=>"111110111",
  34835=>"000000000",
  34836=>"011110110",
  34837=>"000000000",
  34838=>"111111001",
  34839=>"000000000",
  34840=>"111110100",
  34841=>"000010110",
  34842=>"001001101",
  34843=>"111110110",
  34844=>"001000000",
  34845=>"111001000",
  34846=>"100010010",
  34847=>"000000000",
  34848=>"111111111",
  34849=>"001000000",
  34850=>"111111111",
  34851=>"111001001",
  34852=>"111111111",
  34853=>"100100111",
  34854=>"111111111",
  34855=>"011000110",
  34856=>"001000001",
  34857=>"111111111",
  34858=>"111111000",
  34859=>"111111111",
  34860=>"111000000",
  34861=>"100000000",
  34862=>"001001000",
  34863=>"110110110",
  34864=>"000001010",
  34865=>"100101111",
  34866=>"000000000",
  34867=>"000000110",
  34868=>"000000110",
  34869=>"011001000",
  34870=>"100000000",
  34871=>"111101100",
  34872=>"000000000",
  34873=>"111111001",
  34874=>"111111111",
  34875=>"000011111",
  34876=>"100100101",
  34877=>"001111110",
  34878=>"001111111",
  34879=>"111111111",
  34880=>"111111000",
  34881=>"110110010",
  34882=>"111111011",
  34883=>"010000000",
  34884=>"000000010",
  34885=>"000000000",
  34886=>"111111000",
  34887=>"111000000",
  34888=>"111111111",
  34889=>"111010111",
  34890=>"111111010",
  34891=>"111111111",
  34892=>"000000000",
  34893=>"110110100",
  34894=>"111111110",
  34895=>"100000000",
  34896=>"000100100",
  34897=>"111111111",
  34898=>"111100000",
  34899=>"001001011",
  34900=>"000111111",
  34901=>"111111011",
  34902=>"111111000",
  34903=>"011011011",
  34904=>"111111111",
  34905=>"110000000",
  34906=>"111111111",
  34907=>"011011010",
  34908=>"001100100",
  34909=>"000000111",
  34910=>"001000000",
  34911=>"000000000",
  34912=>"000000000",
  34913=>"111111000",
  34914=>"011000101",
  34915=>"000000101",
  34916=>"001001001",
  34917=>"011001001",
  34918=>"111111001",
  34919=>"110111111",
  34920=>"111111111",
  34921=>"000111111",
  34922=>"111111011",
  34923=>"111000000",
  34924=>"111011001",
  34925=>"000001111",
  34926=>"111111111",
  34927=>"111111111",
  34928=>"000000000",
  34929=>"111111011",
  34930=>"000111111",
  34931=>"100100001",
  34932=>"000000000",
  34933=>"000000100",
  34934=>"010010010",
  34935=>"000000000",
  34936=>"111111111",
  34937=>"000000000",
  34938=>"000000110",
  34939=>"111110111",
  34940=>"111101101",
  34941=>"000000000",
  34942=>"000001111",
  34943=>"011000100",
  34944=>"000011010",
  34945=>"011000000",
  34946=>"111111111",
  34947=>"100100110",
  34948=>"111111101",
  34949=>"111111111",
  34950=>"110100000",
  34951=>"111110100",
  34952=>"000000000",
  34953=>"011000000",
  34954=>"100101111",
  34955=>"100000100",
  34956=>"000000000",
  34957=>"111001111",
  34958=>"000100000",
  34959=>"000000000",
  34960=>"111111111",
  34961=>"101111111",
  34962=>"000000000",
  34963=>"001001001",
  34964=>"100100111",
  34965=>"000000000",
  34966=>"111111111",
  34967=>"111000000",
  34968=>"111111111",
  34969=>"110000000",
  34970=>"111001111",
  34971=>"111111110",
  34972=>"111111111",
  34973=>"000111100",
  34974=>"000000101",
  34975=>"000000000",
  34976=>"000000001",
  34977=>"111000000",
  34978=>"111111111",
  34979=>"111111000",
  34980=>"011001001",
  34981=>"011011110",
  34982=>"101100000",
  34983=>"000110110",
  34984=>"011001000",
  34985=>"000110000",
  34986=>"000000000",
  34987=>"001000001",
  34988=>"000000010",
  34989=>"000001001",
  34990=>"111111111",
  34991=>"000000000",
  34992=>"101100110",
  34993=>"000001001",
  34994=>"111111111",
  34995=>"001001000",
  34996=>"000000000",
  34997=>"000110110",
  34998=>"000000000",
  34999=>"111111111",
  35000=>"111111101",
  35001=>"000000111",
  35002=>"111111111",
  35003=>"000100111",
  35004=>"001001001",
  35005=>"111101001",
  35006=>"111001000",
  35007=>"011001111",
  35008=>"001011011",
  35009=>"000000011",
  35010=>"001000000",
  35011=>"111111000",
  35012=>"111111110",
  35013=>"000000000",
  35014=>"111111111",
  35015=>"001101101",
  35016=>"110110111",
  35017=>"111011011",
  35018=>"111111111",
  35019=>"111111111",
  35020=>"000001100",
  35021=>"000000000",
  35022=>"111110111",
  35023=>"001000000",
  35024=>"000000000",
  35025=>"000001000",
  35026=>"000000000",
  35027=>"000000000",
  35028=>"011101001",
  35029=>"000000000",
  35030=>"000011000",
  35031=>"101000000",
  35032=>"111101000",
  35033=>"001000000",
  35034=>"111111111",
  35035=>"000000000",
  35036=>"011000000",
  35037=>"001001000",
  35038=>"111111101",
  35039=>"111010000",
  35040=>"000000000",
  35041=>"100000111",
  35042=>"111111111",
  35043=>"000000000",
  35044=>"111111011",
  35045=>"100000000",
  35046=>"011011111",
  35047=>"001111111",
  35048=>"000000000",
  35049=>"111111111",
  35050=>"000001111",
  35051=>"111111000",
  35052=>"101111111",
  35053=>"000000111",
  35054=>"000000000",
  35055=>"000000000",
  35056=>"011111001",
  35057=>"100110110",
  35058=>"011001101",
  35059=>"111100001",
  35060=>"111111100",
  35061=>"000011001",
  35062=>"010010100",
  35063=>"000000000",
  35064=>"001101111",
  35065=>"011111111",
  35066=>"111100111",
  35067=>"000000000",
  35068=>"011001000",
  35069=>"001001001",
  35070=>"011010000",
  35071=>"010000111",
  35072=>"111101111",
  35073=>"010010001",
  35074=>"000000110",
  35075=>"111100110",
  35076=>"000000000",
  35077=>"001111111",
  35078=>"000000000",
  35079=>"101100111",
  35080=>"101111101",
  35081=>"000111111",
  35082=>"100100110",
  35083=>"110011111",
  35084=>"001101101",
  35085=>"101111111",
  35086=>"001001011",
  35087=>"000011111",
  35088=>"010111111",
  35089=>"111100111",
  35090=>"001001101",
  35091=>"011011001",
  35092=>"011111000",
  35093=>"111111001",
  35094=>"111001001",
  35095=>"001000000",
  35096=>"111111111",
  35097=>"111111011",
  35098=>"000000000",
  35099=>"110110100",
  35100=>"010000000",
  35101=>"000110111",
  35102=>"001111000",
  35103=>"111111111",
  35104=>"111111101",
  35105=>"000000001",
  35106=>"011000000",
  35107=>"111001001",
  35108=>"100100100",
  35109=>"000000100",
  35110=>"111111111",
  35111=>"001011111",
  35112=>"101111000",
  35113=>"111011011",
  35114=>"001000000",
  35115=>"000100111",
  35116=>"001110111",
  35117=>"001011111",
  35118=>"000000000",
  35119=>"001000100",
  35120=>"000000000",
  35121=>"000000001",
  35122=>"111011111",
  35123=>"101111001",
  35124=>"000000001",
  35125=>"001111111",
  35126=>"100100000",
  35127=>"110000000",
  35128=>"111111111",
  35129=>"001000001",
  35130=>"000000000",
  35131=>"000000100",
  35132=>"000000000",
  35133=>"000000000",
  35134=>"111111111",
  35135=>"000010000",
  35136=>"100011011",
  35137=>"000000000",
  35138=>"000000100",
  35139=>"000000000",
  35140=>"111111111",
  35141=>"110110111",
  35142=>"000000000",
  35143=>"100000000",
  35144=>"000010110",
  35145=>"000000000",
  35146=>"111111110",
  35147=>"001000000",
  35148=>"001111001",
  35149=>"001001000",
  35150=>"011000000",
  35151=>"111111000",
  35152=>"100100100",
  35153=>"011000011",
  35154=>"111111100",
  35155=>"111111111",
  35156=>"000111111",
  35157=>"011011111",
  35158=>"100000000",
  35159=>"000000000",
  35160=>"000000001",
  35161=>"111000000",
  35162=>"100100000",
  35163=>"111111111",
  35164=>"111111111",
  35165=>"111111011",
  35166=>"001101100",
  35167=>"111111010",
  35168=>"000000000",
  35169=>"000000001",
  35170=>"001000110",
  35171=>"011001000",
  35172=>"010000001",
  35173=>"101111111",
  35174=>"010000000",
  35175=>"000101000",
  35176=>"101001001",
  35177=>"011111011",
  35178=>"001001111",
  35179=>"000000110",
  35180=>"000001011",
  35181=>"111010010",
  35182=>"000000000",
  35183=>"110100000",
  35184=>"111111111",
  35185=>"111111111",
  35186=>"000000000",
  35187=>"011011111",
  35188=>"000111111",
  35189=>"011001000",
  35190=>"000000000",
  35191=>"000000000",
  35192=>"110100000",
  35193=>"101000110",
  35194=>"011000101",
  35195=>"111011011",
  35196=>"111111111",
  35197=>"111000000",
  35198=>"111111001",
  35199=>"000000000",
  35200=>"110111111",
  35201=>"000000000",
  35202=>"100100000",
  35203=>"000100000",
  35204=>"000000000",
  35205=>"111001111",
  35206=>"111100000",
  35207=>"100100000",
  35208=>"000000000",
  35209=>"110001011",
  35210=>"000000000",
  35211=>"111111111",
  35212=>"111001101",
  35213=>"001101111",
  35214=>"000001000",
  35215=>"000000001",
  35216=>"000100110",
  35217=>"110000000",
  35218=>"111111111",
  35219=>"000000000",
  35220=>"110000000",
  35221=>"000000000",
  35222=>"010011000",
  35223=>"111111111",
  35224=>"111111111",
  35225=>"001111001",
  35226=>"111111111",
  35227=>"111011001",
  35228=>"001101100",
  35229=>"001011111",
  35230=>"000111111",
  35231=>"000000011",
  35232=>"000000000",
  35233=>"110111011",
  35234=>"111111111",
  35235=>"000000111",
  35236=>"111011011",
  35237=>"111111010",
  35238=>"111111111",
  35239=>"000100111",
  35240=>"100100111",
  35241=>"011111111",
  35242=>"000100111",
  35243=>"001100111",
  35244=>"111111111",
  35245=>"101111011",
  35246=>"000000111",
  35247=>"111111111",
  35248=>"011010011",
  35249=>"000000000",
  35250=>"000000000",
  35251=>"001001001",
  35252=>"111101001",
  35253=>"101001000",
  35254=>"001001011",
  35255=>"101111100",
  35256=>"110111000",
  35257=>"000001111",
  35258=>"100100000",
  35259=>"111111111",
  35260=>"111111111",
  35261=>"000000000",
  35262=>"000100100",
  35263=>"011011001",
  35264=>"000000000",
  35265=>"001011001",
  35266=>"000000000",
  35267=>"000000000",
  35268=>"011001000",
  35269=>"111111111",
  35270=>"011101001",
  35271=>"000000111",
  35272=>"011100100",
  35273=>"111111000",
  35274=>"001000100",
  35275=>"000000000",
  35276=>"111111111",
  35277=>"101101101",
  35278=>"011111100",
  35279=>"000000000",
  35280=>"000000100",
  35281=>"111111000",
  35282=>"111111100",
  35283=>"101000111",
  35284=>"000000000",
  35285=>"000000000",
  35286=>"001101111",
  35287=>"100111111",
  35288=>"000000000",
  35289=>"000110100",
  35290=>"000110011",
  35291=>"000000000",
  35292=>"010011011",
  35293=>"101000000",
  35294=>"011010000",
  35295=>"011011001",
  35296=>"100000100",
  35297=>"111111111",
  35298=>"011111111",
  35299=>"111001011",
  35300=>"100101001",
  35301=>"011011011",
  35302=>"000000000",
  35303=>"000000010",
  35304=>"001001000",
  35305=>"000011011",
  35306=>"100001111",
  35307=>"011011110",
  35308=>"111110110",
  35309=>"100110100",
  35310=>"110100100",
  35311=>"011100111",
  35312=>"001001111",
  35313=>"000001011",
  35314=>"000000000",
  35315=>"001111111",
  35316=>"111111111",
  35317=>"011110100",
  35318=>"110000000",
  35319=>"110010100",
  35320=>"000000000",
  35321=>"100100100",
  35322=>"000000000",
  35323=>"001000000",
  35324=>"000010110",
  35325=>"000100111",
  35326=>"001011000",
  35327=>"000000100",
  35328=>"110111100",
  35329=>"000000100",
  35330=>"000100111",
  35331=>"100000000",
  35332=>"000000000",
  35333=>"000000000",
  35334=>"111111111",
  35335=>"000000000",
  35336=>"111011011",
  35337=>"110000000",
  35338=>"000001111",
  35339=>"000000100",
  35340=>"000001001",
  35341=>"010110000",
  35342=>"011001001",
  35343=>"111111111",
  35344=>"101101100",
  35345=>"111111000",
  35346=>"111000000",
  35347=>"011001111",
  35348=>"001001111",
  35349=>"000000000",
  35350=>"000111111",
  35351=>"000000000",
  35352=>"000100100",
  35353=>"011001101",
  35354=>"000011111",
  35355=>"100100000",
  35356=>"000000000",
  35357=>"000111110",
  35358=>"000100110",
  35359=>"001000111",
  35360=>"111111011",
  35361=>"111111111",
  35362=>"000010000",
  35363=>"101000100",
  35364=>"000000000",
  35365=>"000000000",
  35366=>"111111000",
  35367=>"011011001",
  35368=>"000111100",
  35369=>"111111111",
  35370=>"111111111",
  35371=>"101000000",
  35372=>"010111110",
  35373=>"001011111",
  35374=>"110000001",
  35375=>"101100101",
  35376=>"000001000",
  35377=>"111111111",
  35378=>"100111111",
  35379=>"100011111",
  35380=>"110110000",
  35381=>"100000100",
  35382=>"001111111",
  35383=>"101111111",
  35384=>"000001101",
  35385=>"111111101",
  35386=>"000001111",
  35387=>"000000100",
  35388=>"010000111",
  35389=>"001001001",
  35390=>"111100100",
  35391=>"111000010",
  35392=>"101111110",
  35393=>"110000011",
  35394=>"000011011",
  35395=>"011001111",
  35396=>"111111100",
  35397=>"011011111",
  35398=>"111111110",
  35399=>"000000000",
  35400=>"000000100",
  35401=>"001000010",
  35402=>"111110011",
  35403=>"100101001",
  35404=>"111100000",
  35405=>"000001111",
  35406=>"111111111",
  35407=>"011111111",
  35408=>"000000110",
  35409=>"110110000",
  35410=>"111110000",
  35411=>"100111100",
  35412=>"111111111",
  35413=>"001001000",
  35414=>"100000000",
  35415=>"000111111",
  35416=>"000000000",
  35417=>"111111111",
  35418=>"111001111",
  35419=>"110010000",
  35420=>"111111111",
  35421=>"000000000",
  35422=>"111000000",
  35423=>"000111011",
  35424=>"011000000",
  35425=>"111111110",
  35426=>"111111111",
  35427=>"010000000",
  35428=>"111111111",
  35429=>"111111111",
  35430=>"000000001",
  35431=>"111100000",
  35432=>"110111111",
  35433=>"111111111",
  35434=>"011011010",
  35435=>"111110101",
  35436=>"100000000",
  35437=>"000000001",
  35438=>"000000100",
  35439=>"111110010",
  35440=>"110111111",
  35441=>"010000110",
  35442=>"010010010",
  35443=>"101111111",
  35444=>"000000001",
  35445=>"001011001",
  35446=>"111111111",
  35447=>"111111111",
  35448=>"000000111",
  35449=>"000000000",
  35450=>"111100100",
  35451=>"011000000",
  35452=>"000000000",
  35453=>"011011001",
  35454=>"111111000",
  35455=>"000111101",
  35456=>"000110111",
  35457=>"001001011",
  35458=>"111000000",
  35459=>"000000100",
  35460=>"000000010",
  35461=>"000000110",
  35462=>"000000000",
  35463=>"110110000",
  35464=>"000001111",
  35465=>"001000110",
  35466=>"111111001",
  35467=>"111111111",
  35468=>"011111111",
  35469=>"011000000",
  35470=>"110000100",
  35471=>"000111111",
  35472=>"000000000",
  35473=>"000000000",
  35474=>"000100111",
  35475=>"111111001",
  35476=>"010100000",
  35477=>"000000000",
  35478=>"001000000",
  35479=>"000000000",
  35480=>"111111000",
  35481=>"101001111",
  35482=>"000000111",
  35483=>"000000000",
  35484=>"001111011",
  35485=>"111111110",
  35486=>"000000111",
  35487=>"111001000",
  35488=>"111111111",
  35489=>"111100100",
  35490=>"000000100",
  35491=>"000001111",
  35492=>"111111110",
  35493=>"111111111",
  35494=>"000000000",
  35495=>"011010011",
  35496=>"000000000",
  35497=>"111110111",
  35498=>"000111111",
  35499=>"111111110",
  35500=>"111001000",
  35501=>"001000000",
  35502=>"000000100",
  35503=>"111011000",
  35504=>"000000000",
  35505=>"000000011",
  35506=>"000000000",
  35507=>"111111111",
  35508=>"111101000",
  35509=>"101101000",
  35510=>"001011000",
  35511=>"111000011",
  35512=>"000001011",
  35513=>"000000000",
  35514=>"001000000",
  35515=>"100000000",
  35516=>"000011111",
  35517=>"111111001",
  35518=>"100000011",
  35519=>"111111110",
  35520=>"000001000",
  35521=>"110100000",
  35522=>"111111111",
  35523=>"111110000",
  35524=>"000000000",
  35525=>"000000011",
  35526=>"110111111",
  35527=>"000010000",
  35528=>"000010000",
  35529=>"000000010",
  35530=>"010000000",
  35531=>"011111011",
  35532=>"010010111",
  35533=>"010000000",
  35534=>"001001001",
  35535=>"111111000",
  35536=>"010011111",
  35537=>"000000000",
  35538=>"000100111",
  35539=>"001001001",
  35540=>"000000000",
  35541=>"001110000",
  35542=>"011011000",
  35543=>"111111101",
  35544=>"111100000",
  35545=>"000000100",
  35546=>"000000000",
  35547=>"000010010",
  35548=>"100000101",
  35549=>"000000111",
  35550=>"111111000",
  35551=>"111111110",
  35552=>"000000000",
  35553=>"111111010",
  35554=>"010000000",
  35555=>"000000001",
  35556=>"001001011",
  35557=>"000000000",
  35558=>"111100101",
  35559=>"111111111",
  35560=>"000000000",
  35561=>"111111110",
  35562=>"100101111",
  35563=>"111111111",
  35564=>"111111100",
  35565=>"011000000",
  35566=>"111111100",
  35567=>"000000011",
  35568=>"001001010",
  35569=>"111001111",
  35570=>"000001111",
  35571=>"011111011",
  35572=>"000000000",
  35573=>"000000010",
  35574=>"011010000",
  35575=>"110110110",
  35576=>"000001011",
  35577=>"000000000",
  35578=>"111110000",
  35579=>"010000000",
  35580=>"100000011",
  35581=>"101001001",
  35582=>"111111111",
  35583=>"111110111",
  35584=>"000000001",
  35585=>"001010010",
  35586=>"110111111",
  35587=>"111011000",
  35588=>"111111001",
  35589=>"111111111",
  35590=>"111111000",
  35591=>"000000000",
  35592=>"111111000",
  35593=>"000000000",
  35594=>"000000000",
  35595=>"011000111",
  35596=>"110110000",
  35597=>"000000000",
  35598=>"111111000",
  35599=>"000010111",
  35600=>"000000001",
  35601=>"100000000",
  35602=>"000001111",
  35603=>"000000111",
  35604=>"000000000",
  35605=>"110000100",
  35606=>"011011011",
  35607=>"100000111",
  35608=>"001001000",
  35609=>"000000100",
  35610=>"000110111",
  35611=>"111111011",
  35612=>"000000000",
  35613=>"000000000",
  35614=>"000000111",
  35615=>"111111000",
  35616=>"011011011",
  35617=>"111111000",
  35618=>"001000000",
  35619=>"111111001",
  35620=>"100101001",
  35621=>"100110111",
  35622=>"110010110",
  35623=>"111111111",
  35624=>"111110000",
  35625=>"000001011",
  35626=>"000000011",
  35627=>"111101111",
  35628=>"000000000",
  35629=>"000000110",
  35630=>"100000000",
  35631=>"110000000",
  35632=>"110110110",
  35633=>"001001000",
  35634=>"000000000",
  35635=>"001111111",
  35636=>"100100110",
  35637=>"000000110",
  35638=>"011111111",
  35639=>"000000000",
  35640=>"100000000",
  35641=>"111000001",
  35642=>"111101111",
  35643=>"110100100",
  35644=>"000000111",
  35645=>"000000000",
  35646=>"011011000",
  35647=>"010110111",
  35648=>"111111111",
  35649=>"000011010",
  35650=>"000001011",
  35651=>"000010110",
  35652=>"000110110",
  35653=>"111111000",
  35654=>"000000111",
  35655=>"111111000",
  35656=>"000000000",
  35657=>"011110100",
  35658=>"100100000",
  35659=>"110110100",
  35660=>"111111000",
  35661=>"001111000",
  35662=>"111111111",
  35663=>"100111111",
  35664=>"111110000",
  35665=>"111111001",
  35666=>"110110000",
  35667=>"100000000",
  35668=>"111111110",
  35669=>"011001001",
  35670=>"000001111",
  35671=>"111111111",
  35672=>"111111111",
  35673=>"000000000",
  35674=>"000000000",
  35675=>"001111001",
  35676=>"111111111",
  35677=>"011111111",
  35678=>"000000000",
  35679=>"010000011",
  35680=>"111101111",
  35681=>"000111111",
  35682=>"110011011",
  35683=>"001111111",
  35684=>"000000010",
  35685=>"000100010",
  35686=>"000000000",
  35687=>"001000000",
  35688=>"001111001",
  35689=>"111010110",
  35690=>"111111000",
  35691=>"000000001",
  35692=>"011110000",
  35693=>"000000001",
  35694=>"111111111",
  35695=>"010010000",
  35696=>"000100110",
  35697=>"011000000",
  35698=>"111111110",
  35699=>"111111000",
  35700=>"101101111",
  35701=>"000000111",
  35702=>"100100111",
  35703=>"000000111",
  35704=>"011111111",
  35705=>"000111001",
  35706=>"111111111",
  35707=>"111111111",
  35708=>"111111111",
  35709=>"000000110",
  35710=>"000000111",
  35711=>"111111111",
  35712=>"000000000",
  35713=>"111111000",
  35714=>"000000011",
  35715=>"000100111",
  35716=>"100101111",
  35717=>"000000000",
  35718=>"101100111",
  35719=>"001000100",
  35720=>"000111111",
  35721=>"111111100",
  35722=>"001001011",
  35723=>"010000110",
  35724=>"111100111",
  35725=>"010010000",
  35726=>"000000100",
  35727=>"110000000",
  35728=>"110000010",
  35729=>"000001111",
  35730=>"110111111",
  35731=>"000001111",
  35732=>"111111111",
  35733=>"000000001",
  35734=>"111000000",
  35735=>"100100000",
  35736=>"000000001",
  35737=>"101101110",
  35738=>"111111111",
  35739=>"000000111",
  35740=>"000000000",
  35741=>"000000000",
  35742=>"000000000",
  35743=>"100100101",
  35744=>"111000000",
  35745=>"001011010",
  35746=>"000111111",
  35747=>"001111111",
  35748=>"110000111",
  35749=>"000011011",
  35750=>"111000000",
  35751=>"000000111",
  35752=>"000001001",
  35753=>"011000100",
  35754=>"110100111",
  35755=>"000000000",
  35756=>"111110000",
  35757=>"001001101",
  35758=>"010010111",
  35759=>"000000000",
  35760=>"100100000",
  35761=>"000000000",
  35762=>"111100001",
  35763=>"000000000",
  35764=>"000000100",
  35765=>"101000000",
  35766=>"000000001",
  35767=>"111111111",
  35768=>"001001000",
  35769=>"101101000",
  35770=>"100110001",
  35771=>"000000111",
  35772=>"101001000",
  35773=>"011001000",
  35774=>"100100000",
  35775=>"010010010",
  35776=>"000000000",
  35777=>"111011011",
  35778=>"000111011",
  35779=>"000000101",
  35780=>"000011111",
  35781=>"111011011",
  35782=>"111111111",
  35783=>"000000101",
  35784=>"100111000",
  35785=>"111000000",
  35786=>"111111100",
  35787=>"000000000",
  35788=>"000000000",
  35789=>"000000000",
  35790=>"000000010",
  35791=>"111111000",
  35792=>"111111111",
  35793=>"000000000",
  35794=>"111111111",
  35795=>"010000011",
  35796=>"111110011",
  35797=>"000011111",
  35798=>"001000010",
  35799=>"111101000",
  35800=>"111111111",
  35801=>"110110000",
  35802=>"010000001",
  35803=>"111111111",
  35804=>"101000000",
  35805=>"011101111",
  35806=>"001011000",
  35807=>"010010000",
  35808=>"111111110",
  35809=>"111111000",
  35810=>"000000000",
  35811=>"010111001",
  35812=>"110100000",
  35813=>"100000001",
  35814=>"011011000",
  35815=>"000000111",
  35816=>"000001001",
  35817=>"000011001",
  35818=>"110110111",
  35819=>"000000000",
  35820=>"000011011",
  35821=>"111111001",
  35822=>"010010010",
  35823=>"111000001",
  35824=>"111110000",
  35825=>"111000011",
  35826=>"111100001",
  35827=>"000000010",
  35828=>"000000000",
  35829=>"000010011",
  35830=>"000000000",
  35831=>"011001011",
  35832=>"011111011",
  35833=>"000000010",
  35834=>"111111111",
  35835=>"000000100",
  35836=>"001001000",
  35837=>"010000100",
  35838=>"000000000",
  35839=>"111111101",
  35840=>"010000000",
  35841=>"111101111",
  35842=>"111111111",
  35843=>"000000111",
  35844=>"000000000",
  35845=>"110111111",
  35846=>"000000000",
  35847=>"000000000",
  35848=>"100000111",
  35849=>"000000000",
  35850=>"110110110",
  35851=>"111011011",
  35852=>"100000000",
  35853=>"010110111",
  35854=>"000110111",
  35855=>"100100111",
  35856=>"111111111",
  35857=>"111111110",
  35858=>"000000000",
  35859=>"000000000",
  35860=>"000000000",
  35861=>"000011111",
  35862=>"111111110",
  35863=>"111111110",
  35864=>"111110110",
  35865=>"100111111",
  35866=>"000000000",
  35867=>"111110111",
  35868=>"111111111",
  35869=>"111111111",
  35870=>"110111111",
  35871=>"011011001",
  35872=>"111011000",
  35873=>"111110000",
  35874=>"111111111",
  35875=>"111111111",
  35876=>"000000111",
  35877=>"111000111",
  35878=>"100111111",
  35879=>"001000001",
  35880=>"111110000",
  35881=>"000000000",
  35882=>"111100111",
  35883=>"001000011",
  35884=>"000000000",
  35885=>"111111111",
  35886=>"111111000",
  35887=>"111111101",
  35888=>"000000000",
  35889=>"000000000",
  35890=>"000111100",
  35891=>"000000001",
  35892=>"111100000",
  35893=>"101111111",
  35894=>"110100100",
  35895=>"111111000",
  35896=>"000000001",
  35897=>"111111111",
  35898=>"111111111",
  35899=>"111111111",
  35900=>"111111011",
  35901=>"111000000",
  35902=>"000000110",
  35903=>"100100111",
  35904=>"001011001",
  35905=>"000000111",
  35906=>"000000000",
  35907=>"000011111",
  35908=>"111111111",
  35909=>"000001111",
  35910=>"000001011",
  35911=>"111111111",
  35912=>"000110000",
  35913=>"001001111",
  35914=>"110111110",
  35915=>"110111011",
  35916=>"000000000",
  35917=>"110000000",
  35918=>"110110010",
  35919=>"000011000",
  35920=>"000000111",
  35921=>"000000000",
  35922=>"000110110",
  35923=>"101111111",
  35924=>"000000000",
  35925=>"010011001",
  35926=>"110100000",
  35927=>"000000000",
  35928=>"001001111",
  35929=>"000101111",
  35930=>"010110100",
  35931=>"111010010",
  35932=>"001000000",
  35933=>"111111111",
  35934=>"101101111",
  35935=>"000000000",
  35936=>"000000000",
  35937=>"001011010",
  35938=>"100100100",
  35939=>"000000000",
  35940=>"000011011",
  35941=>"011011111",
  35942=>"011001000",
  35943=>"111111111",
  35944=>"001111000",
  35945=>"000010111",
  35946=>"100110111",
  35947=>"110010010",
  35948=>"000000000",
  35949=>"000000000",
  35950=>"011111011",
  35951=>"111111000",
  35952=>"111111111",
  35953=>"010111111",
  35954=>"111111100",
  35955=>"111000000",
  35956=>"000000000",
  35957=>"111111000",
  35958=>"111111111",
  35959=>"000000110",
  35960=>"000000000",
  35961=>"000110100",
  35962=>"000000000",
  35963=>"000000000",
  35964=>"111111111",
  35965=>"000000000",
  35966=>"000000110",
  35967=>"000000000",
  35968=>"000010000",
  35969=>"111111111",
  35970=>"000000011",
  35971=>"110000000",
  35972=>"000000001",
  35973=>"111001000",
  35974=>"000000000",
  35975=>"001001000",
  35976=>"111111111",
  35977=>"111000000",
  35978=>"000000001",
  35979=>"011111111",
  35980=>"111011011",
  35981=>"111111111",
  35982=>"000010000",
  35983=>"000000111",
  35984=>"111111111",
  35985=>"110000000",
  35986=>"111111100",
  35987=>"111000000",
  35988=>"000000100",
  35989=>"110110000",
  35990=>"000000000",
  35991=>"111111111",
  35992=>"100100110",
  35993=>"000000000",
  35994=>"000101100",
  35995=>"000000111",
  35996=>"000000000",
  35997=>"111110111",
  35998=>"010100100",
  35999=>"111001011",
  36000=>"000100000",
  36001=>"111111010",
  36002=>"011001111",
  36003=>"111111111",
  36004=>"000000000",
  36005=>"011111111",
  36006=>"111101101",
  36007=>"111111011",
  36008=>"000001000",
  36009=>"000010111",
  36010=>"010010110",
  36011=>"000000000",
  36012=>"000000000",
  36013=>"110010000",
  36014=>"000000000",
  36015=>"000000000",
  36016=>"000000000",
  36017=>"001011011",
  36018=>"110111111",
  36019=>"000000000",
  36020=>"111001111",
  36021=>"011001000",
  36022=>"110010000",
  36023=>"100100110",
  36024=>"000000100",
  36025=>"111111111",
  36026=>"000000000",
  36027=>"000000000",
  36028=>"000010000",
  36029=>"111111111",
  36030=>"000000001",
  36031=>"001011111",
  36032=>"111111111",
  36033=>"000000011",
  36034=>"111110111",
  36035=>"000000000",
  36036=>"111011111",
  36037=>"000000000",
  36038=>"011001000",
  36039=>"000000001",
  36040=>"000000000",
  36041=>"000000000",
  36042=>"111100100",
  36043=>"010010000",
  36044=>"111111011",
  36045=>"111111111",
  36046=>"111111111",
  36047=>"000000000",
  36048=>"111111100",
  36049=>"111111110",
  36050=>"110000110",
  36051=>"110110000",
  36052=>"111001111",
  36053=>"111110000",
  36054=>"010010000",
  36055=>"101001011",
  36056=>"000000000",
  36057=>"000000111",
  36058=>"111111011",
  36059=>"011011000",
  36060=>"000000000",
  36061=>"110010000",
  36062=>"111011011",
  36063=>"111111000",
  36064=>"000000000",
  36065=>"111000111",
  36066=>"110000000",
  36067=>"000000000",
  36068=>"100101100",
  36069=>"010111111",
  36070=>"110111111",
  36071=>"000000000",
  36072=>"000001000",
  36073=>"000000000",
  36074=>"111110000",
  36075=>"001000010",
  36076=>"111111011",
  36077=>"111000001",
  36078=>"001000000",
  36079=>"000111111",
  36080=>"010111111",
  36081=>"111001100",
  36082=>"011111111",
  36083=>"000000101",
  36084=>"000000000",
  36085=>"001001001",
  36086=>"011011011",
  36087=>"000010000",
  36088=>"111111110",
  36089=>"000011001",
  36090=>"000000000",
  36091=>"000000000",
  36092=>"111111110",
  36093=>"000000000",
  36094=>"000110000",
  36095=>"110111111",
  36096=>"000000000",
  36097=>"000000000",
  36098=>"000010010",
  36099=>"000000000",
  36100=>"101111111",
  36101=>"010010111",
  36102=>"000000110",
  36103=>"000000111",
  36104=>"000000000",
  36105=>"000000000",
  36106=>"000000111",
  36107=>"111111111",
  36108=>"111000000",
  36109=>"111111111",
  36110=>"000001000",
  36111=>"110111111",
  36112=>"000000000",
  36113=>"000000110",
  36114=>"010000001",
  36115=>"000111111",
  36116=>"000000000",
  36117=>"000000000",
  36118=>"111111001",
  36119=>"000101101",
  36120=>"111111110",
  36121=>"111111111",
  36122=>"100000000",
  36123=>"000000000",
  36124=>"111011011",
  36125=>"100000000",
  36126=>"111100000",
  36127=>"111001111",
  36128=>"000000000",
  36129=>"000101101",
  36130=>"111111111",
  36131=>"111111111",
  36132=>"100000000",
  36133=>"000000111",
  36134=>"111110110",
  36135=>"111111111",
  36136=>"000000000",
  36137=>"110110111",
  36138=>"111110000",
  36139=>"000000000",
  36140=>"000000000",
  36141=>"100100000",
  36142=>"000000000",
  36143=>"010000000",
  36144=>"000110110",
  36145=>"110110111",
  36146=>"111011101",
  36147=>"111111111",
  36148=>"000000000",
  36149=>"111111111",
  36150=>"100110100",
  36151=>"111111111",
  36152=>"111011001",
  36153=>"111111111",
  36154=>"000010010",
  36155=>"000011001",
  36156=>"111111111",
  36157=>"001000000",
  36158=>"011011011",
  36159=>"000000000",
  36160=>"111111111",
  36161=>"111001101",
  36162=>"000000000",
  36163=>"111011111",
  36164=>"000000111",
  36165=>"111111111",
  36166=>"111111111",
  36167=>"000000000",
  36168=>"010000000",
  36169=>"001000101",
  36170=>"110000000",
  36171=>"111101001",
  36172=>"111001001",
  36173=>"111011000",
  36174=>"010000001",
  36175=>"111111000",
  36176=>"000000110",
  36177=>"010010001",
  36178=>"000010011",
  36179=>"000000000",
  36180=>"000010010",
  36181=>"111111011",
  36182=>"110000000",
  36183=>"110110000",
  36184=>"000000000",
  36185=>"111111111",
  36186=>"000000000",
  36187=>"000000001",
  36188=>"111111111",
  36189=>"111111000",
  36190=>"111111111",
  36191=>"111111111",
  36192=>"000000000",
  36193=>"111111111",
  36194=>"111101100",
  36195=>"000010010",
  36196=>"110110111",
  36197=>"110000100",
  36198=>"111111111",
  36199=>"000000000",
  36200=>"000000000",
  36201=>"111011011",
  36202=>"111111111",
  36203=>"000000011",
  36204=>"001111111",
  36205=>"001110100",
  36206=>"110110110",
  36207=>"010010110",
  36208=>"011111011",
  36209=>"000000000",
  36210=>"000000011",
  36211=>"111001001",
  36212=>"000000000",
  36213=>"100110110",
  36214=>"000001001",
  36215=>"100100000",
  36216=>"111111111",
  36217=>"000000001",
  36218=>"111111100",
  36219=>"111111100",
  36220=>"010001111",
  36221=>"111111111",
  36222=>"110000000",
  36223=>"000011111",
  36224=>"000000010",
  36225=>"000000011",
  36226=>"111111111",
  36227=>"000000000",
  36228=>"000000000",
  36229=>"111111111",
  36230=>"111111111",
  36231=>"000001001",
  36232=>"111000000",
  36233=>"101111110",
  36234=>"111111100",
  36235=>"010111111",
  36236=>"000000010",
  36237=>"111101111",
  36238=>"101101110",
  36239=>"000000000",
  36240=>"000010000",
  36241=>"000000000",
  36242=>"000000000",
  36243=>"111111111",
  36244=>"000000000",
  36245=>"000000000",
  36246=>"000001111",
  36247=>"100000000",
  36248=>"011011000",
  36249=>"011111111",
  36250=>"000000100",
  36251=>"000000011",
  36252=>"111111011",
  36253=>"010100110",
  36254=>"100100000",
  36255=>"000000000",
  36256=>"011000000",
  36257=>"111111110",
  36258=>"011000010",
  36259=>"011111011",
  36260=>"000000001",
  36261=>"000000000",
  36262=>"111111111",
  36263=>"111111111",
  36264=>"111001000",
  36265=>"111100111",
  36266=>"110000111",
  36267=>"111100100",
  36268=>"110110110",
  36269=>"000000000",
  36270=>"000000000",
  36271=>"000000000",
  36272=>"011111111",
  36273=>"000111111",
  36274=>"111100000",
  36275=>"000000000",
  36276=>"100000000",
  36277=>"000100000",
  36278=>"111111111",
  36279=>"000111111",
  36280=>"000000011",
  36281=>"000000000",
  36282=>"111111111",
  36283=>"001001001",
  36284=>"000001001",
  36285=>"000000001",
  36286=>"111101101",
  36287=>"110100100",
  36288=>"111111111",
  36289=>"000000000",
  36290=>"000000000",
  36291=>"001000000",
  36292=>"001000000",
  36293=>"000000111",
  36294=>"100111111",
  36295=>"000000000",
  36296=>"000110100",
  36297=>"011111110",
  36298=>"000000000",
  36299=>"010111111",
  36300=>"000000000",
  36301=>"000000000",
  36302=>"010011111",
  36303=>"000011011",
  36304=>"000000000",
  36305=>"111001111",
  36306=>"110100000",
  36307=>"000000000",
  36308=>"000001000",
  36309=>"000000000",
  36310=>"110000000",
  36311=>"111111111",
  36312=>"111111111",
  36313=>"000000000",
  36314=>"110100111",
  36315=>"000000000",
  36316=>"010000001",
  36317=>"111111111",
  36318=>"000000000",
  36319=>"111110111",
  36320=>"000000000",
  36321=>"110000000",
  36322=>"100111110",
  36323=>"000111111",
  36324=>"111011000",
  36325=>"000010000",
  36326=>"000000000",
  36327=>"111011000",
  36328=>"111111111",
  36329=>"000000000",
  36330=>"111001001",
  36331=>"111111111",
  36332=>"111100000",
  36333=>"111101001",
  36334=>"111111100",
  36335=>"000000100",
  36336=>"000000000",
  36337=>"000111000",
  36338=>"100110000",
  36339=>"011111011",
  36340=>"100000000",
  36341=>"111111111",
  36342=>"111110111",
  36343=>"000000000",
  36344=>"000011111",
  36345=>"011000110",
  36346=>"111111101",
  36347=>"111001000",
  36348=>"011111111",
  36349=>"000000110",
  36350=>"110000000",
  36351=>"000000000",
  36352=>"111000000",
  36353=>"011000000",
  36354=>"101000000",
  36355=>"110110111",
  36356=>"100110110",
  36357=>"111001111",
  36358=>"000000000",
  36359=>"111111111",
  36360=>"111001000",
  36361=>"000000000",
  36362=>"000000110",
  36363=>"111001000",
  36364=>"100100000",
  36365=>"110101010",
  36366=>"111001100",
  36367=>"000010010",
  36368=>"000001001",
  36369=>"111111111",
  36370=>"111000000",
  36371=>"111010000",
  36372=>"110000000",
  36373=>"111111110",
  36374=>"000111111",
  36375=>"000000000",
  36376=>"110100100",
  36377=>"000110111",
  36378=>"111011000",
  36379=>"111011011",
  36380=>"000000000",
  36381=>"111101100",
  36382=>"001100111",
  36383=>"111110111",
  36384=>"100000000",
  36385=>"000010111",
  36386=>"100000000",
  36387=>"011000000",
  36388=>"000000000",
  36389=>"000110110",
  36390=>"111001111",
  36391=>"100000001",
  36392=>"111100000",
  36393=>"111001001",
  36394=>"001000000",
  36395=>"111001101",
  36396=>"100000000",
  36397=>"100000000",
  36398=>"000110111",
  36399=>"000000111",
  36400=>"111111111",
  36401=>"000000001",
  36402=>"011001011",
  36403=>"011011111",
  36404=>"000000000",
  36405=>"110110110",
  36406=>"111110111",
  36407=>"011000000",
  36408=>"000000000",
  36409=>"000000000",
  36410=>"000000011",
  36411=>"011011000",
  36412=>"111111111",
  36413=>"111111111",
  36414=>"000000001",
  36415=>"111011111",
  36416=>"111111001",
  36417=>"000000000",
  36418=>"011111111",
  36419=>"100000011",
  36420=>"100000000",
  36421=>"000000011",
  36422=>"101000000",
  36423=>"111111111",
  36424=>"011000000",
  36425=>"001101111",
  36426=>"000111111",
  36427=>"001001000",
  36428=>"111111111",
  36429=>"111111000",
  36430=>"111101111",
  36431=>"010000001",
  36432=>"100100111",
  36433=>"000000110",
  36434=>"110000000",
  36435=>"110101101",
  36436=>"000000000",
  36437=>"111000000",
  36438=>"011001111",
  36439=>"000000000",
  36440=>"110011000",
  36441=>"111100100",
  36442=>"000111111",
  36443=>"000001001",
  36444=>"111011111",
  36445=>"000000000",
  36446=>"000001001",
  36447=>"111111101",
  36448=>"100000100",
  36449=>"111011111",
  36450=>"001001010",
  36451=>"000000000",
  36452=>"000000111",
  36453=>"101111111",
  36454=>"000000000",
  36455=>"000000001",
  36456=>"000000000",
  36457=>"011011010",
  36458=>"000000000",
  36459=>"000000000",
  36460=>"111110110",
  36461=>"000000000",
  36462=>"001001101",
  36463=>"000001001",
  36464=>"110111011",
  36465=>"111111011",
  36466=>"011011011",
  36467=>"000000111",
  36468=>"111010000",
  36469=>"111111000",
  36470=>"000000000",
  36471=>"111011111",
  36472=>"000000000",
  36473=>"111101100",
  36474=>"111101000",
  36475=>"001000001",
  36476=>"001001111",
  36477=>"110111011",
  36478=>"111111110",
  36479=>"000000000",
  36480=>"000000000",
  36481=>"111111000",
  36482=>"111000000",
  36483=>"010000011",
  36484=>"110010011",
  36485=>"000000111",
  36486=>"111111111",
  36487=>"110111000",
  36488=>"111111011",
  36489=>"100000011",
  36490=>"110000001",
  36491=>"111111111",
  36492=>"000010111",
  36493=>"000000111",
  36494=>"000000001",
  36495=>"110111111",
  36496=>"111111111",
  36497=>"111111111",
  36498=>"111001000",
  36499=>"110000000",
  36500=>"000111111",
  36501=>"000111111",
  36502=>"000000000",
  36503=>"000000000",
  36504=>"111111111",
  36505=>"011111111",
  36506=>"000000011",
  36507=>"001001001",
  36508=>"001111111",
  36509=>"100000000",
  36510=>"000000000",
  36511=>"000000000",
  36512=>"001000000",
  36513=>"110100000",
  36514=>"101000101",
  36515=>"111001001",
  36516=>"110000000",
  36517=>"100110111",
  36518=>"111001111",
  36519=>"111011010",
  36520=>"111111111",
  36521=>"101000000",
  36522=>"000100111",
  36523=>"000000111",
  36524=>"001111111",
  36525=>"101101111",
  36526=>"111111111",
  36527=>"000000111",
  36528=>"000000000",
  36529=>"011111011",
  36530=>"110111111",
  36531=>"000000000",
  36532=>"000000000",
  36533=>"111000000",
  36534=>"000111000",
  36535=>"000000000",
  36536=>"111001000",
  36537=>"000000000",
  36538=>"101111000",
  36539=>"111111000",
  36540=>"001000111",
  36541=>"000000000",
  36542=>"000000110",
  36543=>"111111000",
  36544=>"001000000",
  36545=>"000000000",
  36546=>"110111101",
  36547=>"101111000",
  36548=>"000000000",
  36549=>"111000000",
  36550=>"100000000",
  36551=>"001001000",
  36552=>"111111111",
  36553=>"000111111",
  36554=>"111101001",
  36555=>"000001111",
  36556=>"000000000",
  36557=>"111000000",
  36558=>"000111111",
  36559=>"111111111",
  36560=>"000000111",
  36561=>"011011111",
  36562=>"101011000",
  36563=>"000000000",
  36564=>"000001111",
  36565=>"000001000",
  36566=>"111111111",
  36567=>"111001101",
  36568=>"000100111",
  36569=>"100100101",
  36570=>"010000011",
  36571=>"011111111",
  36572=>"000000011",
  36573=>"000111111",
  36574=>"000000111",
  36575=>"100110111",
  36576=>"000000000",
  36577=>"011111111",
  36578=>"100111000",
  36579=>"000000000",
  36580=>"111111111",
  36581=>"000100100",
  36582=>"100111111",
  36583=>"111111010",
  36584=>"000000000",
  36585=>"111111011",
  36586=>"111111000",
  36587=>"000000000",
  36588=>"110111011",
  36589=>"001011111",
  36590=>"110111001",
  36591=>"000110110",
  36592=>"000000000",
  36593=>"000000000",
  36594=>"011111011",
  36595=>"111000000",
  36596=>"000000000",
  36597=>"110110011",
  36598=>"111000011",
  36599=>"111111111",
  36600=>"000000110",
  36601=>"111011000",
  36602=>"100000000",
  36603=>"001000000",
  36604=>"111111110",
  36605=>"100000000",
  36606=>"001000100",
  36607=>"000000000",
  36608=>"100100110",
  36609=>"110110100",
  36610=>"000000000",
  36611=>"111001001",
  36612=>"000000000",
  36613=>"000000000",
  36614=>"001001001",
  36615=>"111111100",
  36616=>"111001001",
  36617=>"000000000",
  36618=>"000000000",
  36619=>"000000001",
  36620=>"110110110",
  36621=>"110111111",
  36622=>"110110110",
  36623=>"111111111",
  36624=>"101000000",
  36625=>"000000100",
  36626=>"111111111",
  36627=>"111100100",
  36628=>"111010000",
  36629=>"111111111",
  36630=>"001001101",
  36631=>"001011001",
  36632=>"000000001",
  36633=>"000000111",
  36634=>"000110111",
  36635=>"000000010",
  36636=>"100110110",
  36637=>"111000000",
  36638=>"110110110",
  36639=>"111111111",
  36640=>"000000000",
  36641=>"000000001",
  36642=>"001111111",
  36643=>"000000001",
  36644=>"111111111",
  36645=>"111111111",
  36646=>"000000110",
  36647=>"011011011",
  36648=>"111111111",
  36649=>"000000000",
  36650=>"111000111",
  36651=>"111001000",
  36652=>"111101101",
  36653=>"010000000",
  36654=>"000010000",
  36655=>"001000111",
  36656=>"100100001",
  36657=>"011111111",
  36658=>"111111111",
  36659=>"000000000",
  36660=>"000010010",
  36661=>"111011001",
  36662=>"111000000",
  36663=>"110111111",
  36664=>"100000000",
  36665=>"111001100",
  36666=>"111111111",
  36667=>"111111111",
  36668=>"000000000",
  36669=>"000000001",
  36670=>"000000000",
  36671=>"111111000",
  36672=>"000000000",
  36673=>"111111111",
  36674=>"000100000",
  36675=>"000000111",
  36676=>"000000000",
  36677=>"001100100",
  36678=>"000111111",
  36679=>"000000000",
  36680=>"000000010",
  36681=>"110000000",
  36682=>"100000100",
  36683=>"100110010",
  36684=>"101111001",
  36685=>"010011111",
  36686=>"001001011",
  36687=>"011011111",
  36688=>"111110111",
  36689=>"001111111",
  36690=>"100000111",
  36691=>"111110111",
  36692=>"000000000",
  36693=>"011001011",
  36694=>"100100111",
  36695=>"010011001",
  36696=>"000100110",
  36697=>"111111010",
  36698=>"110000011",
  36699=>"101011111",
  36700=>"000000000",
  36701=>"000000000",
  36702=>"000000000",
  36703=>"011000111",
  36704=>"111001111",
  36705=>"111000000",
  36706=>"000000000",
  36707=>"000000010",
  36708=>"110110001",
  36709=>"111011000",
  36710=>"101000000",
  36711=>"111111111",
  36712=>"010010000",
  36713=>"000000000",
  36714=>"101111111",
  36715=>"111111111",
  36716=>"111111101",
  36717=>"111011011",
  36718=>"001111000",
  36719=>"000000000",
  36720=>"100111111",
  36721=>"000111111",
  36722=>"000000000",
  36723=>"111111111",
  36724=>"000000111",
  36725=>"110111111",
  36726=>"101000000",
  36727=>"111111111",
  36728=>"111001101",
  36729=>"111111000",
  36730=>"111110111",
  36731=>"111110110",
  36732=>"111000000",
  36733=>"000111111",
  36734=>"111111101",
  36735=>"101101111",
  36736=>"011001001",
  36737=>"000000111",
  36738=>"001011111",
  36739=>"011010000",
  36740=>"111100000",
  36741=>"000100100",
  36742=>"001001100",
  36743=>"000000111",
  36744=>"000011111",
  36745=>"000000000",
  36746=>"101111111",
  36747=>"111111110",
  36748=>"111111111",
  36749=>"000000100",
  36750=>"000001100",
  36751=>"111111111",
  36752=>"000000111",
  36753=>"111111000",
  36754=>"100000011",
  36755=>"000100000",
  36756=>"111010100",
  36757=>"000100000",
  36758=>"000000000",
  36759=>"111000000",
  36760=>"111000101",
  36761=>"111111011",
  36762=>"111111111",
  36763=>"111111110",
  36764=>"001000000",
  36765=>"111111110",
  36766=>"000101111",
  36767=>"000000000",
  36768=>"111111111",
  36769=>"001001111",
  36770=>"000000100",
  36771=>"000100111",
  36772=>"000100111",
  36773=>"001000001",
  36774=>"111000000",
  36775=>"111000011",
  36776=>"000000000",
  36777=>"111101111",
  36778=>"000000001",
  36779=>"010010000",
  36780=>"010010000",
  36781=>"101101010",
  36782=>"111111000",
  36783=>"111111111",
  36784=>"111111111",
  36785=>"111111110",
  36786=>"110100000",
  36787=>"000000111",
  36788=>"000011011",
  36789=>"111111000",
  36790=>"000000111",
  36791=>"000000000",
  36792=>"000000101",
  36793=>"101011000",
  36794=>"111011000",
  36795=>"000000000",
  36796=>"000000100",
  36797=>"111111111",
  36798=>"111000100",
  36799=>"010000001",
  36800=>"000000001",
  36801=>"010001111",
  36802=>"111111000",
  36803=>"111111011",
  36804=>"000000111",
  36805=>"011011000",
  36806=>"111000000",
  36807=>"111101000",
  36808=>"111110111",
  36809=>"000110111",
  36810=>"101000000",
  36811=>"000000000",
  36812=>"000000000",
  36813=>"001001001",
  36814=>"100000000",
  36815=>"000000111",
  36816=>"001000111",
  36817=>"000111100",
  36818=>"011111111",
  36819=>"111011000",
  36820=>"111111011",
  36821=>"110111111",
  36822=>"111111110",
  36823=>"111110000",
  36824=>"000101111",
  36825=>"111100000",
  36826=>"000000011",
  36827=>"110110000",
  36828=>"000000000",
  36829=>"111111011",
  36830=>"111011000",
  36831=>"000000100",
  36832=>"110010111",
  36833=>"000000000",
  36834=>"111111111",
  36835=>"111100001",
  36836=>"000000010",
  36837=>"111111111",
  36838=>"010000111",
  36839=>"111111011",
  36840=>"110100111",
  36841=>"000000000",
  36842=>"000000000",
  36843=>"111010100",
  36844=>"000000001",
  36845=>"011001011",
  36846=>"111000110",
  36847=>"110010011",
  36848=>"000000011",
  36849=>"000000000",
  36850=>"111000001",
  36851=>"011000000",
  36852=>"111111000",
  36853=>"001000111",
  36854=>"110111111",
  36855=>"111111101",
  36856=>"010110010",
  36857=>"011111111",
  36858=>"000010000",
  36859=>"000000110",
  36860=>"000000000",
  36861=>"111001000",
  36862=>"000110111",
  36863=>"000000111",
  36864=>"111111111",
  36865=>"001011111",
  36866=>"111111111",
  36867=>"010100100",
  36868=>"001000000",
  36869=>"111011000",
  36870=>"010111111",
  36871=>"000000111",
  36872=>"110000000",
  36873=>"111111000",
  36874=>"110111111",
  36875=>"111111110",
  36876=>"100110110",
  36877=>"011111111",
  36878=>"000000000",
  36879=>"000000000",
  36880=>"001000001",
  36881=>"000110111",
  36882=>"000110000",
  36883=>"110110000",
  36884=>"111111001",
  36885=>"001000000",
  36886=>"100111111",
  36887=>"110100000",
  36888=>"100000000",
  36889=>"000100111",
  36890=>"111000000",
  36891=>"100111111",
  36892=>"000000001",
  36893=>"000000001",
  36894=>"111110110",
  36895=>"000010011",
  36896=>"011000000",
  36897=>"101101000",
  36898=>"110111111",
  36899=>"111000000",
  36900=>"011011111",
  36901=>"111111000",
  36902=>"000000111",
  36903=>"000000001",
  36904=>"111001111",
  36905=>"000111111",
  36906=>"001000001",
  36907=>"011011000",
  36908=>"000111111",
  36909=>"011111111",
  36910=>"100000000",
  36911=>"001011001",
  36912=>"000000000",
  36913=>"000011000",
  36914=>"011011001",
  36915=>"111111000",
  36916=>"101000001",
  36917=>"111101000",
  36918=>"111111000",
  36919=>"001001000",
  36920=>"111111111",
  36921=>"111011011",
  36922=>"010111111",
  36923=>"111000111",
  36924=>"101001101",
  36925=>"000111111",
  36926=>"111111100",
  36927=>"000000001",
  36928=>"011011011",
  36929=>"011001001",
  36930=>"111111111",
  36931=>"010010000",
  36932=>"100111001",
  36933=>"000000000",
  36934=>"000000000",
  36935=>"111111111",
  36936=>"000001000",
  36937=>"000000000",
  36938=>"111000000",
  36939=>"000000000",
  36940=>"111111000",
  36941=>"000000000",
  36942=>"111000000",
  36943=>"000000100",
  36944=>"110111000",
  36945=>"010111111",
  36946=>"111111111",
  36947=>"011111101",
  36948=>"000000001",
  36949=>"111000011",
  36950=>"110000000",
  36951=>"111111111",
  36952=>"011111111",
  36953=>"111111111",
  36954=>"110110111",
  36955=>"010110000",
  36956=>"111001000",
  36957=>"111000000",
  36958=>"100000000",
  36959=>"101101111",
  36960=>"000111111",
  36961=>"111111111",
  36962=>"000111111",
  36963=>"011111000",
  36964=>"111100000",
  36965=>"000000110",
  36966=>"110111011",
  36967=>"000000111",
  36968=>"000000001",
  36969=>"000000000",
  36970=>"000000000",
  36971=>"000010111",
  36972=>"111111111",
  36973=>"000111111",
  36974=>"111001001",
  36975=>"111111111",
  36976=>"111000000",
  36977=>"001000100",
  36978=>"111000110",
  36979=>"100000111",
  36980=>"111111011",
  36981=>"000111110",
  36982=>"000000000",
  36983=>"011110000",
  36984=>"010010000",
  36985=>"111000001",
  36986=>"000001101",
  36987=>"000000000",
  36988=>"001111101",
  36989=>"011111111",
  36990=>"111111010",
  36991=>"110000000",
  36992=>"001000000",
  36993=>"111111101",
  36994=>"111111101",
  36995=>"100100100",
  36996=>"011111111",
  36997=>"011000000",
  36998=>"000100000",
  36999=>"000001101",
  37000=>"000111000",
  37001=>"001011000",
  37002=>"001000000",
  37003=>"100000000",
  37004=>"100001001",
  37005=>"111101000",
  37006=>"101111111",
  37007=>"000000000",
  37008=>"111111000",
  37009=>"110000000",
  37010=>"111100111",
  37011=>"111001000",
  37012=>"000000000",
  37013=>"111001111",
  37014=>"001111111",
  37015=>"000000001",
  37016=>"111000000",
  37017=>"000000111",
  37018=>"000000000",
  37019=>"000000000",
  37020=>"000000000",
  37021=>"110000001",
  37022=>"000101111",
  37023=>"100001000",
  37024=>"000010110",
  37025=>"000010110",
  37026=>"110111110",
  37027=>"011000000",
  37028=>"000100000",
  37029=>"100111111",
  37030=>"010110000",
  37031=>"111100000",
  37032=>"000000000",
  37033=>"001011111",
  37034=>"000000000",
  37035=>"000000000",
  37036=>"111111001",
  37037=>"110110110",
  37038=>"111100111",
  37039=>"000011111",
  37040=>"000000001",
  37041=>"000001111",
  37042=>"000111111",
  37043=>"111100000",
  37044=>"000001111",
  37045=>"000000000",
  37046=>"000000000",
  37047=>"000000000",
  37048=>"111111111",
  37049=>"111000000",
  37050=>"000001101",
  37051=>"000100100",
  37052=>"100100000",
  37053=>"000000000",
  37054=>"111111111",
  37055=>"011111111",
  37056=>"011000101",
  37057=>"000000001",
  37058=>"000100000",
  37059=>"001000001",
  37060=>"000000000",
  37061=>"011000000",
  37062=>"100000000",
  37063=>"011011111",
  37064=>"111101000",
  37065=>"111110111",
  37066=>"000000000",
  37067=>"000000000",
  37068=>"000010011",
  37069=>"000000010",
  37070=>"000000010",
  37071=>"000000000",
  37072=>"110111111",
  37073=>"111011111",
  37074=>"000111111",
  37075=>"011000000",
  37076=>"000000000",
  37077=>"111000000",
  37078=>"111110100",
  37079=>"000000111",
  37080=>"000000111",
  37081=>"111111111",
  37082=>"111000000",
  37083=>"110000110",
  37084=>"001011111",
  37085=>"000010111",
  37086=>"100011000",
  37087=>"111111111",
  37088=>"010000000",
  37089=>"001011111",
  37090=>"111111111",
  37091=>"110111110",
  37092=>"010000001",
  37093=>"000000000",
  37094=>"111111111",
  37095=>"111111111",
  37096=>"000111111",
  37097=>"111111111",
  37098=>"110111111",
  37099=>"111011111",
  37100=>"000000000",
  37101=>"111111111",
  37102=>"000110011",
  37103=>"111011000",
  37104=>"111111000",
  37105=>"111111111",
  37106=>"010111000",
  37107=>"101000100",
  37108=>"000000010",
  37109=>"101100100",
  37110=>"000100111",
  37111=>"111111111",
  37112=>"000000000",
  37113=>"000000011",
  37114=>"000111111",
  37115=>"000001111",
  37116=>"000111111",
  37117=>"111001000",
  37118=>"110110110",
  37119=>"000111111",
  37120=>"100000000",
  37121=>"111111011",
  37122=>"110111111",
  37123=>"001000001",
  37124=>"000111111",
  37125=>"000000011",
  37126=>"000001001",
  37127=>"000000111",
  37128=>"111111110",
  37129=>"010010000",
  37130=>"111011001",
  37131=>"011111111",
  37132=>"100000100",
  37133=>"111100000",
  37134=>"100000000",
  37135=>"000011000",
  37136=>"111111111",
  37137=>"001000000",
  37138=>"000000000",
  37139=>"000000010",
  37140=>"011011010",
  37141=>"000000000",
  37142=>"000011110",
  37143=>"101111011",
  37144=>"111001001",
  37145=>"000000000",
  37146=>"101001001",
  37147=>"001011000",
  37148=>"000000000",
  37149=>"000000000",
  37150=>"000000000",
  37151=>"101101111",
  37152=>"111100000",
  37153=>"111110000",
  37154=>"001111111",
  37155=>"001001111",
  37156=>"000000101",
  37157=>"000000000",
  37158=>"000100000",
  37159=>"011100000",
  37160=>"111101100",
  37161=>"110110000",
  37162=>"100111111",
  37163=>"111111111",
  37164=>"000101000",
  37165=>"101111001",
  37166=>"111000000",
  37167=>"000000111",
  37168=>"001101111",
  37169=>"000001101",
  37170=>"111000100",
  37171=>"111111111",
  37172=>"010010010",
  37173=>"111111101",
  37174=>"000000000",
  37175=>"111111110",
  37176=>"010110000",
  37177=>"111111000",
  37178=>"000000000",
  37179=>"000000000",
  37180=>"000000000",
  37181=>"000010111",
  37182=>"100100111",
  37183=>"111111111",
  37184=>"101000000",
  37185=>"111111111",
  37186=>"001001101",
  37187=>"111000000",
  37188=>"001000000",
  37189=>"000000000",
  37190=>"000000111",
  37191=>"100111111",
  37192=>"000000001",
  37193=>"110000000",
  37194=>"000111110",
  37195=>"111111111",
  37196=>"111111000",
  37197=>"111111111",
  37198=>"000000010",
  37199=>"111101111",
  37200=>"001001000",
  37201=>"000000111",
  37202=>"011001111",
  37203=>"000000111",
  37204=>"100111000",
  37205=>"000000001",
  37206=>"110111111",
  37207=>"101000011",
  37208=>"001001111",
  37209=>"010011000",
  37210=>"100000111",
  37211=>"111000011",
  37212=>"000000000",
  37213=>"000000111",
  37214=>"011111000",
  37215=>"001001101",
  37216=>"001011111",
  37217=>"111011111",
  37218=>"101101001",
  37219=>"000000000",
  37220=>"111111111",
  37221=>"111111101",
  37222=>"100110111",
  37223=>"111000000",
  37224=>"110111101",
  37225=>"000001001",
  37226=>"110110111",
  37227=>"111000000",
  37228=>"000111001",
  37229=>"000000000",
  37230=>"000011111",
  37231=>"000000000",
  37232=>"110001001",
  37233=>"111010011",
  37234=>"001011001",
  37235=>"001111111",
  37236=>"111010000",
  37237=>"101111000",
  37238=>"000111111",
  37239=>"100000110",
  37240=>"000000111",
  37241=>"111011000",
  37242=>"110011000",
  37243=>"111000100",
  37244=>"011011001",
  37245=>"111111111",
  37246=>"111111111",
  37247=>"101101001",
  37248=>"000000100",
  37249=>"001000000",
  37250=>"011011001",
  37251=>"000011001",
  37252=>"111110000",
  37253=>"010000000",
  37254=>"111111001",
  37255=>"001000000",
  37256=>"011111000",
  37257=>"010000111",
  37258=>"010000000",
  37259=>"000000010",
  37260=>"101111111",
  37261=>"110000000",
  37262=>"111111011",
  37263=>"111111111",
  37264=>"111111111",
  37265=>"110000000",
  37266=>"111111111",
  37267=>"001001111",
  37268=>"111111111",
  37269=>"111010000",
  37270=>"100111111",
  37271=>"001001101",
  37272=>"000000001",
  37273=>"111000000",
  37274=>"010111110",
  37275=>"001001101",
  37276=>"110110111",
  37277=>"111100000",
  37278=>"111111111",
  37279=>"111111000",
  37280=>"100000011",
  37281=>"101101000",
  37282=>"111111000",
  37283=>"000100111",
  37284=>"000000000",
  37285=>"111111111",
  37286=>"111001000",
  37287=>"111111111",
  37288=>"000000000",
  37289=>"110111111",
  37290=>"110111111",
  37291=>"111111111",
  37292=>"000100110",
  37293=>"001001111",
  37294=>"110111111",
  37295=>"000000000",
  37296=>"000000000",
  37297=>"010010011",
  37298=>"000101111",
  37299=>"000000000",
  37300=>"111001000",
  37301=>"000101110",
  37302=>"100100001",
  37303=>"111011100",
  37304=>"000000000",
  37305=>"110110111",
  37306=>"111111111",
  37307=>"001001111",
  37308=>"000000000",
  37309=>"100000111",
  37310=>"110000000",
  37311=>"001001011",
  37312=>"110110111",
  37313=>"000000000",
  37314=>"111011000",
  37315=>"111011000",
  37316=>"111110111",
  37317=>"111100100",
  37318=>"111000000",
  37319=>"101111111",
  37320=>"111100000",
  37321=>"001010110",
  37322=>"111111010",
  37323=>"000001001",
  37324=>"000000000",
  37325=>"010000111",
  37326=>"000000000",
  37327=>"111111000",
  37328=>"111011000",
  37329=>"111111100",
  37330=>"001101000",
  37331=>"100001111",
  37332=>"001001001",
  37333=>"111100000",
  37334=>"000110110",
  37335=>"000110010",
  37336=>"000000000",
  37337=>"111100000",
  37338=>"111111111",
  37339=>"000000110",
  37340=>"000000000",
  37341=>"000000000",
  37342=>"001000100",
  37343=>"000001011",
  37344=>"111111000",
  37345=>"011001010",
  37346=>"000001111",
  37347=>"001001001",
  37348=>"111111011",
  37349=>"000000000",
  37350=>"000000111",
  37351=>"110110111",
  37352=>"110000000",
  37353=>"111111000",
  37354=>"110111111",
  37355=>"000100100",
  37356=>"111111100",
  37357=>"101101111",
  37358=>"111110100",
  37359=>"111011001",
  37360=>"000000011",
  37361=>"000000000",
  37362=>"110110110",
  37363=>"110000000",
  37364=>"011001110",
  37365=>"000000000",
  37366=>"111011000",
  37367=>"001101001",
  37368=>"111001010",
  37369=>"011101111",
  37370=>"000111111",
  37371=>"010111001",
  37372=>"111111000",
  37373=>"111111001",
  37374=>"111111111",
  37375=>"111001111",
  37376=>"000111111",
  37377=>"000111111",
  37378=>"111111111",
  37379=>"000000000",
  37380=>"000001001",
  37381=>"100100111",
  37382=>"000000000",
  37383=>"001111111",
  37384=>"110000000",
  37385=>"111000000",
  37386=>"001001000",
  37387=>"000000000",
  37388=>"100100100",
  37389=>"001000000",
  37390=>"000000101",
  37391=>"000000001",
  37392=>"000000111",
  37393=>"110000000",
  37394=>"111111111",
  37395=>"000000000",
  37396=>"000000000",
  37397=>"101000011",
  37398=>"000000000",
  37399=>"011011111",
  37400=>"001001001",
  37401=>"100001001",
  37402=>"111000000",
  37403=>"101110100",
  37404=>"011001000",
  37405=>"110110100",
  37406=>"001011011",
  37407=>"000000001",
  37408=>"000000000",
  37409=>"000000000",
  37410=>"100100000",
  37411=>"000000000",
  37412=>"010110110",
  37413=>"111110000",
  37414=>"001000100",
  37415=>"000000000",
  37416=>"111111111",
  37417=>"000000000",
  37418=>"101111000",
  37419=>"111111111",
  37420=>"100000111",
  37421=>"000000000",
  37422=>"111111111",
  37423=>"000000000",
  37424=>"111111100",
  37425=>"000010001",
  37426=>"001001000",
  37427=>"111110111",
  37428=>"000000000",
  37429=>"100100100",
  37430=>"111111111",
  37431=>"100001101",
  37432=>"010000000",
  37433=>"000001001",
  37434=>"111111100",
  37435=>"000000010",
  37436=>"111111111",
  37437=>"111111110",
  37438=>"000000000",
  37439=>"101101111",
  37440=>"000000000",
  37441=>"110110011",
  37442=>"000111111",
  37443=>"110100000",
  37444=>"111100110",
  37445=>"111100100",
  37446=>"000000111",
  37447=>"000010011",
  37448=>"011011001",
  37449=>"001001001",
  37450=>"111111100",
  37451=>"000001111",
  37452=>"111111111",
  37453=>"111111111",
  37454=>"010010011",
  37455=>"000000000",
  37456=>"100000100",
  37457=>"111110110",
  37458=>"111011011",
  37459=>"101001011",
  37460=>"111101101",
  37461=>"000000000",
  37462=>"011011011",
  37463=>"111000000",
  37464=>"111111111",
  37465=>"111111111",
  37466=>"111111111",
  37467=>"010000100",
  37468=>"000010011",
  37469=>"111000111",
  37470=>"000100000",
  37471=>"000000000",
  37472=>"000000000",
  37473=>"000000000",
  37474=>"100100111",
  37475=>"111111111",
  37476=>"001001111",
  37477=>"000001001",
  37478=>"101000000",
  37479=>"011011111",
  37480=>"111111000",
  37481=>"111111111",
  37482=>"111001111",
  37483=>"111111001",
  37484=>"100100111",
  37485=>"000010000",
  37486=>"110100100",
  37487=>"000000000",
  37488=>"000001000",
  37489=>"000000000",
  37490=>"011011001",
  37491=>"000011001",
  37492=>"000000000",
  37493=>"000000100",
  37494=>"101000000",
  37495=>"000001111",
  37496=>"111111111",
  37497=>"000000111",
  37498=>"000000000",
  37499=>"111111111",
  37500=>"100100110",
  37501=>"111011111",
  37502=>"001001000",
  37503=>"000000000",
  37504=>"000000000",
  37505=>"111111000",
  37506=>"111000000",
  37507=>"111111111",
  37508=>"100110000",
  37509=>"111011111",
  37510=>"111001000",
  37511=>"000001111",
  37512=>"101111001",
  37513=>"000000000",
  37514=>"000000000",
  37515=>"000000000",
  37516=>"011100100",
  37517=>"000000111",
  37518=>"110110111",
  37519=>"001000000",
  37520=>"011011011",
  37521=>"111011011",
  37522=>"111111010",
  37523=>"000001011",
  37524=>"000010011",
  37525=>"110100110",
  37526=>"111111111",
  37527=>"111000000",
  37528=>"110000100",
  37529=>"110010011",
  37530=>"111111100",
  37531=>"000000000",
  37532=>"000000000",
  37533=>"000000000",
  37534=>"000000000",
  37535=>"000000110",
  37536=>"000000000",
  37537=>"110110110",
  37538=>"000110111",
  37539=>"111011101",
  37540=>"000000000",
  37541=>"000000000",
  37542=>"111111111",
  37543=>"000111011",
  37544=>"111111001",
  37545=>"000000000",
  37546=>"000000101",
  37547=>"000000000",
  37548=>"000000000",
  37549=>"111101101",
  37550=>"000000001",
  37551=>"111111000",
  37552=>"000011000",
  37553=>"111101101",
  37554=>"111111111",
  37555=>"111100000",
  37556=>"000100111",
  37557=>"000100000",
  37558=>"111111111",
  37559=>"111110000",
  37560=>"111111111",
  37561=>"111001111",
  37562=>"001001000",
  37563=>"000000000",
  37564=>"111111111",
  37565=>"000100100",
  37566=>"011111000",
  37567=>"000001001",
  37568=>"111111111",
  37569=>"000000000",
  37570=>"111111001",
  37571=>"111111111",
  37572=>"000000000",
  37573=>"000000000",
  37574=>"000000000",
  37575=>"010100110",
  37576=>"000000011",
  37577=>"000000111",
  37578=>"110110100",
  37579=>"011010000",
  37580=>"111110111",
  37581=>"111111111",
  37582=>"111000110",
  37583=>"000000000",
  37584=>"101111111",
  37585=>"001001000",
  37586=>"111110111",
  37587=>"111111111",
  37588=>"100100100",
  37589=>"100111111",
  37590=>"000000000",
  37591=>"111111111",
  37592=>"111110110",
  37593=>"011111111",
  37594=>"111111000",
  37595=>"111111111",
  37596=>"000000111",
  37597=>"010011000",
  37598=>"111010001",
  37599=>"000000001",
  37600=>"000000000",
  37601=>"000000011",
  37602=>"000111110",
  37603=>"111111111",
  37604=>"000000000",
  37605=>"100000100",
  37606=>"111000000",
  37607=>"001000111",
  37608=>"111111111",
  37609=>"001001101",
  37610=>"111000000",
  37611=>"111110111",
  37612=>"000000000",
  37613=>"100100000",
  37614=>"000111111",
  37615=>"000011111",
  37616=>"001000000",
  37617=>"110110110",
  37618=>"111111111",
  37619=>"001000111",
  37620=>"000000000",
  37621=>"100000000",
  37622=>"011010110",
  37623=>"110111111",
  37624=>"000000000",
  37625=>"111111111",
  37626=>"111111000",
  37627=>"111111111",
  37628=>"111111111",
  37629=>"100110110",
  37630=>"011000000",
  37631=>"110110110",
  37632=>"111110000",
  37633=>"111101000",
  37634=>"111011010",
  37635=>"100100000",
  37636=>"111111110",
  37637=>"000000000",
  37638=>"000110100",
  37639=>"111111000",
  37640=>"010000000",
  37641=>"011001001",
  37642=>"111111111",
  37643=>"011111100",
  37644=>"110000110",
  37645=>"111000000",
  37646=>"111010111",
  37647=>"111111110",
  37648=>"011111001",
  37649=>"111101101",
  37650=>"110111111",
  37651=>"110110001",
  37652=>"111001001",
  37653=>"101001111",
  37654=>"000000001",
  37655=>"111110100",
  37656=>"111111110",
  37657=>"000111111",
  37658=>"000000000",
  37659=>"111010110",
  37660=>"110110110",
  37661=>"000000000",
  37662=>"111010000",
  37663=>"000000001",
  37664=>"110100100",
  37665=>"111000000",
  37666=>"010111111",
  37667=>"000000000",
  37668=>"011011001",
  37669=>"001001001",
  37670=>"000001111",
  37671=>"110111000",
  37672=>"000000000",
  37673=>"000000000",
  37674=>"111111101",
  37675=>"001001111",
  37676=>"000000111",
  37677=>"111110000",
  37678=>"000100001",
  37679=>"000000110",
  37680=>"000001001",
  37681=>"111111111",
  37682=>"111111111",
  37683=>"011000111",
  37684=>"111100000",
  37685=>"000000000",
  37686=>"011111111",
  37687=>"000000000",
  37688=>"000000000",
  37689=>"111111111",
  37690=>"011001000",
  37691=>"000000000",
  37692=>"000000111",
  37693=>"100100110",
  37694=>"000111111",
  37695=>"001011111",
  37696=>"000000000",
  37697=>"111111111",
  37698=>"111111111",
  37699=>"111011001",
  37700=>"011000000",
  37701=>"000100111",
  37702=>"000000101",
  37703=>"101100100",
  37704=>"111110110",
  37705=>"000000000",
  37706=>"111111111",
  37707=>"111111111",
  37708=>"001101111",
  37709=>"000000000",
  37710=>"111001100",
  37711=>"110111110",
  37712=>"000100100",
  37713=>"111111111",
  37714=>"000000100",
  37715=>"111111110",
  37716=>"000000000",
  37717=>"001000001",
  37718=>"011011111",
  37719=>"111111111",
  37720=>"111111100",
  37721=>"101000001",
  37722=>"111111000",
  37723=>"000111111",
  37724=>"000000000",
  37725=>"000000000",
  37726=>"111111111",
  37727=>"111111111",
  37728=>"111011011",
  37729=>"111111111",
  37730=>"000000000",
  37731=>"000111011",
  37732=>"100000100",
  37733=>"111111111",
  37734=>"000000000",
  37735=>"100000000",
  37736=>"110010000",
  37737=>"110111110",
  37738=>"111111101",
  37739=>"000111111",
  37740=>"001000000",
  37741=>"000000111",
  37742=>"000011000",
  37743=>"111111111",
  37744=>"000000100",
  37745=>"000110010",
  37746=>"100000000",
  37747=>"000000001",
  37748=>"111110111",
  37749=>"111111111",
  37750=>"000110111",
  37751=>"000000001",
  37752=>"100000000",
  37753=>"000000000",
  37754=>"000000000",
  37755=>"000000000",
  37756=>"000001001",
  37757=>"011000111",
  37758=>"111111110",
  37759=>"000000000",
  37760=>"111111111",
  37761=>"111100110",
  37762=>"111100100",
  37763=>"000011000",
  37764=>"000000000",
  37765=>"011011011",
  37766=>"111111011",
  37767=>"111111111",
  37768=>"110111001",
  37769=>"000001101",
  37770=>"100100100",
  37771=>"111011000",
  37772=>"111000000",
  37773=>"011101001",
  37774=>"111111111",
  37775=>"111111001",
  37776=>"000000110",
  37777=>"000001111",
  37778=>"110111111",
  37779=>"001111111",
  37780=>"111111111",
  37781=>"000001000",
  37782=>"110111111",
  37783=>"100111111",
  37784=>"000000100",
  37785=>"000000000",
  37786=>"111110000",
  37787=>"000000001",
  37788=>"000000000",
  37789=>"111111011",
  37790=>"000000000",
  37791=>"111111111",
  37792=>"111111111",
  37793=>"001001000",
  37794=>"010000000",
  37795=>"000000111",
  37796=>"000000000",
  37797=>"000000000",
  37798=>"111001111",
  37799=>"000000000",
  37800=>"110110000",
  37801=>"110010001",
  37802=>"000000000",
  37803=>"000101111",
  37804=>"111111111",
  37805=>"000000000",
  37806=>"000001000",
  37807=>"111111110",
  37808=>"111111111",
  37809=>"111111110",
  37810=>"111111111",
  37811=>"111111100",
  37812=>"000001011",
  37813=>"111001000",
  37814=>"110111110",
  37815=>"111011111",
  37816=>"110100000",
  37817=>"000010000",
  37818=>"001101111",
  37819=>"111111101",
  37820=>"000000000",
  37821=>"111111111",
  37822=>"011111111",
  37823=>"111110100",
  37824=>"000000100",
  37825=>"000000000",
  37826=>"000000001",
  37827=>"111111000",
  37828=>"111011000",
  37829=>"111110000",
  37830=>"000000000",
  37831=>"000111111",
  37832=>"000000000",
  37833=>"000001111",
  37834=>"111000000",
  37835=>"111111000",
  37836=>"111111111",
  37837=>"000000000",
  37838=>"010010000",
  37839=>"000000110",
  37840=>"010010010",
  37841=>"111100111",
  37842=>"000000000",
  37843=>"111111000",
  37844=>"111101111",
  37845=>"111111000",
  37846=>"100100111",
  37847=>"001011011",
  37848=>"000000000",
  37849=>"000000000",
  37850=>"111111000",
  37851=>"011111001",
  37852=>"000000010",
  37853=>"000111111",
  37854=>"111111110",
  37855=>"011001001",
  37856=>"111111111",
  37857=>"001001000",
  37858=>"001111111",
  37859=>"111111111",
  37860=>"111111111",
  37861=>"111000000",
  37862=>"000000000",
  37863=>"100000110",
  37864=>"111111111",
  37865=>"000111111",
  37866=>"111111111",
  37867=>"111011111",
  37868=>"111111111",
  37869=>"000000100",
  37870=>"000001011",
  37871=>"100000000",
  37872=>"000000000",
  37873=>"111110111",
  37874=>"000000001",
  37875=>"010111111",
  37876=>"000000000",
  37877=>"111111111",
  37878=>"101111111",
  37879=>"100100000",
  37880=>"000000000",
  37881=>"000000000",
  37882=>"111110111",
  37883=>"111110110",
  37884=>"111111111",
  37885=>"011000100",
  37886=>"111111111",
  37887=>"000100100",
  37888=>"010110111",
  37889=>"000010010",
  37890=>"111111000",
  37891=>"111101001",
  37892=>"000000110",
  37893=>"110110111",
  37894=>"011001001",
  37895=>"111111111",
  37896=>"001001011",
  37897=>"000000100",
  37898=>"000111111",
  37899=>"111111111",
  37900=>"000000000",
  37901=>"111000000",
  37902=>"111111110",
  37903=>"110111111",
  37904=>"001000000",
  37905=>"000111111",
  37906=>"111111011",
  37907=>"000000101",
  37908=>"010000000",
  37909=>"111111111",
  37910=>"011111000",
  37911=>"111110110",
  37912=>"000000100",
  37913=>"111111111",
  37914=>"000000100",
  37915=>"000010001",
  37916=>"110111111",
  37917=>"000101101",
  37918=>"000001001",
  37919=>"111101000",
  37920=>"000000000",
  37921=>"000110111",
  37922=>"100100000",
  37923=>"100000000",
  37924=>"000000000",
  37925=>"111111111",
  37926=>"000000000",
  37927=>"111111111",
  37928=>"000000000",
  37929=>"111000000",
  37930=>"111110010",
  37931=>"111100111",
  37932=>"100000000",
  37933=>"000101000",
  37934=>"100100100",
  37935=>"001000000",
  37936=>"000000000",
  37937=>"000000001",
  37938=>"000010000",
  37939=>"110010101",
  37940=>"000000000",
  37941=>"110111110",
  37942=>"111111111",
  37943=>"100100100",
  37944=>"111111111",
  37945=>"000000000",
  37946=>"111000000",
  37947=>"111111111",
  37948=>"000000000",
  37949=>"011011111",
  37950=>"111111111",
  37951=>"011000111",
  37952=>"101111111",
  37953=>"000000000",
  37954=>"111111111",
  37955=>"111111111",
  37956=>"000000001",
  37957=>"111111010",
  37958=>"001001111",
  37959=>"000000000",
  37960=>"001000000",
  37961=>"001001001",
  37962=>"001111111",
  37963=>"111100000",
  37964=>"000000000",
  37965=>"000000000",
  37966=>"000000001",
  37967=>"111111111",
  37968=>"111010010",
  37969=>"111111101",
  37970=>"000000000",
  37971=>"100100110",
  37972=>"000111111",
  37973=>"001011011",
  37974=>"111001001",
  37975=>"110110000",
  37976=>"000000000",
  37977=>"111000101",
  37978=>"111111101",
  37979=>"000000100",
  37980=>"000111111",
  37981=>"000111111",
  37982=>"111111111",
  37983=>"111111111",
  37984=>"001001000",
  37985=>"001000000",
  37986=>"111111111",
  37987=>"000001000",
  37988=>"000000100",
  37989=>"111111111",
  37990=>"111111111",
  37991=>"000010111",
  37992=>"111111111",
  37993=>"111111111",
  37994=>"111101111",
  37995=>"111101111",
  37996=>"111111111",
  37997=>"000000000",
  37998=>"111111111",
  37999=>"000000000",
  38000=>"111111011",
  38001=>"000001000",
  38002=>"000000000",
  38003=>"000001111",
  38004=>"011011011",
  38005=>"100100111",
  38006=>"111111111",
  38007=>"110110100",
  38008=>"000000000",
  38009=>"000110110",
  38010=>"111111000",
  38011=>"000000000",
  38012=>"100100100",
  38013=>"111110110",
  38014=>"000000000",
  38015=>"110000000",
  38016=>"111001011",
  38017=>"101100111",
  38018=>"111111111",
  38019=>"000000000",
  38020=>"111000111",
  38021=>"111100000",
  38022=>"111011111",
  38023=>"111111110",
  38024=>"001111111",
  38025=>"111100101",
  38026=>"000000000",
  38027=>"000011111",
  38028=>"011111111",
  38029=>"000000001",
  38030=>"111111111",
  38031=>"000000000",
  38032=>"000000000",
  38033=>"110111111",
  38034=>"111111111",
  38035=>"111110110",
  38036=>"000110111",
  38037=>"000110111",
  38038=>"111001000",
  38039=>"111011000",
  38040=>"100000000",
  38041=>"111100110",
  38042=>"000110010",
  38043=>"000111010",
  38044=>"111111111",
  38045=>"000101111",
  38046=>"101100111",
  38047=>"111111111",
  38048=>"111111000",
  38049=>"111111111",
  38050=>"111111111",
  38051=>"000000110",
  38052=>"000000000",
  38053=>"000000000",
  38054=>"000111111",
  38055=>"011011010",
  38056=>"000000111",
  38057=>"000000001",
  38058=>"101000000",
  38059=>"110111111",
  38060=>"111111001",
  38061=>"111110010",
  38062=>"000000111",
  38063=>"111111111",
  38064=>"000010111",
  38065=>"111111111",
  38066=>"110111111",
  38067=>"111111100",
  38068=>"000110111",
  38069=>"111001001",
  38070=>"000111111",
  38071=>"001101100",
  38072=>"000000000",
  38073=>"000000000",
  38074=>"010110100",
  38075=>"101111111",
  38076=>"100000000",
  38077=>"100000000",
  38078=>"111111111",
  38079=>"000111111",
  38080=>"000000010",
  38081=>"000000000",
  38082=>"000000000",
  38083=>"000010111",
  38084=>"001111010",
  38085=>"000000000",
  38086=>"000000000",
  38087=>"000000111",
  38088=>"111000000",
  38089=>"000000100",
  38090=>"000000000",
  38091=>"000000000",
  38092=>"101100101",
  38093=>"000000000",
  38094=>"111111111",
  38095=>"111000110",
  38096=>"110110000",
  38097=>"000000000",
  38098=>"000111111",
  38099=>"001000000",
  38100=>"100100000",
  38101=>"111000101",
  38102=>"000000001",
  38103=>"010010000",
  38104=>"000000001",
  38105=>"000100101",
  38106=>"100000000",
  38107=>"111001001",
  38108=>"111111111",
  38109=>"100000000",
  38110=>"000010000",
  38111=>"111100111",
  38112=>"111010000",
  38113=>"000000111",
  38114=>"100100111",
  38115=>"111000000",
  38116=>"110110110",
  38117=>"000000111",
  38118=>"100100100",
  38119=>"111001111",
  38120=>"001111000",
  38121=>"100100001",
  38122=>"111111111",
  38123=>"101001101",
  38124=>"000000000",
  38125=>"000101111",
  38126=>"000000101",
  38127=>"000000000",
  38128=>"100101111",
  38129=>"011001000",
  38130=>"111001101",
  38131=>"011111111",
  38132=>"111111111",
  38133=>"101111111",
  38134=>"000000000",
  38135=>"111101000",
  38136=>"001000000",
  38137=>"001100010",
  38138=>"111010000",
  38139=>"000011000",
  38140=>"000000000",
  38141=>"111110111",
  38142=>"000000000",
  38143=>"100100100",
  38144=>"000000000",
  38145=>"001001111",
  38146=>"111111000",
  38147=>"000000000",
  38148=>"000000111",
  38149=>"000000000",
  38150=>"111111111",
  38151=>"001111000",
  38152=>"000000000",
  38153=>"111100000",
  38154=>"111111111",
  38155=>"110001111",
  38156=>"111101000",
  38157=>"111110110",
  38158=>"011011111",
  38159=>"000111111",
  38160=>"000000000",
  38161=>"010011111",
  38162=>"111111111",
  38163=>"000000100",
  38164=>"000000000",
  38165=>"100010000",
  38166=>"100100100",
  38167=>"100100100",
  38168=>"000000110",
  38169=>"111010111",
  38170=>"101111101",
  38171=>"000111111",
  38172=>"001011011",
  38173=>"000001111",
  38174=>"010111010",
  38175=>"111111111",
  38176=>"000110100",
  38177=>"111000100",
  38178=>"111011111",
  38179=>"111111011",
  38180=>"111111111",
  38181=>"000000000",
  38182=>"000010010",
  38183=>"010000000",
  38184=>"111111111",
  38185=>"111001111",
  38186=>"000000000",
  38187=>"000000000",
  38188=>"111111111",
  38189=>"000010000",
  38190=>"000000000",
  38191=>"101000000",
  38192=>"110110111",
  38193=>"000100111",
  38194=>"111110111",
  38195=>"111111111",
  38196=>"111111111",
  38197=>"000000011",
  38198=>"000000000",
  38199=>"000000000",
  38200=>"000000000",
  38201=>"100100100",
  38202=>"011101111",
  38203=>"101100111",
  38204=>"000000000",
  38205=>"000000111",
  38206=>"000000110",
  38207=>"111111100",
  38208=>"000000000",
  38209=>"000000110",
  38210=>"110111111",
  38211=>"100000000",
  38212=>"001001001",
  38213=>"000100101",
  38214=>"000000111",
  38215=>"000000001",
  38216=>"000111111",
  38217=>"111000000",
  38218=>"000111111",
  38219=>"101101001",
  38220=>"011111111",
  38221=>"111111111",
  38222=>"000000001",
  38223=>"000000110",
  38224=>"000000000",
  38225=>"000000000",
  38226=>"000000000",
  38227=>"111000000",
  38228=>"000000000",
  38229=>"011001001",
  38230=>"000000000",
  38231=>"011111111",
  38232=>"100111001",
  38233=>"001000000",
  38234=>"001001000",
  38235=>"111111111",
  38236=>"001000000",
  38237=>"010000000",
  38238=>"110101000",
  38239=>"000000000",
  38240=>"000000000",
  38241=>"000111111",
  38242=>"000000110",
  38243=>"101101100",
  38244=>"000000001",
  38245=>"000000000",
  38246=>"101100110",
  38247=>"100000010",
  38248=>"111001001",
  38249=>"111111111",
  38250=>"000000000",
  38251=>"001001111",
  38252=>"110110010",
  38253=>"111110100",
  38254=>"100100101",
  38255=>"000000000",
  38256=>"000000010",
  38257=>"000100000",
  38258=>"111111000",
  38259=>"000001001",
  38260=>"111111101",
  38261=>"111111111",
  38262=>"000000000",
  38263=>"000001000",
  38264=>"000000000",
  38265=>"110111111",
  38266=>"111111111",
  38267=>"100000001",
  38268=>"111111111",
  38269=>"111100110",
  38270=>"000000000",
  38271=>"000000000",
  38272=>"001111111",
  38273=>"000000000",
  38274=>"110111111",
  38275=>"000000111",
  38276=>"010000000",
  38277=>"010011011",
  38278=>"110111111",
  38279=>"000000000",
  38280=>"100101000",
  38281=>"110111110",
  38282=>"000000111",
  38283=>"000000000",
  38284=>"111111111",
  38285=>"100100111",
  38286=>"111001011",
  38287=>"111001001",
  38288=>"000011010",
  38289=>"111011111",
  38290=>"110110100",
  38291=>"000000100",
  38292=>"111001000",
  38293=>"000000000",
  38294=>"000000000",
  38295=>"111111111",
  38296=>"010110100",
  38297=>"100000001",
  38298=>"111111100",
  38299=>"111000000",
  38300=>"101101000",
  38301=>"011111010",
  38302=>"000111000",
  38303=>"111111000",
  38304=>"010000000",
  38305=>"000000000",
  38306=>"111101001",
  38307=>"011000000",
  38308=>"111100000",
  38309=>"000000000",
  38310=>"000000000",
  38311=>"000101000",
  38312=>"001000000",
  38313=>"100111111",
  38314=>"111111111",
  38315=>"111100101",
  38316=>"000000000",
  38317=>"000000000",
  38318=>"111110111",
  38319=>"011000111",
  38320=>"111111000",
  38321=>"111110000",
  38322=>"000110111",
  38323=>"111111111",
  38324=>"100110111",
  38325=>"000000000",
  38326=>"000000000",
  38327=>"111111111",
  38328=>"111111000",
  38329=>"111111111",
  38330=>"000110111",
  38331=>"000000000",
  38332=>"111111111",
  38333=>"111111111",
  38334=>"000001000",
  38335=>"100110100",
  38336=>"000000000",
  38337=>"000101000",
  38338=>"111111111",
  38339=>"001111111",
  38340=>"011001001",
  38341=>"000000000",
  38342=>"000000011",
  38343=>"000100111",
  38344=>"000000000",
  38345=>"000000000",
  38346=>"111001000",
  38347=>"011111100",
  38348=>"000000111",
  38349=>"100100111",
  38350=>"111111111",
  38351=>"111111111",
  38352=>"000000000",
  38353=>"000111111",
  38354=>"000000000",
  38355=>"000100100",
  38356=>"100100100",
  38357=>"001001111",
  38358=>"000101111",
  38359=>"000000000",
  38360=>"111111111",
  38361=>"010100100",
  38362=>"100100110",
  38363=>"001001111",
  38364=>"111111111",
  38365=>"001001011",
  38366=>"001000100",
  38367=>"100100001",
  38368=>"000000000",
  38369=>"111111111",
  38370=>"111000000",
  38371=>"000111111",
  38372=>"111111111",
  38373=>"000000000",
  38374=>"000000001",
  38375=>"111000000",
  38376=>"110110010",
  38377=>"000101111",
  38378=>"000000000",
  38379=>"110010011",
  38380=>"111111000",
  38381=>"111111111",
  38382=>"000000000",
  38383=>"001000000",
  38384=>"111101000",
  38385=>"111100000",
  38386=>"110000111",
  38387=>"001001100",
  38388=>"000001001",
  38389=>"100000000",
  38390=>"111100111",
  38391=>"110000100",
  38392=>"000000000",
  38393=>"011001001",
  38394=>"000000000",
  38395=>"101111111",
  38396=>"100111101",
  38397=>"000000000",
  38398=>"100100100",
  38399=>"111111111",
  38400=>"100110111",
  38401=>"001000000",
  38402=>"100000111",
  38403=>"101000000",
  38404=>"111110111",
  38405=>"111111111",
  38406=>"000000101",
  38407=>"111111111",
  38408=>"101111010",
  38409=>"111111111",
  38410=>"000111111",
  38411=>"001001000",
  38412=>"111111111",
  38413=>"011111101",
  38414=>"010110000",
  38415=>"001000001",
  38416=>"001000000",
  38417=>"000000111",
  38418=>"000110111",
  38419=>"000000000",
  38420=>"000000000",
  38421=>"010000000",
  38422=>"100111110",
  38423=>"001011011",
  38424=>"110111101",
  38425=>"001011111",
  38426=>"111111000",
  38427=>"000110111",
  38428=>"111111111",
  38429=>"000000000",
  38430=>"000100000",
  38431=>"110110110",
  38432=>"000000001",
  38433=>"010000000",
  38434=>"111111111",
  38435=>"111011111",
  38436=>"111011011",
  38437=>"000000100",
  38438=>"001001001",
  38439=>"000000011",
  38440=>"111111001",
  38441=>"000011011",
  38442=>"011111111",
  38443=>"111111110",
  38444=>"111110010",
  38445=>"101001000",
  38446=>"101100000",
  38447=>"111111000",
  38448=>"111000001",
  38449=>"000001000",
  38450=>"011010000",
  38451=>"111000000",
  38452=>"110111101",
  38453=>"010000000",
  38454=>"101000101",
  38455=>"000000000",
  38456=>"111001111",
  38457=>"111111111",
  38458=>"111111111",
  38459=>"000111111",
  38460=>"111111111",
  38461=>"000000100",
  38462=>"111110000",
  38463=>"101100000",
  38464=>"011110111",
  38465=>"011001111",
  38466=>"000110010",
  38467=>"110010010",
  38468=>"000000110",
  38469=>"111111011",
  38470=>"000000111",
  38471=>"000000000",
  38472=>"011111111",
  38473=>"111111111",
  38474=>"000111111",
  38475=>"100010111",
  38476=>"111111111",
  38477=>"111000000",
  38478=>"010000000",
  38479=>"101111000",
  38480=>"011111000",
  38481=>"001001111",
  38482=>"000000001",
  38483=>"011011011",
  38484=>"000000000",
  38485=>"111100000",
  38486=>"111101111",
  38487=>"110111110",
  38488=>"111000100",
  38489=>"100111111",
  38490=>"111111011",
  38491=>"000011111",
  38492=>"011000000",
  38493=>"011000000",
  38494=>"000000100",
  38495=>"111111000",
  38496=>"111111111",
  38497=>"111111110",
  38498=>"101101000",
  38499=>"000000011",
  38500=>"111111000",
  38501=>"000000000",
  38502=>"111101000",
  38503=>"000000000",
  38504=>"100111111",
  38505=>"111111111",
  38506=>"000000101",
  38507=>"000000000",
  38508=>"111011111",
  38509=>"011011000",
  38510=>"111111110",
  38511=>"111111110",
  38512=>"011000000",
  38513=>"101101001",
  38514=>"000000101",
  38515=>"000000000",
  38516=>"010011111",
  38517=>"111000000",
  38518=>"010000000",
  38519=>"011111110",
  38520=>"000111111",
  38521=>"111111101",
  38522=>"000000000",
  38523=>"000000000",
  38524=>"110110000",
  38525=>"000000000",
  38526=>"000000000",
  38527=>"011001101",
  38528=>"000000000",
  38529=>"100100100",
  38530=>"000000000",
  38531=>"011111111",
  38532=>"011011001",
  38533=>"000000000",
  38534=>"111110000",
  38535=>"001001111",
  38536=>"001000001",
  38537=>"011000100",
  38538=>"111111000",
  38539=>"111111011",
  38540=>"001101111",
  38541=>"011011000",
  38542=>"011101000",
  38543=>"111110111",
  38544=>"111111011",
  38545=>"000000000",
  38546=>"111111111",
  38547=>"000000000",
  38548=>"100111111",
  38549=>"111111111",
  38550=>"100111111",
  38551=>"101000000",
  38552=>"111000000",
  38553=>"101100110",
  38554=>"000000111",
  38555=>"001001001",
  38556=>"110100000",
  38557=>"111000110",
  38558=>"111111000",
  38559=>"000000000",
  38560=>"111111111",
  38561=>"001001001",
  38562=>"101001011",
  38563=>"010000000",
  38564=>"000000000",
  38565=>"001011110",
  38566=>"111111111",
  38567=>"000110011",
  38568=>"000000000",
  38569=>"000000000",
  38570=>"000000000",
  38571=>"111010000",
  38572=>"011010000",
  38573=>"110110110",
  38574=>"100000010",
  38575=>"000001100",
  38576=>"000000101",
  38577=>"000000001",
  38578=>"011111011",
  38579=>"000001000",
  38580=>"111000000",
  38581=>"000111100",
  38582=>"000000000",
  38583=>"000011001",
  38584=>"100100110",
  38585=>"111111111",
  38586=>"000000111",
  38587=>"111111010",
  38588=>"011010011",
  38589=>"110110111",
  38590=>"110111111",
  38591=>"011011011",
  38592=>"000000000",
  38593=>"000010011",
  38594=>"000000000",
  38595=>"111111001",
  38596=>"111111111",
  38597=>"001000111",
  38598=>"111110100",
  38599=>"111000000",
  38600=>"000000100",
  38601=>"100111111",
  38602=>"110000000",
  38603=>"000000110",
  38604=>"001111111",
  38605=>"001011111",
  38606=>"111111000",
  38607=>"000111111",
  38608=>"000010010",
  38609=>"111111111",
  38610=>"000111111",
  38611=>"000000000",
  38612=>"000000000",
  38613=>"000000000",
  38614=>"111111000",
  38615=>"000000000",
  38616=>"000110111",
  38617=>"000000011",
  38618=>"010011111",
  38619=>"011111111",
  38620=>"000101100",
  38621=>"111001001",
  38622=>"011011111",
  38623=>"100100000",
  38624=>"011011111",
  38625=>"111111111",
  38626=>"111000000",
  38627=>"111111110",
  38628=>"111111110",
  38629=>"000010111",
  38630=>"100100010",
  38631=>"000000000",
  38632=>"111111000",
  38633=>"110100000",
  38634=>"001111101",
  38635=>"111111111",
  38636=>"001000000",
  38637=>"000000000",
  38638=>"110111111",
  38639=>"101001011",
  38640=>"000111111",
  38641=>"011111111",
  38642=>"111110011",
  38643=>"110111111",
  38644=>"001010000",
  38645=>"111111111",
  38646=>"100000010",
  38647=>"100000001",
  38648=>"001111111",
  38649=>"001001000",
  38650=>"111111111",
  38651=>"110000000",
  38652=>"011011110",
  38653=>"110010000",
  38654=>"000000001",
  38655=>"000011111",
  38656=>"110000000",
  38657=>"111111001",
  38658=>"111111111",
  38659=>"000100100",
  38660=>"000000001",
  38661=>"000000000",
  38662=>"111110000",
  38663=>"010000110",
  38664=>"001111111",
  38665=>"000000000",
  38666=>"000111111",
  38667=>"111100110",
  38668=>"001001001",
  38669=>"000000010",
  38670=>"111111111",
  38671=>"111111111",
  38672=>"111111000",
  38673=>"000100110",
  38674=>"111111000",
  38675=>"000000000",
  38676=>"110000111",
  38677=>"111000011",
  38678=>"000111001",
  38679=>"111000101",
  38680=>"100001001",
  38681=>"111111000",
  38682=>"000001000",
  38683=>"000000011",
  38684=>"000100110",
  38685=>"111011000",
  38686=>"110101111",
  38687=>"111111111",
  38688=>"000100000",
  38689=>"000001111",
  38690=>"111111111",
  38691=>"111111110",
  38692=>"000000000",
  38693=>"110011001",
  38694=>"101001000",
  38695=>"111111111",
  38696=>"111111111",
  38697=>"000000111",
  38698=>"111000100",
  38699=>"000101111",
  38700=>"000000000",
  38701=>"110010000",
  38702=>"101011011",
  38703=>"000000000",
  38704=>"000000000",
  38705=>"000011000",
  38706=>"000101110",
  38707=>"011100000",
  38708=>"111001000",
  38709=>"100100100",
  38710=>"111111110",
  38711=>"000000000",
  38712=>"111111111",
  38713=>"000000000",
  38714=>"000101001",
  38715=>"101001111",
  38716=>"110110100",
  38717=>"111111000",
  38718=>"111111001",
  38719=>"000000000",
  38720=>"111111111",
  38721=>"111001010",
  38722=>"011011001",
  38723=>"101101000",
  38724=>"000100111",
  38725=>"011000111",
  38726=>"000000000",
  38727=>"111111000",
  38728=>"001001000",
  38729=>"000111111",
  38730=>"000110100",
  38731=>"001001001",
  38732=>"110111000",
  38733=>"101111111",
  38734=>"000000000",
  38735=>"000001011",
  38736=>"011110000",
  38737=>"000000011",
  38738=>"000001111",
  38739=>"000010111",
  38740=>"000000000",
  38741=>"001001001",
  38742=>"010110111",
  38743=>"100100000",
  38744=>"110000000",
  38745=>"000110000",
  38746=>"111110000",
  38747=>"000101111",
  38748=>"000000101",
  38749=>"111111111",
  38750=>"011111101",
  38751=>"000000000",
  38752=>"000001000",
  38753=>"111000000",
  38754=>"001001000",
  38755=>"111111000",
  38756=>"111110110",
  38757=>"111100100",
  38758=>"111000000",
  38759=>"111111111",
  38760=>"000100100",
  38761=>"000000000",
  38762=>"000000010",
  38763=>"111110110",
  38764=>"000111111",
  38765=>"000000000",
  38766=>"000000000",
  38767=>"000000111",
  38768=>"111111000",
  38769=>"111100000",
  38770=>"000000011",
  38771=>"101001000",
  38772=>"000011111",
  38773=>"100000000",
  38774=>"000000010",
  38775=>"000000011",
  38776=>"000000000",
  38777=>"011011111",
  38778=>"110000000",
  38779=>"000000000",
  38780=>"000111111",
  38781=>"111110110",
  38782=>"111111111",
  38783=>"111111111",
  38784=>"100010110",
  38785=>"111110110",
  38786=>"110111010",
  38787=>"011111111",
  38788=>"001011011",
  38789=>"110000000",
  38790=>"000000110",
  38791=>"000000000",
  38792=>"000000000",
  38793=>"000000000",
  38794=>"111111111",
  38795=>"111001000",
  38796=>"111111111",
  38797=>"100100000",
  38798=>"101001111",
  38799=>"000000010",
  38800=>"000000011",
  38801=>"111111110",
  38802=>"111000000",
  38803=>"000001001",
  38804=>"000001111",
  38805=>"000000000",
  38806=>"111111111",
  38807=>"011000010",
  38808=>"100100100",
  38809=>"111110000",
  38810=>"100000100",
  38811=>"111100111",
  38812=>"000000111",
  38813=>"000000000",
  38814=>"111000100",
  38815=>"000001101",
  38816=>"000000000",
  38817=>"111111111",
  38818=>"101100100",
  38819=>"000000000",
  38820=>"111111000",
  38821=>"111111111",
  38822=>"000001001",
  38823=>"010010000",
  38824=>"000101101",
  38825=>"100111110",
  38826=>"000000000",
  38827=>"111000101",
  38828=>"011011000",
  38829=>"111110010",
  38830=>"000000001",
  38831=>"000011111",
  38832=>"111111000",
  38833=>"111111111",
  38834=>"111111011",
  38835=>"110000000",
  38836=>"011111011",
  38837=>"010111111",
  38838=>"100110010",
  38839=>"111111010",
  38840=>"000101111",
  38841=>"011011111",
  38842=>"111111000",
  38843=>"111011000",
  38844=>"000000001",
  38845=>"111001001",
  38846=>"101000000",
  38847=>"110111111",
  38848=>"100101100",
  38849=>"000111110",
  38850=>"111111111",
  38851=>"000111010",
  38852=>"110110110",
  38853=>"000000100",
  38854=>"111000111",
  38855=>"000000000",
  38856=>"110000000",
  38857=>"101111011",
  38858=>"000001100",
  38859=>"000001000",
  38860=>"000000000",
  38861=>"101000000",
  38862=>"111100110",
  38863=>"000000000",
  38864=>"000000010",
  38865=>"111111111",
  38866=>"000000000",
  38867=>"001000000",
  38868=>"000111111",
  38869=>"111111111",
  38870=>"111111000",
  38871=>"110100011",
  38872=>"101000000",
  38873=>"110111010",
  38874=>"000000111",
  38875=>"001111111",
  38876=>"000000000",
  38877=>"111111111",
  38878=>"000001111",
  38879=>"100100111",
  38880=>"011011111",
  38881=>"000000100",
  38882=>"111000111",
  38883=>"111111111",
  38884=>"101110000",
  38885=>"101111111",
  38886=>"000001111",
  38887=>"010000000",
  38888=>"011110111",
  38889=>"111011011",
  38890=>"000001000",
  38891=>"001000101",
  38892=>"001000111",
  38893=>"011011011",
  38894=>"111000001",
  38895=>"111111111",
  38896=>"100111010",
  38897=>"001111111",
  38898=>"000011001",
  38899=>"000000111",
  38900=>"111111000",
  38901=>"110111010",
  38902=>"111111110",
  38903=>"111110100",
  38904=>"111111000",
  38905=>"001011011",
  38906=>"100100110",
  38907=>"111111110",
  38908=>"110110000",
  38909=>"000000011",
  38910=>"101000000",
  38911=>"111111000",
  38912=>"111111111",
  38913=>"111100110",
  38914=>"000000111",
  38915=>"001001001",
  38916=>"001001111",
  38917=>"000000000",
  38918=>"010111010",
  38919=>"000100111",
  38920=>"001001001",
  38921=>"000000101",
  38922=>"000000000",
  38923=>"000011000",
  38924=>"000000010",
  38925=>"100101111",
  38926=>"000001101",
  38927=>"110111110",
  38928=>"000000111",
  38929=>"000000111",
  38930=>"000001000",
  38931=>"111111111",
  38932=>"000000000",
  38933=>"000010111",
  38934=>"101001111",
  38935=>"110110110",
  38936=>"000101110",
  38937=>"111000000",
  38938=>"000000111",
  38939=>"111111111",
  38940=>"000000000",
  38941=>"111111111",
  38942=>"111111111",
  38943=>"010000000",
  38944=>"000000000",
  38945=>"000000000",
  38946=>"111111111",
  38947=>"101000101",
  38948=>"111111111",
  38949=>"000000111",
  38950=>"111111111",
  38951=>"000101111",
  38952=>"000000001",
  38953=>"000000000",
  38954=>"111011000",
  38955=>"011010010",
  38956=>"000100000",
  38957=>"000000000",
  38958=>"111110010",
  38959=>"111111111",
  38960=>"101111111",
  38961=>"000111111",
  38962=>"000000000",
  38963=>"100000000",
  38964=>"000000000",
  38965=>"100100000",
  38966=>"000000000",
  38967=>"100100111",
  38968=>"111111011",
  38969=>"111111111",
  38970=>"000000000",
  38971=>"000000000",
  38972=>"111100000",
  38973=>"111101111",
  38974=>"000000000",
  38975=>"110001111",
  38976=>"011101000",
  38977=>"000000110",
  38978=>"000000000",
  38979=>"001000000",
  38980=>"110001111",
  38981=>"011010010",
  38982=>"000000001",
  38983=>"111111111",
  38984=>"001011011",
  38985=>"001000001",
  38986=>"111111111",
  38987=>"111111111",
  38988=>"111110111",
  38989=>"000000010",
  38990=>"010000000",
  38991=>"000000000",
  38992=>"110100000",
  38993=>"000111111",
  38994=>"000000000",
  38995=>"011001111",
  38996=>"000000001",
  38997=>"000000010",
  38998=>"100000000",
  38999=>"101111101",
  39000=>"000000000",
  39001=>"111111111",
  39002=>"001000000",
  39003=>"000000000",
  39004=>"000011111",
  39005=>"000000000",
  39006=>"000000000",
  39007=>"110011011",
  39008=>"100000000",
  39009=>"111000110",
  39010=>"100111101",
  39011=>"111111111",
  39012=>"000111111",
  39013=>"111010010",
  39014=>"000111111",
  39015=>"000000010",
  39016=>"000000000",
  39017=>"000000000",
  39018=>"111110010",
  39019=>"000000111",
  39020=>"111100000",
  39021=>"111111111",
  39022=>"111111111",
  39023=>"000000110",
  39024=>"010111111",
  39025=>"011111000",
  39026=>"111111001",
  39027=>"000000010",
  39028=>"111111101",
  39029=>"011011111",
  39030=>"000000111",
  39031=>"000000000",
  39032=>"000000000",
  39033=>"110111111",
  39034=>"010001001",
  39035=>"000000011",
  39036=>"100110100",
  39037=>"000111001",
  39038=>"111111111",
  39039=>"111111011",
  39040=>"000010010",
  39041=>"111111111",
  39042=>"111111000",
  39043=>"000000000",
  39044=>"110111010",
  39045=>"001000000",
  39046=>"000000000",
  39047=>"000000000",
  39048=>"111111111",
  39049=>"000000000",
  39050=>"011111000",
  39051=>"000101000",
  39052=>"110110110",
  39053=>"100010111",
  39054=>"000000000",
  39055=>"000000000",
  39056=>"001000000",
  39057=>"111111111",
  39058=>"000000010",
  39059=>"100000000",
  39060=>"111111110",
  39061=>"000000000",
  39062=>"001111110",
  39063=>"111111111",
  39064=>"000000011",
  39065=>"111111011",
  39066=>"100101111",
  39067=>"000000000",
  39068=>"111001111",
  39069=>"110000100",
  39070=>"001011010",
  39071=>"000000000",
  39072=>"111011111",
  39073=>"111011111",
  39074=>"000011111",
  39075=>"000001000",
  39076=>"000000001",
  39077=>"000000111",
  39078=>"000000000",
  39079=>"111111000",
  39080=>"000000001",
  39081=>"000000000",
  39082=>"100000000",
  39083=>"000000000",
  39084=>"001000011",
  39085=>"011100000",
  39086=>"111111111",
  39087=>"100000000",
  39088=>"001000000",
  39089=>"000000000",
  39090=>"111111111",
  39091=>"111011000",
  39092=>"000000000",
  39093=>"111011001",
  39094=>"111110000",
  39095=>"000000000",
  39096=>"111000110",
  39097=>"110010111",
  39098=>"000010101",
  39099=>"000000010",
  39100=>"001111111",
  39101=>"000000000",
  39102=>"110110000",
  39103=>"000110111",
  39104=>"100100111",
  39105=>"000000111",
  39106=>"101111100",
  39107=>"000000000",
  39108=>"000000000",
  39109=>"100011000",
  39110=>"000000000",
  39111=>"110100000",
  39112=>"000000000",
  39113=>"000000000",
  39114=>"101011111",
  39115=>"000000000",
  39116=>"001101001",
  39117=>"111111111",
  39118=>"000000000",
  39119=>"011001001",
  39120=>"000010000",
  39121=>"111111100",
  39122=>"110111110",
  39123=>"000000000",
  39124=>"101111111",
  39125=>"111110110",
  39126=>"000100111",
  39127=>"000000111",
  39128=>"111111111",
  39129=>"111001000",
  39130=>"000000000",
  39131=>"000010111",
  39132=>"000000000",
  39133=>"111111111",
  39134=>"000111111",
  39135=>"011000000",
  39136=>"000000111",
  39137=>"000010111",
  39138=>"000000101",
  39139=>"111001000",
  39140=>"101111111",
  39141=>"000000000",
  39142=>"110000100",
  39143=>"011001001",
  39144=>"001000000",
  39145=>"010010010",
  39146=>"110111111",
  39147=>"000000011",
  39148=>"000000000",
  39149=>"000000000",
  39150=>"110000000",
  39151=>"000000000",
  39152=>"111111100",
  39153=>"000000001",
  39154=>"111111101",
  39155=>"000000000",
  39156=>"000000000",
  39157=>"110110110",
  39158=>"000010000",
  39159=>"111111111",
  39160=>"000000111",
  39161=>"111111100",
  39162=>"111010011",
  39163=>"000000000",
  39164=>"111111100",
  39165=>"011011001",
  39166=>"111101000",
  39167=>"111111111",
  39168=>"000000000",
  39169=>"000000000",
  39170=>"111111110",
  39171=>"000010000",
  39172=>"001001101",
  39173=>"111011000",
  39174=>"000000000",
  39175=>"111111110",
  39176=>"100000000",
  39177=>"000000100",
  39178=>"000100100",
  39179=>"000000000",
  39180=>"111100000",
  39181=>"111000000",
  39182=>"000011111",
  39183=>"100000000",
  39184=>"100000111",
  39185=>"111111101",
  39186=>"111111111",
  39187=>"001011010",
  39188=>"000001001",
  39189=>"111111111",
  39190=>"000000101",
  39191=>"001101111",
  39192=>"000011111",
  39193=>"011111011",
  39194=>"111111111",
  39195=>"000000000",
  39196=>"000100111",
  39197=>"111111101",
  39198=>"000001001",
  39199=>"000000001",
  39200=>"100111100",
  39201=>"111001000",
  39202=>"000100100",
  39203=>"100101111",
  39204=>"000100111",
  39205=>"000000000",
  39206=>"110111110",
  39207=>"000000000",
  39208=>"111111111",
  39209=>"111111111",
  39210=>"010010111",
  39211=>"000000111",
  39212=>"100100101",
  39213=>"000001001",
  39214=>"111111101",
  39215=>"111111111",
  39216=>"000000000",
  39217=>"110000000",
  39218=>"111111111",
  39219=>"001111111",
  39220=>"111111000",
  39221=>"111000000",
  39222=>"111011111",
  39223=>"111111111",
  39224=>"000000000",
  39225=>"111111111",
  39226=>"111111111",
  39227=>"000000000",
  39228=>"111111111",
  39229=>"011010111",
  39230=>"101111010",
  39231=>"111111111",
  39232=>"011011001",
  39233=>"000000000",
  39234=>"000011011",
  39235=>"101101101",
  39236=>"111111111",
  39237=>"010110111",
  39238=>"000000100",
  39239=>"100111110",
  39240=>"010010110",
  39241=>"000000011",
  39242=>"111011001",
  39243=>"110010111",
  39244=>"000000111",
  39245=>"000000000",
  39246=>"000000000",
  39247=>"110111101",
  39248=>"000001000",
  39249=>"011000000",
  39250=>"111111110",
  39251=>"111111111",
  39252=>"000000000",
  39253=>"111001000",
  39254=>"000000000",
  39255=>"000000111",
  39256=>"111000000",
  39257=>"111111000",
  39258=>"111111000",
  39259=>"000001001",
  39260=>"111010110",
  39261=>"000111111",
  39262=>"111011001",
  39263=>"001001011",
  39264=>"111100101",
  39265=>"001101111",
  39266=>"111111111",
  39267=>"111111111",
  39268=>"111110000",
  39269=>"111111111",
  39270=>"111110110",
  39271=>"110111111",
  39272=>"011001001",
  39273=>"000000110",
  39274=>"100111111",
  39275=>"001001011",
  39276=>"111111011",
  39277=>"010000011",
  39278=>"111111100",
  39279=>"111111111",
  39280=>"111000000",
  39281=>"110011111",
  39282=>"111111000",
  39283=>"000000001",
  39284=>"111111000",
  39285=>"110111111",
  39286=>"111011011",
  39287=>"111111001",
  39288=>"000000000",
  39289=>"000000000",
  39290=>"001010110",
  39291=>"111111111",
  39292=>"111001001",
  39293=>"000000001",
  39294=>"111111101",
  39295=>"111111111",
  39296=>"000100100",
  39297=>"111111111",
  39298=>"100110000",
  39299=>"000000000",
  39300=>"000000100",
  39301=>"111111111",
  39302=>"111110000",
  39303=>"110010011",
  39304=>"111111111",
  39305=>"000011111",
  39306=>"000000111",
  39307=>"000000000",
  39308=>"101111111",
  39309=>"111101111",
  39310=>"000000000",
  39311=>"000011000",
  39312=>"100111000",
  39313=>"111110100",
  39314=>"111111000",
  39315=>"111111110",
  39316=>"111111111",
  39317=>"000010000",
  39318=>"010000000",
  39319=>"001000100",
  39320=>"000011111",
  39321=>"111110000",
  39322=>"111111111",
  39323=>"111000000",
  39324=>"100000000",
  39325=>"000000011",
  39326=>"110110100",
  39327=>"111111111",
  39328=>"011111111",
  39329=>"111111110",
  39330=>"111001100",
  39331=>"000010111",
  39332=>"111111111",
  39333=>"000110111",
  39334=>"011000000",
  39335=>"111000000",
  39336=>"000000000",
  39337=>"000000000",
  39338=>"111111111",
  39339=>"110111110",
  39340=>"000110111",
  39341=>"000000000",
  39342=>"000000000",
  39343=>"111000000",
  39344=>"100100000",
  39345=>"111111111",
  39346=>"000001111",
  39347=>"000000011",
  39348=>"000100111",
  39349=>"011111010",
  39350=>"111111011",
  39351=>"000000001",
  39352=>"000000111",
  39353=>"001010000",
  39354=>"000111111",
  39355=>"000000001",
  39356=>"111111111",
  39357=>"000000110",
  39358=>"000000110",
  39359=>"110100110",
  39360=>"111111111",
  39361=>"000000000",
  39362=>"111111111",
  39363=>"000000000",
  39364=>"111111111",
  39365=>"111111111",
  39366=>"000000000",
  39367=>"000000011",
  39368=>"101000111",
  39369=>"111111001",
  39370=>"100000000",
  39371=>"111111111",
  39372=>"000110110",
  39373=>"111100110",
  39374=>"110111111",
  39375=>"111111111",
  39376=>"000111110",
  39377=>"000000000",
  39378=>"010010111",
  39379=>"111000111",
  39380=>"111111111",
  39381=>"111111111",
  39382=>"000000100",
  39383=>"000000010",
  39384=>"100111111",
  39385=>"111111110",
  39386=>"100100000",
  39387=>"001000000",
  39388=>"000000000",
  39389=>"000110110",
  39390=>"001001000",
  39391=>"001001111",
  39392=>"000000111",
  39393=>"000110100",
  39394=>"000000000",
  39395=>"110000111",
  39396=>"111111111",
  39397=>"000011000",
  39398=>"111111111",
  39399=>"011000100",
  39400=>"000100110",
  39401=>"000000100",
  39402=>"100100100",
  39403=>"000000111",
  39404=>"000000000",
  39405=>"110000000",
  39406=>"111111111",
  39407=>"000110111",
  39408=>"000001001",
  39409=>"110000110",
  39410=>"110111111",
  39411=>"000000000",
  39412=>"101111111",
  39413=>"100100111",
  39414=>"111111101",
  39415=>"111111000",
  39416=>"000000000",
  39417=>"100000001",
  39418=>"000010000",
  39419=>"111111111",
  39420=>"111110110",
  39421=>"110100110",
  39422=>"111101111",
  39423=>"111111000",
  39424=>"000000000",
  39425=>"111111111",
  39426=>"000000000",
  39427=>"000000111",
  39428=>"100100100",
  39429=>"000010011",
  39430=>"111101111",
  39431=>"111111111",
  39432=>"110111111",
  39433=>"001001001",
  39434=>"001001001",
  39435=>"110110111",
  39436=>"001001000",
  39437=>"000010110",
  39438=>"100000000",
  39439=>"100111111",
  39440=>"111111000",
  39441=>"110001111",
  39442=>"000101111",
  39443=>"111111100",
  39444=>"111111000",
  39445=>"001000000",
  39446=>"111000000",
  39447=>"110011000",
  39448=>"111110110",
  39449=>"000000001",
  39450=>"111000101",
  39451=>"111111111",
  39452=>"000000000",
  39453=>"111111001",
  39454=>"001001111",
  39455=>"000000001",
  39456=>"100001000",
  39457=>"111111111",
  39458=>"111110010",
  39459=>"111111110",
  39460=>"111100000",
  39461=>"111011111",
  39462=>"011000000",
  39463=>"111100100",
  39464=>"000000000",
  39465=>"000000000",
  39466=>"011000000",
  39467=>"000000110",
  39468=>"111111111",
  39469=>"111111111",
  39470=>"000011011",
  39471=>"111000000",
  39472=>"000001111",
  39473=>"000000000",
  39474=>"001111111",
  39475=>"000000111",
  39476=>"000000000",
  39477=>"001001000",
  39478=>"111111111",
  39479=>"101011111",
  39480=>"111100101",
  39481=>"011000111",
  39482=>"000000000",
  39483=>"111000000",
  39484=>"000000111",
  39485=>"111101000",
  39486=>"000000000",
  39487=>"111000000",
  39488=>"000000111",
  39489=>"001000101",
  39490=>"111000000",
  39491=>"111111111",
  39492=>"001011111",
  39493=>"111011001",
  39494=>"111111011",
  39495=>"111011000",
  39496=>"000001000",
  39497=>"000000111",
  39498=>"000000100",
  39499=>"111101101",
  39500=>"011111111",
  39501=>"111001001",
  39502=>"110110011",
  39503=>"111111111",
  39504=>"000000000",
  39505=>"000001011",
  39506=>"111111100",
  39507=>"000000000",
  39508=>"001000001",
  39509=>"111111111",
  39510=>"000000111",
  39511=>"011111111",
  39512=>"001000110",
  39513=>"101000111",
  39514=>"111111111",
  39515=>"000000000",
  39516=>"000011000",
  39517=>"000011111",
  39518=>"000000000",
  39519=>"000000000",
  39520=>"000011111",
  39521=>"111111011",
  39522=>"111111111",
  39523=>"111111101",
  39524=>"111110110",
  39525=>"000101111",
  39526=>"111010000",
  39527=>"000100100",
  39528=>"000000000",
  39529=>"111111000",
  39530=>"111001111",
  39531=>"111111111",
  39532=>"000000000",
  39533=>"111111000",
  39534=>"000011011",
  39535=>"111000000",
  39536=>"110001000",
  39537=>"011111001",
  39538=>"111011001",
  39539=>"010010010",
  39540=>"111111111",
  39541=>"111101000",
  39542=>"111111000",
  39543=>"111000000",
  39544=>"000111111",
  39545=>"111000011",
  39546=>"100110110",
  39547=>"111111111",
  39548=>"000100111",
  39549=>"000000000",
  39550=>"000000110",
  39551=>"000011011",
  39552=>"001001000",
  39553=>"000000000",
  39554=>"000000000",
  39555=>"000000001",
  39556=>"000110110",
  39557=>"111000111",
  39558=>"111000111",
  39559=>"111111000",
  39560=>"000000000",
  39561=>"000110010",
  39562=>"111000000",
  39563=>"011000000",
  39564=>"111111110",
  39565=>"000000111",
  39566=>"001000111",
  39567=>"000011101",
  39568=>"111111111",
  39569=>"000000010",
  39570=>"000110110",
  39571=>"101001011",
  39572=>"111111000",
  39573=>"111000000",
  39574=>"101011111",
  39575=>"111111100",
  39576=>"100101000",
  39577=>"111111111",
  39578=>"111000000",
  39579=>"111101101",
  39580=>"111111111",
  39581=>"000111111",
  39582=>"001101101",
  39583=>"001001000",
  39584=>"000000001",
  39585=>"111111111",
  39586=>"111101000",
  39587=>"000000001",
  39588=>"001000111",
  39589=>"000001111",
  39590=>"111111111",
  39591=>"000110100",
  39592=>"011010000",
  39593=>"001001111",
  39594=>"111001111",
  39595=>"111111101",
  39596=>"010000000",
  39597=>"000000101",
  39598=>"111111111",
  39599=>"000000000",
  39600=>"111110000",
  39601=>"000000100",
  39602=>"110111000",
  39603=>"000011111",
  39604=>"000000000",
  39605=>"000000000",
  39606=>"111111000",
  39607=>"111111111",
  39608=>"100111111",
  39609=>"111000000",
  39610=>"100001111",
  39611=>"100001111",
  39612=>"110110111",
  39613=>"111001011",
  39614=>"111110100",
  39615=>"111111111",
  39616=>"000000111",
  39617=>"001001111",
  39618=>"000000111",
  39619=>"111001111",
  39620=>"111111000",
  39621=>"000000000",
  39622=>"000000000",
  39623=>"000101101",
  39624=>"000000000",
  39625=>"000000110",
  39626=>"000100111",
  39627=>"111000000",
  39628=>"011111111",
  39629=>"000000010",
  39630=>"000000011",
  39631=>"000000000",
  39632=>"100111000",
  39633=>"110000000",
  39634=>"111111000",
  39635=>"000000001",
  39636=>"001000000",
  39637=>"110100000",
  39638=>"111111000",
  39639=>"010000111",
  39640=>"111111000",
  39641=>"111111111",
  39642=>"000010010",
  39643=>"000000000",
  39644=>"001011111",
  39645=>"111110000",
  39646=>"110000000",
  39647=>"000000001",
  39648=>"100000110",
  39649=>"000000111",
  39650=>"010111110",
  39651=>"111000000",
  39652=>"000000000",
  39653=>"000000000",
  39654=>"111100000",
  39655=>"100000000",
  39656=>"110110100",
  39657=>"011101111",
  39658=>"101111110",
  39659=>"000110111",
  39660=>"111111111",
  39661=>"011111010",
  39662=>"111111101",
  39663=>"000110100",
  39664=>"000000000",
  39665=>"111111000",
  39666=>"101111111",
  39667=>"000010111",
  39668=>"111111000",
  39669=>"000000000",
  39670=>"111111111",
  39671=>"100000000",
  39672=>"000110111",
  39673=>"000000000",
  39674=>"001001111",
  39675=>"000000000",
  39676=>"000000000",
  39677=>"000000100",
  39678=>"001111100",
  39679=>"111111111",
  39680=>"101111101",
  39681=>"000000000",
  39682=>"111100111",
  39683=>"000000000",
  39684=>"111111111",
  39685=>"111011000",
  39686=>"111101100",
  39687=>"011000101",
  39688=>"000000000",
  39689=>"000000000",
  39690=>"111111111",
  39691=>"111111111",
  39692=>"000001111",
  39693=>"110111110",
  39694=>"110111110",
  39695=>"111000000",
  39696=>"000000100",
  39697=>"011001010",
  39698=>"110010111",
  39699=>"111111100",
  39700=>"111100000",
  39701=>"111111000",
  39702=>"101000001",
  39703=>"111101101",
  39704=>"000100000",
  39705=>"000000000",
  39706=>"000001000",
  39707=>"111000000",
  39708=>"101100111",
  39709=>"001011111",
  39710=>"100110110",
  39711=>"000000000",
  39712=>"111110011",
  39713=>"000010111",
  39714=>"000000000",
  39715=>"000000011",
  39716=>"000000110",
  39717=>"001001000",
  39718=>"000000110",
  39719=>"011111111",
  39720=>"110010000",
  39721=>"000011111",
  39722=>"000000010",
  39723=>"111011110",
  39724=>"000000000",
  39725=>"110110111",
  39726=>"000000000",
  39727=>"000000000",
  39728=>"111111111",
  39729=>"000000000",
  39730=>"000000011",
  39731=>"000000010",
  39732=>"000000111",
  39733=>"000000000",
  39734=>"011010000",
  39735=>"111111100",
  39736=>"111111000",
  39737=>"000000100",
  39738=>"111101100",
  39739=>"111111111",
  39740=>"011111111",
  39741=>"000000000",
  39742=>"110000011",
  39743=>"000000000",
  39744=>"100000101",
  39745=>"111111111",
  39746=>"011000000",
  39747=>"000101111",
  39748=>"111100011",
  39749=>"111011101",
  39750=>"000000000",
  39751=>"001000000",
  39752=>"000000010",
  39753=>"001001000",
  39754=>"000000000",
  39755=>"000000000",
  39756=>"110110000",
  39757=>"111001111",
  39758=>"111000000",
  39759=>"110110000",
  39760=>"110110100",
  39761=>"000000110",
  39762=>"001000000",
  39763=>"000000111",
  39764=>"000100110",
  39765=>"011011011",
  39766=>"110100100",
  39767=>"001001111",
  39768=>"000000000",
  39769=>"111111111",
  39770=>"000011011",
  39771=>"111111111",
  39772=>"000000000",
  39773=>"000000000",
  39774=>"011111000",
  39775=>"000000000",
  39776=>"111111001",
  39777=>"110111111",
  39778=>"100110111",
  39779=>"000000111",
  39780=>"100000000",
  39781=>"000011111",
  39782=>"111111111",
  39783=>"000000000",
  39784=>"001001001",
  39785=>"110010000",
  39786=>"000000111",
  39787=>"000000000",
  39788=>"111111111",
  39789=>"000111111",
  39790=>"011011001",
  39791=>"110000000",
  39792=>"111111111",
  39793=>"110110111",
  39794=>"000000000",
  39795=>"111111000",
  39796=>"111000000",
  39797=>"111000000",
  39798=>"111111111",
  39799=>"000000100",
  39800=>"000000111",
  39801=>"110111111",
  39802=>"000000000",
  39803=>"000000110",
  39804=>"110010010",
  39805=>"111111000",
  39806=>"111111111",
  39807=>"001000000",
  39808=>"000000111",
  39809=>"100000100",
  39810=>"111110110",
  39811=>"111111111",
  39812=>"011111111",
  39813=>"110111111",
  39814=>"000000000",
  39815=>"000000000",
  39816=>"001011010",
  39817=>"111111111",
  39818=>"000000011",
  39819=>"111000000",
  39820=>"001011111",
  39821=>"010110100",
  39822=>"111111111",
  39823=>"000110000",
  39824=>"000111111",
  39825=>"000001111",
  39826=>"111111111",
  39827=>"110110111",
  39828=>"000101010",
  39829=>"000000000",
  39830=>"100100110",
  39831=>"000110111",
  39832=>"101100111",
  39833=>"000000111",
  39834=>"000000000",
  39835=>"000000000",
  39836=>"000110000",
  39837=>"111111111",
  39838=>"000000000",
  39839=>"000000111",
  39840=>"111011000",
  39841=>"111111001",
  39842=>"000000000",
  39843=>"111111111",
  39844=>"000000001",
  39845=>"001011011",
  39846=>"111001111",
  39847=>"111111111",
  39848=>"100111111",
  39849=>"000000000",
  39850=>"111101111",
  39851=>"100000110",
  39852=>"000000000",
  39853=>"000001101",
  39854=>"011010000",
  39855=>"000000000",
  39856=>"111111111",
  39857=>"110110000",
  39858=>"111111111",
  39859=>"011111000",
  39860=>"001000000",
  39861=>"000000000",
  39862=>"111111111",
  39863=>"111101000",
  39864=>"110000000",
  39865=>"111111111",
  39866=>"000011000",
  39867=>"111011111",
  39868=>"101000011",
  39869=>"111111111",
  39870=>"000000001",
  39871=>"100100111",
  39872=>"011011011",
  39873=>"000000111",
  39874=>"000000000",
  39875=>"110110111",
  39876=>"111110111",
  39877=>"000000110",
  39878=>"111111101",
  39879=>"000000011",
  39880=>"100100111",
  39881=>"111100101",
  39882=>"000000001",
  39883=>"000000000",
  39884=>"000000000",
  39885=>"111000000",
  39886=>"100000001",
  39887=>"111111111",
  39888=>"000000000",
  39889=>"111011000",
  39890=>"000100111",
  39891=>"100000111",
  39892=>"101101111",
  39893=>"000000011",
  39894=>"000000000",
  39895=>"111111111",
  39896=>"111110111",
  39897=>"011111111",
  39898=>"111000000",
  39899=>"111100000",
  39900=>"111111000",
  39901=>"001000111",
  39902=>"111111100",
  39903=>"011111111",
  39904=>"110111111",
  39905=>"000000000",
  39906=>"111011000",
  39907=>"111111111",
  39908=>"111000000",
  39909=>"100000011",
  39910=>"000000000",
  39911=>"111111000",
  39912=>"000000000",
  39913=>"000000000",
  39914=>"000000000",
  39915=>"000000000",
  39916=>"000111011",
  39917=>"000001111",
  39918=>"101000000",
  39919=>"100000000",
  39920=>"000000110",
  39921=>"111111111",
  39922=>"111111010",
  39923=>"011001000",
  39924=>"111110110",
  39925=>"011110000",
  39926=>"001001011",
  39927=>"000000000",
  39928=>"111111111",
  39929=>"000000000",
  39930=>"111110010",
  39931=>"111111000",
  39932=>"000000000",
  39933=>"100100100",
  39934=>"111110100",
  39935=>"000000000",
  39936=>"000000000",
  39937=>"111000000",
  39938=>"000000000",
  39939=>"000110110",
  39940=>"000100011",
  39941=>"111111101",
  39942=>"000000000",
  39943=>"111111100",
  39944=>"111111111",
  39945=>"111111101",
  39946=>"000110000",
  39947=>"000000001",
  39948=>"000110111",
  39949=>"001000000",
  39950=>"000000000",
  39951=>"111111000",
  39952=>"111111111",
  39953=>"000111111",
  39954=>"000000100",
  39955=>"000000000",
  39956=>"111111111",
  39957=>"010000000",
  39958=>"111111000",
  39959=>"011011110",
  39960=>"000100100",
  39961=>"101100111",
  39962=>"001000000",
  39963=>"100111110",
  39964=>"001111111",
  39965=>"000000111",
  39966=>"000010000",
  39967=>"111100111",
  39968=>"010000000",
  39969=>"011111110",
  39970=>"000000000",
  39971=>"111101000",
  39972=>"000000000",
  39973=>"111000000",
  39974=>"001001001",
  39975=>"111111111",
  39976=>"111111111",
  39977=>"000000000",
  39978=>"000000000",
  39979=>"001011111",
  39980=>"011111111",
  39981=>"110110000",
  39982=>"000000111",
  39983=>"000110111",
  39984=>"111111011",
  39985=>"111000000",
  39986=>"000000000",
  39987=>"111111000",
  39988=>"000000000",
  39989=>"111111111",
  39990=>"011000001",
  39991=>"111111111",
  39992=>"100000000",
  39993=>"000001000",
  39994=>"000000000",
  39995=>"111000000",
  39996=>"101001111",
  39997=>"000000000",
  39998=>"000000000",
  39999=>"111111111",
  40000=>"001100111",
  40001=>"000000000",
  40002=>"111000000",
  40003=>"100100100",
  40004=>"100000000",
  40005=>"110111111",
  40006=>"001000000",
  40007=>"111111111",
  40008=>"000000011",
  40009=>"101001101",
  40010=>"000000000",
  40011=>"100000000",
  40012=>"000000101",
  40013=>"000000000",
  40014=>"111111111",
  40015=>"000111111",
  40016=>"000000001",
  40017=>"111011000",
  40018=>"000000000",
  40019=>"001111111",
  40020=>"000110000",
  40021=>"110111111",
  40022=>"000000001",
  40023=>"000111111",
  40024=>"111000100",
  40025=>"111000000",
  40026=>"001001000",
  40027=>"001000000",
  40028=>"011011111",
  40029=>"100110110",
  40030=>"000101001",
  40031=>"000000111",
  40032=>"000000000",
  40033=>"000000000",
  40034=>"000000001",
  40035=>"001001111",
  40036=>"111111000",
  40037=>"100100101",
  40038=>"111111000",
  40039=>"111111111",
  40040=>"000001000",
  40041=>"001001111",
  40042=>"000001111",
  40043=>"000101111",
  40044=>"000000000",
  40045=>"111011000",
  40046=>"001000000",
  40047=>"001001001",
  40048=>"010110000",
  40049=>"111111111",
  40050=>"011011011",
  40051=>"011111111",
  40052=>"111111111",
  40053=>"000000011",
  40054=>"000000000",
  40055=>"000111111",
  40056=>"100111101",
  40057=>"111111111",
  40058=>"110000000",
  40059=>"111111011",
  40060=>"100100111",
  40061=>"000110111",
  40062=>"000000000",
  40063=>"000000000",
  40064=>"111001111",
  40065=>"110110100",
  40066=>"000000000",
  40067=>"111111001",
  40068=>"000000000",
  40069=>"111100001",
  40070=>"111111111",
  40071=>"000000000",
  40072=>"111110110",
  40073=>"000000010",
  40074=>"000000100",
  40075=>"000000001",
  40076=>"000000001",
  40077=>"111111110",
  40078=>"111111111",
  40079=>"100000000",
  40080=>"000000000",
  40081=>"000000000",
  40082=>"000000000",
  40083=>"110010111",
  40084=>"110010000",
  40085=>"000000010",
  40086=>"000000000",
  40087=>"000000000",
  40088=>"111001000",
  40089=>"111111111",
  40090=>"000000000",
  40091=>"001000001",
  40092=>"000000011",
  40093=>"000000000",
  40094=>"001101111",
  40095=>"000011000",
  40096=>"111000000",
  40097=>"111100000",
  40098=>"111111010",
  40099=>"111111111",
  40100=>"000000000",
  40101=>"110111111",
  40102=>"111111000",
  40103=>"011011001",
  40104=>"111111111",
  40105=>"111111101",
  40106=>"000111000",
  40107=>"010000010",
  40108=>"001111111",
  40109=>"100011100",
  40110=>"100111111",
  40111=>"111111001",
  40112=>"111111110",
  40113=>"111111111",
  40114=>"111111111",
  40115=>"000000000",
  40116=>"000001001",
  40117=>"000000000",
  40118=>"001011001",
  40119=>"000000000",
  40120=>"100100111",
  40121=>"111111111",
  40122=>"010000011",
  40123=>"001001001",
  40124=>"000000000",
  40125=>"001111111",
  40126=>"111000000",
  40127=>"111111000",
  40128=>"000100101",
  40129=>"111111111",
  40130=>"110110111",
  40131=>"000000000",
  40132=>"010011111",
  40133=>"111000000",
  40134=>"101000000",
  40135=>"000000000",
  40136=>"111101111",
  40137=>"000000000",
  40138=>"000000101",
  40139=>"111110000",
  40140=>"100100000",
  40141=>"000001101",
  40142=>"001111101",
  40143=>"000110110",
  40144=>"001011011",
  40145=>"100111111",
  40146=>"111011000",
  40147=>"000000000",
  40148=>"000000000",
  40149=>"000000000",
  40150=>"100100000",
  40151=>"000000000",
  40152=>"111011000",
  40153=>"100111001",
  40154=>"000000010",
  40155=>"000000000",
  40156=>"111111111",
  40157=>"000100100",
  40158=>"000000000",
  40159=>"000000011",
  40160=>"000001111",
  40161=>"000110011",
  40162=>"000000000",
  40163=>"001000000",
  40164=>"111111111",
  40165=>"100000000",
  40166=>"001010111",
  40167=>"111111000",
  40168=>"000000000",
  40169=>"000000000",
  40170=>"100110100",
  40171=>"000000000",
  40172=>"111111111",
  40173=>"000000010",
  40174=>"000000111",
  40175=>"000000101",
  40176=>"111111111",
  40177=>"000100111",
  40178=>"111100100",
  40179=>"000000000",
  40180=>"111111111",
  40181=>"000000101",
  40182=>"010100000",
  40183=>"000000000",
  40184=>"110110110",
  40185=>"111111111",
  40186=>"101111111",
  40187=>"000000000",
  40188=>"011000000",
  40189=>"101101111",
  40190=>"000110111",
  40191=>"111100000",
  40192=>"000000000",
  40193=>"111111111",
  40194=>"000000000",
  40195=>"000001000",
  40196=>"111111011",
  40197=>"101111111",
  40198=>"000000000",
  40199=>"000000000",
  40200=>"111000000",
  40201=>"000000101",
  40202=>"001001000",
  40203=>"100100000",
  40204=>"001001001",
  40205=>"000010010",
  40206=>"000111111",
  40207=>"000010110",
  40208=>"011000011",
  40209=>"100100000",
  40210=>"010111111",
  40211=>"001101001",
  40212=>"000000000",
  40213=>"111111110",
  40214=>"100100100",
  40215=>"101000000",
  40216=>"111111111",
  40217=>"111111010",
  40218=>"010000001",
  40219=>"101111011",
  40220=>"001001001",
  40221=>"011000000",
  40222=>"111111111",
  40223=>"000110000",
  40224=>"000000000",
  40225=>"000000000",
  40226=>"110111110",
  40227=>"111111111",
  40228=>"101000000",
  40229=>"110111111",
  40230=>"011000000",
  40231=>"000000111",
  40232=>"000000110",
  40233=>"011011111",
  40234=>"000100110",
  40235=>"010011111",
  40236=>"000000000",
  40237=>"100100000",
  40238=>"000000000",
  40239=>"000000001",
  40240=>"101001101",
  40241=>"000000000",
  40242=>"011111111",
  40243=>"000000110",
  40244=>"111111110",
  40245=>"011000000",
  40246=>"000000000",
  40247=>"101000000",
  40248=>"000000000",
  40249=>"111000111",
  40250=>"000111111",
  40251=>"111111000",
  40252=>"110110010",
  40253=>"000000000",
  40254=>"011000010",
  40255=>"111111111",
  40256=>"000000000",
  40257=>"000110000",
  40258=>"000111111",
  40259=>"111111111",
  40260=>"000000100",
  40261=>"111011111",
  40262=>"011000001",
  40263=>"000000000",
  40264=>"111111111",
  40265=>"011001001",
  40266=>"111110110",
  40267=>"000100100",
  40268=>"110011000",
  40269=>"111111011",
  40270=>"001101000",
  40271=>"111100111",
  40272=>"100100100",
  40273=>"000000000",
  40274=>"000000000",
  40275=>"000000000",
  40276=>"000000000",
  40277=>"001011011",
  40278=>"110110011",
  40279=>"111111111",
  40280=>"111111110",
  40281=>"111111111",
  40282=>"000001111",
  40283=>"110111111",
  40284=>"000001000",
  40285=>"000000000",
  40286=>"111111111",
  40287=>"111111111",
  40288=>"111111111",
  40289=>"111111111",
  40290=>"001000001",
  40291=>"101100100",
  40292=>"000001000",
  40293=>"000000000",
  40294=>"111110001",
  40295=>"000000000",
  40296=>"000000000",
  40297=>"110110000",
  40298=>"000000000",
  40299=>"111111101",
  40300=>"000101001",
  40301=>"000000111",
  40302=>"111111111",
  40303=>"000000000",
  40304=>"000111111",
  40305=>"000000000",
  40306=>"000111111",
  40307=>"111111100",
  40308=>"000000100",
  40309=>"111111101",
  40310=>"000000000",
  40311=>"000100110",
  40312=>"111011111",
  40313=>"000100000",
  40314=>"111111111",
  40315=>"111111111",
  40316=>"010111111",
  40317=>"111111111",
  40318=>"011001111",
  40319=>"000000000",
  40320=>"101111111",
  40321=>"111111000",
  40322=>"000111111",
  40323=>"111111111",
  40324=>"100111111",
  40325=>"000000101",
  40326=>"001000000",
  40327=>"110100000",
  40328=>"000000111",
  40329=>"000000110",
  40330=>"110111111",
  40331=>"000000100",
  40332=>"111111111",
  40333=>"111111111",
  40334=>"100100000",
  40335=>"000000000",
  40336=>"011011001",
  40337=>"111111110",
  40338=>"100001100",
  40339=>"001001111",
  40340=>"000000010",
  40341=>"000000000",
  40342=>"011011111",
  40343=>"000000100",
  40344=>"110000000",
  40345=>"011010110",
  40346=>"111110010",
  40347=>"001000000",
  40348=>"110000000",
  40349=>"110111111",
  40350=>"000000000",
  40351=>"111111111",
  40352=>"111111111",
  40353=>"001011111",
  40354=>"100110111",
  40355=>"000000000",
  40356=>"100000000",
  40357=>"000001001",
  40358=>"111111111",
  40359=>"000000000",
  40360=>"111111111",
  40361=>"110111111",
  40362=>"001111111",
  40363=>"010000000",
  40364=>"000001111",
  40365=>"111000001",
  40366=>"000000110",
  40367=>"000100000",
  40368=>"000000000",
  40369=>"000110111",
  40370=>"000000000",
  40371=>"111111111",
  40372=>"111111111",
  40373=>"111110110",
  40374=>"111111111",
  40375=>"000000000",
  40376=>"110000000",
  40377=>"000110111",
  40378=>"010011111",
  40379=>"111111111",
  40380=>"101111111",
  40381=>"111111000",
  40382=>"000000000",
  40383=>"111101101",
  40384=>"110000000",
  40385=>"000000000",
  40386=>"000000000",
  40387=>"111111111",
  40388=>"000000101",
  40389=>"100100101",
  40390=>"000000000",
  40391=>"001000000",
  40392=>"000000000",
  40393=>"011011111",
  40394=>"100101111",
  40395=>"111000000",
  40396=>"000000000",
  40397=>"100111111",
  40398=>"000000000",
  40399=>"000000111",
  40400=>"111000000",
  40401=>"100100000",
  40402=>"000100111",
  40403=>"111111110",
  40404=>"000000000",
  40405=>"000001001",
  40406=>"101111111",
  40407=>"000010011",
  40408=>"100000000",
  40409=>"000111111",
  40410=>"110111111",
  40411=>"111000000",
  40412=>"011011111",
  40413=>"000000100",
  40414=>"011011111",
  40415=>"000000000",
  40416=>"001000000",
  40417=>"000100001",
  40418=>"111111111",
  40419=>"000000111",
  40420=>"111111011",
  40421=>"111010000",
  40422=>"111111111",
  40423=>"000000000",
  40424=>"000000000",
  40425=>"111111111",
  40426=>"111010000",
  40427=>"000000000",
  40428=>"000100100",
  40429=>"000010000",
  40430=>"000111111",
  40431=>"010111111",
  40432=>"100000000",
  40433=>"000111111",
  40434=>"100111111",
  40435=>"001001110",
  40436=>"110111110",
  40437=>"010111111",
  40438=>"111111110",
  40439=>"000000000",
  40440=>"000000100",
  40441=>"001001001",
  40442=>"000000000",
  40443=>"010000100",
  40444=>"000111111",
  40445=>"111111111",
  40446=>"111111111",
  40447=>"111111000",
  40448=>"011011011",
  40449=>"000000011",
  40450=>"111010000",
  40451=>"011111111",
  40452=>"011011011",
  40453=>"111100110",
  40454=>"111111111",
  40455=>"111111111",
  40456=>"001000000",
  40457=>"000100100",
  40458=>"101000000",
  40459=>"001011011",
  40460=>"111110100",
  40461=>"011111111",
  40462=>"101111111",
  40463=>"111000100",
  40464=>"110000000",
  40465=>"011111111",
  40466=>"000000110",
  40467=>"001111111",
  40468=>"000110111",
  40469=>"001011111",
  40470=>"110111111",
  40471=>"111110110",
  40472=>"100000000",
  40473=>"000000000",
  40474=>"111000000",
  40475=>"100000001",
  40476=>"000000000",
  40477=>"000000100",
  40478=>"101111111",
  40479=>"000000111",
  40480=>"000000000",
  40481=>"110111110",
  40482=>"010000000",
  40483=>"111111011",
  40484=>"000000100",
  40485=>"111111001",
  40486=>"000010111",
  40487=>"111001000",
  40488=>"111111100",
  40489=>"000000110",
  40490=>"111101111",
  40491=>"000000000",
  40492=>"000000000",
  40493=>"111111101",
  40494=>"000110110",
  40495=>"111110111",
  40496=>"111111111",
  40497=>"000000000",
  40498=>"111100000",
  40499=>"100000000",
  40500=>"000000000",
  40501=>"000100111",
  40502=>"110110000",
  40503=>"111111000",
  40504=>"001001111",
  40505=>"110111110",
  40506=>"001000000",
  40507=>"000000000",
  40508=>"000000000",
  40509=>"100100110",
  40510=>"111001000",
  40511=>"001000000",
  40512=>"111111011",
  40513=>"000111111",
  40514=>"111111100",
  40515=>"111011011",
  40516=>"000001000",
  40517=>"001001101",
  40518=>"000001000",
  40519=>"000000100",
  40520=>"001001001",
  40521=>"000000111",
  40522=>"100000111",
  40523=>"000000000",
  40524=>"110000000",
  40525=>"001111100",
  40526=>"000000000",
  40527=>"001000000",
  40528=>"111100110",
  40529=>"100110110",
  40530=>"000000000",
  40531=>"111111000",
  40532=>"001001001",
  40533=>"111111000",
  40534=>"001000001",
  40535=>"000000000",
  40536=>"111111001",
  40537=>"000011111",
  40538=>"110010010",
  40539=>"100011011",
  40540=>"000000000",
  40541=>"000000000",
  40542=>"000000111",
  40543=>"110100000",
  40544=>"000000000",
  40545=>"001000000",
  40546=>"000101111",
  40547=>"000000000",
  40548=>"100000011",
  40549=>"011011001",
  40550=>"000110011",
  40551=>"000000001",
  40552=>"110110111",
  40553=>"010000000",
  40554=>"111111111",
  40555=>"111000001",
  40556=>"010000111",
  40557=>"000000100",
  40558=>"000000111",
  40559=>"111001001",
  40560=>"110110111",
  40561=>"000010000",
  40562=>"011011100",
  40563=>"100100100",
  40564=>"111111111",
  40565=>"111111111",
  40566=>"111111111",
  40567=>"101111001",
  40568=>"000000011",
  40569=>"000000000",
  40570=>"000000000",
  40571=>"101000001",
  40572=>"001001001",
  40573=>"000000000",
  40574=>"111001000",
  40575=>"011111111",
  40576=>"000100000",
  40577=>"111001001",
  40578=>"000000000",
  40579=>"100110111",
  40580=>"000000000",
  40581=>"110110000",
  40582=>"000011110",
  40583=>"000000000",
  40584=>"000000000",
  40585=>"000000101",
  40586=>"000000000",
  40587=>"111000001",
  40588=>"000110000",
  40589=>"000000000",
  40590=>"100000000",
  40591=>"101110111",
  40592=>"111111011",
  40593=>"111111111",
  40594=>"000000000",
  40595=>"111001001",
  40596=>"000010110",
  40597=>"100100001",
  40598=>"111111111",
  40599=>"110111110",
  40600=>"000000101",
  40601=>"111010110",
  40602=>"000111111",
  40603=>"111111111",
  40604=>"110111110",
  40605=>"111111000",
  40606=>"111110110",
  40607=>"111101000",
  40608=>"111111111",
  40609=>"000000000",
  40610=>"001000000",
  40611=>"111111101",
  40612=>"011011011",
  40613=>"111101100",
  40614=>"110110000",
  40615=>"000000001",
  40616=>"111000000",
  40617=>"100010010",
  40618=>"001010001",
  40619=>"001001001",
  40620=>"000000000",
  40621=>"000100111",
  40622=>"000010111",
  40623=>"000000000",
  40624=>"111111000",
  40625=>"001000100",
  40626=>"000100000",
  40627=>"000000000",
  40628=>"000000100",
  40629=>"100000000",
  40630=>"111111000",
  40631=>"111111001",
  40632=>"100110000",
  40633=>"000000001",
  40634=>"111000011",
  40635=>"000000111",
  40636=>"111111111",
  40637=>"000000001",
  40638=>"000000000",
  40639=>"000000000",
  40640=>"000000000",
  40641=>"000000000",
  40642=>"000000000",
  40643=>"000000000",
  40644=>"001001111",
  40645=>"000000000",
  40646=>"001001000",
  40647=>"000000001",
  40648=>"010011111",
  40649=>"111111111",
  40650=>"001101000",
  40651=>"000000001",
  40652=>"010010111",
  40653=>"101101001",
  40654=>"010110111",
  40655=>"100000111",
  40656=>"000110110",
  40657=>"110100000",
  40658=>"000000000",
  40659=>"111111101",
  40660=>"000100100",
  40661=>"000000000",
  40662=>"000010000",
  40663=>"000001111",
  40664=>"000010011",
  40665=>"111010010",
  40666=>"011011111",
  40667=>"001000000",
  40668=>"010111111",
  40669=>"000000000",
  40670=>"111111111",
  40671=>"111110100",
  40672=>"111111111",
  40673=>"110111111",
  40674=>"000000000",
  40675=>"111111000",
  40676=>"111111111",
  40677=>"101111110",
  40678=>"111111111",
  40679=>"001000000",
  40680=>"111111111",
  40681=>"111111111",
  40682=>"100111001",
  40683=>"001000100",
  40684=>"110110011",
  40685=>"000010011",
  40686=>"000000101",
  40687=>"111000000",
  40688=>"111111111",
  40689=>"000000001",
  40690=>"011011011",
  40691=>"000011111",
  40692=>"111111111",
  40693=>"001000000",
  40694=>"110110111",
  40695=>"111111000",
  40696=>"000000000",
  40697=>"000000000",
  40698=>"100000111",
  40699=>"000000100",
  40700=>"110111111",
  40701=>"111000000",
  40702=>"111111111",
  40703=>"111111111",
  40704=>"001000010",
  40705=>"111111111",
  40706=>"000000000",
  40707=>"100001001",
  40708=>"111111111",
  40709=>"100100000",
  40710=>"000000000",
  40711=>"111110111",
  40712=>"111001111",
  40713=>"000000000",
  40714=>"111000100",
  40715=>"110100000",
  40716=>"000110100",
  40717=>"110111111",
  40718=>"000000000",
  40719=>"110111111",
  40720=>"111111111",
  40721=>"000000011",
  40722=>"000110111",
  40723=>"100000000",
  40724=>"111111000",
  40725=>"000000000",
  40726=>"110110110",
  40727=>"000001001",
  40728=>"011111001",
  40729=>"000110111",
  40730=>"000000000",
  40731=>"111111011",
  40732=>"111111011",
  40733=>"000000000",
  40734=>"000000000",
  40735=>"111111010",
  40736=>"000000101",
  40737=>"000000000",
  40738=>"111100001",
  40739=>"000100100",
  40740=>"001011001",
  40741=>"000110100",
  40742=>"000000000",
  40743=>"000000000",
  40744=>"000000001",
  40745=>"001110111",
  40746=>"000000000",
  40747=>"011011001",
  40748=>"100000000",
  40749=>"000000111",
  40750=>"010000000",
  40751=>"000000111",
  40752=>"111111011",
  40753=>"111000000",
  40754=>"001000000",
  40755=>"110111111",
  40756=>"000000000",
  40757=>"000000000",
  40758=>"100000001",
  40759=>"011111111",
  40760=>"000000000",
  40761=>"100000100",
  40762=>"100000110",
  40763=>"011000000",
  40764=>"111111111",
  40765=>"000001111",
  40766=>"111111111",
  40767=>"000111111",
  40768=>"000000110",
  40769=>"000000000",
  40770=>"111110000",
  40771=>"000000010",
  40772=>"010000000",
  40773=>"111001000",
  40774=>"011011111",
  40775=>"000000000",
  40776=>"111010011",
  40777=>"111111111",
  40778=>"001001000",
  40779=>"111110000",
  40780=>"110000000",
  40781=>"010011111",
  40782=>"001001001",
  40783=>"001111111",
  40784=>"001100111",
  40785=>"111111111",
  40786=>"111111111",
  40787=>"111111000",
  40788=>"111111111",
  40789=>"010010111",
  40790=>"000000010",
  40791=>"111100000",
  40792=>"101111111",
  40793=>"110100000",
  40794=>"000000000",
  40795=>"011110110",
  40796=>"111111011",
  40797=>"111111011",
  40798=>"000000000",
  40799=>"000000000",
  40800=>"000000010",
  40801=>"000000000",
  40802=>"000010010",
  40803=>"011111111",
  40804=>"111110010",
  40805=>"000110010",
  40806=>"111111111",
  40807=>"000000001",
  40808=>"111100111",
  40809=>"110110010",
  40810=>"111001111",
  40811=>"011111000",
  40812=>"111110111",
  40813=>"110100101",
  40814=>"111111111",
  40815=>"111111010",
  40816=>"111111111",
  40817=>"111111111",
  40818=>"000000000",
  40819=>"111111011",
  40820=>"101000001",
  40821=>"111111110",
  40822=>"111111000",
  40823=>"111111111",
  40824=>"000000001",
  40825=>"111000000",
  40826=>"000000000",
  40827=>"100000000",
  40828=>"000000000",
  40829=>"000000000",
  40830=>"000000111",
  40831=>"111111111",
  40832=>"111000000",
  40833=>"000000000",
  40834=>"110111111",
  40835=>"001001001",
  40836=>"111111111",
  40837=>"110110110",
  40838=>"111111111",
  40839=>"100001011",
  40840=>"000000110",
  40841=>"111001011",
  40842=>"101001001",
  40843=>"000000000",
  40844=>"000011111",
  40845=>"100100101",
  40846=>"111111111",
  40847=>"000000001",
  40848=>"100110111",
  40849=>"110000100",
  40850=>"100110110",
  40851=>"111111111",
  40852=>"101101111",
  40853=>"001100110",
  40854=>"111111111",
  40855=>"000000111",
  40856=>"000000001",
  40857=>"100110111",
  40858=>"111000000",
  40859=>"100000111",
  40860=>"111111111",
  40861=>"000001010",
  40862=>"011011011",
  40863=>"000000111",
  40864=>"111011011",
  40865=>"000111111",
  40866=>"110111111",
  40867=>"011000001",
  40868=>"101110110",
  40869=>"111110000",
  40870=>"000000000",
  40871=>"000111111",
  40872=>"000000000",
  40873=>"000100111",
  40874=>"111100100",
  40875=>"000000000",
  40876=>"000000000",
  40877=>"000110111",
  40878=>"111000000",
  40879=>"000000001",
  40880=>"000000000",
  40881=>"111111111",
  40882=>"000000111",
  40883=>"111011111",
  40884=>"110111111",
  40885=>"000001110",
  40886=>"110101111",
  40887=>"011111111",
  40888=>"000000011",
  40889=>"111111101",
  40890=>"000001011",
  40891=>"100000000",
  40892=>"000000000",
  40893=>"111000100",
  40894=>"000000001",
  40895=>"100010011",
  40896=>"111111111",
  40897=>"000110110",
  40898=>"100110110",
  40899=>"000000000",
  40900=>"111101111",
  40901=>"011111111",
  40902=>"011111111",
  40903=>"000000000",
  40904=>"000000101",
  40905=>"110000001",
  40906=>"000000000",
  40907=>"100010111",
  40908=>"000111111",
  40909=>"010000000",
  40910=>"000000100",
  40911=>"010000000",
  40912=>"110000111",
  40913=>"000001001",
  40914=>"111111111",
  40915=>"111111111",
  40916=>"111111111",
  40917=>"111111100",
  40918=>"111111111",
  40919=>"100001001",
  40920=>"100111011",
  40921=>"111111111",
  40922=>"111011111",
  40923=>"111000010",
  40924=>"101000000",
  40925=>"110111110",
  40926=>"011001000",
  40927=>"111101111",
  40928=>"111111110",
  40929=>"000001001",
  40930=>"111111111",
  40931=>"111111111",
  40932=>"000000111",
  40933=>"111111111",
  40934=>"101111111",
  40935=>"111111111",
  40936=>"010010111",
  40937=>"111111000",
  40938=>"111011000",
  40939=>"000000100",
  40940=>"000111111",
  40941=>"000000001",
  40942=>"001001000",
  40943=>"000111111",
  40944=>"000011001",
  40945=>"000011011",
  40946=>"111111111",
  40947=>"111000110",
  40948=>"011111001",
  40949=>"001011010",
  40950=>"011011011",
  40951=>"000000001",
  40952=>"000111111",
  40953=>"000000000",
  40954=>"111110100",
  40955=>"000000000",
  40956=>"000000001",
  40957=>"110110111",
  40958=>"000111111",
  40959=>"111111111",
  40960=>"001001001",
  40961=>"001000000",
  40962=>"111111111",
  40963=>"000000000",
  40964=>"111011011",
  40965=>"000100100",
  40966=>"010000000",
  40967=>"111111111",
  40968=>"111001000",
  40969=>"000000111",
  40970=>"101011111",
  40971=>"000000001",
  40972=>"110110001",
  40973=>"100111111",
  40974=>"010001111",
  40975=>"110111000",
  40976=>"011111111",
  40977=>"111011111",
  40978=>"000000000",
  40979=>"111111111",
  40980=>"111111111",
  40981=>"010111111",
  40982=>"111111000",
  40983=>"000100111",
  40984=>"000101111",
  40985=>"100110111",
  40986=>"001000000",
  40987=>"010000000",
  40988=>"101100000",
  40989=>"111001001",
  40990=>"101000000",
  40991=>"110111001",
  40992=>"000000000",
  40993=>"110010000",
  40994=>"100110110",
  40995=>"000111110",
  40996=>"000000000",
  40997=>"111111000",
  40998=>"001111111",
  40999=>"000011111",
  41000=>"001011111",
  41001=>"000000000",
  41002=>"000000001",
  41003=>"111111111",
  41004=>"111111001",
  41005=>"111111010",
  41006=>"000000001",
  41007=>"110110000",
  41008=>"000000000",
  41009=>"000000000",
  41010=>"001111110",
  41011=>"000010111",
  41012=>"001000000",
  41013=>"100101001",
  41014=>"000000101",
  41015=>"111011001",
  41016=>"111111111",
  41017=>"000100000",
  41018=>"000000000",
  41019=>"000000111",
  41020=>"101000000",
  41021=>"100111111",
  41022=>"111111000",
  41023=>"000001111",
  41024=>"000001001",
  41025=>"011001000",
  41026=>"111011110",
  41027=>"110010000",
  41028=>"111101001",
  41029=>"110111111",
  41030=>"000000100",
  41031=>"111111111",
  41032=>"001000000",
  41033=>"000000000",
  41034=>"111111001",
  41035=>"111000000",
  41036=>"110111111",
  41037=>"100000000",
  41038=>"110111111",
  41039=>"111111101",
  41040=>"000101100",
  41041=>"111001000",
  41042=>"111111000",
  41043=>"111011001",
  41044=>"111111101",
  41045=>"111111010",
  41046=>"000000000",
  41047=>"111111001",
  41048=>"111110100",
  41049=>"100000111",
  41050=>"000000010",
  41051=>"100000000",
  41052=>"001000111",
  41053=>"000011000",
  41054=>"111000010",
  41055=>"001111111",
  41056=>"000000111",
  41057=>"101000000",
  41058=>"011111111",
  41059=>"101101101",
  41060=>"111111000",
  41061=>"111111111",
  41062=>"000111111",
  41063=>"111111111",
  41064=>"000000111",
  41065=>"001000000",
  41066=>"111111111",
  41067=>"110111110",
  41068=>"111111001",
  41069=>"000000000",
  41070=>"111110111",
  41071=>"111111111",
  41072=>"111111111",
  41073=>"000000011",
  41074=>"000110111",
  41075=>"111111111",
  41076=>"000000000",
  41077=>"000000110",
  41078=>"000000111",
  41079=>"111011111",
  41080=>"111011000",
  41081=>"100000000",
  41082=>"000011111",
  41083=>"111110111",
  41084=>"001101101",
  41085=>"111111111",
  41086=>"111111000",
  41087=>"011000000",
  41088=>"110110111",
  41089=>"111111111",
  41090=>"000101111",
  41091=>"001000000",
  41092=>"000001011",
  41093=>"011011101",
  41094=>"000000000",
  41095=>"000110111",
  41096=>"111111010",
  41097=>"000111100",
  41098=>"001111111",
  41099=>"101111011",
  41100=>"000000111",
  41101=>"000000000",
  41102=>"000000000",
  41103=>"000000000",
  41104=>"001000000",
  41105=>"011000001",
  41106=>"111111111",
  41107=>"011001001",
  41108=>"100000000",
  41109=>"101101111",
  41110=>"011111111",
  41111=>"111001111",
  41112=>"001000111",
  41113=>"001111111",
  41114=>"000000000",
  41115=>"000000000",
  41116=>"111111111",
  41117=>"111001101",
  41118=>"101101111",
  41119=>"000000000",
  41120=>"000000000",
  41121=>"000111111",
  41122=>"000111111",
  41123=>"001000000",
  41124=>"000000111",
  41125=>"111111111",
  41126=>"111000000",
  41127=>"100110111",
  41128=>"111111111",
  41129=>"111000000",
  41130=>"111111000",
  41131=>"001111111",
  41132=>"000000000",
  41133=>"110110110",
  41134=>"011000000",
  41135=>"100100100",
  41136=>"000000000",
  41137=>"100100110",
  41138=>"111111111",
  41139=>"111000000",
  41140=>"000000000",
  41141=>"111000001",
  41142=>"000001111",
  41143=>"000000100",
  41144=>"111011000",
  41145=>"111111111",
  41146=>"000001000",
  41147=>"101111111",
  41148=>"111101110",
  41149=>"110111000",
  41150=>"000000111",
  41151=>"000000000",
  41152=>"100100100",
  41153=>"010100111",
  41154=>"111111111",
  41155=>"100000000",
  41156=>"111110110",
  41157=>"000000000",
  41158=>"001011101",
  41159=>"000001000",
  41160=>"111001001",
  41161=>"100100011",
  41162=>"000110111",
  41163=>"000000000",
  41164=>"000000100",
  41165=>"100111111",
  41166=>"100000000",
  41167=>"000010011",
  41168=>"000000000",
  41169=>"000110111",
  41170=>"100000111",
  41171=>"000000000",
  41172=>"000010111",
  41173=>"000000000",
  41174=>"000001111",
  41175=>"111111111",
  41176=>"000000100",
  41177=>"111111100",
  41178=>"111100000",
  41179=>"100100000",
  41180=>"111110100",
  41181=>"000000111",
  41182=>"011000000",
  41183=>"111111111",
  41184=>"111101001",
  41185=>"011001000",
  41186=>"111111011",
  41187=>"000110011",
  41188=>"000000000",
  41189=>"000010000",
  41190=>"010010111",
  41191=>"111111110",
  41192=>"011000000",
  41193=>"111000011",
  41194=>"000000111",
  41195=>"111011011",
  41196=>"000000000",
  41197=>"000011111",
  41198=>"101111111",
  41199=>"011111001",
  41200=>"011000110",
  41201=>"001000110",
  41202=>"000111111",
  41203=>"001001000",
  41204=>"001001111",
  41205=>"111111111",
  41206=>"000111111",
  41207=>"111111000",
  41208=>"011111111",
  41209=>"100000000",
  41210=>"111111001",
  41211=>"111111111",
  41212=>"101001001",
  41213=>"011011111",
  41214=>"000000000",
  41215=>"001011111",
  41216=>"111111010",
  41217=>"011011001",
  41218=>"111111100",
  41219=>"011110111",
  41220=>"000001000",
  41221=>"110111111",
  41222=>"111111111",
  41223=>"000000000",
  41224=>"111111000",
  41225=>"000000111",
  41226=>"111000000",
  41227=>"110110000",
  41228=>"111101111",
  41229=>"111000000",
  41230=>"101100001",
  41231=>"111110000",
  41232=>"000000000",
  41233=>"101100111",
  41234=>"100111111",
  41235=>"111111111",
  41236=>"011111111",
  41237=>"011001000",
  41238=>"001001000",
  41239=>"110000000",
  41240=>"001000000",
  41241=>"011000000",
  41242=>"010010111",
  41243=>"010000000",
  41244=>"111010000",
  41245=>"111111001",
  41246=>"000000000",
  41247=>"111111111",
  41248=>"111111111",
  41249=>"001000000",
  41250=>"000000000",
  41251=>"111111100",
  41252=>"111111100",
  41253=>"011000111",
  41254=>"000111011",
  41255=>"111000000",
  41256=>"000111111",
  41257=>"000000001",
  41258=>"010110010",
  41259=>"000011111",
  41260=>"111111011",
  41261=>"101111111",
  41262=>"000000101",
  41263=>"110000000",
  41264=>"000001100",
  41265=>"000101101",
  41266=>"000000001",
  41267=>"111111111",
  41268=>"000100111",
  41269=>"001000000",
  41270=>"100100000",
  41271=>"000000000",
  41272=>"000010010",
  41273=>"111111000",
  41274=>"110000010",
  41275=>"000000011",
  41276=>"111111000",
  41277=>"000000111",
  41278=>"101101001",
  41279=>"111111111",
  41280=>"111111000",
  41281=>"000000000",
  41282=>"001000000",
  41283=>"000111111",
  41284=>"111111111",
  41285=>"000111111",
  41286=>"010111111",
  41287=>"000000111",
  41288=>"111001000",
  41289=>"111000000",
  41290=>"000000000",
  41291=>"111100100",
  41292=>"000000100",
  41293=>"000000000",
  41294=>"001100100",
  41295=>"111111111",
  41296=>"000001111",
  41297=>"000000000",
  41298=>"000000000",
  41299=>"100110111",
  41300=>"010000000",
  41301=>"000011000",
  41302=>"111111101",
  41303=>"000111111",
  41304=>"010110010",
  41305=>"000000000",
  41306=>"100000000",
  41307=>"110000000",
  41308=>"000000000",
  41309=>"100111101",
  41310=>"011111111",
  41311=>"000000000",
  41312=>"111111111",
  41313=>"101001101",
  41314=>"110100000",
  41315=>"000001000",
  41316=>"111111110",
  41317=>"111101000",
  41318=>"000001000",
  41319=>"011000000",
  41320=>"111111110",
  41321=>"000000000",
  41322=>"000000010",
  41323=>"001000000",
  41324=>"110110100",
  41325=>"001001000",
  41326=>"000000000",
  41327=>"111111101",
  41328=>"000000100",
  41329=>"011011111",
  41330=>"111010000",
  41331=>"110100000",
  41332=>"111110000",
  41333=>"111011101",
  41334=>"001101001",
  41335=>"110000000",
  41336=>"000111111",
  41337=>"001111011",
  41338=>"000111111",
  41339=>"000000000",
  41340=>"000000000",
  41341=>"001100111",
  41342=>"000000000",
  41343=>"000111111",
  41344=>"100000000",
  41345=>"000000000",
  41346=>"000111111",
  41347=>"000000000",
  41348=>"000000000",
  41349=>"110111111",
  41350=>"000000000",
  41351=>"011011111",
  41352=>"100111111",
  41353=>"100000001",
  41354=>"110110110",
  41355=>"000111111",
  41356=>"101111111",
  41357=>"100110110",
  41358=>"001010110",
  41359=>"111111111",
  41360=>"001000000",
  41361=>"100111111",
  41362=>"000111111",
  41363=>"001011111",
  41364=>"011011010",
  41365=>"000000000",
  41366=>"011011000",
  41367=>"001001000",
  41368=>"000000001",
  41369=>"011000001",
  41370=>"000111111",
  41371=>"111111111",
  41372=>"111111111",
  41373=>"000000011",
  41374=>"001000000",
  41375=>"101111000",
  41376=>"000000000",
  41377=>"111111111",
  41378=>"111111010",
  41379=>"011000000",
  41380=>"000000011",
  41381=>"111010000",
  41382=>"001000000",
  41383=>"101000100",
  41384=>"101000000",
  41385=>"111111100",
  41386=>"001111111",
  41387=>"111111011",
  41388=>"010000000",
  41389=>"011111101",
  41390=>"100000000",
  41391=>"000001011",
  41392=>"000000000",
  41393=>"000000000",
  41394=>"111111111",
  41395=>"000000000",
  41396=>"111111111",
  41397=>"000111111",
  41398=>"111111111",
  41399=>"111010000",
  41400=>"001111111",
  41401=>"000000111",
  41402=>"000000001",
  41403=>"001111111",
  41404=>"000000011",
  41405=>"111111010",
  41406=>"111111111",
  41407=>"000100111",
  41408=>"111111111",
  41409=>"001011011",
  41410=>"111111010",
  41411=>"000000000",
  41412=>"000000000",
  41413=>"001001000",
  41414=>"000111111",
  41415=>"000000000",
  41416=>"001111111",
  41417=>"000101111",
  41418=>"000000000",
  41419=>"000000000",
  41420=>"000000000",
  41421=>"111111111",
  41422=>"000101101",
  41423=>"000000101",
  41424=>"111000101",
  41425=>"000000000",
  41426=>"111111111",
  41427=>"111001001",
  41428=>"111111001",
  41429=>"000000111",
  41430=>"100100000",
  41431=>"111111011",
  41432=>"000000000",
  41433=>"111001001",
  41434=>"000000111",
  41435=>"111111111",
  41436=>"000000000",
  41437=>"000000000",
  41438=>"111111111",
  41439=>"111111111",
  41440=>"001000011",
  41441=>"000000000",
  41442=>"000111111",
  41443=>"001000000",
  41444=>"111111111",
  41445=>"000000000",
  41446=>"001111111",
  41447=>"000000001",
  41448=>"111111110",
  41449=>"110000000",
  41450=>"111111111",
  41451=>"111111111",
  41452=>"001000000",
  41453=>"000000000",
  41454=>"000111111",
  41455=>"011000000",
  41456=>"101100000",
  41457=>"100111111",
  41458=>"111111111",
  41459=>"110000000",
  41460=>"000000000",
  41461=>"000000100",
  41462=>"111111001",
  41463=>"111111000",
  41464=>"000000000",
  41465=>"000000000",
  41466=>"000001111",
  41467=>"011111000",
  41468=>"000111111",
  41469=>"000000001",
  41470=>"101000000",
  41471=>"001000000",
  41472=>"110000110",
  41473=>"000110111",
  41474=>"000000110",
  41475=>"000000000",
  41476=>"111100100",
  41477=>"001000000",
  41478=>"110110000",
  41479=>"000000000",
  41480=>"111000000",
  41481=>"001111001",
  41482=>"000000000",
  41483=>"100100110",
  41484=>"000000000",
  41485=>"011000000",
  41486=>"101001001",
  41487=>"000000000",
  41488=>"110111001",
  41489=>"000011000",
  41490=>"001000000",
  41491=>"000100000",
  41492=>"000000000",
  41493=>"111111111",
  41494=>"110110111",
  41495=>"000000000",
  41496=>"110110000",
  41497=>"000000111",
  41498=>"111111000",
  41499=>"011010111",
  41500=>"000000001",
  41501=>"010010011",
  41502=>"000100100",
  41503=>"110000000",
  41504=>"000001001",
  41505=>"111111111",
  41506=>"111111011",
  41507=>"110111111",
  41508=>"111111111",
  41509=>"111110000",
  41510=>"101111111",
  41511=>"000100110",
  41512=>"111111111",
  41513=>"100000000",
  41514=>"011000000",
  41515=>"111111001",
  41516=>"111111110",
  41517=>"111111111",
  41518=>"001000000",
  41519=>"111000000",
  41520=>"000000000",
  41521=>"010001000",
  41522=>"111111111",
  41523=>"000001011",
  41524=>"000011011",
  41525=>"100010010",
  41526=>"111101111",
  41527=>"000000001",
  41528=>"111111111",
  41529=>"000000000",
  41530=>"000110110",
  41531=>"000000100",
  41532=>"000000000",
  41533=>"011011000",
  41534=>"111000100",
  41535=>"000000000",
  41536=>"001000111",
  41537=>"111111111",
  41538=>"111111111",
  41539=>"110111111",
  41540=>"001001000",
  41541=>"111111000",
  41542=>"110000110",
  41543=>"111111111",
  41544=>"001001111",
  41545=>"000000000",
  41546=>"000000000",
  41547=>"000000100",
  41548=>"111111110",
  41549=>"111111000",
  41550=>"100110111",
  41551=>"111001001",
  41552=>"000111111",
  41553=>"110111111",
  41554=>"100000111",
  41555=>"111111111",
  41556=>"000000000",
  41557=>"100000000",
  41558=>"011111101",
  41559=>"000000000",
  41560=>"011000000",
  41561=>"001101111",
  41562=>"111111001",
  41563=>"111000000",
  41564=>"111111111",
  41565=>"111111000",
  41566=>"111111000",
  41567=>"000000000",
  41568=>"000111111",
  41569=>"000001011",
  41570=>"000000111",
  41571=>"111001001",
  41572=>"000000000",
  41573=>"000000101",
  41574=>"011111111",
  41575=>"100100111",
  41576=>"000000000",
  41577=>"000100111",
  41578=>"000110111",
  41579=>"111111011",
  41580=>"100000011",
  41581=>"110111101",
  41582=>"111111111",
  41583=>"000000000",
  41584=>"011011111",
  41585=>"000001000",
  41586=>"101001000",
  41587=>"010000000",
  41588=>"000000000",
  41589=>"100100100",
  41590=>"011001000",
  41591=>"010000110",
  41592=>"011111111",
  41593=>"001000000",
  41594=>"110110111",
  41595=>"000000000",
  41596=>"001011011",
  41597=>"110111111",
  41598=>"110110101",
  41599=>"011111111",
  41600=>"000000001",
  41601=>"110111111",
  41602=>"001011111",
  41603=>"011011011",
  41604=>"100011000",
  41605=>"000000000",
  41606=>"010111111",
  41607=>"000000010",
  41608=>"111111100",
  41609=>"011000001",
  41610=>"111111111",
  41611=>"111111101",
  41612=>"000101111",
  41613=>"111111111",
  41614=>"000011110",
  41615=>"000100100",
  41616=>"111111111",
  41617=>"000000000",
  41618=>"001111000",
  41619=>"111111111",
  41620=>"000000110",
  41621=>"111100100",
  41622=>"110111111",
  41623=>"000000111",
  41624=>"000000111",
  41625=>"111110111",
  41626=>"110000000",
  41627=>"000000000",
  41628=>"000000001",
  41629=>"001000000",
  41630=>"000111001",
  41631=>"110111101",
  41632=>"101101111",
  41633=>"000000001",
  41634=>"000000000",
  41635=>"000000001",
  41636=>"101101111",
  41637=>"000001111",
  41638=>"111011011",
  41639=>"111111001",
  41640=>"111000000",
  41641=>"100100100",
  41642=>"111000000",
  41643=>"111111111",
  41644=>"010011111",
  41645=>"000000000",
  41646=>"111111111",
  41647=>"000000011",
  41648=>"000000111",
  41649=>"001000001",
  41650=>"010000010",
  41651=>"100110111",
  41652=>"110100101",
  41653=>"000000000",
  41654=>"111010010",
  41655=>"100001111",
  41656=>"110011011",
  41657=>"111111111",
  41658=>"110100000",
  41659=>"111111111",
  41660=>"111111111",
  41661=>"110110000",
  41662=>"111100111",
  41663=>"111111111",
  41664=>"000000000",
  41665=>"100000100",
  41666=>"000000000",
  41667=>"000000000",
  41668=>"111111111",
  41669=>"000000000",
  41670=>"000001001",
  41671=>"000000000",
  41672=>"111110111",
  41673=>"000000100",
  41674=>"001111111",
  41675=>"000000000",
  41676=>"000111111",
  41677=>"011111111",
  41678=>"010111111",
  41679=>"111111111",
  41680=>"111111000",
  41681=>"010000111",
  41682=>"110100111",
  41683=>"110110000",
  41684=>"001001000",
  41685=>"011011011",
  41686=>"111001001",
  41687=>"001000001",
  41688=>"000000000",
  41689=>"111111111",
  41690=>"101100000",
  41691=>"000000000",
  41692=>"010000000",
  41693=>"000000000",
  41694=>"111111000",
  41695=>"111111001",
  41696=>"011111111",
  41697=>"000000000",
  41698=>"010011000",
  41699=>"111111000",
  41700=>"000001001",
  41701=>"101011011",
  41702=>"000000000",
  41703=>"111111001",
  41704=>"111111000",
  41705=>"111001000",
  41706=>"001111111",
  41707=>"111111001",
  41708=>"111111011",
  41709=>"111111111",
  41710=>"110010010",
  41711=>"000001111",
  41712=>"010000111",
  41713=>"100000000",
  41714=>"111111111",
  41715=>"111111110",
  41716=>"000000000",
  41717=>"111111011",
  41718=>"000010000",
  41719=>"000000000",
  41720=>"000000111",
  41721=>"000000000",
  41722=>"000000000",
  41723=>"111111011",
  41724=>"111111111",
  41725=>"000000001",
  41726=>"000000000",
  41727=>"100001000",
  41728=>"000000000",
  41729=>"111111000",
  41730=>"111111111",
  41731=>"000000000",
  41732=>"000101111",
  41733=>"000100000",
  41734=>"000000000",
  41735=>"000000000",
  41736=>"000000100",
  41737=>"110110010",
  41738=>"100111111",
  41739=>"011011001",
  41740=>"111001001",
  41741=>"001011111",
  41742=>"000000000",
  41743=>"000100000",
  41744=>"000001000",
  41745=>"011000000",
  41746=>"000000000",
  41747=>"000110000",
  41748=>"010011101",
  41749=>"010000110",
  41750=>"000001001",
  41751=>"111001000",
  41752=>"110111111",
  41753=>"101100000",
  41754=>"111001000",
  41755=>"000000000",
  41756=>"111011011",
  41757=>"111000000",
  41758=>"111111111",
  41759=>"000000000",
  41760=>"001000000",
  41761=>"000001111",
  41762=>"100000000",
  41763=>"111111111",
  41764=>"000000100",
  41765=>"111111111",
  41766=>"000000000",
  41767=>"011000000",
  41768=>"000100100",
  41769=>"111111011",
  41770=>"001000000",
  41771=>"111111000",
  41772=>"100000000",
  41773=>"010110000",
  41774=>"000001001",
  41775=>"000001001",
  41776=>"000111111",
  41777=>"000001000",
  41778=>"000000000",
  41779=>"110100110",
  41780=>"011000000",
  41781=>"110111111",
  41782=>"000000000",
  41783=>"010000111",
  41784=>"000000000",
  41785=>"001111111",
  41786=>"100110100",
  41787=>"111000000",
  41788=>"001001000",
  41789=>"110110110",
  41790=>"000000110",
  41791=>"000000111",
  41792=>"000000000",
  41793=>"111111111",
  41794=>"000000000",
  41795=>"000000000",
  41796=>"011001011",
  41797=>"111101000",
  41798=>"100000000",
  41799=>"111000001",
  41800=>"000000000",
  41801=>"000000000",
  41802=>"111111111",
  41803=>"111111111",
  41804=>"000000000",
  41805=>"111110111",
  41806=>"110111111",
  41807=>"011001001",
  41808=>"111111000",
  41809=>"100000000",
  41810=>"010111111",
  41811=>"000000100",
  41812=>"111111111",
  41813=>"010000000",
  41814=>"101100100",
  41815=>"111111111",
  41816=>"111110111",
  41817=>"000000111",
  41818=>"011011010",
  41819=>"110100101",
  41820=>"111111111",
  41821=>"000000110",
  41822=>"100000000",
  41823=>"100000000",
  41824=>"100111001",
  41825=>"011000000",
  41826=>"000001000",
  41827=>"000000001",
  41828=>"110000000",
  41829=>"000000000",
  41830=>"011000000",
  41831=>"000000111",
  41832=>"011101001",
  41833=>"000000000",
  41834=>"111111111",
  41835=>"001001011",
  41836=>"001010110",
  41837=>"110111111",
  41838=>"111111111",
  41839=>"000010000",
  41840=>"110000111",
  41841=>"111111000",
  41842=>"111111011",
  41843=>"001000000",
  41844=>"111111111",
  41845=>"110111001",
  41846=>"100000000",
  41847=>"000000000",
  41848=>"111111111",
  41849=>"000000000",
  41850=>"111101100",
  41851=>"000011001",
  41852=>"000000110",
  41853=>"011001000",
  41854=>"100111111",
  41855=>"000000111",
  41856=>"111111110",
  41857=>"111111110",
  41858=>"111111111",
  41859=>"000100110",
  41860=>"111000101",
  41861=>"111111111",
  41862=>"111111111",
  41863=>"000110110",
  41864=>"111111110",
  41865=>"000000000",
  41866=>"110110011",
  41867=>"000000111",
  41868=>"011001001",
  41869=>"000000000",
  41870=>"000100000",
  41871=>"010010111",
  41872=>"111111111",
  41873=>"110000000",
  41874=>"111111111",
  41875=>"110100100",
  41876=>"111111111",
  41877=>"000110000",
  41878=>"000010000",
  41879=>"000000000",
  41880=>"110000001",
  41881=>"000011100",
  41882=>"111110111",
  41883=>"111111100",
  41884=>"100000000",
  41885=>"000011111",
  41886=>"001000000",
  41887=>"000000000",
  41888=>"111111100",
  41889=>"111111111",
  41890=>"000000001",
  41891=>"110100111",
  41892=>"111111100",
  41893=>"000111111",
  41894=>"000001111",
  41895=>"111001000",
  41896=>"100000001",
  41897=>"001001001",
  41898=>"110111100",
  41899=>"111001000",
  41900=>"000000110",
  41901=>"100000000",
  41902=>"000000000",
  41903=>"000000000",
  41904=>"100111111",
  41905=>"000000000",
  41906=>"000100111",
  41907=>"000000000",
  41908=>"110111111",
  41909=>"111111000",
  41910=>"001001111",
  41911=>"111000000",
  41912=>"000000000",
  41913=>"111011000",
  41914=>"010000000",
  41915=>"111110110",
  41916=>"011111000",
  41917=>"100100100",
  41918=>"111111111",
  41919=>"000000000",
  41920=>"111110111",
  41921=>"000000011",
  41922=>"111111111",
  41923=>"001001011",
  41924=>"111100100",
  41925=>"111111111",
  41926=>"001001111",
  41927=>"111011000",
  41928=>"000000000",
  41929=>"111000010",
  41930=>"010000000",
  41931=>"111111111",
  41932=>"000000000",
  41933=>"000000000",
  41934=>"000000000",
  41935=>"000000000",
  41936=>"000000000",
  41937=>"110111111",
  41938=>"000000000",
  41939=>"100000000",
  41940=>"100000000",
  41941=>"111001001",
  41942=>"000111111",
  41943=>"011011111",
  41944=>"000000100",
  41945=>"000111111",
  41946=>"000000100",
  41947=>"000000000",
  41948=>"100000001",
  41949=>"111111111",
  41950=>"001001011",
  41951=>"111001011",
  41952=>"111111111",
  41953=>"110101110",
  41954=>"100000000",
  41955=>"100000000",
  41956=>"000000000",
  41957=>"001001001",
  41958=>"000000000",
  41959=>"100100111",
  41960=>"111111111",
  41961=>"111111000",
  41962=>"101111111",
  41963=>"001001111",
  41964=>"101111111",
  41965=>"000000000",
  41966=>"111111111",
  41967=>"111000000",
  41968=>"111100100",
  41969=>"111111111",
  41970=>"111111111",
  41971=>"111011011",
  41972=>"110100100",
  41973=>"001000000",
  41974=>"111001000",
  41975=>"001001000",
  41976=>"001111000",
  41977=>"100100111",
  41978=>"000000000",
  41979=>"011000000",
  41980=>"001000000",
  41981=>"111110111",
  41982=>"111111111",
  41983=>"000000000",
  41984=>"111111110",
  41985=>"011001111",
  41986=>"001111000",
  41987=>"000100100",
  41988=>"100000000",
  41989=>"001000000",
  41990=>"110000000",
  41991=>"000000111",
  41992=>"111111100",
  41993=>"000000111",
  41994=>"111111111",
  41995=>"111111011",
  41996=>"000001011",
  41997=>"001001111",
  41998=>"100110111",
  41999=>"111111010",
  42000=>"111111110",
  42001=>"000000111",
  42002=>"000111101",
  42003=>"000001111",
  42004=>"111101101",
  42005=>"110110000",
  42006=>"000001111",
  42007=>"001001001",
  42008=>"000000100",
  42009=>"011111111",
  42010=>"111111100",
  42011=>"000000000",
  42012=>"011111110",
  42013=>"111110100",
  42014=>"000000000",
  42015=>"100000000",
  42016=>"100100000",
  42017=>"111111010",
  42018=>"001001111",
  42019=>"000000000",
  42020=>"111111111",
  42021=>"000110111",
  42022=>"000000010",
  42023=>"111111000",
  42024=>"000000000",
  42025=>"111010010",
  42026=>"111111111",
  42027=>"101111111",
  42028=>"111010000",
  42029=>"000001001",
  42030=>"111011110",
  42031=>"111111100",
  42032=>"000000000",
  42033=>"000000000",
  42034=>"000001000",
  42035=>"100101111",
  42036=>"111111100",
  42037=>"000000000",
  42038=>"111111111",
  42039=>"111111111",
  42040=>"000000000",
  42041=>"000011011",
  42042=>"110111111",
  42043=>"010011111",
  42044=>"000000111",
  42045=>"111111111",
  42046=>"110100100",
  42047=>"111111011",
  42048=>"111111000",
  42049=>"000000000",
  42050=>"111111011",
  42051=>"000000011",
  42052=>"110111111",
  42053=>"101000100",
  42054=>"000000000",
  42055=>"000000101",
  42056=>"111111011",
  42057=>"000000000",
  42058=>"110110110",
  42059=>"111111000",
  42060=>"000000000",
  42061=>"110111011",
  42062=>"000000101",
  42063=>"111001111",
  42064=>"000000000",
  42065=>"111111000",
  42066=>"110111110",
  42067=>"001000000",
  42068=>"111111110",
  42069=>"110010000",
  42070=>"100100000",
  42071=>"000000000",
  42072=>"110001001",
  42073=>"111111001",
  42074=>"101101111",
  42075=>"110110110",
  42076=>"000000001",
  42077=>"111111000",
  42078=>"001001101",
  42079=>"000110111",
  42080=>"111000000",
  42081=>"000000000",
  42082=>"111000000",
  42083=>"000000000",
  42084=>"100000000",
  42085=>"000000001",
  42086=>"001111111",
  42087=>"011000111",
  42088=>"010010000",
  42089=>"010010010",
  42090=>"000000010",
  42091=>"000000111",
  42092=>"111111000",
  42093=>"111111111",
  42094=>"101000000",
  42095=>"111111011",
  42096=>"000111111",
  42097=>"000000000",
  42098=>"111111111",
  42099=>"111001111",
  42100=>"111111000",
  42101=>"000111111",
  42102=>"000000000",
  42103=>"000000000",
  42104=>"000000000",
  42105=>"001111111",
  42106=>"001001011",
  42107=>"111111111",
  42108=>"110110110",
  42109=>"111111111",
  42110=>"000000000",
  42111=>"000000000",
  42112=>"111111000",
  42113=>"111111111",
  42114=>"111111011",
  42115=>"111110100",
  42116=>"001001111",
  42117=>"111110000",
  42118=>"101111101",
  42119=>"000000110",
  42120=>"111111111",
  42121=>"111000111",
  42122=>"111000000",
  42123=>"110111111",
  42124=>"000000000",
  42125=>"101000100",
  42126=>"010111111",
  42127=>"111111111",
  42128=>"111001001",
  42129=>"000000000",
  42130=>"111111011",
  42131=>"100000010",
  42132=>"111111000",
  42133=>"100000101",
  42134=>"010000100",
  42135=>"000000000",
  42136=>"000000000",
  42137=>"000000000",
  42138=>"111111000",
  42139=>"000000000",
  42140=>"111111111",
  42141=>"011111111",
  42142=>"111011001",
  42143=>"001001111",
  42144=>"111111111",
  42145=>"000000000",
  42146=>"000000000",
  42147=>"100101101",
  42148=>"000001001",
  42149=>"000000111",
  42150=>"111111111",
  42151=>"111111111",
  42152=>"000000000",
  42153=>"111111010",
  42154=>"111111100",
  42155=>"111111110",
  42156=>"000011111",
  42157=>"111110100",
  42158=>"111111111",
  42159=>"000000000",
  42160=>"000111011",
  42161=>"000001011",
  42162=>"111111111",
  42163=>"111111111",
  42164=>"000001100",
  42165=>"100111110",
  42166=>"110110000",
  42167=>"011001111",
  42168=>"000001000",
  42169=>"001001100",
  42170=>"000111101",
  42171=>"000001111",
  42172=>"010000101",
  42173=>"110110000",
  42174=>"111111110",
  42175=>"000111110",
  42176=>"000000000",
  42177=>"011000111",
  42178=>"000110000",
  42179=>"010110111",
  42180=>"111111100",
  42181=>"000111111",
  42182=>"100101111",
  42183=>"101000101",
  42184=>"111111111",
  42185=>"000000000",
  42186=>"001001000",
  42187=>"010110111",
  42188=>"001001111",
  42189=>"000000000",
  42190=>"000000000",
  42191=>"000000000",
  42192=>"111100000",
  42193=>"001001000",
  42194=>"000000110",
  42195=>"110000000",
  42196=>"000000001",
  42197=>"110110111",
  42198=>"101111111",
  42199=>"111111111",
  42200=>"000000000",
  42201=>"110100000",
  42202=>"000000100",
  42203=>"111111111",
  42204=>"111111110",
  42205=>"000000000",
  42206=>"000000000",
  42207=>"001001111",
  42208=>"111111111",
  42209=>"000000000",
  42210=>"111111111",
  42211=>"000000000",
  42212=>"000000000",
  42213=>"011011011",
  42214=>"111111111",
  42215=>"111100100",
  42216=>"000000000",
  42217=>"000111111",
  42218=>"001001111",
  42219=>"111111111",
  42220=>"000111110",
  42221=>"000000000",
  42222=>"000010111",
  42223=>"111110000",
  42224=>"100100000",
  42225=>"000000111",
  42226=>"000000100",
  42227=>"100100111",
  42228=>"110111011",
  42229=>"000110111",
  42230=>"111111111",
  42231=>"011111111",
  42232=>"000000000",
  42233=>"000000111",
  42234=>"000000000",
  42235=>"000000000",
  42236=>"011000000",
  42237=>"101000000",
  42238=>"111000000",
  42239=>"000000001",
  42240=>"000000000",
  42241=>"001001111",
  42242=>"111111111",
  42243=>"011111110",
  42244=>"000000000",
  42245=>"000110110",
  42246=>"111111000",
  42247=>"000000000",
  42248=>"000000000",
  42249=>"000010000",
  42250=>"000000111",
  42251=>"000000111",
  42252=>"000111110",
  42253=>"111111000",
  42254=>"111111111",
  42255=>"000000000",
  42256=>"000000000",
  42257=>"011111111",
  42258=>"111000000",
  42259=>"000000110",
  42260=>"111101111",
  42261=>"110111111",
  42262=>"111111110",
  42263=>"100110000",
  42264=>"001001000",
  42265=>"111111010",
  42266=>"001000000",
  42267=>"000000111",
  42268=>"111111110",
  42269=>"000010111",
  42270=>"111011001",
  42271=>"000000101",
  42272=>"111101101",
  42273=>"111011000",
  42274=>"000011011",
  42275=>"110111111",
  42276=>"111111011",
  42277=>"111101111",
  42278=>"111111111",
  42279=>"000010111",
  42280=>"111101000",
  42281=>"000000101",
  42282=>"101001000",
  42283=>"111111111",
  42284=>"111110101",
  42285=>"000111111",
  42286=>"000010111",
  42287=>"000000011",
  42288=>"000011111",
  42289=>"000000000",
  42290=>"000000001",
  42291=>"000111111",
  42292=>"000000000",
  42293=>"001011111",
  42294=>"111111111",
  42295=>"111000000",
  42296=>"000010000",
  42297=>"111001011",
  42298=>"111100000",
  42299=>"000000000",
  42300=>"100000000",
  42301=>"000000000",
  42302=>"111100111",
  42303=>"111111111",
  42304=>"000000000",
  42305=>"101101001",
  42306=>"101001101",
  42307=>"000000000",
  42308=>"011111110",
  42309=>"111111111",
  42310=>"000000010",
  42311=>"100111111",
  42312=>"111111111",
  42313=>"111010111",
  42314=>"000000000",
  42315=>"111111111",
  42316=>"001000001",
  42317=>"000000000",
  42318=>"000000000",
  42319=>"100111110",
  42320=>"110001000",
  42321=>"001011000",
  42322=>"001001001",
  42323=>"000000000",
  42324=>"000000000",
  42325=>"011011011",
  42326=>"000000110",
  42327=>"101000110",
  42328=>"001000110",
  42329=>"111111010",
  42330=>"111111111",
  42331=>"111001101",
  42332=>"010000000",
  42333=>"000000000",
  42334=>"000000111",
  42335=>"000001011",
  42336=>"011010000",
  42337=>"100000001",
  42338=>"000011011",
  42339=>"000000000",
  42340=>"011111011",
  42341=>"000000000",
  42342=>"111111111",
  42343=>"111001101",
  42344=>"011111111",
  42345=>"000000111",
  42346=>"000000011",
  42347=>"111111000",
  42348=>"000110110",
  42349=>"000000010",
  42350=>"111111010",
  42351=>"000000000",
  42352=>"000100000",
  42353=>"111001000",
  42354=>"101001111",
  42355=>"000000010",
  42356=>"000000001",
  42357=>"100100000",
  42358=>"000000000",
  42359=>"111111100",
  42360=>"000000000",
  42361=>"000001000",
  42362=>"000000001",
  42363=>"000000001",
  42364=>"111111111",
  42365=>"001000000",
  42366=>"111111111",
  42367=>"111111111",
  42368=>"111101100",
  42369=>"001000000",
  42370=>"111111111",
  42371=>"011000000",
  42372=>"000000110",
  42373=>"010000000",
  42374=>"111111111",
  42375=>"000100111",
  42376=>"101001111",
  42377=>"011011110",
  42378=>"111111111",
  42379=>"110110111",
  42380=>"111111111",
  42381=>"110110110",
  42382=>"111101111",
  42383=>"000000000",
  42384=>"111111010",
  42385=>"001000000",
  42386=>"001111111",
  42387=>"111111001",
  42388=>"000000000",
  42389=>"000001000",
  42390=>"000000101",
  42391=>"111110111",
  42392=>"111111111",
  42393=>"000000001",
  42394=>"111011110",
  42395=>"101000000",
  42396=>"001000000",
  42397=>"111111111",
  42398=>"000100100",
  42399=>"111111000",
  42400=>"000000000",
  42401=>"011011011",
  42402=>"000101111",
  42403=>"111111111",
  42404=>"110111111",
  42405=>"111111111",
  42406=>"000000000",
  42407=>"000000000",
  42408=>"000001000",
  42409=>"101100111",
  42410=>"000000000",
  42411=>"101100000",
  42412=>"000000000",
  42413=>"001110111",
  42414=>"111111111",
  42415=>"000000000",
  42416=>"111111111",
  42417=>"011011111",
  42418=>"000110110",
  42419=>"000000000",
  42420=>"111110010",
  42421=>"110100110",
  42422=>"111111111",
  42423=>"111111111",
  42424=>"111111000",
  42425=>"000000000",
  42426=>"000000101",
  42427=>"111000000",
  42428=>"000000111",
  42429=>"100100111",
  42430=>"111101101",
  42431=>"111111100",
  42432=>"000000000",
  42433=>"000000000",
  42434=>"111111111",
  42435=>"111111000",
  42436=>"100000101",
  42437=>"111110111",
  42438=>"011111110",
  42439=>"111001000",
  42440=>"010000000",
  42441=>"111111111",
  42442=>"111111111",
  42443=>"000000000",
  42444=>"011000000",
  42445=>"111111111",
  42446=>"001000000",
  42447=>"000000110",
  42448=>"001000000",
  42449=>"010000001",
  42450=>"000000101",
  42451=>"000000000",
  42452=>"100010000",
  42453=>"001000000",
  42454=>"000001001",
  42455=>"111110111",
  42456=>"000000000",
  42457=>"111111111",
  42458=>"100100111",
  42459=>"111111111",
  42460=>"000000001",
  42461=>"110110100",
  42462=>"000000111",
  42463=>"000111111",
  42464=>"000001001",
  42465=>"100111011",
  42466=>"111111111",
  42467=>"111111111",
  42468=>"111111111",
  42469=>"000000011",
  42470=>"000000001",
  42471=>"000000000",
  42472=>"111111111",
  42473=>"011010000",
  42474=>"000000000",
  42475=>"011111111",
  42476=>"110110111",
  42477=>"111111001",
  42478=>"000000000",
  42479=>"000000100",
  42480=>"000000111",
  42481=>"111111000",
  42482=>"111111100",
  42483=>"000110000",
  42484=>"000000000",
  42485=>"110000000",
  42486=>"000000000",
  42487=>"000000100",
  42488=>"111111000",
  42489=>"110110001",
  42490=>"111111011",
  42491=>"111111100",
  42492=>"001111111",
  42493=>"000000001",
  42494=>"000000110",
  42495=>"000000000",
  42496=>"000000000",
  42497=>"000000000",
  42498=>"100100000",
  42499=>"111111100",
  42500=>"000110000",
  42501=>"100111110",
  42502=>"000000000",
  42503=>"111000000",
  42504=>"011011001",
  42505=>"000101111",
  42506=>"110000001",
  42507=>"000100101",
  42508=>"000000000",
  42509=>"111111100",
  42510=>"100100100",
  42511=>"000000000",
  42512=>"100000100",
  42513=>"111000000",
  42514=>"111111110",
  42515=>"100100110",
  42516=>"111111111",
  42517=>"001000100",
  42518=>"010000011",
  42519=>"000000100",
  42520=>"011011011",
  42521=>"100000001",
  42522=>"000000001",
  42523=>"000000111",
  42524=>"011111111",
  42525=>"011011011",
  42526=>"111111111",
  42527=>"111111001",
  42528=>"111111010",
  42529=>"010000000",
  42530=>"110100101",
  42531=>"110110111",
  42532=>"000000000",
  42533=>"000000000",
  42534=>"111000000",
  42535=>"000011111",
  42536=>"111110111",
  42537=>"001100111",
  42538=>"000000000",
  42539=>"000010000",
  42540=>"101111000",
  42541=>"111111011",
  42542=>"100100000",
  42543=>"100100000",
  42544=>"111111100",
  42545=>"111111011",
  42546=>"000010011",
  42547=>"010011001",
  42548=>"111001101",
  42549=>"110000000",
  42550=>"010000000",
  42551=>"110100000",
  42552=>"011010011",
  42553=>"111100100",
  42554=>"000000000",
  42555=>"000000000",
  42556=>"110111111",
  42557=>"011011000",
  42558=>"000100111",
  42559=>"000000001",
  42560=>"101100100",
  42561=>"000100000",
  42562=>"010111011",
  42563=>"101101101",
  42564=>"110010011",
  42565=>"111111111",
  42566=>"111001001",
  42567=>"000000000",
  42568=>"110111111",
  42569=>"111101111",
  42570=>"000110111",
  42571=>"111111100",
  42572=>"000011111",
  42573=>"110100111",
  42574=>"110010010",
  42575=>"100100111",
  42576=>"000011001",
  42577=>"101101101",
  42578=>"111111111",
  42579=>"110111001",
  42580=>"111111111",
  42581=>"000010011",
  42582=>"111111110",
  42583=>"010111111",
  42584=>"011010110",
  42585=>"100000000",
  42586=>"111111111",
  42587=>"100000000",
  42588=>"011001011",
  42589=>"000000000",
  42590=>"000000000",
  42591=>"111110100",
  42592=>"101101000",
  42593=>"111111111",
  42594=>"100001000",
  42595=>"111101100",
  42596=>"000110111",
  42597=>"011010000",
  42598=>"001000000",
  42599=>"111010000",
  42600=>"001101100",
  42601=>"111101001",
  42602=>"101101000",
  42603=>"001001001",
  42604=>"000101111",
  42605=>"000000000",
  42606=>"000000010",
  42607=>"111011001",
  42608=>"000000100",
  42609=>"100000100",
  42610=>"111111111",
  42611=>"100100100",
  42612=>"111111111",
  42613=>"010000000",
  42614=>"000000001",
  42615=>"111111110",
  42616=>"000000011",
  42617=>"111111111",
  42618=>"111110110",
  42619=>"000000000",
  42620=>"111111111",
  42621=>"110100110",
  42622=>"110110000",
  42623=>"011011101",
  42624=>"000100000",
  42625=>"000100110",
  42626=>"101111101",
  42627=>"000100100",
  42628=>"001001000",
  42629=>"110101111",
  42630=>"111000000",
  42631=>"011111100",
  42632=>"111110111",
  42633=>"000001001",
  42634=>"001000001",
  42635=>"001001001",
  42636=>"100111011",
  42637=>"100111111",
  42638=>"101111110",
  42639=>"000000000",
  42640=>"000001000",
  42641=>"111001100",
  42642=>"001001111",
  42643=>"000000111",
  42644=>"101101000",
  42645=>"111011011",
  42646=>"000000000",
  42647=>"100100000",
  42648=>"000110000",
  42649=>"111111111",
  42650=>"010000010",
  42651=>"000001000",
  42652=>"011000000",
  42653=>"011011010",
  42654=>"111001001",
  42655=>"100100110",
  42656=>"011000100",
  42657=>"110000000",
  42658=>"001001000",
  42659=>"111110111",
  42660=>"110000110",
  42661=>"000000001",
  42662=>"000000111",
  42663=>"111000000",
  42664=>"111111111",
  42665=>"000000000",
  42666=>"111111011",
  42667=>"001001001",
  42668=>"010001100",
  42669=>"100101101",
  42670=>"110110110",
  42671=>"100000000",
  42672=>"100100000",
  42673=>"000000110",
  42674=>"110110111",
  42675=>"000100001",
  42676=>"010010011",
  42677=>"010111010",
  42678=>"111111111",
  42679=>"111111111",
  42680=>"000000100",
  42681=>"000000000",
  42682=>"110000000",
  42683=>"010000000",
  42684=>"011000001",
  42685=>"000000000",
  42686=>"001001000",
  42687=>"111111111",
  42688=>"000000100",
  42689=>"110110110",
  42690=>"111011111",
  42691=>"000000000",
  42692=>"111111111",
  42693=>"110111111",
  42694=>"111010010",
  42695=>"111111111",
  42696=>"000000000",
  42697=>"110010111",
  42698=>"010000100",
  42699=>"111111111",
  42700=>"111001101",
  42701=>"000110110",
  42702=>"000000000",
  42703=>"000000000",
  42704=>"000111111",
  42705=>"010000111",
  42706=>"011010011",
  42707=>"000000000",
  42708=>"111011000",
  42709=>"101111111",
  42710=>"000000000",
  42711=>"010100000",
  42712=>"111111101",
  42713=>"110110100",
  42714=>"000000100",
  42715=>"111011110",
  42716=>"111111111",
  42717=>"000000000",
  42718=>"111111111",
  42719=>"010000000",
  42720=>"000000000",
  42721=>"101101111",
  42722=>"111001100",
  42723=>"001011111",
  42724=>"000010001",
  42725=>"111110110",
  42726=>"111010010",
  42727=>"111011011",
  42728=>"000110111",
  42729=>"111111111",
  42730=>"111111111",
  42731=>"111000000",
  42732=>"111110000",
  42733=>"000000000",
  42734=>"100101111",
  42735=>"000111110",
  42736=>"000000000",
  42737=>"000000000",
  42738=>"110100000",
  42739=>"010111111",
  42740=>"111111111",
  42741=>"001000000",
  42742=>"001000001",
  42743=>"111111111",
  42744=>"000000000",
  42745=>"011010111",
  42746=>"000000000",
  42747=>"110111000",
  42748=>"111111100",
  42749=>"110110110",
  42750=>"000000100",
  42751=>"010110010",
  42752=>"000000111",
  42753=>"011011010",
  42754=>"110000110",
  42755=>"000000000",
  42756=>"000000000",
  42757=>"000001001",
  42758=>"000000000",
  42759=>"101001111",
  42760=>"010010000",
  42761=>"001000001",
  42762=>"111111111",
  42763=>"000000100",
  42764=>"000000000",
  42765=>"011111111",
  42766=>"000000111",
  42767=>"001001001",
  42768=>"011011011",
  42769=>"000000000",
  42770=>"111000000",
  42771=>"110000000",
  42772=>"110000000",
  42773=>"000000000",
  42774=>"100001000",
  42775=>"111110100",
  42776=>"010000001",
  42777=>"010110111",
  42778=>"011101000",
  42779=>"001000101",
  42780=>"001000000",
  42781=>"001001001",
  42782=>"000000000",
  42783=>"111111000",
  42784=>"001111111",
  42785=>"100111101",
  42786=>"011011111",
  42787=>"000101111",
  42788=>"111011011",
  42789=>"111111111",
  42790=>"001011000",
  42791=>"111011111",
  42792=>"000000010",
  42793=>"000000110",
  42794=>"111111000",
  42795=>"000000000",
  42796=>"000010111",
  42797=>"000010010",
  42798=>"000011101",
  42799=>"000000111",
  42800=>"100001001",
  42801=>"011111111",
  42802=>"111011011",
  42803=>"111111111",
  42804=>"110100000",
  42805=>"001000000",
  42806=>"111100100",
  42807=>"011111111",
  42808=>"101111100",
  42809=>"000000000",
  42810=>"010000000",
  42811=>"111111111",
  42812=>"011011111",
  42813=>"111111111",
  42814=>"010010011",
  42815=>"011000010",
  42816=>"000000100",
  42817=>"111011000",
  42818=>"001001101",
  42819=>"000010100",
  42820=>"000010100",
  42821=>"101100111",
  42822=>"000000011",
  42823=>"111111111",
  42824=>"000000000",
  42825=>"111000000",
  42826=>"111111000",
  42827=>"011001000",
  42828=>"000000000",
  42829=>"110111000",
  42830=>"000111111",
  42831=>"011011010",
  42832=>"111110110",
  42833=>"010011011",
  42834=>"101111111",
  42835=>"011111111",
  42836=>"100100000",
  42837=>"001011011",
  42838=>"101000010",
  42839=>"001000001",
  42840=>"000000100",
  42841=>"111111111",
  42842=>"000111011",
  42843=>"000011111",
  42844=>"000001101",
  42845=>"111111111",
  42846=>"100101111",
  42847=>"110100110",
  42848=>"100000000",
  42849=>"111000000",
  42850=>"000110111",
  42851=>"100111000",
  42852=>"010010100",
  42853=>"110111100",
  42854=>"101101101",
  42855=>"010111111",
  42856=>"100000100",
  42857=>"110111111",
  42858=>"111111111",
  42859=>"001010110",
  42860=>"111111111",
  42861=>"010000000",
  42862=>"000000000",
  42863=>"111011010",
  42864=>"110110110",
  42865=>"000000000",
  42866=>"100000100",
  42867=>"111110110",
  42868=>"010110010",
  42869=>"000000000",
  42870=>"011011111",
  42871=>"101101101",
  42872=>"000111111",
  42873=>"001000000",
  42874=>"111110111",
  42875=>"110111011",
  42876=>"000000000",
  42877=>"110111111",
  42878=>"111000000",
  42879=>"011011011",
  42880=>"000000010",
  42881=>"111100100",
  42882=>"011011011",
  42883=>"011111011",
  42884=>"001001111",
  42885=>"100100110",
  42886=>"111111011",
  42887=>"110111111",
  42888=>"111111111",
  42889=>"100000000",
  42890=>"111011000",
  42891=>"100100101",
  42892=>"111111000",
  42893=>"000000000",
  42894=>"111110111",
  42895=>"111111110",
  42896=>"101111111",
  42897=>"000100110",
  42898=>"000000100",
  42899=>"000000000",
  42900=>"000011111",
  42901=>"011001001",
  42902=>"000000100",
  42903=>"100100000",
  42904=>"000000010",
  42905=>"111111010",
  42906=>"111111111",
  42907=>"000000000",
  42908=>"001001111",
  42909=>"110110100",
  42910=>"010010111",
  42911=>"000000000",
  42912=>"000000000",
  42913=>"000000100",
  42914=>"000000110",
  42915=>"111111010",
  42916=>"000000100",
  42917=>"001111111",
  42918=>"001001000",
  42919=>"111111111",
  42920=>"000100000",
  42921=>"110111100",
  42922=>"000000000",
  42923=>"111111001",
  42924=>"111111001",
  42925=>"101100000",
  42926=>"110000010",
  42927=>"111111111",
  42928=>"001000000",
  42929=>"001001111",
  42930=>"001001100",
  42931=>"011101101",
  42932=>"001000100",
  42933=>"001001111",
  42934=>"000100110",
  42935=>"000100001",
  42936=>"000001111",
  42937=>"111010110",
  42938=>"001001011",
  42939=>"000000000",
  42940=>"001100110",
  42941=>"000110111",
  42942=>"100100100",
  42943=>"110000110",
  42944=>"011011001",
  42945=>"101001001",
  42946=>"111111010",
  42947=>"111010000",
  42948=>"110110100",
  42949=>"001001001",
  42950=>"100000001",
  42951=>"101100100",
  42952=>"011011111",
  42953=>"111111011",
  42954=>"000000000",
  42955=>"100100100",
  42956=>"100001000",
  42957=>"100000000",
  42958=>"111010110",
  42959=>"111111111",
  42960=>"100111101",
  42961=>"100101101",
  42962=>"000100001",
  42963=>"111111110",
  42964=>"000011001",
  42965=>"100110100",
  42966=>"000000101",
  42967=>"111111101",
  42968=>"000000000",
  42969=>"111111110",
  42970=>"010011011",
  42971=>"011010111",
  42972=>"111111110",
  42973=>"101000001",
  42974=>"111011111",
  42975=>"010000000",
  42976=>"101111101",
  42977=>"000100000",
  42978=>"011011111",
  42979=>"111111111",
  42980=>"000100011",
  42981=>"111111011",
  42982=>"100000000",
  42983=>"111111111",
  42984=>"110110111",
  42985=>"111001000",
  42986=>"000011110",
  42987=>"111111100",
  42988=>"101111100",
  42989=>"011011001",
  42990=>"100000001",
  42991=>"111111111",
  42992=>"111011011",
  42993=>"111101101",
  42994=>"000010010",
  42995=>"000100111",
  42996=>"110111001",
  42997=>"000000000",
  42998=>"111111111",
  42999=>"111001000",
  43000=>"100111111",
  43001=>"011000000",
  43002=>"110000000",
  43003=>"000001000",
  43004=>"111110110",
  43005=>"111111110",
  43006=>"111011011",
  43007=>"000000000",
  43008=>"000000000",
  43009=>"100000000",
  43010=>"000100111",
  43011=>"001011111",
  43012=>"000010110",
  43013=>"011010000",
  43014=>"111111110",
  43015=>"000000000",
  43016=>"000111011",
  43017=>"100100000",
  43018=>"111111111",
  43019=>"000000111",
  43020=>"000000000",
  43021=>"110100111",
  43022=>"100010000",
  43023=>"000000000",
  43024=>"011011001",
  43025=>"111111111",
  43026=>"111000000",
  43027=>"000000000",
  43028=>"111111111",
  43029=>"000000000",
  43030=>"111000000",
  43031=>"110111111",
  43032=>"101101111",
  43033=>"000000000",
  43034=>"001000000",
  43035=>"000000000",
  43036=>"100000000",
  43037=>"011111111",
  43038=>"101101001",
  43039=>"110111110",
  43040=>"000001001",
  43041=>"110111110",
  43042=>"111111111",
  43043=>"111111111",
  43044=>"100001111",
  43045=>"111111011",
  43046=>"001001011",
  43047=>"100110111",
  43048=>"001000000",
  43049=>"000100000",
  43050=>"000000000",
  43051=>"110100101",
  43052=>"110100111",
  43053=>"001001101",
  43054=>"111111111",
  43055=>"011111111",
  43056=>"001101000",
  43057=>"111111000",
  43058=>"011011010",
  43059=>"000000000",
  43060=>"011011111",
  43061=>"000000000",
  43062=>"001001001",
  43063=>"000100101",
  43064=>"000110110",
  43065=>"110000000",
  43066=>"111111111",
  43067=>"000110110",
  43068=>"100000000",
  43069=>"111111111",
  43070=>"111111111",
  43071=>"111100000",
  43072=>"111111111",
  43073=>"010010000",
  43074=>"111111111",
  43075=>"111111111",
  43076=>"111100000",
  43077=>"101101111",
  43078=>"111111000",
  43079=>"111111111",
  43080=>"011101001",
  43081=>"111111010",
  43082=>"000000011",
  43083=>"111111001",
  43084=>"001111111",
  43085=>"111111000",
  43086=>"000110111",
  43087=>"111111011",
  43088=>"101101000",
  43089=>"111111010",
  43090=>"000000000",
  43091=>"000000000",
  43092=>"000000000",
  43093=>"110111111",
  43094=>"011000000",
  43095=>"111111111",
  43096=>"000110100",
  43097=>"111111111",
  43098=>"111111111",
  43099=>"101101101",
  43100=>"000100111",
  43101=>"101001011",
  43102=>"000111110",
  43103=>"100111111",
  43104=>"000001001",
  43105=>"111110111",
  43106=>"000001000",
  43107=>"010111110",
  43108=>"011110100",
  43109=>"111111111",
  43110=>"110000001",
  43111=>"001001001",
  43112=>"110110111",
  43113=>"000000000",
  43114=>"000000100",
  43115=>"000010111",
  43116=>"000001011",
  43117=>"101001111",
  43118=>"000000111",
  43119=>"000000000",
  43120=>"100100110",
  43121=>"000010011",
  43122=>"000000001",
  43123=>"000001000",
  43124=>"111111111",
  43125=>"100000101",
  43126=>"111001000",
  43127=>"100000000",
  43128=>"111111001",
  43129=>"000110111",
  43130=>"111111111",
  43131=>"110111111",
  43132=>"100100100",
  43133=>"111111111",
  43134=>"000000000",
  43135=>"111111111",
  43136=>"110000000",
  43137=>"111111111",
  43138=>"001000010",
  43139=>"000111100",
  43140=>"000000000",
  43141=>"111111111",
  43142=>"001110010",
  43143=>"001011111",
  43144=>"111101111",
  43145=>"111111001",
  43146=>"111110100",
  43147=>"111111000",
  43148=>"000000000",
  43149=>"110000000",
  43150=>"000000010",
  43151=>"001111111",
  43152=>"000000000",
  43153=>"000000000",
  43154=>"100100101",
  43155=>"100101000",
  43156=>"110100000",
  43157=>"000000000",
  43158=>"111111011",
  43159=>"111001000",
  43160=>"000000000",
  43161=>"111111111",
  43162=>"001111100",
  43163=>"001011000",
  43164=>"000000000",
  43165=>"011001001",
  43166=>"000000111",
  43167=>"000110110",
  43168=>"000001101",
  43169=>"101000000",
  43170=>"111111000",
  43171=>"111111110",
  43172=>"000000000",
  43173=>"110100100",
  43174=>"000101111",
  43175=>"100000001",
  43176=>"111111111",
  43177=>"000000000",
  43178=>"000000000",
  43179=>"111010000",
  43180=>"111111111",
  43181=>"101111111",
  43182=>"000000000",
  43183=>"000000000",
  43184=>"001000000",
  43185=>"110011001",
  43186=>"000000000",
  43187=>"111111011",
  43188=>"111111111",
  43189=>"111111111",
  43190=>"101000000",
  43191=>"000000000",
  43192=>"111111101",
  43193=>"001000010",
  43194=>"000011010",
  43195=>"111001000",
  43196=>"111111111",
  43197=>"110000000",
  43198=>"000000110",
  43199=>"111011111",
  43200=>"100100100",
  43201=>"101111111",
  43202=>"011111111",
  43203=>"001001000",
  43204=>"111111101",
  43205=>"111110110",
  43206=>"000000000",
  43207=>"101111110",
  43208=>"011011011",
  43209=>"000000000",
  43210=>"100101101",
  43211=>"000000000",
  43212=>"111111010",
  43213=>"111111111",
  43214=>"000000000",
  43215=>"100100100",
  43216=>"111111101",
  43217=>"000000000",
  43218=>"111111001",
  43219=>"000000000",
  43220=>"000011111",
  43221=>"000001011",
  43222=>"000000000",
  43223=>"110100100",
  43224=>"100000100",
  43225=>"000000000",
  43226=>"100000000",
  43227=>"111111100",
  43228=>"111110111",
  43229=>"111111111",
  43230=>"111111111",
  43231=>"111111000",
  43232=>"111111111",
  43233=>"010110110",
  43234=>"110111000",
  43235=>"111111111",
  43236=>"000000000",
  43237=>"111110110",
  43238=>"111111111",
  43239=>"000100000",
  43240=>"000000000",
  43241=>"001101011",
  43242=>"000000000",
  43243=>"000000101",
  43244=>"111111111",
  43245=>"000000000",
  43246=>"000110110",
  43247=>"111111111",
  43248=>"000000000",
  43249=>"100000000",
  43250=>"111111000",
  43251=>"001000011",
  43252=>"100000000",
  43253=>"111111101",
  43254=>"000010010",
  43255=>"000100000",
  43256=>"000000000",
  43257=>"111111111",
  43258=>"111100111",
  43259=>"010000000",
  43260=>"011011111",
  43261=>"111011101",
  43262=>"101000000",
  43263=>"101001111",
  43264=>"111111111",
  43265=>"110100000",
  43266=>"110110000",
  43267=>"110110000",
  43268=>"111111100",
  43269=>"000000000",
  43270=>"001111111",
  43271=>"000010111",
  43272=>"000000000",
  43273=>"000000110",
  43274=>"111111010",
  43275=>"100011000",
  43276=>"111101101",
  43277=>"000000111",
  43278=>"000000000",
  43279=>"000000000",
  43280=>"111100000",
  43281=>"111110111",
  43282=>"111101111",
  43283=>"111111111",
  43284=>"110110100",
  43285=>"000000000",
  43286=>"111111011",
  43287=>"000000000",
  43288=>"001001001",
  43289=>"000001101",
  43290=>"100000000",
  43291=>"111111111",
  43292=>"010111110",
  43293=>"000000100",
  43294=>"111111111",
  43295=>"001111011",
  43296=>"100111001",
  43297=>"000000000",
  43298=>"111011111",
  43299=>"000000000",
  43300=>"100111010",
  43301=>"100100000",
  43302=>"111110100",
  43303=>"000110010",
  43304=>"101001011",
  43305=>"111111011",
  43306=>"001000000",
  43307=>"001011111",
  43308=>"011010010",
  43309=>"011111111",
  43310=>"111111000",
  43311=>"100100000",
  43312=>"001100010",
  43313=>"001001000",
  43314=>"110111111",
  43315=>"000001101",
  43316=>"111111111",
  43317=>"000001011",
  43318=>"110110000",
  43319=>"010011000",
  43320=>"100001011",
  43321=>"000000000",
  43322=>"111111111",
  43323=>"000000000",
  43324=>"110110110",
  43325=>"111001000",
  43326=>"000000000",
  43327=>"100000000",
  43328=>"000001000",
  43329=>"110110000",
  43330=>"000000000",
  43331=>"111111111",
  43332=>"111111110",
  43333=>"000000100",
  43334=>"110110000",
  43335=>"000000000",
  43336=>"111101111",
  43337=>"110111110",
  43338=>"100110100",
  43339=>"111101111",
  43340=>"111110110",
  43341=>"111111100",
  43342=>"001001101",
  43343=>"111101001",
  43344=>"111001001",
  43345=>"000011111",
  43346=>"111111111",
  43347=>"000100111",
  43348=>"000000000",
  43349=>"001001011",
  43350=>"000110111",
  43351=>"000000000",
  43352=>"000110111",
  43353=>"111111111",
  43354=>"110011011",
  43355=>"111111111",
  43356=>"111010110",
  43357=>"100100000",
  43358=>"111111001",
  43359=>"011000000",
  43360=>"101111111",
  43361=>"110000000",
  43362=>"110111111",
  43363=>"000000111",
  43364=>"011011011",
  43365=>"000000000",
  43366=>"001000000",
  43367=>"001000000",
  43368=>"101100111",
  43369=>"110000000",
  43370=>"000000000",
  43371=>"111100111",
  43372=>"011111100",
  43373=>"000000000",
  43374=>"000000010",
  43375=>"011111111",
  43376=>"000000000",
  43377=>"011001001",
  43378=>"000000000",
  43379=>"100100111",
  43380=>"000000000",
  43381=>"001001000",
  43382=>"000000101",
  43383=>"000100001",
  43384=>"000000000",
  43385=>"111001100",
  43386=>"000000000",
  43387=>"111111111",
  43388=>"000000101",
  43389=>"000100111",
  43390=>"111111111",
  43391=>"000000000",
  43392=>"110000001",
  43393=>"101111111",
  43394=>"111111111",
  43395=>"111111111",
  43396=>"100110111",
  43397=>"111111111",
  43398=>"100111111",
  43399=>"111111111",
  43400=>"010000000",
  43401=>"110101111",
  43402=>"000110110",
  43403=>"111110000",
  43404=>"111111111",
  43405=>"100100000",
  43406=>"001000000",
  43407=>"000000111",
  43408=>"000000000",
  43409=>"111111001",
  43410=>"011111000",
  43411=>"110101101",
  43412=>"000000000",
  43413=>"111010000",
  43414=>"100110111",
  43415=>"001001000",
  43416=>"000010010",
  43417=>"000000000",
  43418=>"111111111",
  43419=>"101100100",
  43420=>"000000000",
  43421=>"011111110",
  43422=>"111001001",
  43423=>"000000001",
  43424=>"111111111",
  43425=>"000010011",
  43426=>"000000000",
  43427=>"000001111",
  43428=>"111010111",
  43429=>"000001000",
  43430=>"111011001",
  43431=>"111001000",
  43432=>"000000000",
  43433=>"100110111",
  43434=>"111111100",
  43435=>"000000001",
  43436=>"000000000",
  43437=>"111111111",
  43438=>"000000100",
  43439=>"000011010",
  43440=>"111111111",
  43441=>"110010000",
  43442=>"111111000",
  43443=>"111110111",
  43444=>"000100000",
  43445=>"011000010",
  43446=>"000000000",
  43447=>"111111111",
  43448=>"111111111",
  43449=>"111001001",
  43450=>"000000000",
  43451=>"100000111",
  43452=>"010111111",
  43453=>"001000000",
  43454=>"001000010",
  43455=>"111111011",
  43456=>"000000000",
  43457=>"000000000",
  43458=>"000010000",
  43459=>"111111111",
  43460=>"000000000",
  43461=>"100100111",
  43462=>"000000000",
  43463=>"011011111",
  43464=>"000000000",
  43465=>"111100000",
  43466=>"000000000",
  43467=>"000100110",
  43468=>"111111010",
  43469=>"000000000",
  43470=>"111111001",
  43471=>"000000100",
  43472=>"000110111",
  43473=>"000000001",
  43474=>"001100111",
  43475=>"000000000",
  43476=>"101111111",
  43477=>"000000000",
  43478=>"001011011",
  43479=>"100100100",
  43480=>"000000000",
  43481=>"111111111",
  43482=>"000000001",
  43483=>"010000000",
  43484=>"000000000",
  43485=>"011111011",
  43486=>"000110110",
  43487=>"111100101",
  43488=>"111110110",
  43489=>"111111111",
  43490=>"000111111",
  43491=>"100000011",
  43492=>"000000111",
  43493=>"111000001",
  43494=>"000000000",
  43495=>"110111111",
  43496=>"111111001",
  43497=>"011111111",
  43498=>"000000001",
  43499=>"000000000",
  43500=>"111110000",
  43501=>"101111001",
  43502=>"011111111",
  43503=>"011000000",
  43504=>"000000000",
  43505=>"111111000",
  43506=>"111111111",
  43507=>"011011111",
  43508=>"000100110",
  43509=>"001101100",
  43510=>"000000000",
  43511=>"101000100",
  43512=>"011111111",
  43513=>"101101101",
  43514=>"111001001",
  43515=>"000000000",
  43516=>"011011001",
  43517=>"111111111",
  43518=>"000101001",
  43519=>"110111111",
  43520=>"000000000",
  43521=>"000000101",
  43522=>"111001111",
  43523=>"001100101",
  43524=>"100100111",
  43525=>"111000001",
  43526=>"110111100",
  43527=>"111101101",
  43528=>"100001011",
  43529=>"110000000",
  43530=>"111111111",
  43531=>"111011011",
  43532=>"011000011",
  43533=>"111111001",
  43534=>"001000000",
  43535=>"000000000",
  43536=>"000000000",
  43537=>"000000000",
  43538=>"000000110",
  43539=>"010000111",
  43540=>"111111111",
  43541=>"000000000",
  43542=>"000100100",
  43543=>"111111111",
  43544=>"111111111",
  43545=>"100110110",
  43546=>"011000000",
  43547=>"110110100",
  43548=>"111111111",
  43549=>"000000000",
  43550=>"111011011",
  43551=>"110110000",
  43552=>"000000000",
  43553=>"111111110",
  43554=>"100110111",
  43555=>"111111111",
  43556=>"000000000",
  43557=>"000111110",
  43558=>"110011111",
  43559=>"000000111",
  43560=>"010100000",
  43561=>"000000000",
  43562=>"011111111",
  43563=>"000101111",
  43564=>"001000000",
  43565=>"000001011",
  43566=>"000000000",
  43567=>"111111111",
  43568=>"001000001",
  43569=>"000001011",
  43570=>"101111110",
  43571=>"000000110",
  43572=>"000000010",
  43573=>"001001001",
  43574=>"000111111",
  43575=>"001000000",
  43576=>"000000100",
  43577=>"111000000",
  43578=>"001001111",
  43579=>"000000111",
  43580=>"000000000",
  43581=>"111000000",
  43582=>"110111111",
  43583=>"000000000",
  43584=>"000000000",
  43585=>"010011111",
  43586=>"111111111",
  43587=>"111111000",
  43588=>"000000001",
  43589=>"110110000",
  43590=>"000000111",
  43591=>"000000000",
  43592=>"001000101",
  43593=>"001000111",
  43594=>"000000000",
  43595=>"000000111",
  43596=>"000000110",
  43597=>"111111111",
  43598=>"001111111",
  43599=>"111111001",
  43600=>"000000010",
  43601=>"111000000",
  43602=>"000000000",
  43603=>"000001000",
  43604=>"010111101",
  43605=>"010010111",
  43606=>"011110110",
  43607=>"000001001",
  43608=>"111000110",
  43609=>"000000000",
  43610=>"001101111",
  43611=>"011001000",
  43612=>"100100111",
  43613=>"000111000",
  43614=>"000111111",
  43615=>"110110100",
  43616=>"111011111",
  43617=>"000000000",
  43618=>"111111111",
  43619=>"111111111",
  43620=>"000001101",
  43621=>"111100000",
  43622=>"000000000",
  43623=>"111000000",
  43624=>"000101111",
  43625=>"111100111",
  43626=>"111100100",
  43627=>"000011001",
  43628=>"111111111",
  43629=>"110110100",
  43630=>"001001111",
  43631=>"111011000",
  43632=>"000000000",
  43633=>"111011000",
  43634=>"000110111",
  43635=>"101101000",
  43636=>"000000000",
  43637=>"000000000",
  43638=>"000001111",
  43639=>"110110110",
  43640=>"000101101",
  43641=>"000000000",
  43642=>"000000000",
  43643=>"000000000",
  43644=>"011001011",
  43645=>"000010010",
  43646=>"000000111",
  43647=>"000000110",
  43648=>"100100000",
  43649=>"110100000",
  43650=>"111111110",
  43651=>"111000000",
  43652=>"111111111",
  43653=>"101001111",
  43654=>"000000000",
  43655=>"000000101",
  43656=>"111110110",
  43657=>"000000000",
  43658=>"111111111",
  43659=>"001000000",
  43660=>"111111110",
  43661=>"111111111",
  43662=>"010011000",
  43663=>"111111111",
  43664=>"000000000",
  43665=>"000110111",
  43666=>"000010000",
  43667=>"000000000",
  43668=>"110111111",
  43669=>"000111111",
  43670=>"111011111",
  43671=>"111000110",
  43672=>"000001000",
  43673=>"000100110",
  43674=>"000000000",
  43675=>"000100000",
  43676=>"000000000",
  43677=>"000000000",
  43678=>"111000111",
  43679=>"110100100",
  43680=>"111011101",
  43681=>"111111111",
  43682=>"111111001",
  43683=>"100000100",
  43684=>"011000010",
  43685=>"110111111",
  43686=>"111111111",
  43687=>"000000001",
  43688=>"001000101",
  43689=>"000000000",
  43690=>"100001000",
  43691=>"000000000",
  43692=>"011111111",
  43693=>"100100101",
  43694=>"110100000",
  43695=>"111000011",
  43696=>"001101111",
  43697=>"000001000",
  43698=>"111111110",
  43699=>"111111111",
  43700=>"101101000",
  43701=>"111111111",
  43702=>"000111111",
  43703=>"100100110",
  43704=>"100101000",
  43705=>"100100100",
  43706=>"111111111",
  43707=>"111101101",
  43708=>"001000000",
  43709=>"101000000",
  43710=>"000000000",
  43711=>"100111101",
  43712=>"000000111",
  43713=>"111111111",
  43714=>"000000000",
  43715=>"111111100",
  43716=>"000000000",
  43717=>"000000000",
  43718=>"010110000",
  43719=>"000101111",
  43720=>"000000000",
  43721=>"001000000",
  43722=>"011001000",
  43723=>"001111110",
  43724=>"010000000",
  43725=>"010111000",
  43726=>"000001111",
  43727=>"000000000",
  43728=>"111111110",
  43729=>"001000000",
  43730=>"000000001",
  43731=>"010110010",
  43732=>"000001101",
  43733=>"000000111",
  43734=>"000000000",
  43735=>"010010000",
  43736=>"111111111",
  43737=>"000000000",
  43738=>"110111111",
  43739=>"100111111",
  43740=>"001001111",
  43741=>"010111111",
  43742=>"111111111",
  43743=>"011111110",
  43744=>"111111111",
  43745=>"000010110",
  43746=>"011000000",
  43747=>"000000000",
  43748=>"111111111",
  43749=>"000110110",
  43750=>"000000000",
  43751=>"110110001",
  43752=>"111111111",
  43753=>"000000000",
  43754=>"111111111",
  43755=>"111000000",
  43756=>"011000001",
  43757=>"000000000",
  43758=>"111000000",
  43759=>"011000000",
  43760=>"000000000",
  43761=>"010000000",
  43762=>"001101111",
  43763=>"111111011",
  43764=>"111111111",
  43765=>"011011001",
  43766=>"111110100",
  43767=>"000011000",
  43768=>"000000000",
  43769=>"000010011",
  43770=>"111111011",
  43771=>"000001111",
  43772=>"000100110",
  43773=>"011001111",
  43774=>"000000000",
  43775=>"100000000",
  43776=>"100000000",
  43777=>"000000001",
  43778=>"011011011",
  43779=>"000000011",
  43780=>"011010110",
  43781=>"001111111",
  43782=>"111111111",
  43783=>"000000000",
  43784=>"101101111",
  43785=>"000000000",
  43786=>"000000000",
  43787=>"111111111",
  43788=>"101101001",
  43789=>"100111111",
  43790=>"000111111",
  43791=>"000000011",
  43792=>"111111111",
  43793=>"100111111",
  43794=>"001000000",
  43795=>"000000000",
  43796=>"011111111",
  43797=>"000000000",
  43798=>"010010000",
  43799=>"100111101",
  43800=>"110111111",
  43801=>"000000000",
  43802=>"000000000",
  43803=>"000000000",
  43804=>"111111111",
  43805=>"011000000",
  43806=>"111111110",
  43807=>"001011111",
  43808=>"100111111",
  43809=>"000000001",
  43810=>"110000000",
  43811=>"000000000",
  43812=>"111111111",
  43813=>"110110111",
  43814=>"110110110",
  43815=>"110010000",
  43816=>"000000000",
  43817=>"101000000",
  43818=>"111111111",
  43819=>"000001000",
  43820=>"000000000",
  43821=>"000100110",
  43822=>"000001111",
  43823=>"000100111",
  43824=>"111111000",
  43825=>"000000000",
  43826=>"111000000",
  43827=>"000000000",
  43828=>"111011000",
  43829=>"100000000",
  43830=>"111111111",
  43831=>"000000000",
  43832=>"110000001",
  43833=>"111111111",
  43834=>"111110000",
  43835=>"000000000",
  43836=>"111010000",
  43837=>"111101101",
  43838=>"111101000",
  43839=>"010111110",
  43840=>"100000000",
  43841=>"111101101",
  43842=>"111111111",
  43843=>"000110100",
  43844=>"111111001",
  43845=>"000000000",
  43846=>"111111110",
  43847=>"001001101",
  43848=>"011000000",
  43849=>"111011111",
  43850=>"000000001",
  43851=>"111111111",
  43852=>"111111011",
  43853=>"111000000",
  43854=>"111100000",
  43855=>"101111110",
  43856=>"000000100",
  43857=>"000000000",
  43858=>"000000000",
  43859=>"000010110",
  43860=>"000000111",
  43861=>"111111111",
  43862=>"010111111",
  43863=>"111111011",
  43864=>"000000000",
  43865=>"001101111",
  43866=>"000000000",
  43867=>"001001111",
  43868=>"000000000",
  43869=>"110100100",
  43870=>"010000111",
  43871=>"100000000",
  43872=>"000011111",
  43873=>"010111111",
  43874=>"111110100",
  43875=>"111101001",
  43876=>"000000111",
  43877=>"000000000",
  43878=>"011011000",
  43879=>"000001111",
  43880=>"111110110",
  43881=>"111011111",
  43882=>"000000000",
  43883=>"111001000",
  43884=>"111111111",
  43885=>"111111001",
  43886=>"000000000",
  43887=>"111111111",
  43888=>"111111111",
  43889=>"000000000",
  43890=>"000000111",
  43891=>"110000000",
  43892=>"000100100",
  43893=>"100011111",
  43894=>"011111001",
  43895=>"110111111",
  43896=>"011001000",
  43897=>"000000001",
  43898=>"111111110",
  43899=>"011011111",
  43900=>"111111000",
  43901=>"110000000",
  43902=>"110111111",
  43903=>"000000000",
  43904=>"110111000",
  43905=>"101001111",
  43906=>"101101000",
  43907=>"111111110",
  43908=>"111111111",
  43909=>"111111111",
  43910=>"011000100",
  43911=>"100100110",
  43912=>"001001101",
  43913=>"101111111",
  43914=>"100000000",
  43915=>"001001111",
  43916=>"001111000",
  43917=>"111111110",
  43918=>"000000000",
  43919=>"000000000",
  43920=>"000000000",
  43921=>"000000000",
  43922=>"000010111",
  43923=>"110000000",
  43924=>"111111111",
  43925=>"000000000",
  43926=>"011001001",
  43927=>"000000001",
  43928=>"100100101",
  43929=>"011101000",
  43930=>"110111111",
  43931=>"111111000",
  43932=>"100100000",
  43933=>"011111111",
  43934=>"000111111",
  43935=>"000000011",
  43936=>"000000000",
  43937=>"010001011",
  43938=>"011111010",
  43939=>"000001001",
  43940=>"011010000",
  43941=>"110001000",
  43942=>"000000000",
  43943=>"000010000",
  43944=>"000000000",
  43945=>"111111111",
  43946=>"110000001",
  43947=>"010111111",
  43948=>"000111111",
  43949=>"111010000",
  43950=>"111000110",
  43951=>"110100111",
  43952=>"010010111",
  43953=>"000000111",
  43954=>"111110111",
  43955=>"011011000",
  43956=>"111111111",
  43957=>"100000010",
  43958=>"111110000",
  43959=>"000000000",
  43960=>"000001001",
  43961=>"111110011",
  43962=>"001001000",
  43963=>"010110110",
  43964=>"111001000",
  43965=>"110110110",
  43966=>"000000010",
  43967=>"011111111",
  43968=>"000000000",
  43969=>"001001011",
  43970=>"111000000",
  43971=>"011001000",
  43972=>"011000000",
  43973=>"000000000",
  43974=>"110111111",
  43975=>"111001001",
  43976=>"100111111",
  43977=>"000000100",
  43978=>"000000011",
  43979=>"000000110",
  43980=>"011111000",
  43981=>"101000000",
  43982=>"111111111",
  43983=>"111111111",
  43984=>"000000111",
  43985=>"101100100",
  43986=>"000000000",
  43987=>"001111111",
  43988=>"001001011",
  43989=>"111111111",
  43990=>"000000000",
  43991=>"111101001",
  43992=>"000000000",
  43993=>"100000000",
  43994=>"000000000",
  43995=>"111111111",
  43996=>"000001000",
  43997=>"110110000",
  43998=>"110000100",
  43999=>"000001011",
  44000=>"111111111",
  44001=>"011111100",
  44002=>"000000000",
  44003=>"110010111",
  44004=>"111111001",
  44005=>"000000000",
  44006=>"111111011",
  44007=>"111010000",
  44008=>"000000000",
  44009=>"111111010",
  44010=>"000000000",
  44011=>"111111111",
  44012=>"111111111",
  44013=>"110010000",
  44014=>"110000000",
  44015=>"100000100",
  44016=>"000110110",
  44017=>"000000000",
  44018=>"100000000",
  44019=>"000011111",
  44020=>"111111111",
  44021=>"010000000",
  44022=>"001000100",
  44023=>"000000000",
  44024=>"000000000",
  44025=>"001001101",
  44026=>"101000000",
  44027=>"000000000",
  44028=>"000111111",
  44029=>"000000000",
  44030=>"000010110",
  44031=>"010011110",
  44032=>"000001001",
  44033=>"000110111",
  44034=>"110110111",
  44035=>"111111111",
  44036=>"000100001",
  44037=>"000011011",
  44038=>"001000000",
  44039=>"111111111",
  44040=>"000000110",
  44041=>"111100101",
  44042=>"000000000",
  44043=>"000111001",
  44044=>"100100000",
  44045=>"111100000",
  44046=>"000000000",
  44047=>"011111111",
  44048=>"111111111",
  44049=>"111111111",
  44050=>"111111111",
  44051=>"000001011",
  44052=>"000000000",
  44053=>"111111111",
  44054=>"000010111",
  44055=>"111111111",
  44056=>"111111111",
  44057=>"011011000",
  44058=>"000000000",
  44059=>"111111111",
  44060=>"011000000",
  44061=>"110111000",
  44062=>"000000000",
  44063=>"111010000",
  44064=>"000000000",
  44065=>"111100111",
  44066=>"000000000",
  44067=>"101101100",
  44068=>"111111001",
  44069=>"000001001",
  44070=>"111111111",
  44071=>"000000100",
  44072=>"000000000",
  44073=>"111010000",
  44074=>"001001001",
  44075=>"111111111",
  44076=>"000000000",
  44077=>"111111111",
  44078=>"111111011",
  44079=>"101000111",
  44080=>"000000000",
  44081=>"000000100",
  44082=>"111111111",
  44083=>"100100000",
  44084=>"000000000",
  44085=>"000000000",
  44086=>"000011111",
  44087=>"100111111",
  44088=>"011011101",
  44089=>"011001000",
  44090=>"000000000",
  44091=>"011111111",
  44092=>"000000000",
  44093=>"000001001",
  44094=>"000000000",
  44095=>"011001000",
  44096=>"111000000",
  44097=>"100100110",
  44098=>"111010110",
  44099=>"011001001",
  44100=>"000000000",
  44101=>"000000000",
  44102=>"011111000",
  44103=>"000000000",
  44104=>"011001000",
  44105=>"000000001",
  44106=>"111111111",
  44107=>"100001001",
  44108=>"011000100",
  44109=>"110000101",
  44110=>"000000011",
  44111=>"000010000",
  44112=>"000000000",
  44113=>"000100100",
  44114=>"111011101",
  44115=>"011111111",
  44116=>"000011111",
  44117=>"000000100",
  44118=>"110000000",
  44119=>"000001011",
  44120=>"001001011",
  44121=>"111001001",
  44122=>"111111111",
  44123=>"111111011",
  44124=>"000000000",
  44125=>"000111111",
  44126=>"111111111",
  44127=>"111111111",
  44128=>"000000000",
  44129=>"101111111",
  44130=>"110011011",
  44131=>"111100100",
  44132=>"000000100",
  44133=>"111111111",
  44134=>"101100100",
  44135=>"100000000",
  44136=>"000000000",
  44137=>"000000000",
  44138=>"111011111",
  44139=>"111111111",
  44140=>"100011111",
  44141=>"111111001",
  44142=>"000101111",
  44143=>"010010000",
  44144=>"100000000",
  44145=>"011011000",
  44146=>"000110111",
  44147=>"110100110",
  44148=>"111111111",
  44149=>"000000000",
  44150=>"000000110",
  44151=>"000000000",
  44152=>"000001001",
  44153=>"000000000",
  44154=>"111110100",
  44155=>"001000000",
  44156=>"000010010",
  44157=>"000001001",
  44158=>"000000000",
  44159=>"011111011",
  44160=>"000000000",
  44161=>"001011111",
  44162=>"000000111",
  44163=>"111111111",
  44164=>"111111111",
  44165=>"111000000",
  44166=>"111111111",
  44167=>"111111111",
  44168=>"100000000",
  44169=>"000000000",
  44170=>"000000000",
  44171=>"111111111",
  44172=>"111111101",
  44173=>"000000100",
  44174=>"111111110",
  44175=>"000001001",
  44176=>"000000000",
  44177=>"100011111",
  44178=>"111001011",
  44179=>"001000000",
  44180=>"011011011",
  44181=>"000011001",
  44182=>"000000110",
  44183=>"000000000",
  44184=>"111111001",
  44185=>"111110001",
  44186=>"000000111",
  44187=>"011001000",
  44188=>"111111110",
  44189=>"001011011",
  44190=>"011011001",
  44191=>"111111111",
  44192=>"111000000",
  44193=>"000000000",
  44194=>"000001101",
  44195=>"000000001",
  44196=>"000000100",
  44197=>"011010100",
  44198=>"000000000",
  44199=>"001011011",
  44200=>"001011111",
  44201=>"000000000",
  44202=>"000000000",
  44203=>"011101101",
  44204=>"001000000",
  44205=>"011011011",
  44206=>"111111111",
  44207=>"000000101",
  44208=>"011011000",
  44209=>"110111111",
  44210=>"111111111",
  44211=>"111000001",
  44212=>"000100100",
  44213=>"100111111",
  44214=>"000111111",
  44215=>"000011111",
  44216=>"011001001",
  44217=>"111101000",
  44218=>"000000100",
  44219=>"001011111",
  44220=>"110110010",
  44221=>"001011111",
  44222=>"111111111",
  44223=>"000000101",
  44224=>"000000000",
  44225=>"111111111",
  44226=>"000011111",
  44227=>"011111111",
  44228=>"000100000",
  44229=>"111111111",
  44230=>"111011000",
  44231=>"000000001",
  44232=>"111111011",
  44233=>"000000000",
  44234=>"111111111",
  44235=>"000000000",
  44236=>"011011111",
  44237=>"000100111",
  44238=>"001001011",
  44239=>"000000010",
  44240=>"100110101",
  44241=>"000000000",
  44242=>"111111111",
  44243=>"000000000",
  44244=>"111111100",
  44245=>"001000000",
  44246=>"111111111",
  44247=>"101111111",
  44248=>"001001000",
  44249=>"011011001",
  44250=>"111111011",
  44251=>"000000001",
  44252=>"100000100",
  44253=>"000100100",
  44254=>"000010000",
  44255=>"001011111",
  44256=>"011011011",
  44257=>"111110100",
  44258=>"000000000",
  44259=>"111111111",
  44260=>"011001001",
  44261=>"100110111",
  44262=>"111111111",
  44263=>"100101111",
  44264=>"011011011",
  44265=>"000101000",
  44266=>"001011011",
  44267=>"111111111",
  44268=>"000000000",
  44269=>"000000000",
  44270=>"101111111",
  44271=>"000000000",
  44272=>"111111001",
  44273=>"100000000",
  44274=>"111101111",
  44275=>"000010010",
  44276=>"111111100",
  44277=>"000001000",
  44278=>"010110111",
  44279=>"110010011",
  44280=>"111010000",
  44281=>"110000000",
  44282=>"000100000",
  44283=>"100100100",
  44284=>"000001011",
  44285=>"010111000",
  44286=>"000011011",
  44287=>"001011000",
  44288=>"000011101",
  44289=>"010010011",
  44290=>"111111011",
  44291=>"000000000",
  44292=>"111000000",
  44293=>"000001001",
  44294=>"000000000",
  44295=>"011011111",
  44296=>"000000001",
  44297=>"000000000",
  44298=>"111111011",
  44299=>"001011111",
  44300=>"101000100",
  44301=>"111111111",
  44302=>"110011101",
  44303=>"011111000",
  44304=>"011011011",
  44305=>"000000110",
  44306=>"111111111",
  44307=>"000000001",
  44308=>"100110111",
  44309=>"111001111",
  44310=>"111111011",
  44311=>"111001001",
  44312=>"000000111",
  44313=>"110111100",
  44314=>"000000000",
  44315=>"111111111",
  44316=>"111110100",
  44317=>"100100100",
  44318=>"000000000",
  44319=>"111101001",
  44320=>"101111111",
  44321=>"111111111",
  44322=>"000000111",
  44323=>"111111101",
  44324=>"111111111",
  44325=>"111111101",
  44326=>"101111111",
  44327=>"000011011",
  44328=>"110110111",
  44329=>"000000000",
  44330=>"111001000",
  44331=>"100101111",
  44332=>"111111111",
  44333=>"001101111",
  44334=>"001101001",
  44335=>"000000011",
  44336=>"111011011",
  44337=>"111011111",
  44338=>"000000100",
  44339=>"000000000",
  44340=>"101000111",
  44341=>"000111101",
  44342=>"000000011",
  44343=>"111111111",
  44344=>"111100100",
  44345=>"001000000",
  44346=>"000000111",
  44347=>"010111111",
  44348=>"011001011",
  44349=>"000001001",
  44350=>"111111111",
  44351=>"001011000",
  44352=>"011100000",
  44353=>"000000000",
  44354=>"101011111",
  44355=>"000000000",
  44356=>"001000000",
  44357=>"111111100",
  44358=>"000000000",
  44359=>"000111111",
  44360=>"011111000",
  44361=>"110110110",
  44362=>"101001001",
  44363=>"111111011",
  44364=>"000000000",
  44365=>"000000000",
  44366=>"111111001",
  44367=>"000010000",
  44368=>"100011001",
  44369=>"011111000",
  44370=>"010000000",
  44371=>"000000000",
  44372=>"000100100",
  44373=>"011011011",
  44374=>"000000010",
  44375=>"010110111",
  44376=>"111111111",
  44377=>"111111111",
  44378=>"001000000",
  44379=>"011111111",
  44380=>"000000000",
  44381=>"000000000",
  44382=>"000000011",
  44383=>"111110100",
  44384=>"111111111",
  44385=>"111111111",
  44386=>"000100110",
  44387=>"011111111",
  44388=>"011111111",
  44389=>"000001111",
  44390=>"100100100",
  44391=>"111111011",
  44392=>"110010010",
  44393=>"110110111",
  44394=>"000100100",
  44395=>"000010010",
  44396=>"011011011",
  44397=>"001000100",
  44398=>"111111111",
  44399=>"011000000",
  44400=>"111111111",
  44401=>"111000000",
  44402=>"000000000",
  44403=>"011001000",
  44404=>"111111111",
  44405=>"111111011",
  44406=>"011011111",
  44407=>"111111111",
  44408=>"000000110",
  44409=>"010110110",
  44410=>"000000000",
  44411=>"011011001",
  44412=>"000100000",
  44413=>"111111111",
  44414=>"111111111",
  44415=>"000000000",
  44416=>"111011001",
  44417=>"000000000",
  44418=>"000110001",
  44419=>"001000011",
  44420=>"000000001",
  44421=>"000111111",
  44422=>"000011011",
  44423=>"111001001",
  44424=>"100100100",
  44425=>"000000000",
  44426=>"011111111",
  44427=>"000000110",
  44428=>"111111111",
  44429=>"001001001",
  44430=>"010110000",
  44431=>"000000000",
  44432=>"100000000",
  44433=>"100000100",
  44434=>"111101101",
  44435=>"110110000",
  44436=>"000000000",
  44437=>"000010000",
  44438=>"110100111",
  44439=>"111111111",
  44440=>"000000001",
  44441=>"001011111",
  44442=>"000100100",
  44443=>"011001000",
  44444=>"111111111",
  44445=>"000000000",
  44446=>"000000000",
  44447=>"111111011",
  44448=>"100100100",
  44449=>"110111001",
  44450=>"000011111",
  44451=>"000000110",
  44452=>"111111111",
  44453=>"111000000",
  44454=>"000000000",
  44455=>"111111101",
  44456=>"111111000",
  44457=>"000000000",
  44458=>"000100111",
  44459=>"000000011",
  44460=>"111111111",
  44461=>"111011010",
  44462=>"000011011",
  44463=>"000001001",
  44464=>"010000000",
  44465=>"011011000",
  44466=>"011111111",
  44467=>"111111111",
  44468=>"111111001",
  44469=>"111111111",
  44470=>"111111111",
  44471=>"001000000",
  44472=>"011101101",
  44473=>"111111011",
  44474=>"000100111",
  44475=>"000000000",
  44476=>"111111111",
  44477=>"111110100",
  44478=>"000000111",
  44479=>"010000000",
  44480=>"001000000",
  44481=>"110111111",
  44482=>"000000000",
  44483=>"000011111",
  44484=>"111011000",
  44485=>"001001100",
  44486=>"000000000",
  44487=>"110000111",
  44488=>"000100111",
  44489=>"000111000",
  44490=>"000000000",
  44491=>"000000000",
  44492=>"101111110",
  44493=>"000000000",
  44494=>"011001001",
  44495=>"110100111",
  44496=>"100101111",
  44497=>"011011001",
  44498=>"000000000",
  44499=>"010110110",
  44500=>"000000000",
  44501=>"111001111",
  44502=>"001000000",
  44503=>"000000000",
  44504=>"011111000",
  44505=>"100000000",
  44506=>"101000000",
  44507=>"111111111",
  44508=>"110111111",
  44509=>"001011001",
  44510=>"000011011",
  44511=>"000010010",
  44512=>"010000000",
  44513=>"001000001",
  44514=>"000010000",
  44515=>"100000001",
  44516=>"111111111",
  44517=>"000000111",
  44518=>"000001000",
  44519=>"110100110",
  44520=>"001011001",
  44521=>"111111111",
  44522=>"000010011",
  44523=>"111111111",
  44524=>"001111111",
  44525=>"111101100",
  44526=>"000000000",
  44527=>"000000000",
  44528=>"110111111",
  44529=>"011111111",
  44530=>"011011111",
  44531=>"011011011",
  44532=>"000000000",
  44533=>"110001011",
  44534=>"111111110",
  44535=>"100011011",
  44536=>"110111111",
  44537=>"011011001",
  44538=>"011111111",
  44539=>"101001000",
  44540=>"011010000",
  44541=>"000000000",
  44542=>"011011011",
  44543=>"000000011",
  44544=>"100111111",
  44545=>"111111011",
  44546=>"111100000",
  44547=>"111111111",
  44548=>"001111111",
  44549=>"000000000",
  44550=>"111000000",
  44551=>"000000000",
  44552=>"000101111",
  44553=>"111111000",
  44554=>"111100000",
  44555=>"000000001",
  44556=>"001000000",
  44557=>"000010100",
  44558=>"110100000",
  44559=>"111111111",
  44560=>"111011001",
  44561=>"100111010",
  44562=>"000000000",
  44563=>"001101111",
  44564=>"100000111",
  44565=>"111110111",
  44566=>"010000000",
  44567=>"000001001",
  44568=>"101010010",
  44569=>"111111101",
  44570=>"000011000",
  44571=>"111111010",
  44572=>"011011111",
  44573=>"011000100",
  44574=>"000010000",
  44575=>"000000110",
  44576=>"000000001",
  44577=>"100000000",
  44578=>"001001101",
  44579=>"110111110",
  44580=>"001000000",
  44581=>"000001000",
  44582=>"011010000",
  44583=>"010110111",
  44584=>"111111111",
  44585=>"011011111",
  44586=>"000000000",
  44587=>"110111100",
  44588=>"000000000",
  44589=>"000000000",
  44590=>"110111111",
  44591=>"111001011",
  44592=>"001001001",
  44593=>"000000000",
  44594=>"000000110",
  44595=>"111111111",
  44596=>"000100000",
  44597=>"111101101",
  44598=>"011000001",
  44599=>"000000101",
  44600=>"111111011",
  44601=>"110000000",
  44602=>"111111111",
  44603=>"111111010",
  44604=>"100110111",
  44605=>"111011111",
  44606=>"111111111",
  44607=>"000000000",
  44608=>"101001111",
  44609=>"110000000",
  44610=>"111111000",
  44611=>"111110111",
  44612=>"111001001",
  44613=>"001011111",
  44614=>"000011011",
  44615=>"000000100",
  44616=>"111110110",
  44617=>"000000000",
  44618=>"000000000",
  44619=>"000000111",
  44620=>"110111111",
  44621=>"011011111",
  44622=>"111111000",
  44623=>"000000000",
  44624=>"100000000",
  44625=>"010000000",
  44626=>"000000000",
  44627=>"101101001",
  44628=>"111111111",
  44629=>"010000000",
  44630=>"100000111",
  44631=>"100111111",
  44632=>"001111111",
  44633=>"000110000",
  44634=>"110110110",
  44635=>"111111001",
  44636=>"001100100",
  44637=>"110111111",
  44638=>"000000000",
  44639=>"110000000",
  44640=>"111011001",
  44641=>"111111111",
  44642=>"000000000",
  44643=>"000000000",
  44644=>"000100001",
  44645=>"111010000",
  44646=>"000000110",
  44647=>"000000000",
  44648=>"111010010",
  44649=>"111111110",
  44650=>"111111111",
  44651=>"110111111",
  44652=>"100101101",
  44653=>"000000011",
  44654=>"001000101",
  44655=>"111111111",
  44656=>"111010000",
  44657=>"100000011",
  44658=>"010100100",
  44659=>"000000000",
  44660=>"001000000",
  44661=>"110000000",
  44662=>"110111000",
  44663=>"111111111",
  44664=>"110111111",
  44665=>"001000001",
  44666=>"000011011",
  44667=>"111111111",
  44668=>"000100000",
  44669=>"000111111",
  44670=>"000000000",
  44671=>"000000110",
  44672=>"111111111",
  44673=>"000000001",
  44674=>"000000000",
  44675=>"000000000",
  44676=>"000000100",
  44677=>"111111111",
  44678=>"111111111",
  44679=>"001011000",
  44680=>"000000000",
  44681=>"111111111",
  44682=>"000011111",
  44683=>"001011111",
  44684=>"111111111",
  44685=>"111111111",
  44686=>"100000000",
  44687=>"111111111",
  44688=>"000000000",
  44689=>"000000100",
  44690=>"100001001",
  44691=>"111111111",
  44692=>"000001001",
  44693=>"011111111",
  44694=>"000000000",
  44695=>"000000000",
  44696=>"111011111",
  44697=>"100100111",
  44698=>"000000000",
  44699=>"011011001",
  44700=>"100100100",
  44701=>"111111000",
  44702=>"111000101",
  44703=>"111111111",
  44704=>"111111111",
  44705=>"110000000",
  44706=>"111110100",
  44707=>"111111000",
  44708=>"011111111",
  44709=>"111010011",
  44710=>"000000000",
  44711=>"001011010",
  44712=>"000000000",
  44713=>"000000000",
  44714=>"000100110",
  44715=>"000000000",
  44716=>"110010111",
  44717=>"111111111",
  44718=>"001111111",
  44719=>"000000000",
  44720=>"110011011",
  44721=>"101101101",
  44722=>"011000010",
  44723=>"000000000",
  44724=>"110111000",
  44725=>"100011000",
  44726=>"000010111",
  44727=>"100000000",
  44728=>"100111111",
  44729=>"000000000",
  44730=>"000011000",
  44731=>"110110110",
  44732=>"111111111",
  44733=>"000000111",
  44734=>"000000000",
  44735=>"111111111",
  44736=>"000000000",
  44737=>"011001001",
  44738=>"000000000",
  44739=>"111101111",
  44740=>"000000000",
  44741=>"000000000",
  44742=>"000000110",
  44743=>"111111111",
  44744=>"111111111",
  44745=>"000000111",
  44746=>"101111111",
  44747=>"011001000",
  44748=>"111000110",
  44749=>"000000100",
  44750=>"000011111",
  44751=>"101111111",
  44752=>"000000010",
  44753=>"111111111",
  44754=>"000000000",
  44755=>"001001111",
  44756=>"111111111",
  44757=>"111111000",
  44758=>"000000110",
  44759=>"000100001",
  44760=>"000001011",
  44761=>"111111101",
  44762=>"111111111",
  44763=>"111111000",
  44764=>"111111111",
  44765=>"111111110",
  44766=>"111111111",
  44767=>"001001111",
  44768=>"111111111",
  44769=>"111111111",
  44770=>"001011000",
  44771=>"101000000",
  44772=>"100111111",
  44773=>"111110111",
  44774=>"100000000",
  44775=>"110111111",
  44776=>"000000000",
  44777=>"000111000",
  44778=>"111101000",
  44779=>"011001111",
  44780=>"000000000",
  44781=>"111111111",
  44782=>"000000001",
  44783=>"000000000",
  44784=>"001111111",
  44785=>"000000011",
  44786=>"000000100",
  44787=>"011000110",
  44788=>"111111100",
  44789=>"110000000",
  44790=>"001001111",
  44791=>"000000001",
  44792=>"000000000",
  44793=>"111111111",
  44794=>"111011111",
  44795=>"111111111",
  44796=>"111111011",
  44797=>"111000000",
  44798=>"111000101",
  44799=>"111000000",
  44800=>"011011000",
  44801=>"011011010",
  44802=>"111111111",
  44803=>"000000000",
  44804=>"000001011",
  44805=>"110110011",
  44806=>"000000000",
  44807=>"111000111",
  44808=>"011000000",
  44809=>"000000000",
  44810=>"111111111",
  44811=>"110110000",
  44812=>"000000110",
  44813=>"111011111",
  44814=>"011000010",
  44815=>"000000000",
  44816=>"111111011",
  44817=>"000000000",
  44818=>"101000000",
  44819=>"000000110",
  44820=>"000111111",
  44821=>"011000000",
  44822=>"110100000",
  44823=>"000000000",
  44824=>"110110000",
  44825=>"110110111",
  44826=>"000000000",
  44827=>"110110010",
  44828=>"000000000",
  44829=>"111111101",
  44830=>"101111111",
  44831=>"111111111",
  44832=>"000100110",
  44833=>"111101011",
  44834=>"011000111",
  44835=>"110110000",
  44836=>"010110010",
  44837=>"000000000",
  44838=>"111000000",
  44839=>"110100111",
  44840=>"111111111",
  44841=>"110000000",
  44842=>"111111111",
  44843=>"101111001",
  44844=>"111000101",
  44845=>"111000000",
  44846=>"000000000",
  44847=>"111111111",
  44848=>"000000000",
  44849=>"111011011",
  44850=>"000000100",
  44851=>"010111111",
  44852=>"000000000",
  44853=>"000111111",
  44854=>"111111111",
  44855=>"010111011",
  44856=>"011000000",
  44857=>"111010000",
  44858=>"111011111",
  44859=>"001001010",
  44860=>"011000111",
  44861=>"110100001",
  44862=>"111111111",
  44863=>"111110011",
  44864=>"000111000",
  44865=>"101011000",
  44866=>"111111111",
  44867=>"111111111",
  44868=>"000000000",
  44869=>"100000000",
  44870=>"111111111",
  44871=>"111111111",
  44872=>"111111111",
  44873=>"000000000",
  44874=>"010000000",
  44875=>"000000000",
  44876=>"000000000",
  44877=>"010000000",
  44878=>"111000000",
  44879=>"100111011",
  44880=>"001101011",
  44881=>"000011010",
  44882=>"111000000",
  44883=>"000000111",
  44884=>"001001111",
  44885=>"001000000",
  44886=>"000000000",
  44887=>"000011111",
  44888=>"111111111",
  44889=>"000000000",
  44890=>"111111010",
  44891=>"111110111",
  44892=>"110111111",
  44893=>"100000011",
  44894=>"000000000",
  44895=>"111110110",
  44896=>"001000000",
  44897=>"000100100",
  44898=>"001011010",
  44899=>"000000000",
  44900=>"001001001",
  44901=>"001000000",
  44902=>"000000000",
  44903=>"110000000",
  44904=>"011000000",
  44905=>"000000000",
  44906=>"001111111",
  44907=>"100110100",
  44908=>"111001001",
  44909=>"000011000",
  44910=>"111101111",
  44911=>"111001000",
  44912=>"000110100",
  44913=>"000000000",
  44914=>"011011110",
  44915=>"111111111",
  44916=>"111111111",
  44917=>"000000000",
  44918=>"000000000",
  44919=>"011111111",
  44920=>"000000000",
  44921=>"000000111",
  44922=>"000000011",
  44923=>"111101101",
  44924=>"011011011",
  44925=>"111110111",
  44926=>"011110110",
  44927=>"100000000",
  44928=>"001000000",
  44929=>"011010111",
  44930=>"110111111",
  44931=>"000000000",
  44932=>"100000111",
  44933=>"111111000",
  44934=>"000000011",
  44935=>"010111111",
  44936=>"000010000",
  44937=>"111001000",
  44938=>"011000000",
  44939=>"111001000",
  44940=>"111001011",
  44941=>"110111111",
  44942=>"000000000",
  44943=>"111111111",
  44944=>"000000111",
  44945=>"111000111",
  44946=>"110111111",
  44947=>"100100011",
  44948=>"111111010",
  44949=>"000001000",
  44950=>"100100110",
  44951=>"001100100",
  44952=>"111110000",
  44953=>"001111111",
  44954=>"001110100",
  44955=>"000000000",
  44956=>"111111111",
  44957=>"111111111",
  44958=>"011111100",
  44959=>"001000001",
  44960=>"011011011",
  44961=>"011011011",
  44962=>"111001111",
  44963=>"010000111",
  44964=>"011000111",
  44965=>"111111111",
  44966=>"111111110",
  44967=>"000000001",
  44968=>"111111111",
  44969=>"010010010",
  44970=>"000000000",
  44971=>"000000000",
  44972=>"111001111",
  44973=>"111101000",
  44974=>"011011111",
  44975=>"100110111",
  44976=>"000111111",
  44977=>"111011011",
  44978=>"000000000",
  44979=>"111111111",
  44980=>"110000000",
  44981=>"011111011",
  44982=>"100100111",
  44983=>"110111111",
  44984=>"000000000",
  44985=>"100000000",
  44986=>"111111000",
  44987=>"111111111",
  44988=>"111111111",
  44989=>"000000000",
  44990=>"110000000",
  44991=>"010110110",
  44992=>"000000000",
  44993=>"000000000",
  44994=>"111000000",
  44995=>"000000000",
  44996=>"100110111",
  44997=>"111110110",
  44998=>"010010000",
  44999=>"111111110",
  45000=>"111000000",
  45001=>"001000000",
  45002=>"111110000",
  45003=>"000000000",
  45004=>"010000110",
  45005=>"000000000",
  45006=>"000000000",
  45007=>"000000000",
  45008=>"000000000",
  45009=>"100100010",
  45010=>"000000001",
  45011=>"000000000",
  45012=>"001101111",
  45013=>"110010111",
  45014=>"111111100",
  45015=>"100000100",
  45016=>"111110000",
  45017=>"111000000",
  45018=>"111000000",
  45019=>"111111000",
  45020=>"100100110",
  45021=>"111011001",
  45022=>"000111000",
  45023=>"011001110",
  45024=>"110100000",
  45025=>"001001111",
  45026=>"001000011",
  45027=>"111111111",
  45028=>"111101101",
  45029=>"110110111",
  45030=>"000010000",
  45031=>"110111111",
  45032=>"000000000",
  45033=>"111011111",
  45034=>"111111111",
  45035=>"110110010",
  45036=>"110110000",
  45037=>"100110000",
  45038=>"001111111",
  45039=>"100100110",
  45040=>"000110111",
  45041=>"111101001",
  45042=>"111100111",
  45043=>"000000000",
  45044=>"001000000",
  45045=>"101101111",
  45046=>"001011000",
  45047=>"000000110",
  45048=>"000000000",
  45049=>"001101111",
  45050=>"011000000",
  45051=>"000000000",
  45052=>"100000001",
  45053=>"111000101",
  45054=>"011000010",
  45055=>"000000000",
  45056=>"111111111",
  45057=>"111000111",
  45058=>"101000100",
  45059=>"111111000",
  45060=>"111111111",
  45061=>"101000000",
  45062=>"111111111",
  45063=>"000000001",
  45064=>"111110110",
  45065=>"100111111",
  45066=>"111110111",
  45067=>"111011001",
  45068=>"000110111",
  45069=>"110000011",
  45070=>"100100110",
  45071=>"110111101",
  45072=>"111110110",
  45073=>"111110110",
  45074=>"000111111",
  45075=>"100000000",
  45076=>"001000000",
  45077=>"000000000",
  45078=>"000001011",
  45079=>"000000000",
  45080=>"100000000",
  45081=>"001000100",
  45082=>"111111011",
  45083=>"111111001",
  45084=>"111111000",
  45085=>"000100110",
  45086=>"110100000",
  45087=>"000010000",
  45088=>"000111111",
  45089=>"110111111",
  45090=>"111111111",
  45091=>"001000101",
  45092=>"001000000",
  45093=>"110100100",
  45094=>"100000011",
  45095=>"000000100",
  45096=>"101101001",
  45097=>"000000101",
  45098=>"001000100",
  45099=>"000100100",
  45100=>"111111111",
  45101=>"111111010",
  45102=>"100000100",
  45103=>"000101101",
  45104=>"000000000",
  45105=>"100100000",
  45106=>"111111000",
  45107=>"100000111",
  45108=>"100101000",
  45109=>"000010010",
  45110=>"011000000",
  45111=>"001000000",
  45112=>"000100000",
  45113=>"011011111",
  45114=>"000111111",
  45115=>"110100111",
  45116=>"111000000",
  45117=>"111111111",
  45118=>"011111111",
  45119=>"000000000",
  45120=>"010000001",
  45121=>"111111001",
  45122=>"111001101",
  45123=>"011111111",
  45124=>"000110011",
  45125=>"001001110",
  45126=>"000000000",
  45127=>"000000000",
  45128=>"000000000",
  45129=>"000111111",
  45130=>"111100000",
  45131=>"101111111",
  45132=>"000000000",
  45133=>"111011111",
  45134=>"010011011",
  45135=>"110101001",
  45136=>"000000001",
  45137=>"000111110",
  45138=>"000000011",
  45139=>"111111110",
  45140=>"100100000",
  45141=>"000000001",
  45142=>"111111000",
  45143=>"000000000",
  45144=>"011111111",
  45145=>"111100111",
  45146=>"000000000",
  45147=>"001011011",
  45148=>"101000101",
  45149=>"000000000",
  45150=>"111110111",
  45151=>"100000001",
  45152=>"111111111",
  45153=>"000001111",
  45154=>"101100010",
  45155=>"111111111",
  45156=>"111111110",
  45157=>"110000000",
  45158=>"010000111",
  45159=>"110100100",
  45160=>"111111111",
  45161=>"000000000",
  45162=>"000011010",
  45163=>"001111111",
  45164=>"111111111",
  45165=>"111111111",
  45166=>"011001111",
  45167=>"111111111",
  45168=>"000000010",
  45169=>"000000100",
  45170=>"000000000",
  45171=>"111111000",
  45172=>"010111110",
  45173=>"000110100",
  45174=>"000000000",
  45175=>"111111111",
  45176=>"100101100",
  45177=>"111110100",
  45178=>"111100100",
  45179=>"000000001",
  45180=>"100000000",
  45181=>"000000000",
  45182=>"111100111",
  45183=>"000000000",
  45184=>"111111111",
  45185=>"011011001",
  45186=>"110100001",
  45187=>"100100111",
  45188=>"011001001",
  45189=>"000000000",
  45190=>"110100000",
  45191=>"000000000",
  45192=>"111111111",
  45193=>"111111110",
  45194=>"111111111",
  45195=>"011010110",
  45196=>"001000000",
  45197=>"000000100",
  45198=>"000010011",
  45199=>"111111000",
  45200=>"001000000",
  45201=>"000000000",
  45202=>"000111111",
  45203=>"001001000",
  45204=>"100000000",
  45205=>"000010111",
  45206=>"111111101",
  45207=>"000000000",
  45208=>"101000000",
  45209=>"101001111",
  45210=>"000000111",
  45211=>"110000000",
  45212=>"011111111",
  45213=>"111000000",
  45214=>"110110111",
  45215=>"110111000",
  45216=>"111111111",
  45217=>"110010111",
  45218=>"111111100",
  45219=>"000100111",
  45220=>"000000001",
  45221=>"100111111",
  45222=>"111111000",
  45223=>"011011000",
  45224=>"000110111",
  45225=>"111001111",
  45226=>"001000000",
  45227=>"000000000",
  45228=>"111111000",
  45229=>"000000100",
  45230=>"100000100",
  45231=>"000100111",
  45232=>"000111111",
  45233=>"100110111",
  45234=>"111111111",
  45235=>"111101000",
  45236=>"111000000",
  45237=>"111000001",
  45238=>"000000000",
  45239=>"001101111",
  45240=>"101001101",
  45241=>"111111111",
  45242=>"111100101",
  45243=>"111011001",
  45244=>"000000000",
  45245=>"111111111",
  45246=>"110100000",
  45247=>"000110101",
  45248=>"000000100",
  45249=>"111011010",
  45250=>"000110000",
  45251=>"000000000",
  45252=>"000001001",
  45253=>"000000000",
  45254=>"000001011",
  45255=>"000000000",
  45256=>"110110111",
  45257=>"101000000",
  45258=>"111111001",
  45259=>"000001001",
  45260=>"110000000",
  45261=>"000000000",
  45262=>"010110111",
  45263=>"111110010",
  45264=>"000000100",
  45265=>"111000101",
  45266=>"111000000",
  45267=>"000100000",
  45268=>"000000000",
  45269=>"000001100",
  45270=>"111000000",
  45271=>"100000000",
  45272=>"010000000",
  45273=>"111111111",
  45274=>"111111111",
  45275=>"000000011",
  45276=>"101101100",
  45277=>"000000000",
  45278=>"001001000",
  45279=>"111111111",
  45280=>"100100000",
  45281=>"000000000",
  45282=>"110110110",
  45283=>"000010111",
  45284=>"000000000",
  45285=>"100110111",
  45286=>"011110110",
  45287=>"000000111",
  45288=>"100100111",
  45289=>"111110010",
  45290=>"010111111",
  45291=>"001000000",
  45292=>"111000000",
  45293=>"000000000",
  45294=>"111111101",
  45295=>"101000000",
  45296=>"111111000",
  45297=>"000000111",
  45298=>"001001000",
  45299=>"001000000",
  45300=>"111011111",
  45301=>"011000000",
  45302=>"011000000",
  45303=>"111111110",
  45304=>"111111001",
  45305=>"111111111",
  45306=>"111111011",
  45307=>"000000000",
  45308=>"000001101",
  45309=>"000001000",
  45310=>"000000000",
  45311=>"010110000",
  45312=>"111100100",
  45313=>"011001001",
  45314=>"111110110",
  45315=>"000001111",
  45316=>"111111110",
  45317=>"001111111",
  45318=>"000111111",
  45319=>"011011111",
  45320=>"001111110",
  45321=>"110000000",
  45322=>"100000000",
  45323=>"111111111",
  45324=>"100000100",
  45325=>"000001101",
  45326=>"110111111",
  45327=>"111111000",
  45328=>"000000000",
  45329=>"000000101",
  45330=>"000000000",
  45331=>"000000111",
  45332=>"001111111",
  45333=>"000000111",
  45334=>"000100110",
  45335=>"000011000",
  45336=>"000100100",
  45337=>"111110100",
  45338=>"000000000",
  45339=>"000010000",
  45340=>"110110110",
  45341=>"111101111",
  45342=>"000000000",
  45343=>"000000000",
  45344=>"011111010",
  45345=>"000001001",
  45346=>"011111000",
  45347=>"001111111",
  45348=>"000000111",
  45349=>"000100101",
  45350=>"100111001",
  45351=>"001000000",
  45352=>"111000000",
  45353=>"000101001",
  45354=>"000111111",
  45355=>"000000000",
  45356=>"000010010",
  45357=>"000000000",
  45358=>"111011111",
  45359=>"000000000",
  45360=>"011001000",
  45361=>"000000000",
  45362=>"011001000",
  45363=>"000010011",
  45364=>"010010000",
  45365=>"111111111",
  45366=>"111011111",
  45367=>"000111111",
  45368=>"111011000",
  45369=>"111000000",
  45370=>"111000000",
  45371=>"111000000",
  45372=>"000000000",
  45373=>"000100100",
  45374=>"111111101",
  45375=>"111111111",
  45376=>"111111111",
  45377=>"000100000",
  45378=>"000000111",
  45379=>"000100100",
  45380=>"001001111",
  45381=>"001011111",
  45382=>"111111111",
  45383=>"000111000",
  45384=>"000000000",
  45385=>"111000111",
  45386=>"000001111",
  45387=>"111001000",
  45388=>"011010000",
  45389=>"001011001",
  45390=>"111111000",
  45391=>"100100000",
  45392=>"010011011",
  45393=>"000000000",
  45394=>"111111000",
  45395=>"100101111",
  45396=>"101101001",
  45397=>"011011011",
  45398=>"111111111",
  45399=>"111111111",
  45400=>"100111111",
  45401=>"111000000",
  45402=>"111111111",
  45403=>"101000001",
  45404=>"000000000",
  45405=>"111111111",
  45406=>"111111111",
  45407=>"000000110",
  45408=>"111000000",
  45409=>"000000000",
  45410=>"011000010",
  45411=>"111111001",
  45412=>"000111111",
  45413=>"111111000",
  45414=>"001001000",
  45415=>"010001010",
  45416=>"111000011",
  45417=>"000010100",
  45418=>"111001111",
  45419=>"100100000",
  45420=>"110111111",
  45421=>"011001011",
  45422=>"000000100",
  45423=>"110101101",
  45424=>"001000111",
  45425=>"111111111",
  45426=>"000000111",
  45427=>"100111110",
  45428=>"111111111",
  45429=>"111111111",
  45430=>"111000000",
  45431=>"111111111",
  45432=>"111101000",
  45433=>"111110100",
  45434=>"101111111",
  45435=>"000000000",
  45436=>"001100101",
  45437=>"000000000",
  45438=>"000110000",
  45439=>"001111111",
  45440=>"011011001",
  45441=>"001000001",
  45442=>"100000011",
  45443=>"000000000",
  45444=>"000000000",
  45445=>"000000110",
  45446=>"001000110",
  45447=>"100000000",
  45448=>"111001001",
  45449=>"000000111",
  45450=>"000001000",
  45451=>"000000000",
  45452=>"101000111",
  45453=>"100100110",
  45454=>"111111111",
  45455=>"000000100",
  45456=>"000000000",
  45457=>"011111001",
  45458=>"100100111",
  45459=>"111111001",
  45460=>"111010010",
  45461=>"010011010",
  45462=>"001001001",
  45463=>"110000000",
  45464=>"001000101",
  45465=>"011000001",
  45466=>"000000000",
  45467=>"110101110",
  45468=>"000000000",
  45469=>"000000000",
  45470=>"111001001",
  45471=>"000110011",
  45472=>"011001000",
  45473=>"100000000",
  45474=>"000001110",
  45475=>"000111111",
  45476=>"100000000",
  45477=>"010011001",
  45478=>"111100100",
  45479=>"010000001",
  45480=>"111111111",
  45481=>"011000000",
  45482=>"110111111",
  45483=>"000000000",
  45484=>"111111111",
  45485=>"000010111",
  45486=>"111111111",
  45487=>"001000001",
  45488=>"000000010",
  45489=>"000100000",
  45490=>"110111111",
  45491=>"011001000",
  45492=>"101000100",
  45493=>"010000000",
  45494=>"111111111",
  45495=>"110111111",
  45496=>"001000000",
  45497=>"000000111",
  45498=>"111101111",
  45499=>"000000000",
  45500=>"000000000",
  45501=>"000000000",
  45502=>"111111111",
  45503=>"000000000",
  45504=>"100000111",
  45505=>"111101001",
  45506=>"011111111",
  45507=>"010000110",
  45508=>"000000111",
  45509=>"010000000",
  45510=>"000000111",
  45511=>"000000111",
  45512=>"111100000",
  45513=>"100000000",
  45514=>"001011111",
  45515=>"000000000",
  45516=>"000000000",
  45517=>"111111111",
  45518=>"000000001",
  45519=>"011011111",
  45520=>"111111001",
  45521=>"100000000",
  45522=>"000000000",
  45523=>"000000001",
  45524=>"010000000",
  45525=>"001001001",
  45526=>"000111001",
  45527=>"100110110",
  45528=>"111000000",
  45529=>"001001000",
  45530=>"001000001",
  45531=>"110000000",
  45532=>"000101111",
  45533=>"111111111",
  45534=>"111111001",
  45535=>"100100000",
  45536=>"100000000",
  45537=>"011111111",
  45538=>"001001001",
  45539=>"110001000",
  45540=>"111111001",
  45541=>"000000110",
  45542=>"001001111",
  45543=>"001000101",
  45544=>"010000000",
  45545=>"000000000",
  45546=>"110110000",
  45547=>"101101101",
  45548=>"000010111",
  45549=>"000011011",
  45550=>"111111011",
  45551=>"111110010",
  45552=>"101101101",
  45553=>"000000000",
  45554=>"000000000",
  45555=>"000000000",
  45556=>"100111111",
  45557=>"000000000",
  45558=>"111111000",
  45559=>"001001011",
  45560=>"111111110",
  45561=>"000000011",
  45562=>"111111110",
  45563=>"000000000",
  45564=>"000000000",
  45565=>"000000000",
  45566=>"111000000",
  45567=>"100001101",
  45568=>"000000000",
  45569=>"000000111",
  45570=>"100100101",
  45571=>"111111111",
  45572=>"111111101",
  45573=>"111111000",
  45574=>"001000000",
  45575=>"100100100",
  45576=>"010000111",
  45577=>"100101101",
  45578=>"011000000",
  45579=>"111111000",
  45580=>"111111111",
  45581=>"110110110",
  45582=>"000000101",
  45583=>"011111111",
  45584=>"110110110",
  45585=>"011111111",
  45586=>"000000000",
  45587=>"000000000",
  45588=>"001000111",
  45589=>"111111111",
  45590=>"111111110",
  45591=>"001001001",
  45592=>"111111111",
  45593=>"111101000",
  45594=>"010110000",
  45595=>"001000001",
  45596=>"111100100",
  45597=>"000000101",
  45598=>"000000000",
  45599=>"011010111",
  45600=>"110110100",
  45601=>"011111010",
  45602=>"000000101",
  45603=>"111110111",
  45604=>"010110110",
  45605=>"000011001",
  45606=>"010110010",
  45607=>"011111001",
  45608=>"111101100",
  45609=>"000000000",
  45610=>"011000000",
  45611=>"000000001",
  45612=>"000001111",
  45613=>"110111000",
  45614=>"100001101",
  45615=>"111111111",
  45616=>"110000000",
  45617=>"000001001",
  45618=>"111111111",
  45619=>"000111000",
  45620=>"001000000",
  45621=>"111111011",
  45622=>"111111100",
  45623=>"000001110",
  45624=>"000001111",
  45625=>"000000100",
  45626=>"000001111",
  45627=>"110111111",
  45628=>"000000000",
  45629=>"001000000",
  45630=>"111001000",
  45631=>"000100100",
  45632=>"110110110",
  45633=>"100111111",
  45634=>"000000000",
  45635=>"101100100",
  45636=>"111111011",
  45637=>"011001111",
  45638=>"000000000",
  45639=>"000000101",
  45640=>"101111111",
  45641=>"000000001",
  45642=>"100111111",
  45643=>"111111111",
  45644=>"100100110",
  45645=>"010010000",
  45646=>"000000001",
  45647=>"011000000",
  45648=>"000000000",
  45649=>"100000100",
  45650=>"001101101",
  45651=>"111110110",
  45652=>"001001001",
  45653=>"011011001",
  45654=>"010001001",
  45655=>"001001111",
  45656=>"111001101",
  45657=>"100100111",
  45658=>"111111110",
  45659=>"111111111",
  45660=>"111111111",
  45661=>"010110111",
  45662=>"001101111",
  45663=>"110110110",
  45664=>"111111111",
  45665=>"000001001",
  45666=>"000101101",
  45667=>"000000000",
  45668=>"000000000",
  45669=>"100100000",
  45670=>"000110111",
  45671=>"111100000",
  45672=>"100001111",
  45673=>"111000000",
  45674=>"110011111",
  45675=>"000110110",
  45676=>"000010001",
  45677=>"001000001",
  45678=>"000110100",
  45679=>"111111111",
  45680=>"000111000",
  45681=>"111110110",
  45682=>"101001001",
  45683=>"001001001",
  45684=>"001001111",
  45685=>"111111111",
  45686=>"000000000",
  45687=>"001000100",
  45688=>"001000001",
  45689=>"000100100",
  45690=>"000000000",
  45691=>"000000000",
  45692=>"111111110",
  45693=>"001001001",
  45694=>"001001001",
  45695=>"100101111",
  45696=>"100110111",
  45697=>"011100000",
  45698=>"001011011",
  45699=>"110010000",
  45700=>"011011010",
  45701=>"000000000",
  45702=>"000001001",
  45703=>"010010001",
  45704=>"111011110",
  45705=>"111110110",
  45706=>"000001001",
  45707=>"000000000",
  45708=>"110000101",
  45709=>"111111010",
  45710=>"000000101",
  45711=>"111010111",
  45712=>"100100100",
  45713=>"111111111",
  45714=>"110110000",
  45715=>"111111011",
  45716=>"001001111",
  45717=>"011001001",
  45718=>"110110000",
  45719=>"111110110",
  45720=>"001001000",
  45721=>"111111100",
  45722=>"111001000",
  45723=>"111111111",
  45724=>"001000001",
  45725=>"001111111",
  45726=>"111111000",
  45727=>"000000111",
  45728=>"100100100",
  45729=>"000000000",
  45730=>"011000101",
  45731=>"000111111",
  45732=>"001011001",
  45733=>"011011011",
  45734=>"110110010",
  45735=>"111111000",
  45736=>"001001001",
  45737=>"000010111",
  45738=>"001001000",
  45739=>"000011111",
  45740=>"111100100",
  45741=>"111101100",
  45742=>"111111100",
  45743=>"000000100",
  45744=>"000000001",
  45745=>"110111111",
  45746=>"110111111",
  45747=>"000000000",
  45748=>"111111111",
  45749=>"000000000",
  45750=>"111111111",
  45751=>"111110111",
  45752=>"101101111",
  45753=>"110110110",
  45754=>"001011001",
  45755=>"000001000",
  45756=>"111111111",
  45757=>"001001001",
  45758=>"111111111",
  45759=>"000110110",
  45760=>"010000000",
  45761=>"010000000",
  45762=>"000000000",
  45763=>"000000000",
  45764=>"110111111",
  45765=>"101100111",
  45766=>"000000000",
  45767=>"011111111",
  45768=>"111110110",
  45769=>"000000100",
  45770=>"111111011",
  45771=>"000000000",
  45772=>"000100100",
  45773=>"011111111",
  45774=>"001000000",
  45775=>"011011000",
  45776=>"001001011",
  45777=>"000000000",
  45778=>"001001001",
  45779=>"010010000",
  45780=>"000000000",
  45781=>"100100000",
  45782=>"101100001",
  45783=>"011101101",
  45784=>"110000000",
  45785=>"111111111",
  45786=>"111100000",
  45787=>"111000001",
  45788=>"111111111",
  45789=>"110110111",
  45790=>"000000000",
  45791=>"011001001",
  45792=>"100000000",
  45793=>"110110001",
  45794=>"111111111",
  45795=>"011001000",
  45796=>"001011011",
  45797=>"110111110",
  45798=>"000000000",
  45799=>"111101101",
  45800=>"010011011",
  45801=>"011001001",
  45802=>"101000000",
  45803=>"110000000",
  45804=>"011011001",
  45805=>"000000000",
  45806=>"110111111",
  45807=>"111101000",
  45808=>"000110110",
  45809=>"111111111",
  45810=>"111111111",
  45811=>"000101100",
  45812=>"000000100",
  45813=>"011011011",
  45814=>"011111011",
  45815=>"111111100",
  45816=>"000000000",
  45817=>"000000000",
  45818=>"110111111",
  45819=>"111011011",
  45820=>"111111110",
  45821=>"000000001",
  45822=>"011011000",
  45823=>"111111111",
  45824=>"001101111",
  45825=>"111111111",
  45826=>"011011000",
  45827=>"000100110",
  45828=>"001000100",
  45829=>"000001001",
  45830=>"110110000",
  45831=>"011111111",
  45832=>"110101110",
  45833=>"111000000",
  45834=>"000001000",
  45835=>"000000000",
  45836=>"010000000",
  45837=>"111110110",
  45838=>"111111010",
  45839=>"000100101",
  45840=>"010000000",
  45841=>"010011000",
  45842=>"001001011",
  45843=>"000000000",
  45844=>"000000000",
  45845=>"111111010",
  45846=>"111110110",
  45847=>"000000100",
  45848=>"000000101",
  45849=>"000111111",
  45850=>"110110110",
  45851=>"011011111",
  45852=>"111111011",
  45853=>"110110110",
  45854=>"000001101",
  45855=>"000111111",
  45856=>"001000000",
  45857=>"111111111",
  45858=>"111111011",
  45859=>"100111111",
  45860=>"000000010",
  45861=>"000100000",
  45862=>"011011011",
  45863=>"111011110",
  45864=>"110000000",
  45865=>"010000111",
  45866=>"111111100",
  45867=>"110100100",
  45868=>"011111111",
  45869=>"000000000",
  45870=>"000000000",
  45871=>"011111111",
  45872=>"111111111",
  45873=>"111110111",
  45874=>"000000000",
  45875=>"000000111",
  45876=>"000000000",
  45877=>"111100000",
  45878=>"000000100",
  45879=>"000000100",
  45880=>"000000000",
  45881=>"110100111",
  45882=>"000000111",
  45883=>"010001000",
  45884=>"111100101",
  45885=>"111111100",
  45886=>"000000011",
  45887=>"000001001",
  45888=>"110110000",
  45889=>"111111110",
  45890=>"001001110",
  45891=>"111110110",
  45892=>"000100111",
  45893=>"000100100",
  45894=>"001001001",
  45895=>"111111111",
  45896=>"000000000",
  45897=>"010111111",
  45898=>"111111111",
  45899=>"110110100",
  45900=>"011111100",
  45901=>"000111111",
  45902=>"000000000",
  45903=>"100100110",
  45904=>"011011101",
  45905=>"000001001",
  45906=>"110111111",
  45907=>"000000000",
  45908=>"010000000",
  45909=>"001011011",
  45910=>"000010010",
  45911=>"000111111",
  45912=>"100000000",
  45913=>"111010000",
  45914=>"111010000",
  45915=>"101001101",
  45916=>"110111111",
  45917=>"000000001",
  45918=>"000011011",
  45919=>"111101000",
  45920=>"101101001",
  45921=>"101101101",
  45922=>"100101101",
  45923=>"000000100",
  45924=>"111111011",
  45925=>"001000000",
  45926=>"110000000",
  45927=>"110100000",
  45928=>"110110100",
  45929=>"000100101",
  45930=>"111111110",
  45931=>"110001001",
  45932=>"111111011",
  45933=>"001001000",
  45934=>"000000000",
  45935=>"000111111",
  45936=>"111000011",
  45937=>"000111111",
  45938=>"111111011",
  45939=>"000000000",
  45940=>"011111011",
  45941=>"111111111",
  45942=>"111111111",
  45943=>"111111111",
  45944=>"011011111",
  45945=>"111001001",
  45946=>"000000010",
  45947=>"000010000",
  45948=>"111111010",
  45949=>"000000111",
  45950=>"001001011",
  45951=>"111111111",
  45952=>"111111111",
  45953=>"011001001",
  45954=>"011011001",
  45955=>"000000001",
  45956=>"111111111",
  45957=>"000000000",
  45958=>"110111110",
  45959=>"111111111",
  45960=>"000000000",
  45961=>"101111111",
  45962=>"110111101",
  45963=>"100110110",
  45964=>"110111111",
  45965=>"000000000",
  45966=>"111111110",
  45967=>"011111111",
  45968=>"000000000",
  45969=>"010000000",
  45970=>"000000000",
  45971=>"001001001",
  45972=>"100110110",
  45973=>"011011011",
  45974=>"011001001",
  45975=>"100101001",
  45976=>"000011011",
  45977=>"111110100",
  45978=>"001101111",
  45979=>"111100000",
  45980=>"001001000",
  45981=>"011111001",
  45982=>"000000000",
  45983=>"000111110",
  45984=>"011111011",
  45985=>"001001111",
  45986=>"001110100",
  45987=>"111010100",
  45988=>"101101101",
  45989=>"110111111",
  45990=>"000000110",
  45991=>"000111111",
  45992=>"000000100",
  45993=>"111111001",
  45994=>"000000000",
  45995=>"000001001",
  45996=>"000000000",
  45997=>"001001001",
  45998=>"111110100",
  45999=>"001001011",
  46000=>"111101100",
  46001=>"110110110",
  46002=>"111000000",
  46003=>"000000000",
  46004=>"111100000",
  46005=>"111111111",
  46006=>"100101101",
  46007=>"000000010",
  46008=>"000100101",
  46009=>"010000000",
  46010=>"001000010",
  46011=>"110100000",
  46012=>"010010010",
  46013=>"100000101",
  46014=>"000000000",
  46015=>"111101101",
  46016=>"001000000",
  46017=>"000000000",
  46018=>"000111111",
  46019=>"111111111",
  46020=>"100100100",
  46021=>"000110110",
  46022=>"100001100",
  46023=>"110011011",
  46024=>"000000000",
  46025=>"001001101",
  46026=>"111111111",
  46027=>"011001000",
  46028=>"000000000",
  46029=>"111100100",
  46030=>"000000110",
  46031=>"111111111",
  46032=>"111001001",
  46033=>"000110110",
  46034=>"111110000",
  46035=>"111100111",
  46036=>"100101111",
  46037=>"001000000",
  46038=>"010111111",
  46039=>"000000000",
  46040=>"000111111",
  46041=>"001011010",
  46042=>"110010000",
  46043=>"011000000",
  46044=>"111111111",
  46045=>"000000100",
  46046=>"100110111",
  46047=>"010011011",
  46048=>"010000000",
  46049=>"010111111",
  46050=>"100000101",
  46051=>"111111101",
  46052=>"110010110",
  46053=>"111111111",
  46054=>"000000100",
  46055=>"101101111",
  46056=>"101101100",
  46057=>"000000000",
  46058=>"100110111",
  46059=>"000000000",
  46060=>"100000000",
  46061=>"000000000",
  46062=>"000000101",
  46063=>"000000000",
  46064=>"001011001",
  46065=>"010111110",
  46066=>"111111011",
  46067=>"000000000",
  46068=>"111111110",
  46069=>"011001001",
  46070=>"110100100",
  46071=>"000000000",
  46072=>"000100110",
  46073=>"000000000",
  46074=>"001001000",
  46075=>"000000100",
  46076=>"000000000",
  46077=>"100000100",
  46078=>"110000000",
  46079=>"111101001",
  46080=>"000001111",
  46081=>"111110110",
  46082=>"000000000",
  46083=>"000000101",
  46084=>"001001111",
  46085=>"010111011",
  46086=>"000111010",
  46087=>"101100000",
  46088=>"111111111",
  46089=>"111000000",
  46090=>"111111111",
  46091=>"000000000",
  46092=>"100110000",
  46093=>"001000000",
  46094=>"111111111",
  46095=>"000000000",
  46096=>"000000000",
  46097=>"001100000",
  46098=>"000000000",
  46099=>"110000000",
  46100=>"100000000",
  46101=>"000000000",
  46102=>"111011001",
  46103=>"000011001",
  46104=>"110111111",
  46105=>"000011011",
  46106=>"111111111",
  46107=>"100110100",
  46108=>"111101101",
  46109=>"000000000",
  46110=>"000000001",
  46111=>"001101000",
  46112=>"110110110",
  46113=>"111111111",
  46114=>"000000001",
  46115=>"111111111",
  46116=>"000000000",
  46117=>"000001001",
  46118=>"111111110",
  46119=>"110111000",
  46120=>"111000000",
  46121=>"000000110",
  46122=>"000000001",
  46123=>"001001000",
  46124=>"000100000",
  46125=>"000001110",
  46126=>"000000011",
  46127=>"011011111",
  46128=>"000000001",
  46129=>"000000011",
  46130=>"111000000",
  46131=>"000000111",
  46132=>"110110000",
  46133=>"000000000",
  46134=>"111111111",
  46135=>"110000011",
  46136=>"000000011",
  46137=>"011011011",
  46138=>"000000101",
  46139=>"100000110",
  46140=>"101101111",
  46141=>"111100100",
  46142=>"000000000",
  46143=>"000000101",
  46144=>"000100101",
  46145=>"101111000",
  46146=>"000000000",
  46147=>"000000101",
  46148=>"111111001",
  46149=>"000011011",
  46150=>"000100100",
  46151=>"111111010",
  46152=>"111111001",
  46153=>"111111110",
  46154=>"000001001",
  46155=>"111111111",
  46156=>"011000110",
  46157=>"001111111",
  46158=>"100110110",
  46159=>"111111111",
  46160=>"111111001",
  46161=>"001001001",
  46162=>"000000000",
  46163=>"111011011",
  46164=>"111111111",
  46165=>"100111111",
  46166=>"111100100",
  46167=>"010111111",
  46168=>"000000100",
  46169=>"000000000",
  46170=>"101101111",
  46171=>"100100100",
  46172=>"110110100",
  46173=>"111111111",
  46174=>"000001001",
  46175=>"000011111",
  46176=>"000110110",
  46177=>"000010000",
  46178=>"000000111",
  46179=>"111111111",
  46180=>"001101111",
  46181=>"111000101",
  46182=>"000000111",
  46183=>"100111111",
  46184=>"000100000",
  46185=>"110110000",
  46186=>"010111111",
  46187=>"000001111",
  46188=>"000001001",
  46189=>"000000010",
  46190=>"000000000",
  46191=>"000000111",
  46192=>"110000110",
  46193=>"000101111",
  46194=>"000100100",
  46195=>"000000000",
  46196=>"000000000",
  46197=>"110111111",
  46198=>"000000001",
  46199=>"000000000",
  46200=>"111111111",
  46201=>"001111111",
  46202=>"011001000",
  46203=>"000000000",
  46204=>"011111111",
  46205=>"000000000",
  46206=>"000000000",
  46207=>"001011000",
  46208=>"111111010",
  46209=>"000000000",
  46210=>"000000000",
  46211=>"000000000",
  46212=>"100100010",
  46213=>"000000000",
  46214=>"111011011",
  46215=>"111110000",
  46216=>"001110010",
  46217=>"010111101",
  46218=>"100100000",
  46219=>"000000000",
  46220=>"010110111",
  46221=>"111001111",
  46222=>"010111111",
  46223=>"000011011",
  46224=>"111101100",
  46225=>"000000000",
  46226=>"111001111",
  46227=>"001000101",
  46228=>"000001000",
  46229=>"100110000",
  46230=>"100111000",
  46231=>"000001001",
  46232=>"000000000",
  46233=>"111111111",
  46234=>"000000111",
  46235=>"111111111",
  46236=>"111000000",
  46237=>"110110111",
  46238=>"000110111",
  46239=>"111000000",
  46240=>"000000001",
  46241=>"111111110",
  46242=>"101111011",
  46243=>"111101111",
  46244=>"001001001",
  46245=>"000000000",
  46246=>"111111111",
  46247=>"000001101",
  46248=>"100111111",
  46249=>"111100000",
  46250=>"111111111",
  46251=>"101111000",
  46252=>"011001111",
  46253=>"001001111",
  46254=>"000000001",
  46255=>"010110000",
  46256=>"000111111",
  46257=>"010110100",
  46258=>"001111000",
  46259=>"111111100",
  46260=>"000001011",
  46261=>"000000001",
  46262=>"000100111",
  46263=>"111101000",
  46264=>"111111000",
  46265=>"000110111",
  46266=>"000001001",
  46267=>"110111111",
  46268=>"000100111",
  46269=>"110111010",
  46270=>"010111110",
  46271=>"001000001",
  46272=>"100000110",
  46273=>"111001111",
  46274=>"111111011",
  46275=>"001001111",
  46276=>"111110000",
  46277=>"011000000",
  46278=>"010000011",
  46279=>"010000110",
  46280=>"001000000",
  46281=>"000111111",
  46282=>"010011001",
  46283=>"111001101",
  46284=>"000011000",
  46285=>"111000000",
  46286=>"111111110",
  46287=>"000000000",
  46288=>"100100100",
  46289=>"111010111",
  46290=>"111111111",
  46291=>"111101111",
  46292=>"111000000",
  46293=>"000000000",
  46294=>"000000100",
  46295=>"100110000",
  46296=>"000100111",
  46297=>"000000000",
  46298=>"010111111",
  46299=>"111000100",
  46300=>"000000000",
  46301=>"001101111",
  46302=>"111111111",
  46303=>"010110011",
  46304=>"101100001",
  46305=>"000000111",
  46306=>"111111110",
  46307=>"111111111",
  46308=>"010000000",
  46309=>"001000001",
  46310=>"011010000",
  46311=>"000000111",
  46312=>"000111111",
  46313=>"000000000",
  46314=>"000111111",
  46315=>"110111111",
  46316=>"000000011",
  46317=>"000001111",
  46318=>"111000000",
  46319=>"000110111",
  46320=>"000000000",
  46321=>"110110000",
  46322=>"000001001",
  46323=>"111000000",
  46324=>"000000001",
  46325=>"000100110",
  46326=>"000000000",
  46327=>"001000111",
  46328=>"000000000",
  46329=>"100100111",
  46330=>"000000001",
  46331=>"111111110",
  46332=>"000011000",
  46333=>"100000000",
  46334=>"111111111",
  46335=>"110000111",
  46336=>"000000001",
  46337=>"010010000",
  46338=>"000000000",
  46339=>"111101011",
  46340=>"000000000",
  46341=>"000110011",
  46342=>"111111111",
  46343=>"110100000",
  46344=>"011011111",
  46345=>"001101111",
  46346=>"111101001",
  46347=>"100100010",
  46348=>"000000100",
  46349=>"010000000",
  46350=>"000000101",
  46351=>"111111000",
  46352=>"111110011",
  46353=>"000000001",
  46354=>"000110111",
  46355=>"001000111",
  46356=>"000000111",
  46357=>"000000000",
  46358=>"101101001",
  46359=>"111111111",
  46360=>"111111011",
  46361=>"000111111",
  46362=>"001000000",
  46363=>"000000000",
  46364=>"011011111",
  46365=>"000000001",
  46366=>"111111010",
  46367=>"110110110",
  46368=>"110111011",
  46369=>"111111111",
  46370=>"001011011",
  46371=>"111111001",
  46372=>"000000000",
  46373=>"000000000",
  46374=>"000100110",
  46375=>"000111111",
  46376=>"000000000",
  46377=>"111111111",
  46378=>"111110000",
  46379=>"111111111",
  46380=>"110000000",
  46381=>"000110000",
  46382=>"111010111",
  46383=>"100100000",
  46384=>"000000000",
  46385=>"111111101",
  46386=>"000000011",
  46387=>"001001011",
  46388=>"000000000",
  46389=>"000000110",
  46390=>"100101011",
  46391=>"000000000",
  46392=>"000000000",
  46393=>"000001111",
  46394=>"001000000",
  46395=>"111111010",
  46396=>"111111111",
  46397=>"000000011",
  46398=>"101000000",
  46399=>"111111111",
  46400=>"111111000",
  46401=>"000001001",
  46402=>"111111111",
  46403=>"000000000",
  46404=>"110111111",
  46405=>"000111111",
  46406=>"000111001",
  46407=>"000001000",
  46408=>"000000001",
  46409=>"000111111",
  46410=>"100110110",
  46411=>"000000000",
  46412=>"111010000",
  46413=>"000000110",
  46414=>"000111111",
  46415=>"100111111",
  46416=>"111110111",
  46417=>"000000011",
  46418=>"111111111",
  46419=>"000000000",
  46420=>"010000000",
  46421=>"000101111",
  46422=>"000000001",
  46423=>"000000001",
  46424=>"000101111",
  46425=>"111111111",
  46426=>"000010000",
  46427=>"110100111",
  46428=>"111111111",
  46429=>"000011111",
  46430=>"111111110",
  46431=>"001001011",
  46432=>"100100100",
  46433=>"101101101",
  46434=>"111111100",
  46435=>"000000001",
  46436=>"101001011",
  46437=>"000000000",
  46438=>"111111011",
  46439=>"111011011",
  46440=>"001000001",
  46441=>"111100100",
  46442=>"110110000",
  46443=>"111000000",
  46444=>"101101001",
  46445=>"111011001",
  46446=>"000000000",
  46447=>"111111000",
  46448=>"000000000",
  46449=>"111111111",
  46450=>"111111000",
  46451=>"100100110",
  46452=>"111111111",
  46453=>"110111000",
  46454=>"111100100",
  46455=>"000000001",
  46456=>"100000000",
  46457=>"111101000",
  46458=>"111111000",
  46459=>"111110111",
  46460=>"000000000",
  46461=>"010101111",
  46462=>"010010000",
  46463=>"111111111",
  46464=>"000000000",
  46465=>"111111111",
  46466=>"000111011",
  46467=>"111000000",
  46468=>"000000111",
  46469=>"000000011",
  46470=>"110000000",
  46471=>"111111111",
  46472=>"000000000",
  46473=>"100000000",
  46474=>"111111111",
  46475=>"000111111",
  46476=>"111111111",
  46477=>"110110000",
  46478=>"110111111",
  46479=>"000111111",
  46480=>"001000000",
  46481=>"000000001",
  46482=>"010110010",
  46483=>"111100100",
  46484=>"001001111",
  46485=>"001001000",
  46486=>"001001000",
  46487=>"000011011",
  46488=>"110011011",
  46489=>"111010000",
  46490=>"000000001",
  46491=>"000101111",
  46492=>"111110110",
  46493=>"111000110",
  46494=>"111101000",
  46495=>"111111111",
  46496=>"111111111",
  46497=>"010010000",
  46498=>"111001001",
  46499=>"111111111",
  46500=>"000011101",
  46501=>"111001000",
  46502=>"101000001",
  46503=>"111111000",
  46504=>"000000000",
  46505=>"000000001",
  46506=>"111111111",
  46507=>"011111111",
  46508=>"010000001",
  46509=>"000000000",
  46510=>"111001111",
  46511=>"111111111",
  46512=>"000000100",
  46513=>"000100111",
  46514=>"110111111",
  46515=>"001000000",
  46516=>"000000100",
  46517=>"000011111",
  46518=>"000000000",
  46519=>"100000111",
  46520=>"101011111",
  46521=>"111000000",
  46522=>"010010110",
  46523=>"001100111",
  46524=>"100011111",
  46525=>"111111101",
  46526=>"000000111",
  46527=>"110111011",
  46528=>"001111111",
  46529=>"000000010",
  46530=>"000000000",
  46531=>"111111110",
  46532=>"000001111",
  46533=>"001000111",
  46534=>"110001001",
  46535=>"111000111",
  46536=>"001001000",
  46537=>"000001111",
  46538=>"010111011",
  46539=>"000000000",
  46540=>"000111000",
  46541=>"010000000",
  46542=>"100100110",
  46543=>"001111111",
  46544=>"101110110",
  46545=>"001000000",
  46546=>"001011000",
  46547=>"000000000",
  46548=>"101111111",
  46549=>"111001000",
  46550=>"000000000",
  46551=>"011010000",
  46552=>"000001111",
  46553=>"111110000",
  46554=>"110111111",
  46555=>"000000111",
  46556=>"111111111",
  46557=>"111101101",
  46558=>"001111111",
  46559=>"000000000",
  46560=>"000000000",
  46561=>"000000000",
  46562=>"000111100",
  46563=>"000000011",
  46564=>"000000111",
  46565=>"110001000",
  46566=>"000011111",
  46567=>"111111100",
  46568=>"100111111",
  46569=>"001000111",
  46570=>"000000111",
  46571=>"000110111",
  46572=>"011011000",
  46573=>"000000000",
  46574=>"101001001",
  46575=>"000010001",
  46576=>"000000000",
  46577=>"000000000",
  46578=>"000100100",
  46579=>"001111111",
  46580=>"000000001",
  46581=>"000000000",
  46582=>"001111001",
  46583=>"111011111",
  46584=>"111110110",
  46585=>"001000010",
  46586=>"000000101",
  46587=>"000010000",
  46588=>"111000010",
  46589=>"000000000",
  46590=>"111110000",
  46591=>"000000000",
  46592=>"111000000",
  46593=>"000000000",
  46594=>"111111111",
  46595=>"111111101",
  46596=>"000000110",
  46597=>"111111100",
  46598=>"111000111",
  46599=>"000000000",
  46600=>"000100110",
  46601=>"110000000",
  46602=>"111111111",
  46603=>"011111110",
  46604=>"000100000",
  46605=>"111100111",
  46606=>"000001000",
  46607=>"001111110",
  46608=>"000000011",
  46609=>"111000000",
  46610=>"000000000",
  46611=>"001111111",
  46612=>"100101111",
  46613=>"001001000",
  46614=>"100101111",
  46615=>"100100000",
  46616=>"011101100",
  46617=>"111100000",
  46618=>"011001111",
  46619=>"000111111",
  46620=>"111111011",
  46621=>"111000000",
  46622=>"011101001",
  46623=>"000100111",
  46624=>"000000000",
  46625=>"111101100",
  46626=>"111101001",
  46627=>"000000000",
  46628=>"011111111",
  46629=>"000000001",
  46630=>"100000000",
  46631=>"110110100",
  46632=>"101111111",
  46633=>"000000000",
  46634=>"111111111",
  46635=>"000100100",
  46636=>"100110000",
  46637=>"111011010",
  46638=>"011011000",
  46639=>"111000000",
  46640=>"000000001",
  46641=>"111111011",
  46642=>"000000000",
  46643=>"011011001",
  46644=>"111111000",
  46645=>"000000110",
  46646=>"000011000",
  46647=>"001111111",
  46648=>"011000101",
  46649=>"011000000",
  46650=>"000000111",
  46651=>"000000000",
  46652=>"111111000",
  46653=>"001111001",
  46654=>"001001000",
  46655=>"111111111",
  46656=>"100000001",
  46657=>"000000000",
  46658=>"010111111",
  46659=>"000100000",
  46660=>"000000000",
  46661=>"111111110",
  46662=>"000000000",
  46663=>"000000000",
  46664=>"011001011",
  46665=>"000000000",
  46666=>"000000110",
  46667=>"000111111",
  46668=>"000000011",
  46669=>"111001000",
  46670=>"111000011",
  46671=>"100111111",
  46672=>"001111111",
  46673=>"100000000",
  46674=>"001000000",
  46675=>"110110111",
  46676=>"000000000",
  46677=>"011000111",
  46678=>"000000000",
  46679=>"111111000",
  46680=>"000011011",
  46681=>"111111111",
  46682=>"111111111",
  46683=>"100000000",
  46684=>"010011011",
  46685=>"100000000",
  46686=>"000000001",
  46687=>"101000000",
  46688=>"101001111",
  46689=>"111111111",
  46690=>"000000000",
  46691=>"111001001",
  46692=>"110000000",
  46693=>"111010000",
  46694=>"111111111",
  46695=>"111111111",
  46696=>"010010000",
  46697=>"010011000",
  46698=>"000111111",
  46699=>"000000000",
  46700=>"000001000",
  46701=>"000100110",
  46702=>"000001000",
  46703=>"000000111",
  46704=>"111110111",
  46705=>"000000000",
  46706=>"111001000",
  46707=>"011001000",
  46708=>"001000111",
  46709=>"110110111",
  46710=>"111111111",
  46711=>"011111111",
  46712=>"010111010",
  46713=>"000000111",
  46714=>"000000110",
  46715=>"000000001",
  46716=>"000001011",
  46717=>"111111111",
  46718=>"000000010",
  46719=>"111111111",
  46720=>"000011111",
  46721=>"001111111",
  46722=>"111001000",
  46723=>"000000111",
  46724=>"000000001",
  46725=>"000000000",
  46726=>"110110000",
  46727=>"000000100",
  46728=>"100111111",
  46729=>"101000000",
  46730=>"000000000",
  46731=>"000100111",
  46732=>"010100000",
  46733=>"000010000",
  46734=>"001111111",
  46735=>"111111111",
  46736=>"001111111",
  46737=>"000010000",
  46738=>"100110001",
  46739=>"011000100",
  46740=>"000001000",
  46741=>"000000000",
  46742=>"000000000",
  46743=>"111100000",
  46744=>"010000000",
  46745=>"000000111",
  46746=>"100111110",
  46747=>"111001000",
  46748=>"000000111",
  46749=>"111011011",
  46750=>"001111111",
  46751=>"000011111",
  46752=>"111111111",
  46753=>"100111000",
  46754=>"111101111",
  46755=>"000000111",
  46756=>"100100110",
  46757=>"101111111",
  46758=>"000000000",
  46759=>"000000011",
  46760=>"000011011",
  46761=>"011111111",
  46762=>"111011000",
  46763=>"111110111",
  46764=>"111111111",
  46765=>"001001001",
  46766=>"000111111",
  46767=>"000001000",
  46768=>"000000000",
  46769=>"001001001",
  46770=>"111110111",
  46771=>"111111111",
  46772=>"000001001",
  46773=>"111111111",
  46774=>"011011001",
  46775=>"111111101",
  46776=>"111101111",
  46777=>"000110100",
  46778=>"000000000",
  46779=>"001000100",
  46780=>"111111111",
  46781=>"100101111",
  46782=>"111111110",
  46783=>"000001110",
  46784=>"111111111",
  46785=>"000000010",
  46786=>"000000000",
  46787=>"111111010",
  46788=>"100101111",
  46789=>"111000000",
  46790=>"000000111",
  46791=>"000000000",
  46792=>"111111111",
  46793=>"110111000",
  46794=>"011000000",
  46795=>"100101111",
  46796=>"000100000",
  46797=>"000100100",
  46798=>"011111111",
  46799=>"011000000",
  46800=>"110100111",
  46801=>"100000000",
  46802=>"000110111",
  46803=>"101101011",
  46804=>"001001001",
  46805=>"111111111",
  46806=>"100101000",
  46807=>"000000100",
  46808=>"111101000",
  46809=>"000111000",
  46810=>"111000100",
  46811=>"011111111",
  46812=>"001011111",
  46813=>"001111111",
  46814=>"110111111",
  46815=>"000000000",
  46816=>"000000000",
  46817=>"000100000",
  46818=>"111100100",
  46819=>"000111101",
  46820=>"001000100",
  46821=>"000000001",
  46822=>"000001001",
  46823=>"000100111",
  46824=>"110110111",
  46825=>"011011011",
  46826=>"000011011",
  46827=>"000000000",
  46828=>"000000000",
  46829=>"111000000",
  46830=>"111001011",
  46831=>"110000000",
  46832=>"001111111",
  46833=>"000000001",
  46834=>"000100000",
  46835=>"000000000",
  46836=>"000000000",
  46837=>"100000000",
  46838=>"000000000",
  46839=>"000000000",
  46840=>"001011000",
  46841=>"000000011",
  46842=>"000111110",
  46843=>"000000000",
  46844=>"000000000",
  46845=>"000001111",
  46846=>"000000000",
  46847=>"010000000",
  46848=>"000011111",
  46849=>"001001100",
  46850=>"111000000",
  46851=>"000000100",
  46852=>"001111000",
  46853=>"000001111",
  46854=>"000000011",
  46855=>"000111100",
  46856=>"010000000",
  46857=>"000000000",
  46858=>"001001000",
  46859=>"000000001",
  46860=>"111001001",
  46861=>"111111111",
  46862=>"111111011",
  46863=>"010010000",
  46864=>"000100000",
  46865=>"110000000",
  46866=>"111001111",
  46867=>"100110111",
  46868=>"111111111",
  46869=>"001000000",
  46870=>"111111100",
  46871=>"111111111",
  46872=>"010111111",
  46873=>"111110010",
  46874=>"111111110",
  46875=>"100000111",
  46876=>"001001000",
  46877=>"000000111",
  46878=>"111111111",
  46879=>"100000000",
  46880=>"111000000",
  46881=>"111011011",
  46882=>"000000000",
  46883=>"000001011",
  46884=>"111111111",
  46885=>"111111011",
  46886=>"111111011",
  46887=>"011011000",
  46888=>"111101101",
  46889=>"000000000",
  46890=>"111111000",
  46891=>"000111111",
  46892=>"110110000",
  46893=>"001001000",
  46894=>"000000111",
  46895=>"000000000",
  46896=>"110000000",
  46897=>"000000111",
  46898=>"110110111",
  46899=>"111110110",
  46900=>"000000000",
  46901=>"110100110",
  46902=>"111111000",
  46903=>"111111110",
  46904=>"100000000",
  46905=>"001000101",
  46906=>"111001000",
  46907=>"000110100",
  46908=>"111111111",
  46909=>"111001000",
  46910=>"000000101",
  46911=>"000010010",
  46912=>"000000001",
  46913=>"000100100",
  46914=>"111111011",
  46915=>"111111000",
  46916=>"111111111",
  46917=>"000111111",
  46918=>"111111001",
  46919=>"000000111",
  46920=>"000000000",
  46921=>"000000000",
  46922=>"100000000",
  46923=>"000000000",
  46924=>"111001111",
  46925=>"000000101",
  46926=>"000011010",
  46927=>"000000100",
  46928=>"001011011",
  46929=>"000101000",
  46930=>"000111111",
  46931=>"111100000",
  46932=>"000000000",
  46933=>"000000000",
  46934=>"100000100",
  46935=>"000000000",
  46936=>"010000011",
  46937=>"000000000",
  46938=>"011111111",
  46939=>"000000000",
  46940=>"111011011",
  46941=>"111011111",
  46942=>"011111111",
  46943=>"100001000",
  46944=>"111101100",
  46945=>"111111000",
  46946=>"000000101",
  46947=>"111111000",
  46948=>"010010110",
  46949=>"100000001",
  46950=>"111111111",
  46951=>"000000000",
  46952=>"101001000",
  46953=>"100000000",
  46954=>"111000000",
  46955=>"111111000",
  46956=>"110110000",
  46957=>"000110110",
  46958=>"111111100",
  46959=>"111001000",
  46960=>"011011111",
  46961=>"111110111",
  46962=>"100000010",
  46963=>"001000100",
  46964=>"000000000",
  46965=>"000000000",
  46966=>"001111000",
  46967=>"001000000",
  46968=>"111111010",
  46969=>"000110111",
  46970=>"000000011",
  46971=>"100000001",
  46972=>"000100100",
  46973=>"100100000",
  46974=>"111111000",
  46975=>"111111000",
  46976=>"111111111",
  46977=>"000000000",
  46978=>"011111111",
  46979=>"001001011",
  46980=>"011011000",
  46981=>"000001000",
  46982=>"011010111",
  46983=>"100111110",
  46984=>"000001011",
  46985=>"100000000",
  46986=>"111111001",
  46987=>"111110000",
  46988=>"000111000",
  46989=>"101101111",
  46990=>"111111111",
  46991=>"000000000",
  46992=>"011111111",
  46993=>"100100101",
  46994=>"000000000",
  46995=>"111111111",
  46996=>"011011110",
  46997=>"000000000",
  46998=>"000111111",
  46999=>"100100100",
  47000=>"011111111",
  47001=>"011000000",
  47002=>"000111000",
  47003=>"111011000",
  47004=>"001011111",
  47005=>"100100110",
  47006=>"000010111",
  47007=>"000111111",
  47008=>"000100111",
  47009=>"110110111",
  47010=>"000111111",
  47011=>"011111111",
  47012=>"000000000",
  47013=>"000111111",
  47014=>"000000111",
  47015=>"000000010",
  47016=>"000000000",
  47017=>"010111111",
  47018=>"111100000",
  47019=>"000000111",
  47020=>"000000000",
  47021=>"000000001",
  47022=>"011000000",
  47023=>"000111111",
  47024=>"000000000",
  47025=>"100110000",
  47026=>"000000011",
  47027=>"000111001",
  47028=>"000001000",
  47029=>"100000000",
  47030=>"100111000",
  47031=>"111111011",
  47032=>"000000000",
  47033=>"000000000",
  47034=>"000000000",
  47035=>"101101000",
  47036=>"101101000",
  47037=>"001101101",
  47038=>"111111000",
  47039=>"111111110",
  47040=>"000000110",
  47041=>"000000000",
  47042=>"111111111",
  47043=>"111111100",
  47044=>"110111111",
  47045=>"011111111",
  47046=>"011011000",
  47047=>"111111000",
  47048=>"000001000",
  47049=>"000000011",
  47050=>"011111000",
  47051=>"000000000",
  47052=>"111011000",
  47053=>"010110100",
  47054=>"111001000",
  47055=>"100101101",
  47056=>"100000000",
  47057=>"001000111",
  47058=>"111111111",
  47059=>"111111111",
  47060=>"000011111",
  47061=>"111111111",
  47062=>"011111000",
  47063=>"000000100",
  47064=>"111111111",
  47065=>"111011000",
  47066=>"110111111",
  47067=>"000000001",
  47068=>"011011101",
  47069=>"101000000",
  47070=>"000000000",
  47071=>"100100000",
  47072=>"111111111",
  47073=>"001000001",
  47074=>"111111111",
  47075=>"111111111",
  47076=>"010011011",
  47077=>"111100000",
  47078=>"001000010",
  47079=>"111111111",
  47080=>"110111001",
  47081=>"111111111",
  47082=>"111000111",
  47083=>"000000000",
  47084=>"110111111",
  47085=>"001001011",
  47086=>"000000011",
  47087=>"100000000",
  47088=>"000010001",
  47089=>"011011111",
  47090=>"111111101",
  47091=>"000110101",
  47092=>"011111001",
  47093=>"011001111",
  47094=>"000111001",
  47095=>"111111111",
  47096=>"000111111",
  47097=>"011111001",
  47098=>"110110110",
  47099=>"111011011",
  47100=>"000000111",
  47101=>"101110110",
  47102=>"001000000",
  47103=>"000000100",
  47104=>"110011011",
  47105=>"000001001",
  47106=>"001001001",
  47107=>"111111111",
  47108=>"000010111",
  47109=>"111110110",
  47110=>"000001101",
  47111=>"000001101",
  47112=>"111101101",
  47113=>"000000000",
  47114=>"000101101",
  47115=>"011111111",
  47116=>"100101000",
  47117=>"010000110",
  47118=>"011001101",
  47119=>"011101101",
  47120=>"101001000",
  47121=>"011011101",
  47122=>"000100001",
  47123=>"001001000",
  47124=>"001001101",
  47125=>"101101111",
  47126=>"100110111",
  47127=>"100001001",
  47128=>"111111111",
  47129=>"010010000",
  47130=>"001101101",
  47131=>"000001001",
  47132=>"000000010",
  47133=>"111011011",
  47134=>"011010001",
  47135=>"000000000",
  47136=>"110110110",
  47137=>"110010000",
  47138=>"110110010",
  47139=>"111101101",
  47140=>"000001000",
  47141=>"110110110",
  47142=>"110101101",
  47143=>"011000001",
  47144=>"000001110",
  47145=>"100101101",
  47146=>"001011011",
  47147=>"101100100",
  47148=>"001001001",
  47149=>"010110111",
  47150=>"010000000",
  47151=>"110110110",
  47152=>"001001000",
  47153=>"001001001",
  47154=>"000100100",
  47155=>"000000010",
  47156=>"110110110",
  47157=>"110110110",
  47158=>"001001111",
  47159=>"001111101",
  47160=>"110000001",
  47161=>"000001111",
  47162=>"001001001",
  47163=>"010000111",
  47164=>"101101100",
  47165=>"010000001",
  47166=>"011000000",
  47167=>"111101001",
  47168=>"001000000",
  47169=>"100000110",
  47170=>"001000000",
  47171=>"101001001",
  47172=>"001001001",
  47173=>"000000100",
  47174=>"101101101",
  47175=>"111111111",
  47176=>"001101001",
  47177=>"000000000",
  47178=>"100100000",
  47179=>"110010010",
  47180=>"010000001",
  47181=>"011000011",
  47182=>"111110010",
  47183=>"011000000",
  47184=>"000101001",
  47185=>"101111111",
  47186=>"001100110",
  47187=>"010010000",
  47188=>"000000000",
  47189=>"111111010",
  47190=>"000000000",
  47191=>"010010000",
  47192=>"000000000",
  47193=>"101001000",
  47194=>"101101111",
  47195=>"000000000",
  47196=>"000000101",
  47197=>"101000000",
  47198=>"011011001",
  47199=>"001001011",
  47200=>"010010010",
  47201=>"111101101",
  47202=>"001001000",
  47203=>"111111111",
  47204=>"000111100",
  47205=>"110100000",
  47206=>"000010000",
  47207=>"001111011",
  47208=>"011001011",
  47209=>"001101111",
  47210=>"101101101",
  47211=>"001000100",
  47212=>"011011010",
  47213=>"111111101",
  47214=>"110010010",
  47215=>"101111111",
  47216=>"110110010",
  47217=>"110010001",
  47218=>"110110010",
  47219=>"001000100",
  47220=>"001001001",
  47221=>"000000000",
  47222=>"100000100",
  47223=>"100000111",
  47224=>"111000010",
  47225=>"110110110",
  47226=>"000101000",
  47227=>"001001001",
  47228=>"110110110",
  47229=>"011111001",
  47230=>"000001000",
  47231=>"110001001",
  47232=>"101101101",
  47233=>"110010111",
  47234=>"100010000",
  47235=>"010010000",
  47236=>"111101000",
  47237=>"000001000",
  47238=>"101000110",
  47239=>"110011111",
  47240=>"001000100",
  47241=>"000000101",
  47242=>"011011000",
  47243=>"011000000",
  47244=>"001001001",
  47245=>"011111111",
  47246=>"110100100",
  47247=>"010010010",
  47248=>"100000000",
  47249=>"010110110",
  47250=>"001001111",
  47251=>"011000010",
  47252=>"010010011",
  47253=>"000000000",
  47254=>"101001001",
  47255=>"101101101",
  47256=>"001001101",
  47257=>"111011011",
  47258=>"010010001",
  47259=>"001001000",
  47260=>"001001001",
  47261=>"111110110",
  47262=>"111011111",
  47263=>"010010111",
  47264=>"111001101",
  47265=>"010110110",
  47266=>"010010000",
  47267=>"101111111",
  47268=>"110010001",
  47269=>"000000000",
  47270=>"001001001",
  47271=>"011011011",
  47272=>"101101101",
  47273=>"011001000",
  47274=>"001001000",
  47275=>"100110010",
  47276=>"001111111",
  47277=>"000000000",
  47278=>"110110010",
  47279=>"110110110",
  47280=>"000000010",
  47281=>"010010110",
  47282=>"111111110",
  47283=>"000000010",
  47284=>"110010000",
  47285=>"010000011",
  47286=>"010001101",
  47287=>"000001111",
  47288=>"000000010",
  47289=>"001000010",
  47290=>"010010000",
  47291=>"110010011",
  47292=>"101000100",
  47293=>"110110000",
  47294=>"110110000",
  47295=>"110110110",
  47296=>"111111001",
  47297=>"000000001",
  47298=>"111110111",
  47299=>"001000000",
  47300=>"111011011",
  47301=>"100100101",
  47302=>"110111011",
  47303=>"110110110",
  47304=>"001000000",
  47305=>"111110110",
  47306=>"001011001",
  47307=>"111111010",
  47308=>"010110110",
  47309=>"110100100",
  47310=>"000100110",
  47311=>"010010000",
  47312=>"001001001",
  47313=>"111111111",
  47314=>"000000000",
  47315=>"101001000",
  47316=>"110110111",
  47317=>"010010010",
  47318=>"101101101",
  47319=>"001001001",
  47320=>"110010011",
  47321=>"000001001",
  47322=>"101101101",
  47323=>"111011010",
  47324=>"110110110",
  47325=>"001101001",
  47326=>"110000111",
  47327=>"001001001",
  47328=>"101001100",
  47329=>"111100100",
  47330=>"111101101",
  47331=>"000000001",
  47332=>"000000000",
  47333=>"000101111",
  47334=>"011011000",
  47335=>"111111001",
  47336=>"101001000",
  47337=>"110000001",
  47338=>"111111111",
  47339=>"101101101",
  47340=>"010110110",
  47341=>"111111111",
  47342=>"010010100",
  47343=>"001001001",
  47344=>"110111110",
  47345=>"001011001",
  47346=>"101100110",
  47347=>"110110001",
  47348=>"001000101",
  47349=>"100100100",
  47350=>"000000000",
  47351=>"000000111",
  47352=>"000000111",
  47353=>"000111111",
  47354=>"111111111",
  47355=>"110110000",
  47356=>"011011011",
  47357=>"001001001",
  47358=>"011101101",
  47359=>"001111101",
  47360=>"001001001",
  47361=>"000000001",
  47362=>"010000100",
  47363=>"110000010",
  47364=>"000000000",
  47365=>"101101110",
  47366=>"001010000",
  47367=>"110110001",
  47368=>"010110010",
  47369=>"100100100",
  47370=>"000101111",
  47371=>"010011001",
  47372=>"100100100",
  47373=>"110110100",
  47374=>"010011000",
  47375=>"000111111",
  47376=>"001001001",
  47377=>"010110111",
  47378=>"001101101",
  47379=>"001001011",
  47380=>"001101111",
  47381=>"001001001",
  47382=>"001000000",
  47383=>"010010010",
  47384=>"010010010",
  47385=>"000000111",
  47386=>"100001011",
  47387=>"000101001",
  47388=>"110001001",
  47389=>"000000110",
  47390=>"000001001",
  47391=>"010010110",
  47392=>"011101001",
  47393=>"000111110",
  47394=>"100000111",
  47395=>"000001000",
  47396=>"101101001",
  47397=>"001101011",
  47398=>"010111111",
  47399=>"110110101",
  47400=>"101111111",
  47401=>"010010000",
  47402=>"110110110",
  47403=>"001001101",
  47404=>"000110110",
  47405=>"000000011",
  47406=>"001001011",
  47407=>"111101000",
  47408=>"111111111",
  47409=>"000111101",
  47410=>"111110111",
  47411=>"101101001",
  47412=>"000001110",
  47413=>"111110110",
  47414=>"101101101",
  47415=>"101001001",
  47416=>"011010110",
  47417=>"101101101",
  47418=>"011000000",
  47419=>"111101111",
  47420=>"000000000",
  47421=>"110100000",
  47422=>"000001000",
  47423=>"000000101",
  47424=>"101100101",
  47425=>"000000110",
  47426=>"110110001",
  47427=>"000010000",
  47428=>"101001110",
  47429=>"001100000",
  47430=>"001001000",
  47431=>"110110010",
  47432=>"100000100",
  47433=>"001001001",
  47434=>"001011110",
  47435=>"101001001",
  47436=>"001001001",
  47437=>"101001110",
  47438=>"001000000",
  47439=>"110110100",
  47440=>"001000000",
  47441=>"000000101",
  47442=>"110110110",
  47443=>"100110010",
  47444=>"111111101",
  47445=>"011011001",
  47446=>"011010010",
  47447=>"111010000",
  47448=>"000011011",
  47449=>"000001001",
  47450=>"000110110",
  47451=>"110111010",
  47452=>"001001100",
  47453=>"111111111",
  47454=>"101110110",
  47455=>"001011011",
  47456=>"100001001",
  47457=>"100000000",
  47458=>"100100000",
  47459=>"000000000",
  47460=>"110111111",
  47461=>"000000000",
  47462=>"001101111",
  47463=>"111011001",
  47464=>"110000000",
  47465=>"111111001",
  47466=>"000110010",
  47467=>"001010110",
  47468=>"001001001",
  47469=>"110110110",
  47470=>"101101000",
  47471=>"000000000",
  47472=>"000000001",
  47473=>"001001010",
  47474=>"111111111",
  47475=>"011010010",
  47476=>"001001001",
  47477=>"000100100",
  47478=>"011001000",
  47479=>"011011011",
  47480=>"000000000",
  47481=>"001111111",
  47482=>"111011000",
  47483=>"001000000",
  47484=>"101111000",
  47485=>"000010010",
  47486=>"001001011",
  47487=>"000000000",
  47488=>"000011000",
  47489=>"011111111",
  47490=>"001001001",
  47491=>"001001001",
  47492=>"011111100",
  47493=>"010010110",
  47494=>"001101010",
  47495=>"000011111",
  47496=>"000000000",
  47497=>"000111101",
  47498=>"000000000",
  47499=>"011001101",
  47500=>"001001001",
  47501=>"011011011",
  47502=>"010101111",
  47503=>"001100001",
  47504=>"100100100",
  47505=>"000000111",
  47506=>"111011110",
  47507=>"000001001",
  47508=>"000000001",
  47509=>"000000001",
  47510=>"000000100",
  47511=>"111111111",
  47512=>"111111101",
  47513=>"001000010",
  47514=>"111101001",
  47515=>"011001011",
  47516=>"000100000",
  47517=>"010111001",
  47518=>"110110110",
  47519=>"111011000",
  47520=>"000100000",
  47521=>"011011010",
  47522=>"110010001",
  47523=>"101101100",
  47524=>"110111111",
  47525=>"110111111",
  47526=>"001101111",
  47527=>"100111010",
  47528=>"000000101",
  47529=>"101101001",
  47530=>"000000000",
  47531=>"010010010",
  47532=>"000000000",
  47533=>"001001111",
  47534=>"001011111",
  47535=>"010010111",
  47536=>"101101111",
  47537=>"001000000",
  47538=>"000001111",
  47539=>"001001101",
  47540=>"111110110",
  47541=>"110010000",
  47542=>"000000000",
  47543=>"000111111",
  47544=>"111001001",
  47545=>"011000011",
  47546=>"001000000",
  47547=>"000100100",
  47548=>"111000000",
  47549=>"011110001",
  47550=>"111111111",
  47551=>"010010000",
  47552=>"110110000",
  47553=>"000110111",
  47554=>"111111111",
  47555=>"001000000",
  47556=>"001101001",
  47557=>"001001101",
  47558=>"010000000",
  47559=>"011011010",
  47560=>"000000001",
  47561=>"001000001",
  47562=>"101001001",
  47563=>"000001111",
  47564=>"000000110",
  47565=>"110110111",
  47566=>"000010110",
  47567=>"101111000",
  47568=>"000000010",
  47569=>"010011011",
  47570=>"000010010",
  47571=>"111111111",
  47572=>"000100100",
  47573=>"000010110",
  47574=>"101001101",
  47575=>"011011010",
  47576=>"110010000",
  47577=>"001000000",
  47578=>"101011000",
  47579=>"100100000",
  47580=>"001111111",
  47581=>"110010000",
  47582=>"111110100",
  47583=>"010000001",
  47584=>"101011011",
  47585=>"001000001",
  47586=>"000100111",
  47587=>"000001100",
  47588=>"010010110",
  47589=>"001101101",
  47590=>"100100110",
  47591=>"101101101",
  47592=>"010010010",
  47593=>"000100111",
  47594=>"001001001",
  47595=>"100110000",
  47596=>"111001101",
  47597=>"010010011",
  47598=>"111111111",
  47599=>"011001001",
  47600=>"010011000",
  47601=>"110010011",
  47602=>"101111100",
  47603=>"111100100",
  47604=>"110110010",
  47605=>"001101001",
  47606=>"000000010",
  47607=>"100000000",
  47608=>"010000100",
  47609=>"101000001",
  47610=>"001001001",
  47611=>"001001001",
  47612=>"000101111",
  47613=>"111011001",
  47614=>"111110000",
  47615=>"101000000",
  47616=>"011001000",
  47617=>"110110111",
  47618=>"000000111",
  47619=>"101000000",
  47620=>"111010000",
  47621=>"000000100",
  47622=>"111111111",
  47623=>"000000111",
  47624=>"111111111",
  47625=>"101001101",
  47626=>"111000001",
  47627=>"111001011",
  47628=>"110110110",
  47629=>"010010000",
  47630=>"000000110",
  47631=>"001101000",
  47632=>"000000000",
  47633=>"011111111",
  47634=>"011001101",
  47635=>"010110010",
  47636=>"111111111",
  47637=>"110101001",
  47638=>"000000000",
  47639=>"111111001",
  47640=>"100000000",
  47641=>"100110111",
  47642=>"111111111",
  47643=>"111110111",
  47644=>"111111111",
  47645=>"011111111",
  47646=>"000000000",
  47647=>"000111010",
  47648=>"000010111",
  47649=>"000000011",
  47650=>"011111010",
  47651=>"111111111",
  47652=>"000000000",
  47653=>"000001111",
  47654=>"111111001",
  47655=>"111011111",
  47656=>"001001111",
  47657=>"101100100",
  47658=>"001001111",
  47659=>"110111110",
  47660=>"000111010",
  47661=>"010111010",
  47662=>"100100100",
  47663=>"000100000",
  47664=>"111111111",
  47665=>"011111011",
  47666=>"101111011",
  47667=>"000000000",
  47668=>"001001001",
  47669=>"111010010",
  47670=>"000100111",
  47671=>"100000000",
  47672=>"000100010",
  47673=>"000001111",
  47674=>"111111011",
  47675=>"000000111",
  47676=>"000000000",
  47677=>"001000000",
  47678=>"000000110",
  47679=>"000000001",
  47680=>"010110110",
  47681=>"101101111",
  47682=>"111111111",
  47683=>"010010000",
  47684=>"001001000",
  47685=>"111110110",
  47686=>"000000111",
  47687=>"100100101",
  47688=>"011111001",
  47689=>"000000001",
  47690=>"110110000",
  47691=>"110110110",
  47692=>"000001111",
  47693=>"110101000",
  47694=>"100000000",
  47695=>"000001011",
  47696=>"111100000",
  47697=>"000000111",
  47698=>"000000011",
  47699=>"111111010",
  47700=>"000000000",
  47701=>"000000110",
  47702=>"111111110",
  47703=>"011011000",
  47704=>"001001111",
  47705=>"100000101",
  47706=>"000000111",
  47707=>"000011011",
  47708=>"111111111",
  47709=>"000000101",
  47710=>"100000110",
  47711=>"110000110",
  47712=>"001111111",
  47713=>"000000000",
  47714=>"110110111",
  47715=>"001001001",
  47716=>"110110000",
  47717=>"000000000",
  47718=>"000000111",
  47719=>"110100000",
  47720=>"111111111",
  47721=>"100000000",
  47722=>"110110111",
  47723=>"111111100",
  47724=>"110111111",
  47725=>"000000000",
  47726=>"000000000",
  47727=>"010010000",
  47728=>"001001111",
  47729=>"001001100",
  47730=>"100110011",
  47731=>"111111111",
  47732=>"110010000",
  47733=>"111111000",
  47734=>"000000001",
  47735=>"011111111",
  47736=>"001001000",
  47737=>"010110010",
  47738=>"111100000",
  47739=>"000000001",
  47740=>"001001110",
  47741=>"101000000",
  47742=>"100100110",
  47743=>"110111100",
  47744=>"111100100",
  47745=>"010010010",
  47746=>"110110110",
  47747=>"011011011",
  47748=>"000111100",
  47749=>"100000101",
  47750=>"000010000",
  47751=>"011111000",
  47752=>"111111111",
  47753=>"111100100",
  47754=>"111111111",
  47755=>"110111000",
  47756=>"001001001",
  47757=>"000000000",
  47758=>"010000000",
  47759=>"111111111",
  47760=>"000000101",
  47761=>"001000000",
  47762=>"010110100",
  47763=>"111111111",
  47764=>"110000000",
  47765=>"011010010",
  47766=>"110100100",
  47767=>"000000111",
  47768=>"000000000",
  47769=>"000000100",
  47770=>"010111111",
  47771=>"101111111",
  47772=>"111110010",
  47773=>"100000000",
  47774=>"011000000",
  47775=>"111000000",
  47776=>"010000000",
  47777=>"000000111",
  47778=>"111111101",
  47779=>"010111111",
  47780=>"111111111",
  47781=>"000000000",
  47782=>"001101001",
  47783=>"000000000",
  47784=>"111111111",
  47785=>"000000000",
  47786=>"100000000",
  47787=>"100100101",
  47788=>"111011010",
  47789=>"110110001",
  47790=>"000101110",
  47791=>"000000000",
  47792=>"010111111",
  47793=>"111111000",
  47794=>"011111111",
  47795=>"101101101",
  47796=>"110110000",
  47797=>"000000000",
  47798=>"111111111",
  47799=>"111110010",
  47800=>"000000111",
  47801=>"111111111",
  47802=>"111001000",
  47803=>"110111011",
  47804=>"000000000",
  47805=>"110111010",
  47806=>"111101100",
  47807=>"110000000",
  47808=>"111111111",
  47809=>"011111100",
  47810=>"010000000",
  47811=>"000001011",
  47812=>"101111111",
  47813=>"000000000",
  47814=>"111000000",
  47815=>"000010010",
  47816=>"110110000",
  47817=>"111111111",
  47818=>"111001000",
  47819=>"111111111",
  47820=>"000010000",
  47821=>"101001000",
  47822=>"000111111",
  47823=>"000010010",
  47824=>"000000000",
  47825=>"100000101",
  47826=>"001001001",
  47827=>"100100000",
  47828=>"011011000",
  47829=>"111110110",
  47830=>"101100100",
  47831=>"001000000",
  47832=>"110110110",
  47833=>"000111111",
  47834=>"111111111",
  47835=>"000010011",
  47836=>"100000000",
  47837=>"001101000",
  47838=>"111111000",
  47839=>"110000000",
  47840=>"111101101",
  47841=>"000000000",
  47842=>"111111111",
  47843=>"111110000",
  47844=>"010000000",
  47845=>"000000000",
  47846=>"110110010",
  47847=>"010000110",
  47848=>"111111010",
  47849=>"010110000",
  47850=>"000011000",
  47851=>"110111010",
  47852=>"001101101",
  47853=>"000111111",
  47854=>"111100100",
  47855=>"111101111",
  47856=>"110100110",
  47857=>"111111011",
  47858=>"000000000",
  47859=>"001011000",
  47860=>"111111111",
  47861=>"011010000",
  47862=>"001100010",
  47863=>"011011011",
  47864=>"111111111",
  47865=>"101111001",
  47866=>"000000001",
  47867=>"101000000",
  47868=>"111111001",
  47869=>"000000100",
  47870=>"110000000",
  47871=>"111111110",
  47872=>"000000000",
  47873=>"000000000",
  47874=>"000000011",
  47875=>"000000111",
  47876=>"000010110",
  47877=>"111111111",
  47878=>"001000111",
  47879=>"000111111",
  47880=>"000000000",
  47881=>"111101001",
  47882=>"111100111",
  47883=>"110111110",
  47884=>"001001111",
  47885=>"100000000",
  47886=>"000010111",
  47887=>"000000000",
  47888=>"000000000",
  47889=>"111111010",
  47890=>"000000001",
  47891=>"011000000",
  47892=>"000100110",
  47893=>"001111111",
  47894=>"111111101",
  47895=>"000000000",
  47896=>"001101101",
  47897=>"010111100",
  47898=>"000000010",
  47899=>"010111000",
  47900=>"000001111",
  47901=>"111111111",
  47902=>"000000000",
  47903=>"011100111",
  47904=>"111110000",
  47905=>"000100100",
  47906=>"111110000",
  47907=>"111111111",
  47908=>"111111111",
  47909=>"010000000",
  47910=>"011111011",
  47911=>"111111111",
  47912=>"000000000",
  47913=>"000000000",
  47914=>"111011000",
  47915=>"000000000",
  47916=>"000000001",
  47917=>"000111001",
  47918=>"111111111",
  47919=>"000000011",
  47920=>"011111000",
  47921=>"010010000",
  47922=>"101001101",
  47923=>"000000011",
  47924=>"000000000",
  47925=>"101001001",
  47926=>"100110100",
  47927=>"011001111",
  47928=>"110100000",
  47929=>"000000101",
  47930=>"111001001",
  47931=>"111011000",
  47932=>"000000000",
  47933=>"000000000",
  47934=>"111011000",
  47935=>"011010011",
  47936=>"011100000",
  47937=>"000000000",
  47938=>"111111111",
  47939=>"111111000",
  47940=>"000000000",
  47941=>"000000000",
  47942=>"111111110",
  47943=>"000001000",
  47944=>"001001001",
  47945=>"010100111",
  47946=>"110111110",
  47947=>"101000000",
  47948=>"011000000",
  47949=>"111110000",
  47950=>"001001111",
  47951=>"001001111",
  47952=>"111001111",
  47953=>"111111110",
  47954=>"111111000",
  47955=>"111111111",
  47956=>"011011011",
  47957=>"011011001",
  47958=>"000001111",
  47959=>"000000001",
  47960=>"010011011",
  47961=>"001001111",
  47962=>"000001011",
  47963=>"110100110",
  47964=>"110100100",
  47965=>"001111100",
  47966=>"111111111",
  47967=>"111111111",
  47968=>"100100000",
  47969=>"000000000",
  47970=>"100100000",
  47971=>"101001001",
  47972=>"111001000",
  47973=>"000000000",
  47974=>"001111111",
  47975=>"000001101",
  47976=>"001000000",
  47977=>"010111111",
  47978=>"011011000",
  47979=>"001001001",
  47980=>"110110100",
  47981=>"001000111",
  47982=>"111111000",
  47983=>"001001001",
  47984=>"000000000",
  47985=>"111111110",
  47986=>"001001000",
  47987=>"000001001",
  47988=>"000000000",
  47989=>"011111000",
  47990=>"100000000",
  47991=>"110111000",
  47992=>"101001000",
  47993=>"000000001",
  47994=>"111001000",
  47995=>"001000000",
  47996=>"111000000",
  47997=>"111111111",
  47998=>"000000000",
  47999=>"101000101",
  48000=>"011011001",
  48001=>"111110110",
  48002=>"111111111",
  48003=>"000000000",
  48004=>"000010111",
  48005=>"101111111",
  48006=>"110110110",
  48007=>"111111111",
  48008=>"111111111",
  48009=>"000000000",
  48010=>"000000000",
  48011=>"100101111",
  48012=>"000000101",
  48013=>"111111101",
  48014=>"111100100",
  48015=>"100100100",
  48016=>"000111111",
  48017=>"000000010",
  48018=>"111101101",
  48019=>"111110000",
  48020=>"111001111",
  48021=>"010010000",
  48022=>"001001001",
  48023=>"010000000",
  48024=>"111111111",
  48025=>"111111110",
  48026=>"000101000",
  48027=>"111000100",
  48028=>"111111110",
  48029=>"011011111",
  48030=>"001011001",
  48031=>"111111111",
  48032=>"111110110",
  48033=>"011000000",
  48034=>"001000000",
  48035=>"100100000",
  48036=>"001001000",
  48037=>"101000000",
  48038=>"001001111",
  48039=>"011000000",
  48040=>"111111001",
  48041=>"000000000",
  48042=>"010111111",
  48043=>"000000100",
  48044=>"111111111",
  48045=>"011010000",
  48046=>"111111111",
  48047=>"010000111",
  48048=>"000100111",
  48049=>"111111110",
  48050=>"000000000",
  48051=>"011000000",
  48052=>"001101111",
  48053=>"000001101",
  48054=>"000000000",
  48055=>"110110000",
  48056=>"000100100",
  48057=>"111111011",
  48058=>"000000000",
  48059=>"000000001",
  48060=>"000000001",
  48061=>"111111000",
  48062=>"111100000",
  48063=>"000000000",
  48064=>"011111000",
  48065=>"001001011",
  48066=>"000000001",
  48067=>"000000111",
  48068=>"001000100",
  48069=>"001011111",
  48070=>"000000100",
  48071=>"000000000",
  48072=>"001000000",
  48073=>"111000000",
  48074=>"100100100",
  48075=>"001001111",
  48076=>"111000000",
  48077=>"000000010",
  48078=>"000000000",
  48079=>"011011011",
  48080=>"101101000",
  48081=>"001011011",
  48082=>"000110000",
  48083=>"000000010",
  48084=>"000000000",
  48085=>"111101110",
  48086=>"000000000",
  48087=>"011111011",
  48088=>"001101110",
  48089=>"001000111",
  48090=>"111011011",
  48091=>"010000000",
  48092=>"111101111",
  48093=>"000001001",
  48094=>"001001111",
  48095=>"110110111",
  48096=>"000001001",
  48097=>"000000000",
  48098=>"011000011",
  48099=>"000000000",
  48100=>"001000110",
  48101=>"111111111",
  48102=>"100100111",
  48103=>"100000000",
  48104=>"001101001",
  48105=>"110111111",
  48106=>"100111111",
  48107=>"000000101",
  48108=>"000000111",
  48109=>"000000000",
  48110=>"001001001",
  48111=>"000101111",
  48112=>"001001011",
  48113=>"100000000",
  48114=>"111111111",
  48115=>"000000000",
  48116=>"111111111",
  48117=>"001000101",
  48118=>"110111110",
  48119=>"010010010",
  48120=>"011000000",
  48121=>"000000001",
  48122=>"000110110",
  48123=>"000001001",
  48124=>"000000000",
  48125=>"110111110",
  48126=>"000010000",
  48127=>"100111111",
  48128=>"111000000",
  48129=>"111000000",
  48130=>"101101100",
  48131=>"111111000",
  48132=>"111111111",
  48133=>"001111001",
  48134=>"111001111",
  48135=>"111000000",
  48136=>"001111100",
  48137=>"000000111",
  48138=>"000000000",
  48139=>"011010000",
  48140=>"110000000",
  48141=>"111111000",
  48142=>"111111001",
  48143=>"000000001",
  48144=>"000001111",
  48145=>"111111011",
  48146=>"000111111",
  48147=>"111111111",
  48148=>"101101000",
  48149=>"000000111",
  48150=>"111111111",
  48151=>"111100000",
  48152=>"111011000",
  48153=>"001011111",
  48154=>"111000011",
  48155=>"011001100",
  48156=>"000000110",
  48157=>"000101111",
  48158=>"111101000",
  48159=>"111111000",
  48160=>"100111011",
  48161=>"100100000",
  48162=>"001111000",
  48163=>"100100111",
  48164=>"111110110",
  48165=>"111111111",
  48166=>"110110110",
  48167=>"111111000",
  48168=>"000011111",
  48169=>"000000111",
  48170=>"011001101",
  48171=>"111111111",
  48172=>"000000111",
  48173=>"010000000",
  48174=>"000000111",
  48175=>"111111111",
  48176=>"100001001",
  48177=>"000111111",
  48178=>"000000000",
  48179=>"111111000",
  48180=>"000111110",
  48181=>"000000000",
  48182=>"111111111",
  48183=>"110110000",
  48184=>"111111001",
  48185=>"001001000",
  48186=>"000000000",
  48187=>"000000000",
  48188=>"111000111",
  48189=>"110000111",
  48190=>"110100000",
  48191=>"111111101",
  48192=>"111111111",
  48193=>"000111110",
  48194=>"001000011",
  48195=>"111111100",
  48196=>"000000000",
  48197=>"000000111",
  48198=>"100000000",
  48199=>"111111111",
  48200=>"000001000",
  48201=>"111000000",
  48202=>"111001111",
  48203=>"111111011",
  48204=>"111001111",
  48205=>"111000000",
  48206=>"111111000",
  48207=>"111011000",
  48208=>"100000000",
  48209=>"000011111",
  48210=>"011000000",
  48211=>"011011001",
  48212=>"111111111",
  48213=>"000000000",
  48214=>"111000000",
  48215=>"110111111",
  48216=>"000000110",
  48217=>"111101000",
  48218=>"111000000",
  48219=>"110101000",
  48220=>"000000000",
  48221=>"000011001",
  48222=>"001111111",
  48223=>"000000000",
  48224=>"111111000",
  48225=>"000111111",
  48226=>"000000100",
  48227=>"100110100",
  48228=>"011000000",
  48229=>"101111101",
  48230=>"100001111",
  48231=>"111111111",
  48232=>"000000111",
  48233=>"111111111",
  48234=>"111000000",
  48235=>"000001101",
  48236=>"001000110",
  48237=>"000000001",
  48238=>"110111111",
  48239=>"111000000",
  48240=>"100000110",
  48241=>"000000000",
  48242=>"011110111",
  48243=>"000000111",
  48244=>"001001111",
  48245=>"001111111",
  48246=>"010000000",
  48247=>"000001111",
  48248=>"000111111",
  48249=>"000111111",
  48250=>"000000011",
  48251=>"000101111",
  48252=>"010111011",
  48253=>"111111111",
  48254=>"111111101",
  48255=>"000000011",
  48256=>"000000000",
  48257=>"111101000",
  48258=>"100000000",
  48259=>"000100000",
  48260=>"111111100",
  48261=>"111001111",
  48262=>"000000000",
  48263=>"000000000",
  48264=>"001000000",
  48265=>"000000001",
  48266=>"110100100",
  48267=>"101000111",
  48268=>"000000000",
  48269=>"111100000",
  48270=>"000111111",
  48271=>"101111100",
  48272=>"000100111",
  48273=>"000010111",
  48274=>"000000001",
  48275=>"010000000",
  48276=>"111111000",
  48277=>"000100111",
  48278=>"111111000",
  48279=>"111100000",
  48280=>"111111001",
  48281=>"000000001",
  48282=>"000101001",
  48283=>"100111000",
  48284=>"001011001",
  48285=>"000000111",
  48286=>"111111111",
  48287=>"001000111",
  48288=>"111001000",
  48289=>"100000000",
  48290=>"000000000",
  48291=>"111010000",
  48292=>"100000000",
  48293=>"111111111",
  48294=>"110000000",
  48295=>"000111111",
  48296=>"100100101",
  48297=>"000000000",
  48298=>"111001000",
  48299=>"000000000",
  48300=>"001011111",
  48301=>"111111000",
  48302=>"100111111",
  48303=>"110110010",
  48304=>"111110100",
  48305=>"110000001",
  48306=>"110111110",
  48307=>"111111000",
  48308=>"111111011",
  48309=>"111000000",
  48310=>"000000000",
  48311=>"010010000",
  48312=>"000000101",
  48313=>"011011000",
  48314=>"100000010",
  48315=>"111000000",
  48316=>"000000000",
  48317=>"100000110",
  48318=>"110111111",
  48319=>"000001111",
  48320=>"111111000",
  48321=>"111111000",
  48322=>"111111111",
  48323=>"000111000",
  48324=>"000111111",
  48325=>"000111111",
  48326=>"110111011",
  48327=>"111111011",
  48328=>"000000000",
  48329=>"111100000",
  48330=>"000000110",
  48331=>"000000111",
  48332=>"000000101",
  48333=>"000010000",
  48334=>"111101101",
  48335=>"111111101",
  48336=>"000000000",
  48337=>"101000111",
  48338=>"000000000",
  48339=>"001111001",
  48340=>"111100111",
  48341=>"101001101",
  48342=>"011001001",
  48343=>"000001001",
  48344=>"111111000",
  48345=>"001000101",
  48346=>"111111111",
  48347=>"001000000",
  48348=>"111001001",
  48349=>"110000111",
  48350=>"000000000",
  48351=>"000100110",
  48352=>"000000000",
  48353=>"111011010",
  48354=>"111111111",
  48355=>"000000000",
  48356=>"000000000",
  48357=>"001000000",
  48358=>"111111100",
  48359=>"000100100",
  48360=>"011001000",
  48361=>"111111111",
  48362=>"001111111",
  48363=>"001001000",
  48364=>"011111111",
  48365=>"111111101",
  48366=>"000000111",
  48367=>"111111000",
  48368=>"000111101",
  48369=>"110100000",
  48370=>"111001111",
  48371=>"110000000",
  48372=>"001001100",
  48373=>"000000000",
  48374=>"000100110",
  48375=>"111111100",
  48376=>"111001001",
  48377=>"000011001",
  48378=>"111100100",
  48379=>"000000000",
  48380=>"000100111",
  48381=>"110011010",
  48382=>"011000000",
  48383=>"011111101",
  48384=>"001001111",
  48385=>"011000000",
  48386=>"000001000",
  48387=>"000000000",
  48388=>"000100100",
  48389=>"100100110",
  48390=>"111000000",
  48391=>"001000000",
  48392=>"001001111",
  48393=>"000000000",
  48394=>"111111000",
  48395=>"001000000",
  48396=>"100000110",
  48397=>"111110001",
  48398=>"111111000",
  48399=>"000100100",
  48400=>"000100000",
  48401=>"111111000",
  48402=>"011001011",
  48403=>"111010000",
  48404=>"011011000",
  48405=>"111100000",
  48406=>"100100101",
  48407=>"001011001",
  48408=>"111111000",
  48409=>"000000000",
  48410=>"000111000",
  48411=>"100100000",
  48412=>"000000000",
  48413=>"100111111",
  48414=>"000000000",
  48415=>"110000111",
  48416=>"111100001",
  48417=>"110000111",
  48418=>"111111111",
  48419=>"000001101",
  48420=>"110110000",
  48421=>"111001000",
  48422=>"111100000",
  48423=>"000000111",
  48424=>"110010001",
  48425=>"000000000",
  48426=>"110111011",
  48427=>"111111000",
  48428=>"111111001",
  48429=>"000011111",
  48430=>"100000000",
  48431=>"111111000",
  48432=>"000011011",
  48433=>"110111111",
  48434=>"111111111",
  48435=>"000000000",
  48436=>"111111000",
  48437=>"111011000",
  48438=>"000000000",
  48439=>"000000010",
  48440=>"011111111",
  48441=>"111000000",
  48442=>"111000000",
  48443=>"111110111",
  48444=>"111111001",
  48445=>"011011111",
  48446=>"111111001",
  48447=>"000111111",
  48448=>"000000000",
  48449=>"111000000",
  48450=>"001111100",
  48451=>"010111111",
  48452=>"111111000",
  48453=>"111111111",
  48454=>"001000000",
  48455=>"111001111",
  48456=>"000011111",
  48457=>"111000000",
  48458=>"011001000",
  48459=>"000000110",
  48460=>"000000011",
  48461=>"000001100",
  48462=>"111100000",
  48463=>"000000111",
  48464=>"001001000",
  48465=>"111001001",
  48466=>"001000000",
  48467=>"111111111",
  48468=>"000000000",
  48469=>"001001001",
  48470=>"000010111",
  48471=>"100100110",
  48472=>"011000000",
  48473=>"100000000",
  48474=>"110100000",
  48475=>"101000000",
  48476=>"000010111",
  48477=>"000000010",
  48478=>"000000111",
  48479=>"110111110",
  48480=>"111111000",
  48481=>"000010111",
  48482=>"111100000",
  48483=>"101000000",
  48484=>"000111111",
  48485=>"000000111",
  48486=>"000000000",
  48487=>"000111111",
  48488=>"000000000",
  48489=>"111001001",
  48490=>"010000000",
  48491=>"110110000",
  48492=>"111011111",
  48493=>"111100111",
  48494=>"001000000",
  48495=>"000000000",
  48496=>"001100000",
  48497=>"000000001",
  48498=>"111111111",
  48499=>"000001011",
  48500=>"111000000",
  48501=>"000000111",
  48502=>"000000000",
  48503=>"000000001",
  48504=>"111001001",
  48505=>"010110110",
  48506=>"110000000",
  48507=>"000011111",
  48508=>"111111000",
  48509=>"111000000",
  48510=>"000111000",
  48511=>"000000100",
  48512=>"000110000",
  48513=>"000011000",
  48514=>"100100110",
  48515=>"100100100",
  48516=>"111100000",
  48517=>"110110000",
  48518=>"100100000",
  48519=>"110000000",
  48520=>"111111111",
  48521=>"111111000",
  48522=>"010001001",
  48523=>"111111111",
  48524=>"001000000",
  48525=>"000110011",
  48526=>"011111111",
  48527=>"001011000",
  48528=>"000000010",
  48529=>"111111100",
  48530=>"010111111",
  48531=>"110100100",
  48532=>"110100000",
  48533=>"000111000",
  48534=>"110000000",
  48535=>"110111000",
  48536=>"000000000",
  48537=>"000000011",
  48538=>"111111111",
  48539=>"111111111",
  48540=>"001000000",
  48541=>"000000000",
  48542=>"000111111",
  48543=>"111111000",
  48544=>"001111111",
  48545=>"000111111",
  48546=>"111101101",
  48547=>"101001111",
  48548=>"001000100",
  48549=>"000000000",
  48550=>"000100000",
  48551=>"011111011",
  48552=>"001001011",
  48553=>"000010111",
  48554=>"111111100",
  48555=>"111111111",
  48556=>"000000000",
  48557=>"000101101",
  48558=>"000000111",
  48559=>"000000001",
  48560=>"000111110",
  48561=>"000000000",
  48562=>"100100100",
  48563=>"000100111",
  48564=>"000000011",
  48565=>"101000000",
  48566=>"001001100",
  48567=>"111000000",
  48568=>"111111000",
  48569=>"011111000",
  48570=>"000000100",
  48571=>"001001111",
  48572=>"000001101",
  48573=>"001000100",
  48574=>"000000000",
  48575=>"110110000",
  48576=>"111000000",
  48577=>"000000000",
  48578=>"000111000",
  48579=>"000000111",
  48580=>"000000100",
  48581=>"000000101",
  48582=>"111111000",
  48583=>"011111111",
  48584=>"011000001",
  48585=>"101000000",
  48586=>"111101111",
  48587=>"000110011",
  48588=>"111010000",
  48589=>"111100000",
  48590=>"011000000",
  48591=>"111000001",
  48592=>"111111101",
  48593=>"110011111",
  48594=>"111111000",
  48595=>"101111111",
  48596=>"000000001",
  48597=>"110111111",
  48598=>"000000111",
  48599=>"000000000",
  48600=>"100111111",
  48601=>"111111001",
  48602=>"000000000",
  48603=>"100000100",
  48604=>"111111011",
  48605=>"111000000",
  48606=>"111111000",
  48607=>"111111111",
  48608=>"000000001",
  48609=>"111011000",
  48610=>"100110111",
  48611=>"000000001",
  48612=>"111111110",
  48613=>"000000111",
  48614=>"000000110",
  48615=>"101101000",
  48616=>"111000000",
  48617=>"000011111",
  48618=>"111110001",
  48619=>"111111011",
  48620=>"100000000",
  48621=>"111111001",
  48622=>"000010000",
  48623=>"111111110",
  48624=>"111000110",
  48625=>"011111101",
  48626=>"111111101",
  48627=>"110010010",
  48628=>"111111111",
  48629=>"110111111",
  48630=>"001111111",
  48631=>"000111010",
  48632=>"111100000",
  48633=>"011001101",
  48634=>"110001001",
  48635=>"000000000",
  48636=>"000000111",
  48637=>"111111011",
  48638=>"111111111",
  48639=>"001000000",
  48640=>"111110011",
  48641=>"011000000",
  48642=>"111100100",
  48643=>"000110110",
  48644=>"110100000",
  48645=>"000111010",
  48646=>"000000000",
  48647=>"111001001",
  48648=>"111111000",
  48649=>"000000000",
  48650=>"000000000",
  48651=>"010110111",
  48652=>"000110110",
  48653=>"011011000",
  48654=>"001000000",
  48655=>"000000000",
  48656=>"111111111",
  48657=>"000000000",
  48658=>"000001101",
  48659=>"100100000",
  48660=>"111111010",
  48661=>"000000000",
  48662=>"000000000",
  48663=>"111111111",
  48664=>"110110100",
  48665=>"001001000",
  48666=>"111111101",
  48667=>"011001001",
  48668=>"110111110",
  48669=>"000100000",
  48670=>"111111111",
  48671=>"111111011",
  48672=>"110110000",
  48673=>"011001111",
  48674=>"000000000",
  48675=>"000100000",
  48676=>"000010000",
  48677=>"111111111",
  48678=>"000000111",
  48679=>"100000000",
  48680=>"000000000",
  48681=>"000000000",
  48682=>"111111011",
  48683=>"111111111",
  48684=>"111111111",
  48685=>"101111001",
  48686=>"001001001",
  48687=>"111000111",
  48688=>"111111111",
  48689=>"000111000",
  48690=>"000010110",
  48691=>"011111011",
  48692=>"001001101",
  48693=>"000000000",
  48694=>"000000100",
  48695=>"000001111",
  48696=>"111111111",
  48697=>"000000000",
  48698=>"000000000",
  48699=>"000000000",
  48700=>"111111111",
  48701=>"001001001",
  48702=>"000000000",
  48703=>"001001111",
  48704=>"111111101",
  48705=>"000001111",
  48706=>"100001100",
  48707=>"111100111",
  48708=>"000000000",
  48709=>"111111111",
  48710=>"111111111",
  48711=>"110000000",
  48712=>"111110110",
  48713=>"111111111",
  48714=>"111111111",
  48715=>"110011111",
  48716=>"111111110",
  48717=>"111111111",
  48718=>"000000000",
  48719=>"111111111",
  48720=>"000110111",
  48721=>"000000000",
  48722=>"111111111",
  48723=>"000000000",
  48724=>"110111111",
  48725=>"100000000",
  48726=>"111100111",
  48727=>"010110111",
  48728=>"111111101",
  48729=>"101101101",
  48730=>"111000000",
  48731=>"010110110",
  48732=>"000000011",
  48733=>"111111111",
  48734=>"110110100",
  48735=>"111111111",
  48736=>"000000111",
  48737=>"101001000",
  48738=>"111111110",
  48739=>"000000001",
  48740=>"000000000",
  48741=>"111111111",
  48742=>"001110100",
  48743=>"000000000",
  48744=>"111111000",
  48745=>"111111000",
  48746=>"100100101",
  48747=>"010000000",
  48748=>"110000000",
  48749=>"111111111",
  48750=>"110111111",
  48751=>"000000100",
  48752=>"001001111",
  48753=>"000001011",
  48754=>"111110100",
  48755=>"100100000",
  48756=>"000000000",
  48757=>"111110011",
  48758=>"000100111",
  48759=>"000000000",
  48760=>"000000000",
  48761=>"111101000",
  48762=>"011000000",
  48763=>"100000111",
  48764=>"110110110",
  48765=>"000000001",
  48766=>"001000000",
  48767=>"000000000",
  48768=>"111111000",
  48769=>"111101000",
  48770=>"111110111",
  48771=>"000000000",
  48772=>"111111101",
  48773=>"111111111",
  48774=>"000000000",
  48775=>"111111111",
  48776=>"001000000",
  48777=>"101101111",
  48778=>"000000000",
  48779=>"111111111",
  48780=>"001000000",
  48781=>"100110110",
  48782=>"000000111",
  48783=>"010000100",
  48784=>"111111111",
  48785=>"100000000",
  48786=>"111111111",
  48787=>"000011111",
  48788=>"111000111",
  48789=>"111110110",
  48790=>"111111111",
  48791=>"111111111",
  48792=>"000000000",
  48793=>"111111110",
  48794=>"000000000",
  48795=>"010111111",
  48796=>"111111001",
  48797=>"000000000",
  48798=>"000100100",
  48799=>"101001000",
  48800=>"000000100",
  48801=>"011001001",
  48802=>"011111111",
  48803=>"000010000",
  48804=>"000000000",
  48805=>"000000000",
  48806=>"011011001",
  48807=>"011011011",
  48808=>"111000000",
  48809=>"001001001",
  48810=>"000000111",
  48811=>"111111111",
  48812=>"111111111",
  48813=>"101100001",
  48814=>"001100110",
  48815=>"100000111",
  48816=>"000111111",
  48817=>"000000000",
  48818=>"010111010",
  48819=>"000000000",
  48820=>"011001101",
  48821=>"000000000",
  48822=>"000001001",
  48823=>"001101111",
  48824=>"111100000",
  48825=>"000111000",
  48826=>"000110100",
  48827=>"100100100",
  48828=>"111111111",
  48829=>"100100000",
  48830=>"010000000",
  48831=>"000000000",
  48832=>"001111011",
  48833=>"000000101",
  48834=>"000111010",
  48835=>"111111111",
  48836=>"000000111",
  48837=>"101000000",
  48838=>"011010111",
  48839=>"111111111",
  48840=>"000000000",
  48841=>"111101000",
  48842=>"111111001",
  48843=>"110000000",
  48844=>"111101001",
  48845=>"000100110",
  48846=>"111100111",
  48847=>"111110010",
  48848=>"000000000",
  48849=>"111111111",
  48850=>"000000000",
  48851=>"111111111",
  48852=>"000000000",
  48853=>"111111111",
  48854=>"111111111",
  48855=>"111000111",
  48856=>"000000101",
  48857=>"110111110",
  48858=>"000001000",
  48859=>"000000000",
  48860=>"111101111",
  48861=>"110110111",
  48862=>"000000000",
  48863=>"111000111",
  48864=>"111111111",
  48865=>"000011000",
  48866=>"111100111",
  48867=>"111000000",
  48868=>"001100100",
  48869=>"000000000",
  48870=>"000000000",
  48871=>"111000000",
  48872=>"111011011",
  48873=>"110110111",
  48874=>"000000100",
  48875=>"011001111",
  48876=>"000000011",
  48877=>"111111111",
  48878=>"111111111",
  48879=>"111111111",
  48880=>"000000000",
  48881=>"101001000",
  48882=>"111111100",
  48883=>"000000000",
  48884=>"011000111",
  48885=>"111111111",
  48886=>"100100100",
  48887=>"111011001",
  48888=>"111111111",
  48889=>"000110000",
  48890=>"000110000",
  48891=>"111111111",
  48892=>"111011001",
  48893=>"111110110",
  48894=>"000000101",
  48895=>"110111111",
  48896=>"000011111",
  48897=>"111111011",
  48898=>"000000001",
  48899=>"011001000",
  48900=>"111100100",
  48901=>"000000000",
  48902=>"111111111",
  48903=>"111000111",
  48904=>"001001100",
  48905=>"000000111",
  48906=>"000000000",
  48907=>"000000000",
  48908=>"111111111",
  48909=>"100000010",
  48910=>"101111111",
  48911=>"111111000",
  48912=>"000111111",
  48913=>"001011111",
  48914=>"111111010",
  48915=>"000000001",
  48916=>"000100100",
  48917=>"000000001",
  48918=>"111110100",
  48919=>"000000000",
  48920=>"000000000",
  48921=>"011000000",
  48922=>"111111001",
  48923=>"111110000",
  48924=>"011011001",
  48925=>"111111111",
  48926=>"000111111",
  48927=>"000000111",
  48928=>"000000000",
  48929=>"001001000",
  48930=>"001011000",
  48931=>"000000000",
  48932=>"111000000",
  48933=>"011000110",
  48934=>"000000001",
  48935=>"000000000",
  48936=>"000110000",
  48937=>"000000000",
  48938=>"000000000",
  48939=>"000000000",
  48940=>"110010000",
  48941=>"011111111",
  48942=>"000000000",
  48943=>"000000011",
  48944=>"000010110",
  48945=>"000000000",
  48946=>"111111111",
  48947=>"100000000",
  48948=>"000000000",
  48949=>"111001010",
  48950=>"000000000",
  48951=>"001000000",
  48952=>"111111111",
  48953=>"111111111",
  48954=>"010010111",
  48955=>"111111100",
  48956=>"100111111",
  48957=>"000000111",
  48958=>"010011000",
  48959=>"000000110",
  48960=>"111111111",
  48961=>"111001001",
  48962=>"000010000",
  48963=>"000000000",
  48964=>"111111000",
  48965=>"111011111",
  48966=>"011111111",
  48967=>"001101000",
  48968=>"000000000",
  48969=>"110000000",
  48970=>"000000000",
  48971=>"111111111",
  48972=>"001000111",
  48973=>"111000001",
  48974=>"111111111",
  48975=>"111011011",
  48976=>"111111111",
  48977=>"111111111",
  48978=>"000000111",
  48979=>"010000000",
  48980=>"000100000",
  48981=>"011011011",
  48982=>"000000000",
  48983=>"000000000",
  48984=>"000000000",
  48985=>"000000000",
  48986=>"100000000",
  48987=>"001101101",
  48988=>"111011001",
  48989=>"001000000",
  48990=>"000000000",
  48991=>"000111111",
  48992=>"000000011",
  48993=>"111011111",
  48994=>"111111110",
  48995=>"100001011",
  48996=>"100101100",
  48997=>"000000001",
  48998=>"000001001",
  48999=>"100100100",
  49000=>"111111111",
  49001=>"000001001",
  49002=>"000010000",
  49003=>"111001000",
  49004=>"110010110",
  49005=>"000010111",
  49006=>"000000000",
  49007=>"000000000",
  49008=>"010111111",
  49009=>"000011001",
  49010=>"001000000",
  49011=>"001000000",
  49012=>"111111000",
  49013=>"111111110",
  49014=>"111111111",
  49015=>"111000000",
  49016=>"111111000",
  49017=>"101001000",
  49018=>"000000000",
  49019=>"101111111",
  49020=>"111111010",
  49021=>"111000000",
  49022=>"111111111",
  49023=>"111111111",
  49024=>"000000000",
  49025=>"011001101",
  49026=>"111111111",
  49027=>"000011000",
  49028=>"001101111",
  49029=>"110000000",
  49030=>"011111001",
  49031=>"011000000",
  49032=>"000011111",
  49033=>"111111111",
  49034=>"111111111",
  49035=>"000010000",
  49036=>"111111111",
  49037=>"000000000",
  49038=>"000000010",
  49039=>"000000001",
  49040=>"010000110",
  49041=>"100000100",
  49042=>"111111011",
  49043=>"011111111",
  49044=>"100100111",
  49045=>"000000000",
  49046=>"111111110",
  49047=>"000000000",
  49048=>"001101111",
  49049=>"000000100",
  49050=>"011111101",
  49051=>"011110000",
  49052=>"111110100",
  49053=>"000000000",
  49054=>"000000000",
  49055=>"000000000",
  49056=>"000000000",
  49057=>"111110111",
  49058=>"000100111",
  49059=>"111111111",
  49060=>"100100111",
  49061=>"000000000",
  49062=>"000000010",
  49063=>"111111001",
  49064=>"111000101",
  49065=>"000000000",
  49066=>"100100101",
  49067=>"000100100",
  49068=>"000000000",
  49069=>"111001111",
  49070=>"000000000",
  49071=>"000010000",
  49072=>"100110100",
  49073=>"111111000",
  49074=>"000110000",
  49075=>"111100110",
  49076=>"100111110",
  49077=>"111111111",
  49078=>"111111111",
  49079=>"001011111",
  49080=>"111111011",
  49081=>"011111111",
  49082=>"000000000",
  49083=>"000110000",
  49084=>"111111111",
  49085=>"100100111",
  49086=>"000000000",
  49087=>"101101101",
  49088=>"000000000",
  49089=>"000000000",
  49090=>"011001000",
  49091=>"111111000",
  49092=>"001000100",
  49093=>"111111011",
  49094=>"111000000",
  49095=>"100000111",
  49096=>"001111100",
  49097=>"001000000",
  49098=>"111111111",
  49099=>"111111111",
  49100=>"000011001",
  49101=>"111100101",
  49102=>"001000101",
  49103=>"000000000",
  49104=>"111101111",
  49105=>"000111111",
  49106=>"000100001",
  49107=>"000011000",
  49108=>"000000110",
  49109=>"000000000",
  49110=>"000000110",
  49111=>"000001011",
  49112=>"111111111",
  49113=>"000000100",
  49114=>"000110111",
  49115=>"111111111",
  49116=>"001000000",
  49117=>"000000000",
  49118=>"111111111",
  49119=>"000110111",
  49120=>"011011011",
  49121=>"000001001",
  49122=>"000110110",
  49123=>"111101111",
  49124=>"111101111",
  49125=>"000000111",
  49126=>"100000000",
  49127=>"111111111",
  49128=>"000001000",
  49129=>"000011010",
  49130=>"001001011",
  49131=>"001001111",
  49132=>"111011011",
  49133=>"001001001",
  49134=>"111011000",
  49135=>"000000101",
  49136=>"000000000",
  49137=>"101000000",
  49138=>"000000000",
  49139=>"111001111",
  49140=>"010100000",
  49141=>"000000000",
  49142=>"001011111",
  49143=>"111011111",
  49144=>"000001111",
  49145=>"111110001",
  49146=>"110110110",
  49147=>"111111111",
  49148=>"101000110",
  49149=>"111101111",
  49150=>"111111101",
  49151=>"000110100",
  49152=>"101111111",
  49153=>"111000000",
  49154=>"100111111",
  49155=>"011000000",
  49156=>"000000000",
  49157=>"110111011",
  49158=>"010000000",
  49159=>"111111111",
  49160=>"000000000",
  49161=>"101101111",
  49162=>"000000001",
  49163=>"000000010",
  49164=>"011000000",
  49165=>"111111111",
  49166=>"001011111",
  49167=>"000000000",
  49168=>"000000011",
  49169=>"111011000",
  49170=>"111111111",
  49171=>"111111000",
  49172=>"100000101",
  49173=>"000110110",
  49174=>"000000000",
  49175=>"001011111",
  49176=>"001000000",
  49177=>"111111111",
  49178=>"001000000",
  49179=>"000100100",
  49180=>"100101000",
  49181=>"111100111",
  49182=>"111110000",
  49183=>"000000101",
  49184=>"000111101",
  49185=>"001100000",
  49186=>"011111111",
  49187=>"000000101",
  49188=>"000000000",
  49189=>"111111111",
  49190=>"000000000",
  49191=>"100101111",
  49192=>"111111111",
  49193=>"100111000",
  49194=>"100111111",
  49195=>"000000000",
  49196=>"000001111",
  49197=>"111111011",
  49198=>"000000000",
  49199=>"000010111",
  49200=>"000010011",
  49201=>"000000000",
  49202=>"100100100",
  49203=>"111000000",
  49204=>"101111010",
  49205=>"111010000",
  49206=>"001100101",
  49207=>"111111110",
  49208=>"000111111",
  49209=>"001000100",
  49210=>"000000000",
  49211=>"110000000",
  49212=>"111000000",
  49213=>"011011000",
  49214=>"010010010",
  49215=>"111111111",
  49216=>"000101111",
  49217=>"001001111",
  49218=>"000111111",
  49219=>"111101111",
  49220=>"001011111",
  49221=>"000000000",
  49222=>"000000111",
  49223=>"111111111",
  49224=>"111000000",
  49225=>"000000111",
  49226=>"000000000",
  49227=>"011011000",
  49228=>"000000000",
  49229=>"000100000",
  49230=>"100111111",
  49231=>"101111111",
  49232=>"000000111",
  49233=>"111111111",
  49234=>"000111111",
  49235=>"000001001",
  49236=>"111111001",
  49237=>"000000111",
  49238=>"010000101",
  49239=>"000000000",
  49240=>"101001101",
  49241=>"111100101",
  49242=>"000000000",
  49243=>"000000001",
  49244=>"000000101",
  49245=>"111000000",
  49246=>"111110000",
  49247=>"110000000",
  49248=>"000000111",
  49249=>"010111111",
  49250=>"100000000",
  49251=>"001000110",
  49252=>"111010000",
  49253=>"000001000",
  49254=>"111111111",
  49255=>"001000000",
  49256=>"001111111",
  49257=>"111000000",
  49258=>"111101000",
  49259=>"000000000",
  49260=>"111011010",
  49261=>"000000111",
  49262=>"100100111",
  49263=>"000000111",
  49264=>"011010111",
  49265=>"001001101",
  49266=>"000010010",
  49267=>"000000000",
  49268=>"111110000",
  49269=>"100000000",
  49270=>"000100000",
  49271=>"000111111",
  49272=>"111000000",
  49273=>"000000000",
  49274=>"110000000",
  49275=>"000100111",
  49276=>"111111110",
  49277=>"000111111",
  49278=>"000101101",
  49279=>"010010000",
  49280=>"001000000",
  49281=>"000000001",
  49282=>"111111111",
  49283=>"001111011",
  49284=>"000111111",
  49285=>"111111111",
  49286=>"000001001",
  49287=>"000000111",
  49288=>"111110110",
  49289=>"100111110",
  49290=>"000000000",
  49291=>"000000000",
  49292=>"001111111",
  49293=>"010111111",
  49294=>"111111111",
  49295=>"111111111",
  49296=>"111111111",
  49297=>"010000000",
  49298=>"000000000",
  49299=>"111011000",
  49300=>"111100000",
  49301=>"000000000",
  49302=>"111000000",
  49303=>"100110000",
  49304=>"001001001",
  49305=>"101000100",
  49306=>"101000000",
  49307=>"010000000",
  49308=>"110110101",
  49309=>"111001001",
  49310=>"100100111",
  49311=>"000000101",
  49312=>"000000100",
  49313=>"001000000",
  49314=>"011000100",
  49315=>"111111111",
  49316=>"101001001",
  49317=>"111111110",
  49318=>"011000000",
  49319=>"011111111",
  49320=>"001000000",
  49321=>"000000000",
  49322=>"000000000",
  49323=>"110111111",
  49324=>"000111001",
  49325=>"001000100",
  49326=>"100111101",
  49327=>"011111000",
  49328=>"001000000",
  49329=>"111110111",
  49330=>"010010110",
  49331=>"111000000",
  49332=>"111111111",
  49333=>"000000000",
  49334=>"111010000",
  49335=>"000000000",
  49336=>"100110111",
  49337=>"111000000",
  49338=>"111100000",
  49339=>"000000000",
  49340=>"001000000",
  49341=>"000000111",
  49342=>"000101111",
  49343=>"001111000",
  49344=>"110110000",
  49345=>"111000000",
  49346=>"000100110",
  49347=>"000000000",
  49348=>"111111111",
  49349=>"111111111",
  49350=>"111111111",
  49351=>"000000000",
  49352=>"001111111",
  49353=>"001011000",
  49354=>"100001111",
  49355=>"000100000",
  49356=>"111011000",
  49357=>"000000000",
  49358=>"100000000",
  49359=>"101000000",
  49360=>"000000000",
  49361=>"011111111",
  49362=>"111000111",
  49363=>"000000000",
  49364=>"000000111",
  49365=>"111111111",
  49366=>"111001000",
  49367=>"000000000",
  49368=>"111111111",
  49369=>"111111111",
  49370=>"000000000",
  49371=>"000111111",
  49372=>"000100100",
  49373=>"000000000",
  49374=>"000000000",
  49375=>"000001000",
  49376=>"000000100",
  49377=>"111111000",
  49378=>"101000001",
  49379=>"111000101",
  49380=>"111011000",
  49381=>"000000001",
  49382=>"000110111",
  49383=>"000000111",
  49384=>"111111111",
  49385=>"111001000",
  49386=>"000000101",
  49387=>"000001001",
  49388=>"000000000",
  49389=>"000001101",
  49390=>"111101111",
  49391=>"000000000",
  49392=>"110111111",
  49393=>"111001001",
  49394=>"101101011",
  49395=>"001001111",
  49396=>"000000000",
  49397=>"000001011",
  49398=>"111001011",
  49399=>"001001101",
  49400=>"000001001",
  49401=>"111111100",
  49402=>"111000000",
  49403=>"011111111",
  49404=>"000111111",
  49405=>"000010000",
  49406=>"000010110",
  49407=>"000000001",
  49408=>"111111100",
  49409=>"111010000",
  49410=>"111111011",
  49411=>"011111111",
  49412=>"101111111",
  49413=>"000000011",
  49414=>"101100000",
  49415=>"000000000",
  49416=>"000000000",
  49417=>"111111111",
  49418=>"011111111",
  49419=>"101000101",
  49420=>"111101111",
  49421=>"000000000",
  49422=>"110101101",
  49423=>"111010000",
  49424=>"000000000",
  49425=>"000111111",
  49426=>"110000110",
  49427=>"000000111",
  49428=>"111111111",
  49429=>"111000001",
  49430=>"111011000",
  49431=>"000000001",
  49432=>"000010110",
  49433=>"001011111",
  49434=>"000000000",
  49435=>"111111000",
  49436=>"111111001",
  49437=>"111111111",
  49438=>"000000000",
  49439=>"000100100",
  49440=>"001001111",
  49441=>"000000011",
  49442=>"010111111",
  49443=>"000000100",
  49444=>"111100000",
  49445=>"111111111",
  49446=>"111111110",
  49447=>"110000000",
  49448=>"001000110",
  49449=>"000000111",
  49450=>"111111000",
  49451=>"000000110",
  49452=>"100001000",
  49453=>"111111011",
  49454=>"000000000",
  49455=>"011110000",
  49456=>"111111111",
  49457=>"000010000",
  49458=>"110000000",
  49459=>"111000000",
  49460=>"111111100",
  49461=>"111000000",
  49462=>"000000000",
  49463=>"100111101",
  49464=>"111111000",
  49465=>"000000111",
  49466=>"000000100",
  49467=>"111111010",
  49468=>"111110110",
  49469=>"001000100",
  49470=>"000110101",
  49471=>"111111000",
  49472=>"111111100",
  49473=>"000000000",
  49474=>"000000000",
  49475=>"000000000",
  49476=>"111101000",
  49477=>"001001111",
  49478=>"000000000",
  49479=>"000000001",
  49480=>"000010011",
  49481=>"000000100",
  49482=>"001000111",
  49483=>"110100000",
  49484=>"000000000",
  49485=>"000110000",
  49486=>"000000000",
  49487=>"000100100",
  49488=>"110111000",
  49489=>"000000100",
  49490=>"100000000",
  49491=>"000110000",
  49492=>"111111111",
  49493=>"111000000",
  49494=>"111100000",
  49495=>"000000000",
  49496=>"000000000",
  49497=>"000001000",
  49498=>"010111110",
  49499=>"000101111",
  49500=>"000000000",
  49501=>"011011111",
  49502=>"000011111",
  49503=>"000011111",
  49504=>"000111111",
  49505=>"111110000",
  49506=>"111011011",
  49507=>"001000000",
  49508=>"111111111",
  49509=>"110110000",
  49510=>"000000110",
  49511=>"111111110",
  49512=>"011011001",
  49513=>"111000000",
  49514=>"111111001",
  49515=>"000101110",
  49516=>"010000000",
  49517=>"111101001",
  49518=>"000000000",
  49519=>"011011110",
  49520=>"000000000",
  49521=>"111001000",
  49522=>"111011011",
  49523=>"001001110",
  49524=>"101111111",
  49525=>"000000000",
  49526=>"111101101",
  49527=>"011111000",
  49528=>"011111110",
  49529=>"011000000",
  49530=>"000000000",
  49531=>"011111111",
  49532=>"000100111",
  49533=>"010110100",
  49534=>"110111111",
  49535=>"000000000",
  49536=>"110001000",
  49537=>"011111110",
  49538=>"001001000",
  49539=>"000000000",
  49540=>"110000000",
  49541=>"000000000",
  49542=>"000000000",
  49543=>"111100101",
  49544=>"000000111",
  49545=>"000000001",
  49546=>"010111111",
  49547=>"111111000",
  49548=>"111111111",
  49549=>"011011011",
  49550=>"101011111",
  49551=>"011111111",
  49552=>"000011111",
  49553=>"000111111",
  49554=>"111001111",
  49555=>"111001001",
  49556=>"111111111",
  49557=>"111011000",
  49558=>"000000000",
  49559=>"011111110",
  49560=>"000000111",
  49561=>"110100110",
  49562=>"001001111",
  49563=>"001000000",
  49564=>"010111111",
  49565=>"000010011",
  49566=>"111000011",
  49567=>"000000000",
  49568=>"000000000",
  49569=>"010110110",
  49570=>"111111101",
  49571=>"000000000",
  49572=>"001111111",
  49573=>"000000000",
  49574=>"000110111",
  49575=>"000000111",
  49576=>"000000000",
  49577=>"000000000",
  49578=>"001001000",
  49579=>"111111111",
  49580=>"111111000",
  49581=>"000111111",
  49582=>"000001111",
  49583=>"111111111",
  49584=>"100000000",
  49585=>"101000000",
  49586=>"111111100",
  49587=>"111111111",
  49588=>"110100111",
  49589=>"011110111",
  49590=>"101111111",
  49591=>"000000000",
  49592=>"000000010",
  49593=>"001100100",
  49594=>"111000000",
  49595=>"000001000",
  49596=>"000001011",
  49597=>"111111110",
  49598=>"000000000",
  49599=>"011011011",
  49600=>"111000101",
  49601=>"000110110",
  49602=>"111111111",
  49603=>"000111111",
  49604=>"000110001",
  49605=>"001001011",
  49606=>"001111111",
  49607=>"011000101",
  49608=>"001111001",
  49609=>"000111111",
  49610=>"010000000",
  49611=>"111111001",
  49612=>"100100110",
  49613=>"000111111",
  49614=>"000000000",
  49615=>"110110110",
  49616=>"111111111",
  49617=>"111001000",
  49618=>"011000000",
  49619=>"111111110",
  49620=>"111111111",
  49621=>"000101101",
  49622=>"111111111",
  49623=>"100000100",
  49624=>"000010000",
  49625=>"110111111",
  49626=>"011011000",
  49627=>"000111111",
  49628=>"001001011",
  49629=>"000000100",
  49630=>"111000000",
  49631=>"001011001",
  49632=>"111111110",
  49633=>"000001000",
  49634=>"101111111",
  49635=>"000000101",
  49636=>"000000111",
  49637=>"111110110",
  49638=>"100000111",
  49639=>"000000000",
  49640=>"011111111",
  49641=>"000000000",
  49642=>"111000001",
  49643=>"100000000",
  49644=>"100000000",
  49645=>"000000001",
  49646=>"011111111",
  49647=>"111111110",
  49648=>"111111110",
  49649=>"111111111",
  49650=>"111111111",
  49651=>"111101101",
  49652=>"000111111",
  49653=>"000000000",
  49654=>"000111111",
  49655=>"111000000",
  49656=>"111111010",
  49657=>"110100011",
  49658=>"000000011",
  49659=>"000100111",
  49660=>"011011111",
  49661=>"000000100",
  49662=>"111111000",
  49663=>"000000000",
  49664=>"000000000",
  49665=>"000000000",
  49666=>"000000000",
  49667=>"111111100",
  49668=>"100010110",
  49669=>"111111100",
  49670=>"100000000",
  49671=>"111111111",
  49672=>"000111000",
  49673=>"000000000",
  49674=>"111110000",
  49675=>"100100000",
  49676=>"010011011",
  49677=>"000000000",
  49678=>"111100111",
  49679=>"111101111",
  49680=>"111000011",
  49681=>"000001000",
  49682=>"111111101",
  49683=>"111111111",
  49684=>"110111111",
  49685=>"000000000",
  49686=>"111000001",
  49687=>"111111111",
  49688=>"111011101",
  49689=>"111100100",
  49690=>"000000111",
  49691=>"100000000",
  49692=>"111111101",
  49693=>"110100000",
  49694=>"100100110",
  49695=>"111101000",
  49696=>"000000000",
  49697=>"100000000",
  49698=>"111111111",
  49699=>"000010010",
  49700=>"110000000",
  49701=>"111111111",
  49702=>"000000100",
  49703=>"111111111",
  49704=>"000000000",
  49705=>"000011011",
  49706=>"111111111",
  49707=>"001111111",
  49708=>"110111111",
  49709=>"000000000",
  49710=>"111101111",
  49711=>"111111111",
  49712=>"000000000",
  49713=>"111111111",
  49714=>"001110110",
  49715=>"011001001",
  49716=>"000000000",
  49717=>"000000000",
  49718=>"100000000",
  49719=>"000000111",
  49720=>"100100111",
  49721=>"100000110",
  49722=>"000000000",
  49723=>"010110010",
  49724=>"000111111",
  49725=>"000011111",
  49726=>"111111111",
  49727=>"111111111",
  49728=>"111111111",
  49729=>"011111100",
  49730=>"110111111",
  49731=>"000000000",
  49732=>"111111111",
  49733=>"011111111",
  49734=>"001101000",
  49735=>"000000000",
  49736=>"110110110",
  49737=>"111111111",
  49738=>"000000000",
  49739=>"111111011",
  49740=>"000000110",
  49741=>"000000000",
  49742=>"111100100",
  49743=>"111111111",
  49744=>"100111110",
  49745=>"111111010",
  49746=>"000000011",
  49747=>"000000000",
  49748=>"000000110",
  49749=>"001111111",
  49750=>"001000000",
  49751=>"000000000",
  49752=>"110110110",
  49753=>"000000000",
  49754=>"000000000",
  49755=>"110110111",
  49756=>"000010000",
  49757=>"111000000",
  49758=>"111111111",
  49759=>"111110111",
  49760=>"000000000",
  49761=>"110111111",
  49762=>"111001001",
  49763=>"111111111",
  49764=>"000000000",
  49765=>"000000100",
  49766=>"111111100",
  49767=>"111111111",
  49768=>"000001001",
  49769=>"000000000",
  49770=>"000000111",
  49771=>"000011000",
  49772=>"111011111",
  49773=>"111111111",
  49774=>"001001000",
  49775=>"000000000",
  49776=>"001001011",
  49777=>"000000010",
  49778=>"111010000",
  49779=>"100000010",
  49780=>"111111111",
  49781=>"000000000",
  49782=>"110110111",
  49783=>"000100100",
  49784=>"000000000",
  49785=>"111000000",
  49786=>"000000000",
  49787=>"001001111",
  49788=>"011011001",
  49789=>"000000000",
  49790=>"111111111",
  49791=>"111111111",
  49792=>"111111111",
  49793=>"000000000",
  49794=>"111001101",
  49795=>"001010010",
  49796=>"000000011",
  49797=>"000011111",
  49798=>"001000110",
  49799=>"111110111",
  49800=>"000000000",
  49801=>"000000000",
  49802=>"111111000",
  49803=>"000000000",
  49804=>"011011111",
  49805=>"000110111",
  49806=>"111111111",
  49807=>"111111011",
  49808=>"000000001",
  49809=>"011110000",
  49810=>"111111111",
  49811=>"100000000",
  49812=>"100000000",
  49813=>"011001001",
  49814=>"100000000",
  49815=>"000000000",
  49816=>"111111110",
  49817=>"111111111",
  49818=>"111111111",
  49819=>"100000100",
  49820=>"110111111",
  49821=>"000000000",
  49822=>"111111101",
  49823=>"000000000",
  49824=>"111110000",
  49825=>"111111111",
  49826=>"000000010",
  49827=>"111111111",
  49828=>"000000000",
  49829=>"100100001",
  49830=>"110111010",
  49831=>"111111111",
  49832=>"111111111",
  49833=>"000000101",
  49834=>"111111111",
  49835=>"001111000",
  49836=>"111111000",
  49837=>"000100111",
  49838=>"111101111",
  49839=>"000000000",
  49840=>"000000000",
  49841=>"011011000",
  49842=>"010011010",
  49843=>"111111111",
  49844=>"011101111",
  49845=>"101111101",
  49846=>"000000000",
  49847=>"101000111",
  49848=>"101111111",
  49849=>"000000000",
  49850=>"000000111",
  49851=>"001000101",
  49852=>"110111011",
  49853=>"000000110",
  49854=>"111111111",
  49855=>"000000000",
  49856=>"111000000",
  49857=>"111110111",
  49858=>"011000000",
  49859=>"000001001",
  49860=>"111111111",
  49861=>"111111111",
  49862=>"111111111",
  49863=>"000000000",
  49864=>"100111101",
  49865=>"010100000",
  49866=>"111111111",
  49867=>"001000000",
  49868=>"110111101",
  49869=>"100100110",
  49870=>"111111111",
  49871=>"111000000",
  49872=>"111100111",
  49873=>"000000000",
  49874=>"001001001",
  49875=>"100100000",
  49876=>"101000000",
  49877=>"111111111",
  49878=>"011111111",
  49879=>"111111111",
  49880=>"001000001",
  49881=>"100101000",
  49882=>"110110111",
  49883=>"001001000",
  49884=>"100000000",
  49885=>"000000010",
  49886=>"111111100",
  49887=>"011011111",
  49888=>"111111111",
  49889=>"000111110",
  49890=>"110111111",
  49891=>"111111101",
  49892=>"000000001",
  49893=>"000100000",
  49894=>"000000000",
  49895=>"111111111",
  49896=>"111001000",
  49897=>"000001000",
  49898=>"100100000",
  49899=>"000000000",
  49900=>"111111111",
  49901=>"111111111",
  49902=>"001001000",
  49903=>"111111111",
  49904=>"000000000",
  49905=>"110111111",
  49906=>"000000000",
  49907=>"000000000",
  49908=>"011010011",
  49909=>"110100110",
  49910=>"100000100",
  49911=>"000000000",
  49912=>"101111000",
  49913=>"111001001",
  49914=>"000000000",
  49915=>"000000000",
  49916=>"111111111",
  49917=>"111111111",
  49918=>"111111000",
  49919=>"000000001",
  49920=>"000101100",
  49921=>"111111111",
  49922=>"000000000",
  49923=>"000000111",
  49924=>"111000010",
  49925=>"111101000",
  49926=>"111111111",
  49927=>"111011111",
  49928=>"111111101",
  49929=>"111011011",
  49930=>"111101111",
  49931=>"000000000",
  49932=>"100000000",
  49933=>"000000001",
  49934=>"111111000",
  49935=>"000000000",
  49936=>"010000000",
  49937=>"111001000",
  49938=>"111111111",
  49939=>"111111111",
  49940=>"000000000",
  49941=>"111111111",
  49942=>"110110110",
  49943=>"000000000",
  49944=>"000000000",
  49945=>"000000000",
  49946=>"000000000",
  49947=>"110000001",
  49948=>"101001001",
  49949=>"111111111",
  49950=>"111111111",
  49951=>"111101000",
  49952=>"110110111",
  49953=>"111111110",
  49954=>"000110111",
  49955=>"111111110",
  49956=>"111111111",
  49957=>"110000000",
  49958=>"001000000",
  49959=>"001100111",
  49960=>"100000111",
  49961=>"000000000",
  49962=>"000000000",
  49963=>"000100110",
  49964=>"011000000",
  49965=>"110111111",
  49966=>"111011111",
  49967=>"111111101",
  49968=>"001111000",
  49969=>"011111111",
  49970=>"011111011",
  49971=>"111111111",
  49972=>"110000000",
  49973=>"000000000",
  49974=>"111111101",
  49975=>"111111111",
  49976=>"000000000",
  49977=>"111111111",
  49978=>"110111000",
  49979=>"111111111",
  49980=>"011001001",
  49981=>"111100000",
  49982=>"000000000",
  49983=>"000000000",
  49984=>"111000111",
  49985=>"000000000",
  49986=>"000000000",
  49987=>"000000000",
  49988=>"111111111",
  49989=>"000000110",
  49990=>"100111000",
  49991=>"000000000",
  49992=>"111111111",
  49993=>"100111111",
  49994=>"000000000",
  49995=>"111011111",
  49996=>"000000111",
  49997=>"000000000",
  49998=>"100000001",
  49999=>"111001000",
  50000=>"111011001",
  50001=>"001000000",
  50002=>"000000001",
  50003=>"010000000",
  50004=>"111110100",
  50005=>"101000000",
  50006=>"000000000",
  50007=>"101000000",
  50008=>"000000000",
  50009=>"000000000",
  50010=>"000100111",
  50011=>"000000000",
  50012=>"111111111",
  50013=>"000000000",
  50014=>"000000000",
  50015=>"000000000",
  50016=>"111111111",
  50017=>"111111011",
  50018=>"010000000",
  50019=>"011011001",
  50020=>"001001111",
  50021=>"000000000",
  50022=>"000000000",
  50023=>"111110000",
  50024=>"111111111",
  50025=>"000000000",
  50026=>"000000000",
  50027=>"111111111",
  50028=>"010011011",
  50029=>"001000000",
  50030=>"111000000",
  50031=>"111000111",
  50032=>"100100111",
  50033=>"111111111",
  50034=>"000000011",
  50035=>"000000000",
  50036=>"111111111",
  50037=>"000000001",
  50038=>"111101101",
  50039=>"111111000",
  50040=>"111111001",
  50041=>"001001001",
  50042=>"100100000",
  50043=>"111111000",
  50044=>"001000101",
  50045=>"111111111",
  50046=>"111001001",
  50047=>"111101000",
  50048=>"001000000",
  50049=>"111111101",
  50050=>"110100111",
  50051=>"111111000",
  50052=>"000010011",
  50053=>"011011011",
  50054=>"111001001",
  50055=>"000000001",
  50056=>"111111111",
  50057=>"011011011",
  50058=>"111000000",
  50059=>"011011011",
  50060=>"111110000",
  50061=>"100110010",
  50062=>"000000000",
  50063=>"011111111",
  50064=>"011111011",
  50065=>"000000001",
  50066=>"000000000",
  50067=>"100101101",
  50068=>"111111111",
  50069=>"000000100",
  50070=>"111110110",
  50071=>"011111111",
  50072=>"111110000",
  50073=>"111111100",
  50074=>"101111110",
  50075=>"101101000",
  50076=>"100000111",
  50077=>"000000000",
  50078=>"001000001",
  50079=>"000111110",
  50080=>"000000000",
  50081=>"100100110",
  50082=>"101001111",
  50083=>"000000001",
  50084=>"100000000",
  50085=>"000000000",
  50086=>"000001111",
  50087=>"000000000",
  50088=>"001001110",
  50089=>"011010111",
  50090=>"000000000",
  50091=>"110100000",
  50092=>"001011000",
  50093=>"000000000",
  50094=>"111111110",
  50095=>"111111011",
  50096=>"111111011",
  50097=>"000000000",
  50098=>"000000000",
  50099=>"111100000",
  50100=>"110110110",
  50101=>"000000000",
  50102=>"000010011",
  50103=>"111101111",
  50104=>"111111111",
  50105=>"111111111",
  50106=>"000000100",
  50107=>"100100110",
  50108=>"111111111",
  50109=>"111111111",
  50110=>"011110110",
  50111=>"111111111",
  50112=>"110111111",
  50113=>"110000110",
  50114=>"111111111",
  50115=>"100111011",
  50116=>"100100000",
  50117=>"001011111",
  50118=>"001100100",
  50119=>"000011111",
  50120=>"111111000",
  50121=>"111111111",
  50122=>"000000111",
  50123=>"000000000",
  50124=>"111100000",
  50125=>"000000100",
  50126=>"001001001",
  50127=>"000000000",
  50128=>"111111011",
  50129=>"000000000",
  50130=>"000000000",
  50131=>"100111111",
  50132=>"110110111",
  50133=>"000000100",
  50134=>"111111011",
  50135=>"000100100",
  50136=>"111100000",
  50137=>"110000000",
  50138=>"110110111",
  50139=>"000011111",
  50140=>"101100100",
  50141=>"001000111",
  50142=>"000000010",
  50143=>"110100100",
  50144=>"111111111",
  50145=>"000000111",
  50146=>"110111111",
  50147=>"110110111",
  50148=>"111011111",
  50149=>"000000000",
  50150=>"001000000",
  50151=>"011001101",
  50152=>"111111100",
  50153=>"000000000",
  50154=>"000000000",
  50155=>"111001001",
  50156=>"111111111",
  50157=>"001001111",
  50158=>"000000011",
  50159=>"111100100",
  50160=>"111111000",
  50161=>"000000000",
  50162=>"111111101",
  50163=>"100111111",
  50164=>"111111001",
  50165=>"111111101",
  50166=>"111000000",
  50167=>"000000000",
  50168=>"111111111",
  50169=>"011001000",
  50170=>"110110000",
  50171=>"111001000",
  50172=>"111111111",
  50173=>"101101111",
  50174=>"011001000",
  50175=>"000000000",
  50176=>"001111111",
  50177=>"000000000",
  50178=>"000011111",
  50179=>"000011111",
  50180=>"111111111",
  50181=>"000000010",
  50182=>"111111100",
  50183=>"111000000",
  50184=>"000000000",
  50185=>"110001000",
  50186=>"111000001",
  50187=>"010110111",
  50188=>"011111110",
  50189=>"111111000",
  50190=>"000000000",
  50191=>"001111110",
  50192=>"000110111",
  50193=>"011111111",
  50194=>"111101000",
  50195=>"111011000",
  50196=>"000110000",
  50197=>"000000111",
  50198=>"000000000",
  50199=>"111111111",
  50200=>"110111000",
  50201=>"001000111",
  50202=>"111001000",
  50203=>"011111111",
  50204=>"111111111",
  50205=>"000110111",
  50206=>"001001101",
  50207=>"100110111",
  50208=>"000011011",
  50209=>"111000000",
  50210=>"111111000",
  50211=>"111000000",
  50212=>"000000000",
  50213=>"111111111",
  50214=>"111111111",
  50215=>"100100111",
  50216=>"111111111",
  50217=>"111000000",
  50218=>"111111111",
  50219=>"111111011",
  50220=>"000000111",
  50221=>"111001000",
  50222=>"000000111",
  50223=>"000000000",
  50224=>"000001111",
  50225=>"111001000",
  50226=>"111111000",
  50227=>"101000000",
  50228=>"001001000",
  50229=>"011011011",
  50230=>"111111111",
  50231=>"000001111",
  50232=>"111111111",
  50233=>"000000000",
  50234=>"000110110",
  50235=>"000101000",
  50236=>"111111010",
  50237=>"000000001",
  50238=>"111111110",
  50239=>"000000011",
  50240=>"000000100",
  50241=>"001001111",
  50242=>"000000000",
  50243=>"100100111",
  50244=>"011000000",
  50245=>"001001011",
  50246=>"000000000",
  50247=>"001000000",
  50248=>"000000000",
  50249=>"000100000",
  50250=>"111111000",
  50251=>"101000001",
  50252=>"000111111",
  50253=>"000000100",
  50254=>"000011000",
  50255=>"111111111",
  50256=>"110000000",
  50257=>"111110000",
  50258=>"111111000",
  50259=>"110110000",
  50260=>"000000000",
  50261=>"110000000",
  50262=>"000000100",
  50263=>"000000000",
  50264=>"111111010",
  50265=>"100000000",
  50266=>"000000000",
  50267=>"111110100",
  50268=>"000000111",
  50269=>"111111111",
  50270=>"000000000",
  50271=>"000000011",
  50272=>"111111000",
  50273=>"111111111",
  50274=>"000111111",
  50275=>"111111001",
  50276=>"110110000",
  50277=>"111111000",
  50278=>"000000000",
  50279=>"111111111",
  50280=>"000000010",
  50281=>"110000101",
  50282=>"111000111",
  50283=>"000000000",
  50284=>"111011011",
  50285=>"111000000",
  50286=>"111111111",
  50287=>"110011000",
  50288=>"100000000",
  50289=>"000000001",
  50290=>"000000111",
  50291=>"000000000",
  50292=>"111111100",
  50293=>"000000000",
  50294=>"111111111",
  50295=>"111101011",
  50296=>"000000000",
  50297=>"101100100",
  50298=>"010000000",
  50299=>"011001111",
  50300=>"110110000",
  50301=>"000111111",
  50302=>"111101001",
  50303=>"000000000",
  50304=>"111000000",
  50305=>"000000111",
  50306=>"000000000",
  50307=>"111111011",
  50308=>"001000011",
  50309=>"111011100",
  50310=>"111111111",
  50311=>"100100110",
  50312=>"111111110",
  50313=>"100000000",
  50314=>"111111000",
  50315=>"111111111",
  50316=>"000001000",
  50317=>"111111111",
  50318=>"111111000",
  50319=>"000000000",
  50320=>"100100100",
  50321=>"010000000",
  50322=>"000000000",
  50323=>"000000000",
  50324=>"010111111",
  50325=>"000000111",
  50326=>"000000000",
  50327=>"101001000",
  50328=>"000000111",
  50329=>"011111110",
  50330=>"111111111",
  50331=>"000010011",
  50332=>"000000001",
  50333=>"101110000",
  50334=>"000110111",
  50335=>"000111000",
  50336=>"111111111",
  50337=>"001000100",
  50338=>"111111111",
  50339=>"111100000",
  50340=>"000001000",
  50341=>"001001000",
  50342=>"011111000",
  50343=>"000000000",
  50344=>"111100100",
  50345=>"110000000",
  50346=>"000000111",
  50347=>"000000001",
  50348=>"110111111",
  50349=>"101100000",
  50350=>"001000111",
  50351=>"111000000",
  50352=>"000001111",
  50353=>"111100100",
  50354=>"011111011",
  50355=>"000000000",
  50356=>"111011001",
  50357=>"101000000",
  50358=>"000000000",
  50359=>"000111111",
  50360=>"101111111",
  50361=>"000010000",
  50362=>"000000000",
  50363=>"000000111",
  50364=>"111111111",
  50365=>"000000111",
  50366=>"000111111",
  50367=>"000000111",
  50368=>"000100111",
  50369=>"000000000",
  50370=>"011111111",
  50371=>"111000000",
  50372=>"000000000",
  50373=>"000111111",
  50374=>"110011000",
  50375=>"000000000",
  50376=>"000000011",
  50377=>"000010111",
  50378=>"100100111",
  50379=>"100011001",
  50380=>"111110110",
  50381=>"000000101",
  50382=>"111111001",
  50383=>"011111100",
  50384=>"001000000",
  50385=>"110111011",
  50386=>"000000000",
  50387=>"111000010",
  50388=>"000000000",
  50389=>"111110111",
  50390=>"111111111",
  50391=>"000001111",
  50392=>"111000111",
  50393=>"111111111",
  50394=>"011111000",
  50395=>"111100100",
  50396=>"111110000",
  50397=>"011010111",
  50398=>"000000000",
  50399=>"011111111",
  50400=>"111111011",
  50401=>"111111111",
  50402=>"111011000",
  50403=>"000000111",
  50404=>"000110110",
  50405=>"111011011",
  50406=>"111111000",
  50407=>"001001111",
  50408=>"000000001",
  50409=>"110111011",
  50410=>"101001000",
  50411=>"000100000",
  50412=>"001011111",
  50413=>"111110000",
  50414=>"000000001",
  50415=>"011000000",
  50416=>"101000000",
  50417=>"000000001",
  50418=>"000111111",
  50419=>"001000001",
  50420=>"001111111",
  50421=>"111111110",
  50422=>"000000111",
  50423=>"111000001",
  50424=>"111000000",
  50425=>"111000000",
  50426=>"001000000",
  50427=>"111111111",
  50428=>"000000110",
  50429=>"011011111",
  50430=>"111000101",
  50431=>"001000000",
  50432=>"001101101",
  50433=>"111111000",
  50434=>"001001111",
  50435=>"111111111",
  50436=>"111101000",
  50437=>"001111111",
  50438=>"100000101",
  50439=>"000001111",
  50440=>"111011000",
  50441=>"111110111",
  50442=>"111111111",
  50443=>"000111111",
  50444=>"111111111",
  50445=>"000000000",
  50446=>"000101100",
  50447=>"000111111",
  50448=>"111111100",
  50449=>"000000000",
  50450=>"000000011",
  50451=>"010111111",
  50452=>"100110111",
  50453=>"000111111",
  50454=>"000000000",
  50455=>"010000100",
  50456=>"000000001",
  50457=>"010000000",
  50458=>"111001000",
  50459=>"000000000",
  50460=>"110111011",
  50461=>"000000000",
  50462=>"111111111",
  50463=>"000000101",
  50464=>"010010110",
  50465=>"111010000",
  50466=>"000000000",
  50467=>"111111110",
  50468=>"000000100",
  50469=>"001000000",
  50470=>"010000000",
  50471=>"000000111",
  50472=>"110110111",
  50473=>"000000000",
  50474=>"100100111",
  50475=>"010010111",
  50476=>"111001111",
  50477=>"100100001",
  50478=>"111111110",
  50479=>"000000000",
  50480=>"111100100",
  50481=>"111000000",
  50482=>"111100100",
  50483=>"111111000",
  50484=>"000111111",
  50485=>"000111111",
  50486=>"000001111",
  50487=>"111000000",
  50488=>"111111011",
  50489=>"111000000",
  50490=>"000000000",
  50491=>"001101000",
  50492=>"111111111",
  50493=>"000000111",
  50494=>"000000000",
  50495=>"000000000",
  50496=>"000000000",
  50497=>"111100000",
  50498=>"000000100",
  50499=>"000000111",
  50500=>"110111110",
  50501=>"111111111",
  50502=>"110111111",
  50503=>"111111100",
  50504=>"111111111",
  50505=>"000000000",
  50506=>"100000000",
  50507=>"001001000",
  50508=>"000000001",
  50509=>"000000000",
  50510=>"000000000",
  50511=>"001011011",
  50512=>"111011111",
  50513=>"000000000",
  50514=>"111111111",
  50515=>"111111111",
  50516=>"000011000",
  50517=>"011011011",
  50518=>"000000000",
  50519=>"111100000",
  50520=>"001011111",
  50521=>"001111111",
  50522=>"111111000",
  50523=>"000000111",
  50524=>"011001111",
  50525=>"000000100",
  50526=>"111001000",
  50527=>"000010011",
  50528=>"000000000",
  50529=>"000000001",
  50530=>"000110110",
  50531=>"111111111",
  50532=>"000111111",
  50533=>"000100111",
  50534=>"001000000",
  50535=>"000111111",
  50536=>"111001001",
  50537=>"111111111",
  50538=>"111000000",
  50539=>"001011111",
  50540=>"001001100",
  50541=>"000000000",
  50542=>"000000100",
  50543=>"101111100",
  50544=>"001111011",
  50545=>"011111111",
  50546=>"110000000",
  50547=>"001000000",
  50548=>"000000110",
  50549=>"100000000",
  50550=>"111000110",
  50551=>"111111100",
  50552=>"000000000",
  50553=>"000000000",
  50554=>"000000000",
  50555=>"111010001",
  50556=>"000000000",
  50557=>"000000000",
  50558=>"101111111",
  50559=>"000111111",
  50560=>"111001000",
  50561=>"000111001",
  50562=>"100100100",
  50563=>"111100100",
  50564=>"111000000",
  50565=>"111111111",
  50566=>"111111000",
  50567=>"111111000",
  50568=>"000111111",
  50569=>"111111111",
  50570=>"000000000",
  50571=>"110111111",
  50572=>"101101111",
  50573=>"110111111",
  50574=>"001001000",
  50575=>"000000000",
  50576=>"000000000",
  50577=>"100000000",
  50578=>"111000000",
  50579=>"100100110",
  50580=>"000000111",
  50581=>"000000000",
  50582=>"100100000",
  50583=>"111111100",
  50584=>"000000000",
  50585=>"000000000",
  50586=>"111111001",
  50587=>"010111111",
  50588=>"001111111",
  50589=>"100001101",
  50590=>"010111111",
  50591=>"000000001",
  50592=>"110011100",
  50593=>"011000000",
  50594=>"111000000",
  50595=>"110110000",
  50596=>"000000110",
  50597=>"111000000",
  50598=>"100100000",
  50599=>"010110010",
  50600=>"000001001",
  50601=>"000000000",
  50602=>"000000000",
  50603=>"000000000",
  50604=>"000000000",
  50605=>"111111111",
  50606=>"111101100",
  50607=>"000000000",
  50608=>"000000000",
  50609=>"010011001",
  50610=>"111111000",
  50611=>"000000000",
  50612=>"000000000",
  50613=>"111111000",
  50614=>"111111110",
  50615=>"011111000",
  50616=>"111010000",
  50617=>"000001001",
  50618=>"111010001",
  50619=>"000100111",
  50620=>"000011111",
  50621=>"101111111",
  50622=>"110111111",
  50623=>"011110111",
  50624=>"100000000",
  50625=>"111111110",
  50626=>"111110111",
  50627=>"111011000",
  50628=>"001000000",
  50629=>"111000011",
  50630=>"000000111",
  50631=>"000100000",
  50632=>"111111111",
  50633=>"100000000",
  50634=>"100000000",
  50635=>"111000111",
  50636=>"000000000",
  50637=>"111111111",
  50638=>"000000011",
  50639=>"011000100",
  50640=>"000000000",
  50641=>"001111001",
  50642=>"111011011",
  50643=>"111111111",
  50644=>"000000111",
  50645=>"000000000",
  50646=>"000000000",
  50647=>"110111001",
  50648=>"111111110",
  50649=>"000101000",
  50650=>"000010000",
  50651=>"100000100",
  50652=>"000000100",
  50653=>"000000000",
  50654=>"010000000",
  50655=>"110111111",
  50656=>"100000000",
  50657=>"110000000",
  50658=>"000000000",
  50659=>"100111111",
  50660=>"000000000",
  50661=>"111111111",
  50662=>"000110110",
  50663=>"000001000",
  50664=>"000000001",
  50665=>"111111110",
  50666=>"000011111",
  50667=>"111011000",
  50668=>"000011111",
  50669=>"110011001",
  50670=>"000000000",
  50671=>"000100110",
  50672=>"111111000",
  50673=>"111111111",
  50674=>"111111111",
  50675=>"000101111",
  50676=>"000011111",
  50677=>"000011001",
  50678=>"001000000",
  50679=>"111111000",
  50680=>"111111100",
  50681=>"001001011",
  50682=>"111110110",
  50683=>"100000100",
  50684=>"010111111",
  50685=>"000001001",
  50686=>"000000000",
  50687=>"000000000",
  50688=>"111100000",
  50689=>"110110110",
  50690=>"111011111",
  50691=>"111111010",
  50692=>"111111111",
  50693=>"000010000",
  50694=>"000111111",
  50695=>"111101101",
  50696=>"000000000",
  50697=>"000000111",
  50698=>"111111010",
  50699=>"111000000",
  50700=>"111111111",
  50701=>"000000000",
  50702=>"001101111",
  50703=>"000000000",
  50704=>"111001000",
  50705=>"010000000",
  50706=>"111111011",
  50707=>"000000000",
  50708=>"101110110",
  50709=>"111111111",
  50710=>"100111111",
  50711=>"011011001",
  50712=>"001011000",
  50713=>"101001011",
  50714=>"111111111",
  50715=>"100000000",
  50716=>"100100000",
  50717=>"111111111",
  50718=>"100000111",
  50719=>"010010010",
  50720=>"111010000",
  50721=>"110110110",
  50722=>"110110100",
  50723=>"111111000",
  50724=>"000101101",
  50725=>"000000000",
  50726=>"111111111",
  50727=>"000000110",
  50728=>"111111101",
  50729=>"010011001",
  50730=>"111111111",
  50731=>"110111010",
  50732=>"000000100",
  50733=>"110110000",
  50734=>"111001100",
  50735=>"111111111",
  50736=>"000000000",
  50737=>"000000111",
  50738=>"001000111",
  50739=>"000000000",
  50740=>"111111111",
  50741=>"100000000",
  50742=>"001001001",
  50743=>"000000011",
  50744=>"111111001",
  50745=>"000000010",
  50746=>"111111111",
  50747=>"110000000",
  50748=>"100101111",
  50749=>"001001001",
  50750=>"111111101",
  50751=>"001000000",
  50752=>"001000000",
  50753=>"111101001",
  50754=>"001001001",
  50755=>"000000110",
  50756=>"101011001",
  50757=>"000000111",
  50758=>"110010010",
  50759=>"000000000",
  50760=>"111111100",
  50761=>"110110111",
  50762=>"111111101",
  50763=>"000000001",
  50764=>"011011111",
  50765=>"001011000",
  50766=>"000000000",
  50767=>"111000000",
  50768=>"000110111",
  50769=>"111111000",
  50770=>"000000001",
  50771=>"000100101",
  50772=>"011011000",
  50773=>"010111111",
  50774=>"001111100",
  50775=>"111111111",
  50776=>"000000111",
  50777=>"101000000",
  50778=>"111111111",
  50779=>"001110110",
  50780=>"000000111",
  50781=>"000000000",
  50782=>"000000000",
  50783=>"000100000",
  50784=>"111001111",
  50785=>"000010000",
  50786=>"111111111",
  50787=>"111111000",
  50788=>"010010000",
  50789=>"011111111",
  50790=>"011000000",
  50791=>"001000000",
  50792=>"000000111",
  50793=>"111111001",
  50794=>"111111011",
  50795=>"110110010",
  50796=>"110111111",
  50797=>"111111111",
  50798=>"111001101",
  50799=>"000000000",
  50800=>"011000000",
  50801=>"001001111",
  50802=>"001001000",
  50803=>"011000010",
  50804=>"001111111",
  50805=>"111111110",
  50806=>"011001000",
  50807=>"011011011",
  50808=>"111111101",
  50809=>"000000000",
  50810=>"110000010",
  50811=>"001000000",
  50812=>"100100101",
  50813=>"000000000",
  50814=>"111111011",
  50815=>"110100000",
  50816=>"110000000",
  50817=>"100100011",
  50818=>"110000000",
  50819=>"010000000",
  50820=>"010000000",
  50821=>"111111101",
  50822=>"000000001",
  50823=>"110000000",
  50824=>"010110010",
  50825=>"000000000",
  50826=>"000010011",
  50827=>"000000000",
  50828=>"000000000",
  50829=>"000001111",
  50830=>"101111111",
  50831=>"000000000",
  50832=>"111101101",
  50833=>"000000000",
  50834=>"000111001",
  50835=>"000000000",
  50836=>"111111111",
  50837=>"000000000",
  50838=>"010000000",
  50839=>"101000100",
  50840=>"000000101",
  50841=>"111111111",
  50842=>"111111111",
  50843=>"111110000",
  50844=>"101000000",
  50845=>"111000000",
  50846=>"111011011",
  50847=>"001001001",
  50848=>"110111111",
  50849=>"010110000",
  50850=>"000000000",
  50851=>"000000111",
  50852=>"001000111",
  50853=>"010000000",
  50854=>"000100001",
  50855=>"001001101",
  50856=>"111111011",
  50857=>"001001001",
  50858=>"110111110",
  50859=>"000000001",
  50860=>"001000000",
  50861=>"100011111",
  50862=>"000000000",
  50863=>"100000000",
  50864=>"000100111",
  50865=>"111100100",
  50866=>"111111111",
  50867=>"000000101",
  50868=>"011011111",
  50869=>"111111111",
  50870=>"000000101",
  50871=>"011000000",
  50872=>"000000101",
  50873=>"101111111",
  50874=>"000110111",
  50875=>"110110111",
  50876=>"000110000",
  50877=>"111110110",
  50878=>"000000000",
  50879=>"110110000",
  50880=>"000000101",
  50881=>"111001000",
  50882=>"110000000",
  50883=>"001000001",
  50884=>"000000000",
  50885=>"000000000",
  50886=>"111111111",
  50887=>"110000000",
  50888=>"000000000",
  50889=>"001000000",
  50890=>"111100000",
  50891=>"110111110",
  50892=>"000000000",
  50893=>"000000100",
  50894=>"111111110",
  50895=>"000100000",
  50896=>"000000110",
  50897=>"000000000",
  50898=>"111000111",
  50899=>"000000010",
  50900=>"000000100",
  50901=>"000000111",
  50902=>"000000000",
  50903=>"111111111",
  50904=>"000000000",
  50905=>"000011111",
  50906=>"111111111",
  50907=>"000000000",
  50908=>"110110111",
  50909=>"111111111",
  50910=>"000000000",
  50911=>"000000000",
  50912=>"111001000",
  50913=>"000000000",
  50914=>"000000010",
  50915=>"010001111",
  50916=>"000001000",
  50917=>"100111101",
  50918=>"001000100",
  50919=>"000000000",
  50920=>"011111011",
  50921=>"111111110",
  50922=>"000000001",
  50923=>"001000000",
  50924=>"000000111",
  50925=>"000000000",
  50926=>"100100110",
  50927=>"110110011",
  50928=>"000000000",
  50929=>"101101001",
  50930=>"100000100",
  50931=>"110110110",
  50932=>"000000001",
  50933=>"010111011",
  50934=>"000000000",
  50935=>"001000000",
  50936=>"000001101",
  50937=>"000001011",
  50938=>"011111000",
  50939=>"111101000",
  50940=>"110110110",
  50941=>"111010110",
  50942=>"000000000",
  50943=>"000110111",
  50944=>"111011010",
  50945=>"111111111",
  50946=>"000000000",
  50947=>"011111000",
  50948=>"000000111",
  50949=>"000001001",
  50950=>"011001111",
  50951=>"111101111",
  50952=>"100111111",
  50953=>"000000000",
  50954=>"001000000",
  50955=>"111111111",
  50956=>"011011111",
  50957=>"010011111",
  50958=>"000000000",
  50959=>"010111001",
  50960=>"000000011",
  50961=>"110000000",
  50962=>"111111101",
  50963=>"001111111",
  50964=>"111111111",
  50965=>"101101000",
  50966=>"000000100",
  50967=>"111111111",
  50968=>"000000001",
  50969=>"111111111",
  50970=>"110010000",
  50971=>"001000000",
  50972=>"111111110",
  50973=>"000000100",
  50974=>"000001000",
  50975=>"111000000",
  50976=>"000100110",
  50977=>"000000000",
  50978=>"110111011",
  50979=>"111000000",
  50980=>"100111111",
  50981=>"110110110",
  50982=>"011000000",
  50983=>"000000001",
  50984=>"100000100",
  50985=>"111000000",
  50986=>"010110111",
  50987=>"000000110",
  50988=>"100101100",
  50989=>"111111110",
  50990=>"001011111",
  50991=>"000000000",
  50992=>"111011000",
  50993=>"111111110",
  50994=>"001111111",
  50995=>"111111111",
  50996=>"111001111",
  50997=>"000000000",
  50998=>"000000000",
  50999=>"000000111",
  51000=>"011000000",
  51001=>"101000101",
  51002=>"000000000",
  51003=>"111000111",
  51004=>"011011001",
  51005=>"100101111",
  51006=>"010011011",
  51007=>"000011111",
  51008=>"000000000",
  51009=>"111111010",
  51010=>"000000101",
  51011=>"111110110",
  51012=>"000000000",
  51013=>"000100100",
  51014=>"000000111",
  51015=>"111111111",
  51016=>"111111111",
  51017=>"000000000",
  51018=>"000000000",
  51019=>"111111111",
  51020=>"000000000",
  51021=>"000000000",
  51022=>"011111111",
  51023=>"000000000",
  51024=>"100011011",
  51025=>"000000000",
  51026=>"000000000",
  51027=>"000000100",
  51028=>"110100100",
  51029=>"011011011",
  51030=>"000000100",
  51031=>"001000111",
  51032=>"111111111",
  51033=>"110010110",
  51034=>"111101111",
  51035=>"110010000",
  51036=>"000000111",
  51037=>"000000000",
  51038=>"110110110",
  51039=>"000000111",
  51040=>"000000000",
  51041=>"000000000",
  51042=>"110000000",
  51043=>"000000000",
  51044=>"000000001",
  51045=>"110111111",
  51046=>"000010000",
  51047=>"001001000",
  51048=>"001011011",
  51049=>"000000111",
  51050=>"001001111",
  51051=>"111010001",
  51052=>"000100101",
  51053=>"000110011",
  51054=>"000000000",
  51055=>"111111111",
  51056=>"111110111",
  51057=>"001111111",
  51058=>"010000111",
  51059=>"000000100",
  51060=>"000000101",
  51061=>"001001111",
  51062=>"000000000",
  51063=>"000000000",
  51064=>"111011111",
  51065=>"111111110",
  51066=>"000110111",
  51067=>"111111111",
  51068=>"000000001",
  51069=>"000000111",
  51070=>"100111000",
  51071=>"000000000",
  51072=>"100000100",
  51073=>"100000100",
  51074=>"111111111",
  51075=>"000011011",
  51076=>"000000100",
  51077=>"000110111",
  51078=>"000000000",
  51079=>"001011000",
  51080=>"111111111",
  51081=>"111101001",
  51082=>"100000000",
  51083=>"111011010",
  51084=>"111111101",
  51085=>"100100111",
  51086=>"111111000",
  51087=>"000000111",
  51088=>"000000000",
  51089=>"111111111",
  51090=>"000000000",
  51091=>"001001111",
  51092=>"111111111",
  51093=>"000000000",
  51094=>"100100000",
  51095=>"000000000",
  51096=>"111001000",
  51097=>"000000111",
  51098=>"110100000",
  51099=>"000001111",
  51100=>"000001101",
  51101=>"010000000",
  51102=>"000000000",
  51103=>"111111111",
  51104=>"000000011",
  51105=>"111011111",
  51106=>"000011000",
  51107=>"000000111",
  51108=>"000000100",
  51109=>"111000100",
  51110=>"111001111",
  51111=>"111111011",
  51112=>"000000000",
  51113=>"101111111",
  51114=>"111111111",
  51115=>"111001101",
  51116=>"010011000",
  51117=>"011001000",
  51118=>"000000000",
  51119=>"000000000",
  51120=>"000111001",
  51121=>"000000000",
  51122=>"001011111",
  51123=>"111111111",
  51124=>"000100111",
  51125=>"110101000",
  51126=>"111111111",
  51127=>"000101110",
  51128=>"000000100",
  51129=>"010111111",
  51130=>"111001001",
  51131=>"111111111",
  51132=>"101001001",
  51133=>"001000000",
  51134=>"000000000",
  51135=>"101101111",
  51136=>"001000111",
  51137=>"000000010",
  51138=>"110110000",
  51139=>"101101100",
  51140=>"111011111",
  51141=>"111111111",
  51142=>"000000000",
  51143=>"111111010",
  51144=>"111001000",
  51145=>"000011111",
  51146=>"000000000",
  51147=>"100000110",
  51148=>"100000001",
  51149=>"000010111",
  51150=>"111101101",
  51151=>"010111111",
  51152=>"001000000",
  51153=>"100110111",
  51154=>"000000101",
  51155=>"111101101",
  51156=>"111111111",
  51157=>"001101001",
  51158=>"000001001",
  51159=>"011101111",
  51160=>"000000000",
  51161=>"011011000",
  51162=>"111111111",
  51163=>"111111110",
  51164=>"110111111",
  51165=>"111101111",
  51166=>"111111100",
  51167=>"100000100",
  51168=>"001000000",
  51169=>"000001011",
  51170=>"000111111",
  51171=>"000000000",
  51172=>"111111111",
  51173=>"101001000",
  51174=>"111111111",
  51175=>"000000000",
  51176=>"010010000",
  51177=>"111111111",
  51178=>"000000000",
  51179=>"111111010",
  51180=>"000000000",
  51181=>"111111000",
  51182=>"110000000",
  51183=>"110111111",
  51184=>"000110111",
  51185=>"000000000",
  51186=>"000000001",
  51187=>"010011010",
  51188=>"000000111",
  51189=>"000000000",
  51190=>"000001101",
  51191=>"000100100",
  51192=>"100000000",
  51193=>"000000000",
  51194=>"001001111",
  51195=>"001000000",
  51196=>"111001011",
  51197=>"000000001",
  51198=>"010111111",
  51199=>"001011111",
  51200=>"100000101",
  51201=>"101011000",
  51202=>"101000000",
  51203=>"011000000",
  51204=>"000010111",
  51205=>"111111111",
  51206=>"001000011",
  51207=>"111111111",
  51208=>"000110111",
  51209=>"011111111",
  51210=>"010001111",
  51211=>"000000110",
  51212=>"111110000",
  51213=>"111100100",
  51214=>"000110000",
  51215=>"111111011",
  51216=>"111001001",
  51217=>"000000111",
  51218=>"011111111",
  51219=>"010010111",
  51220=>"011001011",
  51221=>"000000111",
  51222=>"000000111",
  51223=>"000000000",
  51224=>"111111000",
  51225=>"111001001",
  51226=>"000000111",
  51227=>"000000000",
  51228=>"111111010",
  51229=>"110000001",
  51230=>"000110000",
  51231=>"000000000",
  51232=>"010011000",
  51233=>"111111111",
  51234=>"111111000",
  51235=>"111000011",
  51236=>"000000000",
  51237=>"111000000",
  51238=>"000011111",
  51239=>"111000001",
  51240=>"100000001",
  51241=>"001001111",
  51242=>"101000101",
  51243=>"111110110",
  51244=>"110110111",
  51245=>"111111101",
  51246=>"100110111",
  51247=>"001101111",
  51248=>"000000100",
  51249=>"101000000",
  51250=>"100000000",
  51251=>"011010010",
  51252=>"000111011",
  51253=>"100001001",
  51254=>"111001000",
  51255=>"111111111",
  51256=>"000100000",
  51257=>"111111111",
  51258=>"000000001",
  51259=>"000000000",
  51260=>"111111101",
  51261=>"001000000",
  51262=>"000100110",
  51263=>"110100000",
  51264=>"011111000",
  51265=>"111111000",
  51266=>"001011111",
  51267=>"011000000",
  51268=>"001000100",
  51269=>"110000000",
  51270=>"000000000",
  51271=>"000000000",
  51272=>"011111101",
  51273=>"000000111",
  51274=>"100111111",
  51275=>"001110110",
  51276=>"110000000",
  51277=>"110100110",
  51278=>"011001011",
  51279=>"111111111",
  51280=>"110111101",
  51281=>"100000111",
  51282=>"000000001",
  51283=>"011001100",
  51284=>"111111111",
  51285=>"000010110",
  51286=>"101000100",
  51287=>"110000001",
  51288=>"000000101",
  51289=>"100000000",
  51290=>"000000001",
  51291=>"000000111",
  51292=>"111111111",
  51293=>"000111111",
  51294=>"111000000",
  51295=>"111111111",
  51296=>"000000000",
  51297=>"000000011",
  51298=>"111111110",
  51299=>"000001000",
  51300=>"001000000",
  51301=>"010111000",
  51302=>"111000111",
  51303=>"010000111",
  51304=>"111000010",
  51305=>"111111100",
  51306=>"001011111",
  51307=>"000011001",
  51308=>"000110100",
  51309=>"000000110",
  51310=>"111111111",
  51311=>"000110111",
  51312=>"100000000",
  51313=>"000000111",
  51314=>"000000000",
  51315=>"111111101",
  51316=>"011011011",
  51317=>"000000000",
  51318=>"011111000",
  51319=>"111111000",
  51320=>"000011000",
  51321=>"111000000",
  51322=>"111000000",
  51323=>"111111111",
  51324=>"110000000",
  51325=>"111011111",
  51326=>"000000110",
  51327=>"010111101",
  51328=>"111000000",
  51329=>"111111000",
  51330=>"111000000",
  51331=>"111101000",
  51332=>"001111111",
  51333=>"111101111",
  51334=>"011100000",
  51335=>"000000110",
  51336=>"110000000",
  51337=>"111010110",
  51338=>"000000000",
  51339=>"111111111",
  51340=>"111110101",
  51341=>"011011101",
  51342=>"101111111",
  51343=>"110111100",
  51344=>"000000001",
  51345=>"110111111",
  51346=>"011000010",
  51347=>"000010110",
  51348=>"111001000",
  51349=>"000011111",
  51350=>"000101111",
  51351=>"111000000",
  51352=>"000001111",
  51353=>"111111111",
  51354=>"000000000",
  51355=>"000111010",
  51356=>"000000101",
  51357=>"001000000",
  51358=>"111111111",
  51359=>"000011111",
  51360=>"000011000",
  51361=>"110011001",
  51362=>"111000010",
  51363=>"000000111",
  51364=>"000000000",
  51365=>"000000011",
  51366=>"111010000",
  51367=>"000100100",
  51368=>"111111111",
  51369=>"101111111",
  51370=>"010000000",
  51371=>"110001000",
  51372=>"101001000",
  51373=>"111110000",
  51374=>"100000000",
  51375=>"000000100",
  51376=>"111111111",
  51377=>"000000000",
  51378=>"110111010",
  51379=>"000001000",
  51380=>"000000000",
  51381=>"111111110",
  51382=>"000000000",
  51383=>"111111111",
  51384=>"111111111",
  51385=>"111111111",
  51386=>"000000001",
  51387=>"011111111",
  51388=>"111111111",
  51389=>"000111111",
  51390=>"111000001",
  51391=>"011111111",
  51392=>"100000110",
  51393=>"111111000",
  51394=>"010111111",
  51395=>"010111111",
  51396=>"000111000",
  51397=>"000110000",
  51398=>"111000000",
  51399=>"111111111",
  51400=>"011111111",
  51401=>"111111111",
  51402=>"111101111",
  51403=>"000000101",
  51404=>"111100001",
  51405=>"000000000",
  51406=>"001000000",
  51407=>"111000000",
  51408=>"111111111",
  51409=>"000000110",
  51410=>"000011111",
  51411=>"000000101",
  51412=>"111110100",
  51413=>"110000110",
  51414=>"111101001",
  51415=>"111111110",
  51416=>"001010000",
  51417=>"111111111",
  51418=>"000000111",
  51419=>"001111111",
  51420=>"011010000",
  51421=>"101110000",
  51422=>"000010111",
  51423=>"011111111",
  51424=>"111111111",
  51425=>"001111010",
  51426=>"010111000",
  51427=>"011001110",
  51428=>"111111111",
  51429=>"100000111",
  51430=>"111111111",
  51431=>"000110110",
  51432=>"000000111",
  51433=>"111111001",
  51434=>"001000000",
  51435=>"000000000",
  51436=>"111111111",
  51437=>"001000000",
  51438=>"000000001",
  51439=>"111000000",
  51440=>"001000010",
  51441=>"000000111",
  51442=>"000000000",
  51443=>"000000000",
  51444=>"011111111",
  51445=>"111111110",
  51446=>"000101111",
  51447=>"111000000",
  51448=>"111111111",
  51449=>"011111000",
  51450=>"111000111",
  51451=>"100101101",
  51452=>"000000000",
  51453=>"110010000",
  51454=>"010000011",
  51455=>"000000000",
  51456=>"001000000",
  51457=>"001000000",
  51458=>"111111000",
  51459=>"110110100",
  51460=>"000000011",
  51461=>"101001100",
  51462=>"000110111",
  51463=>"001001000",
  51464=>"011000110",
  51465=>"110100100",
  51466=>"000000101",
  51467=>"111111000",
  51468=>"000001101",
  51469=>"100110100",
  51470=>"110110110",
  51471=>"111101111",
  51472=>"010111111",
  51473=>"000000000",
  51474=>"110100100",
  51475=>"000000001",
  51476=>"000000111",
  51477=>"010111111",
  51478=>"110110110",
  51479=>"000110111",
  51480=>"000001001",
  51481=>"111110110",
  51482=>"000100000",
  51483=>"000111111",
  51484=>"100100100",
  51485=>"111111110",
  51486=>"000001111",
  51487=>"000100000",
  51488=>"100101011",
  51489=>"111111011",
  51490=>"001000000",
  51491=>"000001111",
  51492=>"000000000",
  51493=>"000001110",
  51494=>"101000000",
  51495=>"000010111",
  51496=>"110111110",
  51497=>"000000000",
  51498=>"000000000",
  51499=>"000000000",
  51500=>"000000010",
  51501=>"111110110",
  51502=>"000000000",
  51503=>"000001000",
  51504=>"111111111",
  51505=>"011011101",
  51506=>"111110110",
  51507=>"000001001",
  51508=>"111000101",
  51509=>"111010100",
  51510=>"011011010",
  51511=>"111001010",
  51512=>"000000110",
  51513=>"000010111",
  51514=>"000000111",
  51515=>"100000000",
  51516=>"111111011",
  51517=>"111000000",
  51518=>"000000000",
  51519=>"000000000",
  51520=>"000000110",
  51521=>"111000000",
  51522=>"001010000",
  51523=>"111100000",
  51524=>"000110010",
  51525=>"011111111",
  51526=>"100111111",
  51527=>"000000000",
  51528=>"010110110",
  51529=>"000000000",
  51530=>"100001111",
  51531=>"011111111",
  51532=>"000110111",
  51533=>"011010111",
  51534=>"000000111",
  51535=>"000000000",
  51536=>"010111001",
  51537=>"001001011",
  51538=>"000000000",
  51539=>"000000000",
  51540=>"110000000",
  51541=>"111001001",
  51542=>"100111111",
  51543=>"111100000",
  51544=>"111100111",
  51545=>"000000000",
  51546=>"111110000",
  51547=>"111111111",
  51548=>"000000000",
  51549=>"011111010",
  51550=>"101001111",
  51551=>"110111011",
  51552=>"110000111",
  51553=>"111100000",
  51554=>"000011001",
  51555=>"111111111",
  51556=>"100111001",
  51557=>"111001111",
  51558=>"111000000",
  51559=>"011000000",
  51560=>"110110110",
  51561=>"101111011",
  51562=>"111111111",
  51563=>"111111110",
  51564=>"000000100",
  51565=>"000011101",
  51566=>"110111111",
  51567=>"000000111",
  51568=>"000010010",
  51569=>"110111111",
  51570=>"000000000",
  51571=>"111111010",
  51572=>"000111101",
  51573=>"000001011",
  51574=>"011110111",
  51575=>"100000000",
  51576=>"111111100",
  51577=>"111111110",
  51578=>"001001101",
  51579=>"000000001",
  51580=>"111111111",
  51581=>"111111110",
  51582=>"000000001",
  51583=>"111111111",
  51584=>"110110110",
  51585=>"000000000",
  51586=>"111001000",
  51587=>"000000011",
  51588=>"000000000",
  51589=>"101100101",
  51590=>"111011010",
  51591=>"101000000",
  51592=>"001001000",
  51593=>"000000001",
  51594=>"000001111",
  51595=>"000111100",
  51596=>"111111111",
  51597=>"000111000",
  51598=>"110110110",
  51599=>"100101111",
  51600=>"000000000",
  51601=>"001000110",
  51602=>"111101000",
  51603=>"111110110",
  51604=>"111111111",
  51605=>"000111111",
  51606=>"111011111",
  51607=>"110100000",
  51608=>"000000000",
  51609=>"011111111",
  51610=>"111111111",
  51611=>"000000111",
  51612=>"111111111",
  51613=>"000000000",
  51614=>"100000000",
  51615=>"000011111",
  51616=>"000000111",
  51617=>"000100011",
  51618=>"111111111",
  51619=>"000000001",
  51620=>"110111000",
  51621=>"000000000",
  51622=>"000000000",
  51623=>"010000000",
  51624=>"000011000",
  51625=>"011111111",
  51626=>"001011011",
  51627=>"111000000",
  51628=>"000000000",
  51629=>"111001111",
  51630=>"111111111",
  51631=>"010011111",
  51632=>"111111111",
  51633=>"111110010",
  51634=>"111000000",
  51635=>"011000111",
  51636=>"111011000",
  51637=>"000000000",
  51638=>"010011001",
  51639=>"000001001",
  51640=>"111000000",
  51641=>"011111111",
  51642=>"111111111",
  51643=>"101000000",
  51644=>"000111000",
  51645=>"011001000",
  51646=>"100101011",
  51647=>"100100000",
  51648=>"111111101",
  51649=>"001111001",
  51650=>"000001001",
  51651=>"111111111",
  51652=>"111000000",
  51653=>"111000000",
  51654=>"111111000",
  51655=>"100000100",
  51656=>"000100010",
  51657=>"000000010",
  51658=>"000000000",
  51659=>"000110111",
  51660=>"000000000",
  51661=>"000000000",
  51662=>"011011000",
  51663=>"111111111",
  51664=>"111111011",
  51665=>"011011000",
  51666=>"000000010",
  51667=>"111111010",
  51668=>"000000000",
  51669=>"000000000",
  51670=>"011111111",
  51671=>"000001000",
  51672=>"111111111",
  51673=>"111111000",
  51674=>"000000000",
  51675=>"000010111",
  51676=>"000000000",
  51677=>"111111000",
  51678=>"010010000",
  51679=>"001000110",
  51680=>"001111111",
  51681=>"000100111",
  51682=>"000100001",
  51683=>"000111111",
  51684=>"010110010",
  51685=>"101000000",
  51686=>"000000111",
  51687=>"111111111",
  51688=>"101001111",
  51689=>"011111111",
  51690=>"000011111",
  51691=>"001011000",
  51692=>"010110111",
  51693=>"011011001",
  51694=>"000000111",
  51695=>"000111111",
  51696=>"111100000",
  51697=>"111111111",
  51698=>"111011011",
  51699=>"000111110",
  51700=>"011000000",
  51701=>"111111111",
  51702=>"100111111",
  51703=>"000001111",
  51704=>"000000000",
  51705=>"001001000",
  51706=>"111111110",
  51707=>"111000000",
  51708=>"000010010",
  51709=>"000111111",
  51710=>"111001000",
  51711=>"111101000",
  51712=>"110100000",
  51713=>"000000001",
  51714=>"111000111",
  51715=>"111111111",
  51716=>"110000000",
  51717=>"001001011",
  51718=>"111111000",
  51719=>"000000000",
  51720=>"000000000",
  51721=>"000000100",
  51722=>"100000000",
  51723=>"001000000",
  51724=>"110111111",
  51725=>"111111111",
  51726=>"000000000",
  51727=>"111000000",
  51728=>"111001000",
  51729=>"110110111",
  51730=>"011011000",
  51731=>"111111110",
  51732=>"000000111",
  51733=>"110110111",
  51734=>"111111111",
  51735=>"110100100",
  51736=>"111000000",
  51737=>"100111100",
  51738=>"000000001",
  51739=>"111101100",
  51740=>"111111111",
  51741=>"000000000",
  51742=>"111011111",
  51743=>"111111110",
  51744=>"011111111",
  51745=>"000000010",
  51746=>"000001000",
  51747=>"111111111",
  51748=>"100000000",
  51749=>"000111111",
  51750=>"010000001",
  51751=>"111000000",
  51752=>"000000011",
  51753=>"000000000",
  51754=>"000000000",
  51755=>"111111111",
  51756=>"000000011",
  51757=>"000000101",
  51758=>"010010000",
  51759=>"111111111",
  51760=>"000000111",
  51761=>"000000000",
  51762=>"001001111",
  51763=>"000000111",
  51764=>"111111000",
  51765=>"111110000",
  51766=>"111111111",
  51767=>"001100101",
  51768=>"000000000",
  51769=>"000000011",
  51770=>"000110111",
  51771=>"011111111",
  51772=>"001000001",
  51773=>"110100100",
  51774=>"111111111",
  51775=>"000000000",
  51776=>"110111111",
  51777=>"000000100",
  51778=>"000000000",
  51779=>"000000111",
  51780=>"110000000",
  51781=>"111110100",
  51782=>"000000111",
  51783=>"111111111",
  51784=>"111111111",
  51785=>"001111111",
  51786=>"111110110",
  51787=>"000000000",
  51788=>"000111111",
  51789=>"111111100",
  51790=>"100100110",
  51791=>"001001011",
  51792=>"000000000",
  51793=>"010010011",
  51794=>"111001011",
  51795=>"110000000",
  51796=>"000000000",
  51797=>"000000000",
  51798=>"000000000",
  51799=>"101111111",
  51800=>"111001000",
  51801=>"111001001",
  51802=>"110000110",
  51803=>"110111011",
  51804=>"111111111",
  51805=>"101000111",
  51806=>"000000000",
  51807=>"000011111",
  51808=>"000111111",
  51809=>"011111111",
  51810=>"111111111",
  51811=>"000000000",
  51812=>"000000000",
  51813=>"010011011",
  51814=>"000111111",
  51815=>"000000000",
  51816=>"111111111",
  51817=>"111111111",
  51818=>"000000000",
  51819=>"111111110",
  51820=>"111111100",
  51821=>"000000010",
  51822=>"000100111",
  51823=>"111111100",
  51824=>"111110000",
  51825=>"000000110",
  51826=>"111111011",
  51827=>"111111100",
  51828=>"111111000",
  51829=>"100111000",
  51830=>"100100110",
  51831=>"000000000",
  51832=>"001011111",
  51833=>"000010000",
  51834=>"000000000",
  51835=>"100111111",
  51836=>"111111000",
  51837=>"000000000",
  51838=>"100000000",
  51839=>"110110000",
  51840=>"111111111",
  51841=>"111111111",
  51842=>"100000000",
  51843=>"000001001",
  51844=>"001001111",
  51845=>"111100100",
  51846=>"100011111",
  51847=>"111111111",
  51848=>"111101001",
  51849=>"111111111",
  51850=>"011010000",
  51851=>"111000000",
  51852=>"001111111",
  51853=>"000000001",
  51854=>"011000111",
  51855=>"111111111",
  51856=>"101101111",
  51857=>"100000000",
  51858=>"000000001",
  51859=>"000110110",
  51860=>"000000000",
  51861=>"111000011",
  51862=>"000111111",
  51863=>"000000011",
  51864=>"111101111",
  51865=>"111111111",
  51866=>"000000000",
  51867=>"111111000",
  51868=>"110100000",
  51869=>"111111011",
  51870=>"111000000",
  51871=>"000000000",
  51872=>"110110000",
  51873=>"000001111",
  51874=>"010011000",
  51875=>"111111111",
  51876=>"000011111",
  51877=>"111111111",
  51878=>"111100101",
  51879=>"011011000",
  51880=>"111111111",
  51881=>"000000000",
  51882=>"000000000",
  51883=>"000011111",
  51884=>"000000101",
  51885=>"100000000",
  51886=>"001001000",
  51887=>"001101000",
  51888=>"011011111",
  51889=>"010111011",
  51890=>"111010011",
  51891=>"000000000",
  51892=>"111010000",
  51893=>"000000000",
  51894=>"000111100",
  51895=>"110111111",
  51896=>"000000000",
  51897=>"000011000",
  51898=>"111000000",
  51899=>"111000110",
  51900=>"000000010",
  51901=>"111110000",
  51902=>"111010000",
  51903=>"000000000",
  51904=>"111111000",
  51905=>"000000000",
  51906=>"001000000",
  51907=>"000000010",
  51908=>"001111111",
  51909=>"000000111",
  51910=>"011000000",
  51911=>"111001001",
  51912=>"111000000",
  51913=>"011111111",
  51914=>"111101011",
  51915=>"100000000",
  51916=>"000111111",
  51917=>"100000000",
  51918=>"111010000",
  51919=>"100110111",
  51920=>"111111110",
  51921=>"111111111",
  51922=>"000000100",
  51923=>"100100100",
  51924=>"000000000",
  51925=>"000000000",
  51926=>"000111111",
  51927=>"111111111",
  51928=>"000011111",
  51929=>"000000011",
  51930=>"111000100",
  51931=>"000000000",
  51932=>"101111111",
  51933=>"000000000",
  51934=>"000111111",
  51935=>"000000000",
  51936=>"111001000",
  51937=>"010111111",
  51938=>"010111111",
  51939=>"011110010",
  51940=>"111111000",
  51941=>"111111111",
  51942=>"110011000",
  51943=>"111111110",
  51944=>"000111000",
  51945=>"111100010",
  51946=>"111100000",
  51947=>"000000000",
  51948=>"111000000",
  51949=>"000000111",
  51950=>"111010100",
  51951=>"100001011",
  51952=>"100111000",
  51953=>"000000000",
  51954=>"111111111",
  51955=>"111000000",
  51956=>"111111111",
  51957=>"000011111",
  51958=>"011000000",
  51959=>"100111111",
  51960=>"010111111",
  51961=>"001111111",
  51962=>"000000000",
  51963=>"111001101",
  51964=>"111111011",
  51965=>"111111011",
  51966=>"111110111",
  51967=>"100000000",
  51968=>"000000000",
  51969=>"001001001",
  51970=>"000000111",
  51971=>"111111110",
  51972=>"111111111",
  51973=>"100000100",
  51974=>"111111111",
  51975=>"000100111",
  51976=>"000000001",
  51977=>"111111010",
  51978=>"011000100",
  51979=>"111111100",
  51980=>"001001101",
  51981=>"111111100",
  51982=>"000000000",
  51983=>"000000111",
  51984=>"001101111",
  51985=>"000111111",
  51986=>"111111111",
  51987=>"000000000",
  51988=>"110111111",
  51989=>"000111111",
  51990=>"011011000",
  51991=>"000000001",
  51992=>"000000000",
  51993=>"111000110",
  51994=>"111011000",
  51995=>"111100100",
  51996=>"110110011",
  51997=>"010000000",
  51998=>"000000100",
  51999=>"100000111",
  52000=>"000010011",
  52001=>"000000111",
  52002=>"110100000",
  52003=>"111111111",
  52004=>"001001001",
  52005=>"111100100",
  52006=>"111111111",
  52007=>"000100111",
  52008=>"111110111",
  52009=>"110100000",
  52010=>"001000101",
  52011=>"101110100",
  52012=>"000100010",
  52013=>"111111011",
  52014=>"110010010",
  52015=>"000000000",
  52016=>"110000011",
  52017=>"111000000",
  52018=>"000000000",
  52019=>"111110100",
  52020=>"110000000",
  52021=>"010000000",
  52022=>"111000000",
  52023=>"000111111",
  52024=>"000000000",
  52025=>"000000001",
  52026=>"101000000",
  52027=>"000000111",
  52028=>"010111111",
  52029=>"011000000",
  52030=>"001000001",
  52031=>"000001111",
  52032=>"000000010",
  52033=>"000000011",
  52034=>"010111010",
  52035=>"111011000",
  52036=>"000011000",
  52037=>"000000000",
  52038=>"111111010",
  52039=>"001000000",
  52040=>"001000011",
  52041=>"000000111",
  52042=>"000000100",
  52043=>"100001101",
  52044=>"111111111",
  52045=>"111111001",
  52046=>"011111111",
  52047=>"001001000",
  52048=>"111111111",
  52049=>"000000111",
  52050=>"000000001",
  52051=>"111111111",
  52052=>"000000111",
  52053=>"011000000",
  52054=>"111111111",
  52055=>"000001111",
  52056=>"011100001",
  52057=>"001001101",
  52058=>"000000000",
  52059=>"111011110",
  52060=>"111111111",
  52061=>"111100101",
  52062=>"011000100",
  52063=>"111111000",
  52064=>"111111000",
  52065=>"000000000",
  52066=>"000000111",
  52067=>"101111111",
  52068=>"110111000",
  52069=>"100000000",
  52070=>"010110111",
  52071=>"000000000",
  52072=>"011011011",
  52073=>"111011111",
  52074=>"111111000",
  52075=>"011111111",
  52076=>"111111010",
  52077=>"100100100",
  52078=>"111001000",
  52079=>"011000000",
  52080=>"000000111",
  52081=>"111000000",
  52082=>"001111011",
  52083=>"111111000",
  52084=>"110000000",
  52085=>"000000000",
  52086=>"111111110",
  52087=>"010000000",
  52088=>"111001001",
  52089=>"000111111",
  52090=>"111111111",
  52091=>"000000000",
  52092=>"000101111",
  52093=>"000000000",
  52094=>"001010110",
  52095=>"111111111",
  52096=>"000000000",
  52097=>"111111111",
  52098=>"011001001",
  52099=>"111000000",
  52100=>"000010111",
  52101=>"000000000",
  52102=>"111111111",
  52103=>"000000001",
  52104=>"110100100",
  52105=>"100110111",
  52106=>"001000101",
  52107=>"000000111",
  52108=>"111101101",
  52109=>"001011011",
  52110=>"010011000",
  52111=>"010000100",
  52112=>"000000111",
  52113=>"111000000",
  52114=>"000000111",
  52115=>"000100111",
  52116=>"111101111",
  52117=>"000000000",
  52118=>"001001001",
  52119=>"000000111",
  52120=>"000010110",
  52121=>"110001011",
  52122=>"111111000",
  52123=>"000000000",
  52124=>"000000111",
  52125=>"111111111",
  52126=>"000000000",
  52127=>"011111111",
  52128=>"010000000",
  52129=>"111011010",
  52130=>"001000001",
  52131=>"110000100",
  52132=>"111111110",
  52133=>"111010111",
  52134=>"001000000",
  52135=>"000011111",
  52136=>"000000000",
  52137=>"011011111",
  52138=>"111111111",
  52139=>"001000000",
  52140=>"000000000",
  52141=>"111111110",
  52142=>"000000000",
  52143=>"100101101",
  52144=>"000000000",
  52145=>"000010000",
  52146=>"000000001",
  52147=>"111100000",
  52148=>"111000000",
  52149=>"001000001",
  52150=>"001000011",
  52151=>"110110000",
  52152=>"111100110",
  52153=>"011001111",
  52154=>"110000000",
  52155=>"111111111",
  52156=>"111111001",
  52157=>"111011000",
  52158=>"010111111",
  52159=>"001111001",
  52160=>"000010011",
  52161=>"100111111",
  52162=>"000000000",
  52163=>"111111111",
  52164=>"111111000",
  52165=>"111101111",
  52166=>"111111111",
  52167=>"111111101",
  52168=>"001000000",
  52169=>"000000100",
  52170=>"000000101",
  52171=>"011000000",
  52172=>"000000000",
  52173=>"001011011",
  52174=>"111000001",
  52175=>"000000000",
  52176=>"000000111",
  52177=>"111110011",
  52178=>"111111011",
  52179=>"111110000",
  52180=>"101101011",
  52181=>"111110000",
  52182=>"000000101",
  52183=>"011111111",
  52184=>"101000000",
  52185=>"000100111",
  52186=>"001001111",
  52187=>"111111110",
  52188=>"000000111",
  52189=>"001101101",
  52190=>"001000001",
  52191=>"110100000",
  52192=>"001000000",
  52193=>"000000000",
  52194=>"100111000",
  52195=>"000000000",
  52196=>"111111111",
  52197=>"000000000",
  52198=>"101000000",
  52199=>"000000111",
  52200=>"000000000",
  52201=>"110111000",
  52202=>"110000000",
  52203=>"011111001",
  52204=>"111111000",
  52205=>"000000111",
  52206=>"000000000",
  52207=>"111000000",
  52208=>"000000000",
  52209=>"111000001",
  52210=>"011111111",
  52211=>"000000000",
  52212=>"111111111",
  52213=>"000000000",
  52214=>"111111111",
  52215=>"000000000",
  52216=>"111000000",
  52217=>"101101111",
  52218=>"000000000",
  52219=>"111111111",
  52220=>"111000111",
  52221=>"000111111",
  52222=>"000111110",
  52223=>"111111111",
  52224=>"000011111",
  52225=>"011010010",
  52226=>"111111111",
  52227=>"011000000",
  52228=>"111111011",
  52229=>"000000000",
  52230=>"000101111",
  52231=>"111111111",
  52232=>"001111111",
  52233=>"001000000",
  52234=>"111111111",
  52235=>"111111111",
  52236=>"100100100",
  52237=>"001011111",
  52238=>"111111111",
  52239=>"000000000",
  52240=>"010110011",
  52241=>"111111111",
  52242=>"000111111",
  52243=>"110000000",
  52244=>"000111110",
  52245=>"000000111",
  52246=>"000000001",
  52247=>"000001111",
  52248=>"100011111",
  52249=>"010111000",
  52250=>"101000000",
  52251=>"000000000",
  52252=>"000101111",
  52253=>"111111111",
  52254=>"100001001",
  52255=>"010111111",
  52256=>"111111111",
  52257=>"110000000",
  52258=>"100100110",
  52259=>"110000000",
  52260=>"111111111",
  52261=>"101000000",
  52262=>"111110111",
  52263=>"100000000",
  52264=>"101101111",
  52265=>"000000100",
  52266=>"001000000",
  52267=>"001101000",
  52268=>"000001111",
  52269=>"000000000",
  52270=>"000000001",
  52271=>"111111111",
  52272=>"000000000",
  52273=>"111111111",
  52274=>"011111011",
  52275=>"000100100",
  52276=>"000000000",
  52277=>"000001100",
  52278=>"000111111",
  52279=>"001010100",
  52280=>"111111111",
  52281=>"000000000",
  52282=>"000000000",
  52283=>"001000000",
  52284=>"101101101",
  52285=>"000000000",
  52286=>"000000100",
  52287=>"000000000",
  52288=>"001001000",
  52289=>"000000000",
  52290=>"101101000",
  52291=>"000100111",
  52292=>"111111111",
  52293=>"001000011",
  52294=>"000000111",
  52295=>"000000000",
  52296=>"000001001",
  52297=>"001000000",
  52298=>"111111111",
  52299=>"111111111",
  52300=>"100100100",
  52301=>"000111110",
  52302=>"000000000",
  52303=>"001001111",
  52304=>"000000000",
  52305=>"111111111",
  52306=>"100111000",
  52307=>"011111111",
  52308=>"000000000",
  52309=>"000000001",
  52310=>"100101110",
  52311=>"111111111",
  52312=>"111111111",
  52313=>"000000000",
  52314=>"111111111",
  52315=>"000101101",
  52316=>"111101110",
  52317=>"110000001",
  52318=>"111111000",
  52319=>"000000110",
  52320=>"100000000",
  52321=>"001001001",
  52322=>"000000000",
  52323=>"111111111",
  52324=>"111010000",
  52325=>"101001000",
  52326=>"000000001",
  52327=>"000000101",
  52328=>"100000100",
  52329=>"111111111",
  52330=>"000100110",
  52331=>"111001111",
  52332=>"010111111",
  52333=>"000111100",
  52334=>"111110111",
  52335=>"110110111",
  52336=>"111101000",
  52337=>"000001000",
  52338=>"000001001",
  52339=>"111111001",
  52340=>"000000000",
  52341=>"000100111",
  52342=>"111111111",
  52343=>"111000000",
  52344=>"000000000",
  52345=>"111111001",
  52346=>"000000000",
  52347=>"001101111",
  52348=>"000000000",
  52349=>"000000000",
  52350=>"111111100",
  52351=>"000000000",
  52352=>"111000000",
  52353=>"111111001",
  52354=>"000000000",
  52355=>"111111001",
  52356=>"011111111",
  52357=>"000000000",
  52358=>"100000000",
  52359=>"011000000",
  52360=>"001110111",
  52361=>"010000000",
  52362=>"000000000",
  52363=>"111111111",
  52364=>"111101101",
  52365=>"000110010",
  52366=>"001001000",
  52367=>"000000000",
  52368=>"000001111",
  52369=>"111111111",
  52370=>"001111111",
  52371=>"000000000",
  52372=>"000011010",
  52373=>"111111111",
  52374=>"101111000",
  52375=>"111000111",
  52376=>"000000000",
  52377=>"000000000",
  52378=>"111111110",
  52379=>"111111011",
  52380=>"100100111",
  52381=>"110111000",
  52382=>"111111011",
  52383=>"111100000",
  52384=>"000000000",
  52385=>"110000001",
  52386=>"000000110",
  52387=>"000000000",
  52388=>"001000100",
  52389=>"000000011",
  52390=>"010111111",
  52391=>"110110000",
  52392=>"011011000",
  52393=>"000000000",
  52394=>"111111111",
  52395=>"110000001",
  52396=>"000111111",
  52397=>"100111111",
  52398=>"111111111",
  52399=>"111111111",
  52400=>"000000010",
  52401=>"000000000",
  52402=>"111111111",
  52403=>"111111000",
  52404=>"111111111",
  52405=>"111111000",
  52406=>"000000000",
  52407=>"111111111",
  52408=>"000000000",
  52409=>"000000000",
  52410=>"001000111",
  52411=>"111100111",
  52412=>"001000100",
  52413=>"111111111",
  52414=>"101111111",
  52415=>"110001001",
  52416=>"000111111",
  52417=>"000000000",
  52418=>"111101100",
  52419=>"000000000",
  52420=>"000000000",
  52421=>"000000000",
  52422=>"111110110",
  52423=>"111111111",
  52424=>"111011000",
  52425=>"000000111",
  52426=>"000000000",
  52427=>"111111111",
  52428=>"100111100",
  52429=>"000100111",
  52430=>"110000000",
  52431=>"110111111",
  52432=>"001000111",
  52433=>"000000011",
  52434=>"111110111",
  52435=>"000000000",
  52436=>"110111101",
  52437=>"011101111",
  52438=>"111000000",
  52439=>"011011100",
  52440=>"000101111",
  52441=>"101111000",
  52442=>"000000000",
  52443=>"001111111",
  52444=>"000111111",
  52445=>"000001001",
  52446=>"000011111",
  52447=>"111111010",
  52448=>"111111111",
  52449=>"000000010",
  52450=>"000000000",
  52451=>"100110000",
  52452=>"010111111",
  52453=>"111111010",
  52454=>"000111111",
  52455=>"111111111",
  52456=>"000000100",
  52457=>"000000111",
  52458=>"100000000",
  52459=>"001000000",
  52460=>"101000000",
  52461=>"110000000",
  52462=>"100110111",
  52463=>"000000000",
  52464=>"110111010",
  52465=>"000001111",
  52466=>"111001111",
  52467=>"101001111",
  52468=>"111111111",
  52469=>"100011101",
  52470=>"111111111",
  52471=>"000000100",
  52472=>"101001111",
  52473=>"111111001",
  52474=>"000000000",
  52475=>"000000000",
  52476=>"011001001",
  52477=>"010000100",
  52478=>"000000000",
  52479=>"011000000",
  52480=>"001111111",
  52481=>"110110110",
  52482=>"111110000",
  52483=>"111111001",
  52484=>"000101000",
  52485=>"000001011",
  52486=>"000100100",
  52487=>"001111100",
  52488=>"000000000",
  52489=>"001000000",
  52490=>"001111111",
  52491=>"111111110",
  52492=>"111111111",
  52493=>"000010111",
  52494=>"000000111",
  52495=>"111000000",
  52496=>"111111111",
  52497=>"100100111",
  52498=>"000000000",
  52499=>"000010000",
  52500=>"111100000",
  52501=>"001111111",
  52502=>"000100111",
  52503=>"000111111",
  52504=>"010000010",
  52505=>"111111100",
  52506=>"111000000",
  52507=>"111111111",
  52508=>"111110100",
  52509=>"100100000",
  52510=>"111111111",
  52511=>"111111111",
  52512=>"100001011",
  52513=>"000000000",
  52514=>"110000111",
  52515=>"000000100",
  52516=>"000000000",
  52517=>"011000000",
  52518=>"101100111",
  52519=>"000000000",
  52520=>"000100111",
  52521=>"000000000",
  52522=>"111000000",
  52523=>"010000001",
  52524=>"111001000",
  52525=>"111111111",
  52526=>"000000111",
  52527=>"011010010",
  52528=>"001000010",
  52529=>"111111100",
  52530=>"011110000",
  52531=>"000000000",
  52532=>"000000000",
  52533=>"001000000",
  52534=>"111111001",
  52535=>"111000111",
  52536=>"010010000",
  52537=>"111000000",
  52538=>"000000110",
  52539=>"111111000",
  52540=>"000000110",
  52541=>"000000000",
  52542=>"011000100",
  52543=>"111111011",
  52544=>"010000000",
  52545=>"000000110",
  52546=>"100000000",
  52547=>"001000000",
  52548=>"100011000",
  52549=>"101111111",
  52550=>"000000000",
  52551=>"100100100",
  52552=>"111111111",
  52553=>"111111110",
  52554=>"110111111",
  52555=>"000000011",
  52556=>"000100001",
  52557=>"111000000",
  52558=>"001000000",
  52559=>"111111101",
  52560=>"000111111",
  52561=>"000000111",
  52562=>"010111111",
  52563=>"000000111",
  52564=>"000110111",
  52565=>"011011001",
  52566=>"000000011",
  52567=>"000000000",
  52568=>"111111100",
  52569=>"111111111",
  52570=>"111111011",
  52571=>"111111111",
  52572=>"000000000",
  52573=>"000000110",
  52574=>"111101000",
  52575=>"000010011",
  52576=>"111110100",
  52577=>"011111111",
  52578=>"000100000",
  52579=>"111111111",
  52580=>"000100101",
  52581=>"111001001",
  52582=>"000111000",
  52583=>"001001010",
  52584=>"000000000",
  52585=>"000100101",
  52586=>"110000100",
  52587=>"000001000",
  52588=>"011011010",
  52589=>"000000111",
  52590=>"001000000",
  52591=>"110110001",
  52592=>"111111111",
  52593=>"111111111",
  52594=>"001001001",
  52595=>"110110111",
  52596=>"100111110",
  52597=>"111111111",
  52598=>"110111111",
  52599=>"001000110",
  52600=>"111000000",
  52601=>"000100111",
  52602=>"111010000",
  52603=>"001000000",
  52604=>"111111000",
  52605=>"000000010",
  52606=>"101101111",
  52607=>"100111101",
  52608=>"001011011",
  52609=>"111111111",
  52610=>"000000001",
  52611=>"111111111",
  52612=>"000000000",
  52613=>"000000000",
  52614=>"111110110",
  52615=>"000000000",
  52616=>"111000000",
  52617=>"000000011",
  52618=>"111111011",
  52619=>"010000010",
  52620=>"101111111",
  52621=>"100100101",
  52622=>"001011100",
  52623=>"000111111",
  52624=>"111111001",
  52625=>"000000110",
  52626=>"110110110",
  52627=>"000000011",
  52628=>"111111111",
  52629=>"000000000",
  52630=>"111000111",
  52631=>"110010000",
  52632=>"111111111",
  52633=>"000000011",
  52634=>"111111010",
  52635=>"110010000",
  52636=>"000000010",
  52637=>"001001100",
  52638=>"111111111",
  52639=>"111111100",
  52640=>"111111111",
  52641=>"011000000",
  52642=>"000001000",
  52643=>"111111000",
  52644=>"000001111",
  52645=>"000000000",
  52646=>"000000010",
  52647=>"000000000",
  52648=>"111100011",
  52649=>"101110000",
  52650=>"100100100",
  52651=>"111111111",
  52652=>"010000100",
  52653=>"000000000",
  52654=>"000000000",
  52655=>"110111111",
  52656=>"100111111",
  52657=>"111111111",
  52658=>"100100000",
  52659=>"000111111",
  52660=>"000000111",
  52661=>"100100111",
  52662=>"101111111",
  52663=>"000010011",
  52664=>"001011000",
  52665=>"111111111",
  52666=>"111111010",
  52667=>"000000000",
  52668=>"000000000",
  52669=>"111111000",
  52670=>"010000010",
  52671=>"000000000",
  52672=>"111000000",
  52673=>"000000001",
  52674=>"000000000",
  52675=>"100100000",
  52676=>"110100000",
  52677=>"100111001",
  52678=>"111000000",
  52679=>"011000000",
  52680=>"000111111",
  52681=>"000111111",
  52682=>"001000000",
  52683=>"100000101",
  52684=>"000000111",
  52685=>"111111000",
  52686=>"101111111",
  52687=>"000001000",
  52688=>"000000000",
  52689=>"110000000",
  52690=>"000111111",
  52691=>"111111111",
  52692=>"111111111",
  52693=>"111111111",
  52694=>"111111111",
  52695=>"110000001",
  52696=>"111111110",
  52697=>"000000000",
  52698=>"111000011",
  52699=>"000100101",
  52700=>"000000111",
  52701=>"000000000",
  52702=>"100000111",
  52703=>"111111110",
  52704=>"110110111",
  52705=>"001001000",
  52706=>"111111100",
  52707=>"111111110",
  52708=>"011001011",
  52709=>"011011111",
  52710=>"111111011",
  52711=>"111100000",
  52712=>"111010010",
  52713=>"100100101",
  52714=>"000000000",
  52715=>"000000000",
  52716=>"100000000",
  52717=>"010110110",
  52718=>"111111111",
  52719=>"111111111",
  52720=>"000000000",
  52721=>"000100101",
  52722=>"001000000",
  52723=>"000000000",
  52724=>"000100000",
  52725=>"000000000",
  52726=>"111110100",
  52727=>"111011111",
  52728=>"001111001",
  52729=>"000001001",
  52730=>"101101100",
  52731=>"111111111",
  52732=>"000000111",
  52733=>"000000011",
  52734=>"000001000",
  52735=>"111111111",
  52736=>"000100100",
  52737=>"000110000",
  52738=>"100000000",
  52739=>"000000000",
  52740=>"111001000",
  52741=>"110000000",
  52742=>"000011111",
  52743=>"111111111",
  52744=>"111111010",
  52745=>"111010000",
  52746=>"001001001",
  52747=>"000000001",
  52748=>"110100001",
  52749=>"100000000",
  52750=>"011000100",
  52751=>"000000000",
  52752=>"111000100",
  52753=>"000000000",
  52754=>"111111111",
  52755=>"000000000",
  52756=>"000000111",
  52757=>"000000100",
  52758=>"011001000",
  52759=>"111001111",
  52760=>"000100000",
  52761=>"001001000",
  52762=>"100000000",
  52763=>"000001000",
  52764=>"111111001",
  52765=>"110000111",
  52766=>"111111000",
  52767=>"000011111",
  52768=>"110111111",
  52769=>"000000000",
  52770=>"111111111",
  52771=>"111100000",
  52772=>"101101101",
  52773=>"000001000",
  52774=>"110000000",
  52775=>"000001000",
  52776=>"111111011",
  52777=>"100100111",
  52778=>"001011111",
  52779=>"111101001",
  52780=>"111111111",
  52781=>"000000000",
  52782=>"011010011",
  52783=>"000000011",
  52784=>"000111100",
  52785=>"111111111",
  52786=>"001111111",
  52787=>"010100000",
  52788=>"000000000",
  52789=>"111010010",
  52790=>"111111001",
  52791=>"001000000",
  52792=>"111101000",
  52793=>"000000110",
  52794=>"001011011",
  52795=>"111111111",
  52796=>"100000000",
  52797=>"111110111",
  52798=>"111110110",
  52799=>"000000000",
  52800=>"110111111",
  52801=>"001001000",
  52802=>"110000000",
  52803=>"000100100",
  52804=>"111111111",
  52805=>"111111001",
  52806=>"000001111",
  52807=>"111111111",
  52808=>"011100000",
  52809=>"000000111",
  52810=>"011001101",
  52811=>"011111111",
  52812=>"000101111",
  52813=>"000100100",
  52814=>"111111010",
  52815=>"110110000",
  52816=>"000010111",
  52817=>"000100000",
  52818=>"111111011",
  52819=>"001001001",
  52820=>"011011110",
  52821=>"111111111",
  52822=>"111100000",
  52823=>"111111111",
  52824=>"111111111",
  52825=>"000000111",
  52826=>"000000111",
  52827=>"111111110",
  52828=>"011111101",
  52829=>"000000000",
  52830=>"111111111",
  52831=>"100100000",
  52832=>"111111111",
  52833=>"011000000",
  52834=>"001111011",
  52835=>"000000000",
  52836=>"101000111",
  52837=>"011111111",
  52838=>"000100000",
  52839=>"111011001",
  52840=>"110111111",
  52841=>"111111111",
  52842=>"010111111",
  52843=>"000010010",
  52844=>"101001001",
  52845=>"000000000",
  52846=>"001101001",
  52847=>"000000011",
  52848=>"000000010",
  52849=>"000000000",
  52850=>"110110100",
  52851=>"000110111",
  52852=>"001001111",
  52853=>"001001000",
  52854=>"000000000",
  52855=>"011101111",
  52856=>"111111111",
  52857=>"001000000",
  52858=>"000000111",
  52859=>"111111111",
  52860=>"100110111",
  52861=>"110111001",
  52862=>"000000101",
  52863=>"111111111",
  52864=>"000000111",
  52865=>"010000100",
  52866=>"111111111",
  52867=>"000000000",
  52868=>"000000000",
  52869=>"111111111",
  52870=>"000000000",
  52871=>"001001001",
  52872=>"111000000",
  52873=>"111110100",
  52874=>"011111111",
  52875=>"000100000",
  52876=>"000100101",
  52877=>"001000001",
  52878=>"111000000",
  52879=>"000000000",
  52880=>"100000000",
  52881=>"111111111",
  52882=>"101110110",
  52883=>"011010010",
  52884=>"110111111",
  52885=>"011111000",
  52886=>"100000000",
  52887=>"000000000",
  52888=>"000001001",
  52889=>"000000111",
  52890=>"000111111",
  52891=>"000001111",
  52892=>"111111111",
  52893=>"111111001",
  52894=>"110110001",
  52895=>"000001001",
  52896=>"111010111",
  52897=>"011101000",
  52898=>"111001000",
  52899=>"000011011",
  52900=>"011000010",
  52901=>"110111111",
  52902=>"111111111",
  52903=>"111110100",
  52904=>"000001000",
  52905=>"111111111",
  52906=>"010000000",
  52907=>"111111010",
  52908=>"000000001",
  52909=>"000110000",
  52910=>"111000111",
  52911=>"000100111",
  52912=>"000100111",
  52913=>"000100100",
  52914=>"010111111",
  52915=>"000001111",
  52916=>"110110000",
  52917=>"110111111",
  52918=>"000000000",
  52919=>"000000000",
  52920=>"111111011",
  52921=>"001000000",
  52922=>"001000000",
  52923=>"000000000",
  52924=>"010111110",
  52925=>"000000000",
  52926=>"111000000",
  52927=>"000001001",
  52928=>"000000000",
  52929=>"111001001",
  52930=>"100000000",
  52931=>"111001101",
  52932=>"100001001",
  52933=>"000000001",
  52934=>"000000111",
  52935=>"000001101",
  52936=>"100100110",
  52937=>"000001000",
  52938=>"000010011",
  52939=>"000100111",
  52940=>"000000000",
  52941=>"111111110",
  52942=>"010010100",
  52943=>"011110100",
  52944=>"110100010",
  52945=>"000000000",
  52946=>"100100110",
  52947=>"000001011",
  52948=>"100100001",
  52949=>"111011011",
  52950=>"110100000",
  52951=>"111101001",
  52952=>"100000000",
  52953=>"111111111",
  52954=>"111111111",
  52955=>"111111111",
  52956=>"101001011",
  52957=>"111110110",
  52958=>"000000011",
  52959=>"000000111",
  52960=>"000000000",
  52961=>"110000010",
  52962=>"110000000",
  52963=>"111111111",
  52964=>"111000100",
  52965=>"110111011",
  52966=>"000000000",
  52967=>"111101111",
  52968=>"000000000",
  52969=>"000000001",
  52970=>"000000000",
  52971=>"000000010",
  52972=>"000000010",
  52973=>"100000000",
  52974=>"000000000",
  52975=>"111011000",
  52976=>"100111001",
  52977=>"011011111",
  52978=>"000110111",
  52979=>"000100000",
  52980=>"111111111",
  52981=>"000001000",
  52982=>"110111111",
  52983=>"100100110",
  52984=>"101000011",
  52985=>"011011111",
  52986=>"011001011",
  52987=>"000000101",
  52988=>"111011001",
  52989=>"110110110",
  52990=>"111111111",
  52991=>"000001111",
  52992=>"111111111",
  52993=>"111010000",
  52994=>"011010110",
  52995=>"000111111",
  52996=>"001001001",
  52997=>"100000000",
  52998=>"000001001",
  52999=>"000000000",
  53000=>"101101111",
  53001=>"000000111",
  53002=>"000000000",
  53003=>"100000000",
  53004=>"110110110",
  53005=>"000000111",
  53006=>"110110010",
  53007=>"000000000",
  53008=>"111100100",
  53009=>"111111111",
  53010=>"100100110",
  53011=>"011011000",
  53012=>"110111011",
  53013=>"000100001",
  53014=>"001001001",
  53015=>"000000000",
  53016=>"000001011",
  53017=>"000000000",
  53018=>"000000000",
  53019=>"110110111",
  53020=>"100000100",
  53021=>"000101001",
  53022=>"001001000",
  53023=>"110111111",
  53024=>"111101001",
  53025=>"000001111",
  53026=>"000110010",
  53027=>"000010001",
  53028=>"111111110",
  53029=>"000000000",
  53030=>"100000000",
  53031=>"010000000",
  53032=>"000000000",
  53033=>"111111111",
  53034=>"110111111",
  53035=>"000110111",
  53036=>"000110101",
  53037=>"111111111",
  53038=>"000111010",
  53039=>"110111111",
  53040=>"110001001",
  53041=>"011111111",
  53042=>"111111111",
  53043=>"111111011",
  53044=>"111111010",
  53045=>"111111111",
  53046=>"111000111",
  53047=>"001111111",
  53048=>"111100000",
  53049=>"000000000",
  53050=>"111111111",
  53051=>"000010010",
  53052=>"000000000",
  53053=>"001000001",
  53054=>"111111011",
  53055=>"000000111",
  53056=>"000100111",
  53057=>"100100110",
  53058=>"000000001",
  53059=>"000000000",
  53060=>"111111000",
  53061=>"111001000",
  53062=>"111111111",
  53063=>"000000000",
  53064=>"111110111",
  53065=>"000000000",
  53066=>"100100100",
  53067=>"110111101",
  53068=>"000000000",
  53069=>"100110000",
  53070=>"100101111",
  53071=>"111110000",
  53072=>"111111111",
  53073=>"000000100",
  53074=>"000000000",
  53075=>"011010110",
  53076=>"101000000",
  53077=>"011011111",
  53078=>"100000000",
  53079=>"000000000",
  53080=>"000100111",
  53081=>"100100001",
  53082=>"111111011",
  53083=>"000000110",
  53084=>"000000101",
  53085=>"011001001",
  53086=>"111111000",
  53087=>"111111110",
  53088=>"110000000",
  53089=>"111100110",
  53090=>"111101100",
  53091=>"000000100",
  53092=>"111011000",
  53093=>"111110100",
  53094=>"110000011",
  53095=>"111111111",
  53096=>"010110100",
  53097=>"100000000",
  53098=>"011001101",
  53099=>"000011101",
  53100=>"000001011",
  53101=>"000010100",
  53102=>"011011011",
  53103=>"001001001",
  53104=>"100100001",
  53105=>"111111111",
  53106=>"000000011",
  53107=>"111111111",
  53108=>"111111111",
  53109=>"100000000",
  53110=>"111101001",
  53111=>"000100111",
  53112=>"110111111",
  53113=>"111000000",
  53114=>"000000000",
  53115=>"111100000",
  53116=>"111111111",
  53117=>"000000000",
  53118=>"111000110",
  53119=>"111111011",
  53120=>"100001011",
  53121=>"000111101",
  53122=>"111000001",
  53123=>"011011011",
  53124=>"111100111",
  53125=>"111100000",
  53126=>"110110110",
  53127=>"100110000",
  53128=>"011110110",
  53129=>"000011111",
  53130=>"111111011",
  53131=>"000000110",
  53132=>"000000000",
  53133=>"000110000",
  53134=>"111110000",
  53135=>"111000111",
  53136=>"100000111",
  53137=>"111111111",
  53138=>"000100111",
  53139=>"000000000",
  53140=>"101110111",
  53141=>"110000000",
  53142=>"011011011",
  53143=>"111011000",
  53144=>"000001111",
  53145=>"010111111",
  53146=>"111111111",
  53147=>"100100000",
  53148=>"000000000",
  53149=>"111111011",
  53150=>"111100100",
  53151=>"111111111",
  53152=>"000000000",
  53153=>"011000110",
  53154=>"010011000",
  53155=>"111111000",
  53156=>"000110111",
  53157=>"111100000",
  53158=>"000101111",
  53159=>"000010011",
  53160=>"000000000",
  53161=>"110000100",
  53162=>"000000000",
  53163=>"110111111",
  53164=>"011001001",
  53165=>"111111011",
  53166=>"111111111",
  53167=>"111000000",
  53168=>"000100111",
  53169=>"111111111",
  53170=>"000000000",
  53171=>"000111111",
  53172=>"111110000",
  53173=>"110100110",
  53174=>"110000000",
  53175=>"100100000",
  53176=>"000000000",
  53177=>"000110000",
  53178=>"111111111",
  53179=>"000111111",
  53180=>"000000000",
  53181=>"001001111",
  53182=>"000000000",
  53183=>"011010000",
  53184=>"111111011",
  53185=>"000000000",
  53186=>"111111111",
  53187=>"111111111",
  53188=>"111111110",
  53189=>"000000001",
  53190=>"111111111",
  53191=>"100100000",
  53192=>"100100101",
  53193=>"000000000",
  53194=>"000000001",
  53195=>"000000000",
  53196=>"000001000",
  53197=>"111111111",
  53198=>"000000000",
  53199=>"110110111",
  53200=>"011000111",
  53201=>"000000000",
  53202=>"110110111",
  53203=>"111111010",
  53204=>"010010011",
  53205=>"000000000",
  53206=>"111101101",
  53207=>"011011010",
  53208=>"000000001",
  53209=>"110000110",
  53210=>"000000001",
  53211=>"100000011",
  53212=>"000000010",
  53213=>"000100100",
  53214=>"111111100",
  53215=>"010000010",
  53216=>"110111111",
  53217=>"000000000",
  53218=>"111111111",
  53219=>"111000000",
  53220=>"011010001",
  53221=>"111000111",
  53222=>"110111111",
  53223=>"110000000",
  53224=>"110100111",
  53225=>"101100100",
  53226=>"111011000",
  53227=>"000000000",
  53228=>"101101111",
  53229=>"000101101",
  53230=>"111111111",
  53231=>"111110000",
  53232=>"000000000",
  53233=>"011111111",
  53234=>"000111000",
  53235=>"000111111",
  53236=>"100110000",
  53237=>"011000000",
  53238=>"111111111",
  53239=>"000100110",
  53240=>"000100111",
  53241=>"100110110",
  53242=>"111111111",
  53243=>"111111100",
  53244=>"110111010",
  53245=>"000000111",
  53246=>"100111111",
  53247=>"000000000",
  53248=>"111111111",
  53249=>"001001000",
  53250=>"000000000",
  53251=>"001000000",
  53252=>"110110110",
  53253=>"101100000",
  53254=>"000001111",
  53255=>"000000000",
  53256=>"111100000",
  53257=>"000111111",
  53258=>"111111110",
  53259=>"010011000",
  53260=>"111111111",
  53261=>"111001000",
  53262=>"010011100",
  53263=>"001011001",
  53264=>"001000001",
  53265=>"011111110",
  53266=>"100100100",
  53267=>"111111111",
  53268=>"001111111",
  53269=>"010010010",
  53270=>"111111111",
  53271=>"011011010",
  53272=>"110010010",
  53273=>"110111111",
  53274=>"111111111",
  53275=>"011011011",
  53276=>"101111111",
  53277=>"011010000",
  53278=>"111111111",
  53279=>"111101111",
  53280=>"000000001",
  53281=>"111111111",
  53282=>"111000000",
  53283=>"000001110",
  53284=>"111111000",
  53285=>"000000010",
  53286=>"110110100",
  53287=>"100100000",
  53288=>"111111000",
  53289=>"000001011",
  53290=>"111111000",
  53291=>"111010001",
  53292=>"000011000",
  53293=>"000000000",
  53294=>"001001111",
  53295=>"111111011",
  53296=>"000000110",
  53297=>"000000111",
  53298=>"111101001",
  53299=>"111111111",
  53300=>"000000000",
  53301=>"001001101",
  53302=>"001000000",
  53303=>"110111111",
  53304=>"001001101",
  53305=>"000000000",
  53306=>"001000000",
  53307=>"011011000",
  53308=>"000000000",
  53309=>"111111111",
  53310=>"001011111",
  53311=>"111111011",
  53312=>"000000000",
  53313=>"100100101",
  53314=>"000000000",
  53315=>"001000111",
  53316=>"011000011",
  53317=>"111110001",
  53318=>"111111000",
  53319=>"111111000",
  53320=>"000000000",
  53321=>"000100000",
  53322=>"101111111",
  53323=>"111001001",
  53324=>"111111111",
  53325=>"000000000",
  53326=>"000011010",
  53327=>"000000001",
  53328=>"111111011",
  53329=>"000000000",
  53330=>"101000000",
  53331=>"110110000",
  53332=>"000001111",
  53333=>"111111111",
  53334=>"000011001",
  53335=>"110111111",
  53336=>"111110111",
  53337=>"000000000",
  53338=>"111111100",
  53339=>"011011111",
  53340=>"000000010",
  53341=>"111111111",
  53342=>"111111111",
  53343=>"111111111",
  53344=>"111111110",
  53345=>"111111110",
  53346=>"000000011",
  53347=>"111111111",
  53348=>"000000000",
  53349=>"001000101",
  53350=>"011011011",
  53351=>"111000000",
  53352=>"000000000",
  53353=>"000000111",
  53354=>"010000100",
  53355=>"111111001",
  53356=>"001111111",
  53357=>"000000000",
  53358=>"011001101",
  53359=>"111111110",
  53360=>"000010000",
  53361=>"000000000",
  53362=>"111111011",
  53363=>"100101111",
  53364=>"000001001",
  53365=>"011001101",
  53366=>"011000011",
  53367=>"001000001",
  53368=>"000000000",
  53369=>"011111000",
  53370=>"000001100",
  53371=>"010000000",
  53372=>"011011001",
  53373=>"000001111",
  53374=>"000000000",
  53375=>"000000000",
  53376=>"111111111",
  53377=>"000000100",
  53378=>"000000011",
  53379=>"011011011",
  53380=>"111111111",
  53381=>"000000111",
  53382=>"000001111",
  53383=>"000010111",
  53384=>"000000000",
  53385=>"100000100",
  53386=>"111111111",
  53387=>"111111111",
  53388=>"111111000",
  53389=>"111111111",
  53390=>"111111100",
  53391=>"000000100",
  53392=>"110000001",
  53393=>"000000010",
  53394=>"000101111",
  53395=>"111111100",
  53396=>"000000000",
  53397=>"111011111",
  53398=>"111111111",
  53399=>"000000000",
  53400=>"111111110",
  53401=>"111111001",
  53402=>"000000000",
  53403=>"000000100",
  53404=>"001011001",
  53405=>"100101000",
  53406=>"001011001",
  53407=>"000111111",
  53408=>"111111111",
  53409=>"011001000",
  53410=>"111000000",
  53411=>"111111100",
  53412=>"001100100",
  53413=>"111110111",
  53414=>"010111111",
  53415=>"110010110",
  53416=>"000001111",
  53417=>"111111111",
  53418=>"111000000",
  53419=>"111111000",
  53420=>"111011001",
  53421=>"011001111",
  53422=>"000000000",
  53423=>"000000000",
  53424=>"000000111",
  53425=>"011001111",
  53426=>"110110110",
  53427=>"000000000",
  53428=>"101101111",
  53429=>"101111011",
  53430=>"000001011",
  53431=>"000000000",
  53432=>"000000000",
  53433=>"110110110",
  53434=>"101100100",
  53435=>"000000110",
  53436=>"000000000",
  53437=>"000000010",
  53438=>"100111000",
  53439=>"000001001",
  53440=>"000000011",
  53441=>"001011000",
  53442=>"000010111",
  53443=>"111011000",
  53444=>"111111100",
  53445=>"111111111",
  53446=>"000001011",
  53447=>"001101100",
  53448=>"101111111",
  53449=>"000111111",
  53450=>"001001001",
  53451=>"100100000",
  53452=>"111111000",
  53453=>"111111111",
  53454=>"100000000",
  53455=>"000001001",
  53456=>"111111000",
  53457=>"000000000",
  53458=>"111000000",
  53459=>"000000111",
  53460=>"000000111",
  53461=>"110110111",
  53462=>"111001011",
  53463=>"111111011",
  53464=>"111001111",
  53465=>"100100100",
  53466=>"000011000",
  53467=>"000000001",
  53468=>"111111001",
  53469=>"001011111",
  53470=>"010000000",
  53471=>"011001111",
  53472=>"111111111",
  53473=>"000000111",
  53474=>"000000000",
  53475=>"111100100",
  53476=>"100100111",
  53477=>"100100000",
  53478=>"001001001",
  53479=>"111111111",
  53480=>"110111000",
  53481=>"111111111",
  53482=>"110111111",
  53483=>"010000000",
  53484=>"000001111",
  53485=>"000000000",
  53486=>"111110000",
  53487=>"000000000",
  53488=>"111111000",
  53489=>"111000000",
  53490=>"110110100",
  53491=>"111111110",
  53492=>"001001111",
  53493=>"111111111",
  53494=>"000000111",
  53495=>"000011011",
  53496=>"000000000",
  53497=>"011001000",
  53498=>"111111111",
  53499=>"101100000",
  53500=>"111111111",
  53501=>"100100100",
  53502=>"011001111",
  53503=>"001101001",
  53504=>"111111111",
  53505=>"110000000",
  53506=>"111111111",
  53507=>"000000000",
  53508=>"100100000",
  53509=>"101111100",
  53510=>"101111111",
  53511=>"001000101",
  53512=>"111111111",
  53513=>"111111111",
  53514=>"111011000",
  53515=>"111111111",
  53516=>"111111111",
  53517=>"000000000",
  53518=>"110110110",
  53519=>"000000000",
  53520=>"111111111",
  53521=>"001000000",
  53522=>"000000011",
  53523=>"101100101",
  53524=>"010000000",
  53525=>"000000001",
  53526=>"111010010",
  53527=>"001000101",
  53528=>"110110110",
  53529=>"000000000",
  53530=>"011011111",
  53531=>"111001000",
  53532=>"001001001",
  53533=>"100000000",
  53534=>"111111111",
  53535=>"101111110",
  53536=>"111001001",
  53537=>"000000000",
  53538=>"010000000",
  53539=>"111111000",
  53540=>"111101100",
  53541=>"000000000",
  53542=>"001001011",
  53543=>"111110010",
  53544=>"111111011",
  53545=>"111011111",
  53546=>"110110110",
  53547=>"000011011",
  53548=>"111111111",
  53549=>"010010010",
  53550=>"000000000",
  53551=>"000000001",
  53552=>"110011101",
  53553=>"101111111",
  53554=>"000000000",
  53555=>"111111111",
  53556=>"000000000",
  53557=>"000111111",
  53558=>"111000000",
  53559=>"101111110",
  53560=>"011000000",
  53561=>"000000000",
  53562=>"000000000",
  53563=>"001101101",
  53564=>"111111111",
  53565=>"111000100",
  53566=>"101111111",
  53567=>"111111111",
  53568=>"111111111",
  53569=>"111011111",
  53570=>"000010111",
  53571=>"000001111",
  53572=>"011001111",
  53573=>"110001111",
  53574=>"000001111",
  53575=>"111111101",
  53576=>"011011111",
  53577=>"111000000",
  53578=>"000000000",
  53579=>"110111010",
  53580=>"001001000",
  53581=>"000000000",
  53582=>"001000101",
  53583=>"110110111",
  53584=>"111100101",
  53585=>"000001111",
  53586=>"000000000",
  53587=>"111111100",
  53588=>"000000000",
  53589=>"100100111",
  53590=>"011000000",
  53591=>"111000000",
  53592=>"111000000",
  53593=>"000000000",
  53594=>"010111000",
  53595=>"000111001",
  53596=>"110111011",
  53597=>"111111111",
  53598=>"110010000",
  53599=>"001000000",
  53600=>"000000000",
  53601=>"111111000",
  53602=>"111110111",
  53603=>"111111101",
  53604=>"111011011",
  53605=>"000000000",
  53606=>"000000111",
  53607=>"111011010",
  53608=>"111111001",
  53609=>"001001001",
  53610=>"010111110",
  53611=>"000000000",
  53612=>"000000000",
  53613=>"101111111",
  53614=>"000000110",
  53615=>"100000110",
  53616=>"111111111",
  53617=>"111111111",
  53618=>"000011111",
  53619=>"011011110",
  53620=>"011000000",
  53621=>"101000111",
  53622=>"101000101",
  53623=>"010101100",
  53624=>"000000100",
  53625=>"111111111",
  53626=>"000010111",
  53627=>"111000101",
  53628=>"011011100",
  53629=>"000000001",
  53630=>"001011111",
  53631=>"100000000",
  53632=>"111111111",
  53633=>"111111000",
  53634=>"111111111",
  53635=>"000000010",
  53636=>"111111001",
  53637=>"001101111",
  53638=>"110000000",
  53639=>"111011010",
  53640=>"010111111",
  53641=>"111011111",
  53642=>"111111111",
  53643=>"011001000",
  53644=>"111111111",
  53645=>"011011010",
  53646=>"000000000",
  53647=>"000000000",
  53648=>"111111111",
  53649=>"000111110",
  53650=>"000111111",
  53651=>"111111111",
  53652=>"000000000",
  53653=>"000000000",
  53654=>"000000110",
  53655=>"011001001",
  53656=>"001000111",
  53657=>"111101001",
  53658=>"011000100",
  53659=>"111111000",
  53660=>"111111111",
  53661=>"111111110",
  53662=>"101000000",
  53663=>"000001001",
  53664=>"111001101",
  53665=>"001001111",
  53666=>"000110000",
  53667=>"111111111",
  53668=>"111111101",
  53669=>"111111110",
  53670=>"100010111",
  53671=>"111111000",
  53672=>"100000000",
  53673=>"010010000",
  53674=>"101111111",
  53675=>"001110110",
  53676=>"110000000",
  53677=>"001111111",
  53678=>"001001000",
  53679=>"000000100",
  53680=>"000000000",
  53681=>"111111111",
  53682=>"100100100",
  53683=>"000011111",
  53684=>"001000000",
  53685=>"000100000",
  53686=>"111111111",
  53687=>"110110111",
  53688=>"000000000",
  53689=>"000001000",
  53690=>"001100101",
  53691=>"111111111",
  53692=>"000000000",
  53693=>"100111111",
  53694=>"101000000",
  53695=>"000000011",
  53696=>"011000000",
  53697=>"000010000",
  53698=>"111111111",
  53699=>"111111011",
  53700=>"110110111",
  53701=>"100110111",
  53702=>"011111000",
  53703=>"000100000",
  53704=>"111111100",
  53705=>"011001011",
  53706=>"111111111",
  53707=>"000000000",
  53708=>"111000111",
  53709=>"111110110",
  53710=>"110000000",
  53711=>"000000100",
  53712=>"111111110",
  53713=>"100110110",
  53714=>"000000000",
  53715=>"111111111",
  53716=>"010011110",
  53717=>"111000001",
  53718=>"000111111",
  53719=>"011010000",
  53720=>"000000000",
  53721=>"001001011",
  53722=>"000001111",
  53723=>"000010011",
  53724=>"100000100",
  53725=>"111111100",
  53726=>"000111111",
  53727=>"110111110",
  53728=>"000000011",
  53729=>"000000000",
  53730=>"000000110",
  53731=>"001110000",
  53732=>"111111111",
  53733=>"001111111",
  53734=>"000011010",
  53735=>"000000111",
  53736=>"100111100",
  53737=>"111111111",
  53738=>"101001110",
  53739=>"000000111",
  53740=>"000000000",
  53741=>"001000100",
  53742=>"101111111",
  53743=>"000000000",
  53744=>"000100001",
  53745=>"111111111",
  53746=>"100000000",
  53747=>"111110010",
  53748=>"100110110",
  53749=>"000000000",
  53750=>"111111110",
  53751=>"000110000",
  53752=>"000000111",
  53753=>"110100100",
  53754=>"110110100",
  53755=>"111111111",
  53756=>"000000000",
  53757=>"110010000",
  53758=>"000000000",
  53759=>"000000000",
  53760=>"111111111",
  53761=>"000110100",
  53762=>"000000000",
  53763=>"000000000",
  53764=>"100000000",
  53765=>"000000000",
  53766=>"001111001",
  53767=>"000000000",
  53768=>"111111011",
  53769=>"111111011",
  53770=>"011111010",
  53771=>"110100010",
  53772=>"101111111",
  53773=>"110111110",
  53774=>"000000000",
  53775=>"000000000",
  53776=>"111111111",
  53777=>"000000000",
  53778=>"000000000",
  53779=>"000000000",
  53780=>"111000100",
  53781=>"100100111",
  53782=>"000000010",
  53783=>"010011000",
  53784=>"000000000",
  53785=>"110110100",
  53786=>"000000000",
  53787=>"011001000",
  53788=>"000001000",
  53789=>"111110110",
  53790=>"110110110",
  53791=>"111000000",
  53792=>"110000000",
  53793=>"111000000",
  53794=>"100000000",
  53795=>"110000000",
  53796=>"111111111",
  53797=>"111111111",
  53798=>"111111110",
  53799=>"010111011",
  53800=>"000000000",
  53801=>"000000000",
  53802=>"000000000",
  53803=>"100111111",
  53804=>"111111111",
  53805=>"000000000",
  53806=>"111011010",
  53807=>"000000000",
  53808=>"000000000",
  53809=>"110111111",
  53810=>"010111111",
  53811=>"111111111",
  53812=>"100100000",
  53813=>"000000001",
  53814=>"000000000",
  53815=>"111111100",
  53816=>"111111000",
  53817=>"011001011",
  53818=>"111111111",
  53819=>"110110110",
  53820=>"000000000",
  53821=>"011111000",
  53822=>"010010000",
  53823=>"111100000",
  53824=>"000000000",
  53825=>"111111110",
  53826=>"101100000",
  53827=>"111011000",
  53828=>"110111111",
  53829=>"000010000",
  53830=>"000000100",
  53831=>"011111111",
  53832=>"111111011",
  53833=>"111111101",
  53834=>"011001000",
  53835=>"110000000",
  53836=>"000010010",
  53837=>"000000000",
  53838=>"000000111",
  53839=>"111111111",
  53840=>"111111111",
  53841=>"000000000",
  53842=>"000000000",
  53843=>"000000001",
  53844=>"000111000",
  53845=>"011111100",
  53846=>"110100101",
  53847=>"111011111",
  53848=>"000000000",
  53849=>"000011000",
  53850=>"111111111",
  53851=>"111001011",
  53852=>"000000001",
  53853=>"111111000",
  53854=>"000000010",
  53855=>"110110110",
  53856=>"000000000",
  53857=>"111100000",
  53858=>"000000000",
  53859=>"000000000",
  53860=>"000000000",
  53861=>"110000000",
  53862=>"111111111",
  53863=>"111000000",
  53864=>"000000000",
  53865=>"111111111",
  53866=>"100101111",
  53867=>"111111000",
  53868=>"000100000",
  53869=>"111111111",
  53870=>"000000000",
  53871=>"000000010",
  53872=>"000000000",
  53873=>"000000000",
  53874=>"100110111",
  53875=>"000011111",
  53876=>"000000100",
  53877=>"111001000",
  53878=>"110111111",
  53879=>"000010110",
  53880=>"000000000",
  53881=>"000000010",
  53882=>"000000000",
  53883=>"111111000",
  53884=>"000000000",
  53885=>"000000000",
  53886=>"000000000",
  53887=>"000000000",
  53888=>"001001101",
  53889=>"111111111",
  53890=>"000111101",
  53891=>"000000000",
  53892=>"111011001",
  53893=>"111111111",
  53894=>"111101001",
  53895=>"000000000",
  53896=>"000000000",
  53897=>"111001001",
  53898=>"111111111",
  53899=>"101100111",
  53900=>"111111111",
  53901=>"111111110",
  53902=>"111110100",
  53903=>"111111111",
  53904=>"011111111",
  53905=>"100100000",
  53906=>"000000000",
  53907=>"111111100",
  53908=>"000000000",
  53909=>"110100111",
  53910=>"000000000",
  53911=>"000000000",
  53912=>"010000000",
  53913=>"111111111",
  53914=>"000000000",
  53915=>"111111111",
  53916=>"000000000",
  53917=>"010000000",
  53918=>"011011000",
  53919=>"011111000",
  53920=>"111111110",
  53921=>"000000000",
  53922=>"111111111",
  53923=>"111111100",
  53924=>"000110000",
  53925=>"000110100",
  53926=>"111111111",
  53927=>"111011001",
  53928=>"000000000",
  53929=>"000000010",
  53930=>"000100101",
  53931=>"111111111",
  53932=>"000000000",
  53933=>"011011001",
  53934=>"100100111",
  53935=>"011001000",
  53936=>"000111111",
  53937=>"111111011",
  53938=>"101111111",
  53939=>"111100111",
  53940=>"110111111",
  53941=>"000000000",
  53942=>"111111110",
  53943=>"111111111",
  53944=>"111011111",
  53945=>"000000000",
  53946=>"000000000",
  53947=>"000001111",
  53948=>"000000000",
  53949=>"101001000",
  53950=>"111000000",
  53951=>"111111111",
  53952=>"110000000",
  53953=>"111111111",
  53954=>"000000000",
  53955=>"000000000",
  53956=>"000000000",
  53957=>"000000000",
  53958=>"000001111",
  53959=>"111111111",
  53960=>"110110000",
  53961=>"111110100",
  53962=>"100000000",
  53963=>"001111111",
  53964=>"000011011",
  53965=>"000001110",
  53966=>"100111000",
  53967=>"000000001",
  53968=>"000000000",
  53969=>"001101101",
  53970=>"000000000",
  53971=>"000000000",
  53972=>"110111111",
  53973=>"111111000",
  53974=>"000000000",
  53975=>"001100110",
  53976=>"111111111",
  53977=>"111111111",
  53978=>"111001000",
  53979=>"000010111",
  53980=>"101100000",
  53981=>"101101111",
  53982=>"000111111",
  53983=>"000000000",
  53984=>"000010000",
  53985=>"000100111",
  53986=>"110111000",
  53987=>"100100111",
  53988=>"111101000",
  53989=>"100100110",
  53990=>"111111000",
  53991=>"110111111",
  53992=>"110010011",
  53993=>"010010000",
  53994=>"000000000",
  53995=>"110111110",
  53996=>"111001011",
  53997=>"000000000",
  53998=>"000000010",
  53999=>"001000000",
  54000=>"100000000",
  54001=>"111111111",
  54002=>"111111111",
  54003=>"010000000",
  54004=>"000010000",
  54005=>"111111011",
  54006=>"000000011",
  54007=>"111111000",
  54008=>"000000000",
  54009=>"111111100",
  54010=>"000111111",
  54011=>"010011000",
  54012=>"001101111",
  54013=>"001000100",
  54014=>"111111111",
  54015=>"000000001",
  54016=>"000000000",
  54017=>"110011011",
  54018=>"000000111",
  54019=>"010111111",
  54020=>"111111100",
  54021=>"111111101",
  54022=>"000000000",
  54023=>"000000000",
  54024=>"011000000",
  54025=>"111111111",
  54026=>"000000000",
  54027=>"100011111",
  54028=>"011011000",
  54029=>"000000000",
  54030=>"000000000",
  54031=>"111000000",
  54032=>"000000000",
  54033=>"000000101",
  54034=>"000000000",
  54035=>"000000000",
  54036=>"111100010",
  54037=>"111111110",
  54038=>"011011011",
  54039=>"111111111",
  54040=>"111111111",
  54041=>"111111111",
  54042=>"111111111",
  54043=>"111111101",
  54044=>"111111111",
  54045=>"111101111",
  54046=>"000000000",
  54047=>"110111111",
  54048=>"000000001",
  54049=>"000000101",
  54050=>"011011011",
  54051=>"000000000",
  54052=>"000000000",
  54053=>"000000000",
  54054=>"110000001",
  54055=>"000000100",
  54056=>"111110110",
  54057=>"111111111",
  54058=>"000000100",
  54059=>"001101100",
  54060=>"111100110",
  54061=>"110111111",
  54062=>"000100101",
  54063=>"000000000",
  54064=>"000000000",
  54065=>"111111000",
  54066=>"111111110",
  54067=>"111101111",
  54068=>"000000000",
  54069=>"000000011",
  54070=>"011111000",
  54071=>"001111111",
  54072=>"000000000",
  54073=>"000000111",
  54074=>"000100111",
  54075=>"000000000",
  54076=>"011111111",
  54077=>"000000100",
  54078=>"011001011",
  54079=>"111011111",
  54080=>"000000000",
  54081=>"000000000",
  54082=>"111110111",
  54083=>"111100111",
  54084=>"011001011",
  54085=>"111111011",
  54086=>"110111111",
  54087=>"000000111",
  54088=>"110110000",
  54089=>"000110110",
  54090=>"001011100",
  54091=>"110011000",
  54092=>"000100000",
  54093=>"000111111",
  54094=>"001001111",
  54095=>"000110111",
  54096=>"000000100",
  54097=>"000000001",
  54098=>"110010000",
  54099=>"000000000",
  54100=>"111000110",
  54101=>"000000001",
  54102=>"110111011",
  54103=>"011111101",
  54104=>"111111110",
  54105=>"000111111",
  54106=>"111111011",
  54107=>"000000000",
  54108=>"111111111",
  54109=>"000000000",
  54110=>"000000100",
  54111=>"111111110",
  54112=>"111110100",
  54113=>"000000000",
  54114=>"100110111",
  54115=>"000001101",
  54116=>"001011111",
  54117=>"000000000",
  54118=>"111000000",
  54119=>"001001000",
  54120=>"011010000",
  54121=>"000000010",
  54122=>"000000000",
  54123=>"111010010",
  54124=>"000000011",
  54125=>"010010000",
  54126=>"111011011",
  54127=>"111111111",
  54128=>"100100111",
  54129=>"000000000",
  54130=>"111111110",
  54131=>"011111110",
  54132=>"001111111",
  54133=>"111000000",
  54134=>"000000000",
  54135=>"000000000",
  54136=>"011011111",
  54137=>"111111111",
  54138=>"111111111",
  54139=>"000100000",
  54140=>"000000000",
  54141=>"111111111",
  54142=>"111111111",
  54143=>"000000000",
  54144=>"000000111",
  54145=>"111011000",
  54146=>"001011010",
  54147=>"101101111",
  54148=>"111110000",
  54149=>"111000000",
  54150=>"000000000",
  54151=>"000000000",
  54152=>"111111111",
  54153=>"100000000",
  54154=>"100110110",
  54155=>"000001000",
  54156=>"000000000",
  54157=>"111111000",
  54158=>"110100000",
  54159=>"000000000",
  54160=>"000000011",
  54161=>"111111011",
  54162=>"000000100",
  54163=>"111111011",
  54164=>"111111110",
  54165=>"000000000",
  54166=>"110100100",
  54167=>"000000000",
  54168=>"011111111",
  54169=>"000000000",
  54170=>"001000000",
  54171=>"111001001",
  54172=>"100111111",
  54173=>"111111111",
  54174=>"000001000",
  54175=>"000000000",
  54176=>"111001000",
  54177=>"001001001",
  54178=>"000000000",
  54179=>"001111111",
  54180=>"001110110",
  54181=>"010110000",
  54182=>"111111111",
  54183=>"111111111",
  54184=>"111100100",
  54185=>"000000000",
  54186=>"000000111",
  54187=>"101001001",
  54188=>"000000111",
  54189=>"111000000",
  54190=>"010010000",
  54191=>"111111111",
  54192=>"011111010",
  54193=>"111011011",
  54194=>"000000000",
  54195=>"000001000",
  54196=>"001011010",
  54197=>"000000000",
  54198=>"000000100",
  54199=>"111111111",
  54200=>"000010000",
  54201=>"011101110",
  54202=>"000100000",
  54203=>"111000001",
  54204=>"110111111",
  54205=>"111111111",
  54206=>"000000000",
  54207=>"011010010",
  54208=>"000000000",
  54209=>"000000000",
  54210=>"000000000",
  54211=>"011111111",
  54212=>"111110000",
  54213=>"100000000",
  54214=>"000011111",
  54215=>"000111111",
  54216=>"000000000",
  54217=>"000000000",
  54218=>"001101100",
  54219=>"111111111",
  54220=>"000000000",
  54221=>"000000000",
  54222=>"000111010",
  54223=>"111111111",
  54224=>"000000000",
  54225=>"000000000",
  54226=>"111111111",
  54227=>"111011011",
  54228=>"111111110",
  54229=>"000000000",
  54230=>"000000000",
  54231=>"000000100",
  54232=>"011111100",
  54233=>"110111011",
  54234=>"001111111",
  54235=>"110110111",
  54236=>"101100101",
  54237=>"111111111",
  54238=>"110110110",
  54239=>"111111011",
  54240=>"000000000",
  54241=>"111110111",
  54242=>"000000000",
  54243=>"111111111",
  54244=>"000110111",
  54245=>"111111111",
  54246=>"100100100",
  54247=>"001111100",
  54248=>"100110110",
  54249=>"111111100",
  54250=>"111111111",
  54251=>"000000000",
  54252=>"000000001",
  54253=>"000100110",
  54254=>"000000011",
  54255=>"111111000",
  54256=>"000000010",
  54257=>"110110000",
  54258=>"000011001",
  54259=>"010110000",
  54260=>"110111111",
  54261=>"000100110",
  54262=>"000000000",
  54263=>"100110110",
  54264=>"000000000",
  54265=>"000010000",
  54266=>"000001111",
  54267=>"000000000",
  54268=>"000010011",
  54269=>"111111111",
  54270=>"000000000",
  54271=>"111111000",
  54272=>"001011011",
  54273=>"001101000",
  54274=>"001000101",
  54275=>"000000000",
  54276=>"011100100",
  54277=>"111111011",
  54278=>"000000000",
  54279=>"111100100",
  54280=>"011111011",
  54281=>"000000101",
  54282=>"001001000",
  54283=>"111110010",
  54284=>"000000110",
  54285=>"100000000",
  54286=>"110110000",
  54287=>"001001001",
  54288=>"000001011",
  54289=>"000000111",
  54290=>"000100011",
  54291=>"000000000",
  54292=>"111000000",
  54293=>"100100110",
  54294=>"001000000",
  54295=>"001111110",
  54296=>"101101111",
  54297=>"111111101",
  54298=>"101111111",
  54299=>"110111111",
  54300=>"011000000",
  54301=>"000000000",
  54302=>"100111011",
  54303=>"000000000",
  54304=>"111000000",
  54305=>"001000001",
  54306=>"000100100",
  54307=>"000000110",
  54308=>"000000111",
  54309=>"111111000",
  54310=>"111110111",
  54311=>"111000000",
  54312=>"000111111",
  54313=>"111111111",
  54314=>"111111000",
  54315=>"111111000",
  54316=>"111111111",
  54317=>"100000000",
  54318=>"110001001",
  54319=>"001011011",
  54320=>"111000000",
  54321=>"000000001",
  54322=>"100111100",
  54323=>"111000000",
  54324=>"100000101",
  54325=>"111111101",
  54326=>"001001001",
  54327=>"001001101",
  54328=>"000000110",
  54329=>"000000000",
  54330=>"000111111",
  54331=>"000000000",
  54332=>"100000111",
  54333=>"000000100",
  54334=>"110000000",
  54335=>"111111110",
  54336=>"000001001",
  54337=>"101100000",
  54338=>"000011111",
  54339=>"000000000",
  54340=>"111000000",
  54341=>"001011001",
  54342=>"000000000",
  54343=>"110011000",
  54344=>"111111111",
  54345=>"111000111",
  54346=>"111111111",
  54347=>"000000000",
  54348=>"111111111",
  54349=>"000000011",
  54350=>"111100000",
  54351=>"111111111",
  54352=>"000000001",
  54353=>"000000000",
  54354=>"000000000",
  54355=>"111001100",
  54356=>"111111111",
  54357=>"000000000",
  54358=>"000000000",
  54359=>"111111111",
  54360=>"000000000",
  54361=>"111000000",
  54362=>"111111111",
  54363=>"110100100",
  54364=>"011111100",
  54365=>"111111111",
  54366=>"001000110",
  54367=>"111111110",
  54368=>"011000111",
  54369=>"000000000",
  54370=>"000001011",
  54371=>"001011011",
  54372=>"111111000",
  54373=>"011001001",
  54374=>"000100111",
  54375=>"011011111",
  54376=>"111111111",
  54377=>"111111111",
  54378=>"001111111",
  54379=>"100111000",
  54380=>"111011100",
  54381=>"111111010",
  54382=>"000000100",
  54383=>"110111110",
  54384=>"011111001",
  54385=>"000000000",
  54386=>"111111111",
  54387=>"110111111",
  54388=>"111111111",
  54389=>"100101110",
  54390=>"000000110",
  54391=>"111111111",
  54392=>"100000000",
  54393=>"000000000",
  54394=>"111000100",
  54395=>"000000000",
  54396=>"111110100",
  54397=>"011111111",
  54398=>"011000000",
  54399=>"111111111",
  54400=>"000000011",
  54401=>"111111111",
  54402=>"111000001",
  54403=>"101110111",
  54404=>"000000000",
  54405=>"111000000",
  54406=>"000011110",
  54407=>"111111110",
  54408=>"001001001",
  54409=>"100100000",
  54410=>"001000000",
  54411=>"001000000",
  54412=>"111111111",
  54413=>"000000111",
  54414=>"101111111",
  54415=>"111111000",
  54416=>"111111000",
  54417=>"011001000",
  54418=>"110111111",
  54419=>"111000000",
  54420=>"111111111",
  54421=>"000110100",
  54422=>"000111111",
  54423=>"110111000",
  54424=>"000000000",
  54425=>"111111000",
  54426=>"001001000",
  54427=>"000000000",
  54428=>"000001111",
  54429=>"011011111",
  54430=>"100000000",
  54431=>"000111011",
  54432=>"111000000",
  54433=>"010111111",
  54434=>"011111110",
  54435=>"000001111",
  54436=>"110000111",
  54437=>"000000000",
  54438=>"111000101",
  54439=>"000100111",
  54440=>"111111111",
  54441=>"000000000",
  54442=>"011011000",
  54443=>"111111111",
  54444=>"111111001",
  54445=>"100100110",
  54446=>"100110000",
  54447=>"000000000",
  54448=>"111111100",
  54449=>"100111110",
  54450=>"010111111",
  54451=>"111001000",
  54452=>"110111111",
  54453=>"000011011",
  54454=>"000001101",
  54455=>"001001011",
  54456=>"000000000",
  54457=>"101000001",
  54458=>"111000111",
  54459=>"111001001",
  54460=>"000000000",
  54461=>"011011111",
  54462=>"001000000",
  54463=>"000000000",
  54464=>"111111111",
  54465=>"111111111",
  54466=>"000000000",
  54467=>"110100000",
  54468=>"111110000",
  54469=>"000000000",
  54470=>"000000000",
  54471=>"000000000",
  54472=>"111111111",
  54473=>"011001000",
  54474=>"000001000",
  54475=>"010111111",
  54476=>"000000001",
  54477=>"000110111",
  54478=>"000000000",
  54479=>"011000000",
  54480=>"011101111",
  54481=>"111011000",
  54482=>"011011111",
  54483=>"000000111",
  54484=>"111111111",
  54485=>"000000000",
  54486=>"001000000",
  54487=>"000011110",
  54488=>"000000010",
  54489=>"011011000",
  54490=>"110110110",
  54491=>"111111111",
  54492=>"111111111",
  54493=>"111000000",
  54494=>"111111111",
  54495=>"001000100",
  54496=>"000000000",
  54497=>"000010000",
  54498=>"000011000",
  54499=>"111111001",
  54500=>"111111111",
  54501=>"000011011",
  54502=>"111111000",
  54503=>"000000000",
  54504=>"111111110",
  54505=>"000000000",
  54506=>"111111111",
  54507=>"000000000",
  54508=>"000000000",
  54509=>"000000011",
  54510=>"000000000",
  54511=>"001001000",
  54512=>"001100100",
  54513=>"111111111",
  54514=>"000111001",
  54515=>"100100100",
  54516=>"001011111",
  54517=>"100111011",
  54518=>"000000000",
  54519=>"111111010",
  54520=>"001011000",
  54521=>"000111001",
  54522=>"000000000",
  54523=>"011111111",
  54524=>"110100100",
  54525=>"111001000",
  54526=>"000000000",
  54527=>"000000000",
  54528=>"110110010",
  54529=>"100101101",
  54530=>"011011011",
  54531=>"000000000",
  54532=>"110111110",
  54533=>"000111111",
  54534=>"111101111",
  54535=>"001101111",
  54536=>"100110110",
  54537=>"000000000",
  54538=>"111111000",
  54539=>"101000000",
  54540=>"111111110",
  54541=>"011001111",
  54542=>"000000000",
  54543=>"000000100",
  54544=>"001000000",
  54545=>"111111111",
  54546=>"110000000",
  54547=>"001111011",
  54548=>"001000000",
  54549=>"000011111",
  54550=>"100101111",
  54551=>"000000000",
  54552=>"111111110",
  54553=>"111111111",
  54554=>"000000000",
  54555=>"000110110",
  54556=>"111111111",
  54557=>"000000000",
  54558=>"000000000",
  54559=>"111111110",
  54560=>"000000001",
  54561=>"011111010",
  54562=>"111111111",
  54563=>"101000001",
  54564=>"110111011",
  54565=>"000011111",
  54566=>"100000011",
  54567=>"000000000",
  54568=>"111111111",
  54569=>"011001001",
  54570=>"111000000",
  54571=>"111100110",
  54572=>"000000001",
  54573=>"100000100",
  54574=>"000000000",
  54575=>"000000000",
  54576=>"110111111",
  54577=>"000000000",
  54578=>"000000000",
  54579=>"000110010",
  54580=>"000000100",
  54581=>"111111000",
  54582=>"000000000",
  54583=>"000000100",
  54584=>"101001000",
  54585=>"111000000",
  54586=>"110100000",
  54587=>"000000001",
  54588=>"000000000",
  54589=>"011000000",
  54590=>"111111000",
  54591=>"111111000",
  54592=>"111101111",
  54593=>"000011111",
  54594=>"111000001",
  54595=>"111101000",
  54596=>"000000000",
  54597=>"001101000",
  54598=>"010000111",
  54599=>"111000101",
  54600=>"110111111",
  54601=>"000111111",
  54602=>"111111101",
  54603=>"110111110",
  54604=>"111111111",
  54605=>"111111011",
  54606=>"000000111",
  54607=>"000110110",
  54608=>"000101000",
  54609=>"111000110",
  54610=>"000000111",
  54611=>"000000000",
  54612=>"000000000",
  54613=>"000000011",
  54614=>"100000011",
  54615=>"001111111",
  54616=>"011111111",
  54617=>"111111001",
  54618=>"110101101",
  54619=>"000000000",
  54620=>"001001001",
  54621=>"010111111",
  54622=>"111000000",
  54623=>"100000000",
  54624=>"111111111",
  54625=>"111011111",
  54626=>"110111111",
  54627=>"100000001",
  54628=>"000000000",
  54629=>"000101101",
  54630=>"100000000",
  54631=>"001000000",
  54632=>"111101101",
  54633=>"000011111",
  54634=>"111100110",
  54635=>"111000001",
  54636=>"011111000",
  54637=>"110000100",
  54638=>"111000001",
  54639=>"011010000",
  54640=>"000100111",
  54641=>"000000011",
  54642=>"101000001",
  54643=>"110111001",
  54644=>"011011000",
  54645=>"001000100",
  54646=>"111111110",
  54647=>"000000111",
  54648=>"011000101",
  54649=>"011111010",
  54650=>"000000100",
  54651=>"001000000",
  54652=>"011111111",
  54653=>"111111111",
  54654=>"011111000",
  54655=>"111111000",
  54656=>"000011111",
  54657=>"111001011",
  54658=>"110110000",
  54659=>"000000011",
  54660=>"000000000",
  54661=>"110111111",
  54662=>"000100101",
  54663=>"111011011",
  54664=>"000000000",
  54665=>"011011111",
  54666=>"110110111",
  54667=>"000000001",
  54668=>"100100000",
  54669=>"101111111",
  54670=>"111111110",
  54671=>"111111111",
  54672=>"000000111",
  54673=>"011111100",
  54674=>"000000011",
  54675=>"000000000",
  54676=>"000000000",
  54677=>"000000000",
  54678=>"000000000",
  54679=>"111101101",
  54680=>"000000000",
  54681=>"000111111",
  54682=>"111111101",
  54683=>"000000100",
  54684=>"000000000",
  54685=>"000000100",
  54686=>"101000000",
  54687=>"000000010",
  54688=>"000000011",
  54689=>"001000101",
  54690=>"101001000",
  54691=>"000010010",
  54692=>"001001101",
  54693=>"000010111",
  54694=>"000000110",
  54695=>"111111111",
  54696=>"100000000",
  54697=>"000000000",
  54698=>"101111101",
  54699=>"111101111",
  54700=>"011111111",
  54701=>"000000000",
  54702=>"000000000",
  54703=>"111111110",
  54704=>"001111111",
  54705=>"000010011",
  54706=>"101100111",
  54707=>"000000000",
  54708=>"000000111",
  54709=>"000000000",
  54710=>"011111000",
  54711=>"111111111",
  54712=>"111111000",
  54713=>"000000000",
  54714=>"000010000",
  54715=>"000000000",
  54716=>"001111111",
  54717=>"111111110",
  54718=>"111011000",
  54719=>"110100100",
  54720=>"000000010",
  54721=>"111111001",
  54722=>"001011111",
  54723=>"111110000",
  54724=>"000000100",
  54725=>"010000000",
  54726=>"101000100",
  54727=>"111111111",
  54728=>"111111101",
  54729=>"000000000",
  54730=>"101000000",
  54731=>"111111111",
  54732=>"111001000",
  54733=>"000001001",
  54734=>"010011111",
  54735=>"010111110",
  54736=>"111011111",
  54737=>"100000101",
  54738=>"010010001",
  54739=>"000000000",
  54740=>"110110000",
  54741=>"111111000",
  54742=>"111110000",
  54743=>"000000000",
  54744=>"111111110",
  54745=>"000000000",
  54746=>"001001111",
  54747=>"010000011",
  54748=>"000000000",
  54749=>"000000000",
  54750=>"000100110",
  54751=>"111111111",
  54752=>"100101000",
  54753=>"111111111",
  54754=>"111001011",
  54755=>"000000000",
  54756=>"111111011",
  54757=>"101101101",
  54758=>"000111111",
  54759=>"000000111",
  54760=>"111111111",
  54761=>"110111001",
  54762=>"010000100",
  54763=>"111111111",
  54764=>"001111111",
  54765=>"001001101",
  54766=>"111100100",
  54767=>"111011000",
  54768=>"111001000",
  54769=>"000000000",
  54770=>"000000000",
  54771=>"000000100",
  54772=>"000000011",
  54773=>"000000011",
  54774=>"110111111",
  54775=>"100000000",
  54776=>"111111000",
  54777=>"000000000",
  54778=>"111111010",
  54779=>"000000000",
  54780=>"011111111",
  54781=>"000000000",
  54782=>"001011111",
  54783=>"111110111",
  54784=>"110000110",
  54785=>"010011111",
  54786=>"000000000",
  54787=>"110111010",
  54788=>"001000011",
  54789=>"010000000",
  54790=>"110110000",
  54791=>"111101000",
  54792=>"011111011",
  54793=>"111111111",
  54794=>"001100111",
  54795=>"111100100",
  54796=>"000000000",
  54797=>"111000000",
  54798=>"001111111",
  54799=>"111001011",
  54800=>"111111110",
  54801=>"111111101",
  54802=>"111111101",
  54803=>"111111111",
  54804=>"000000101",
  54805=>"111111000",
  54806=>"110110111",
  54807=>"111111111",
  54808=>"100110111",
  54809=>"011011011",
  54810=>"001001001",
  54811=>"000000000",
  54812=>"111111111",
  54813=>"110110110",
  54814=>"110100100",
  54815=>"100000000",
  54816=>"001000000",
  54817=>"000000011",
  54818=>"000000000",
  54819=>"111110110",
  54820=>"001011000",
  54821=>"111111100",
  54822=>"000000000",
  54823=>"111111000",
  54824=>"000000111",
  54825=>"000010000",
  54826=>"011010110",
  54827=>"110111110",
  54828=>"000000111",
  54829=>"000000001",
  54830=>"010010010",
  54831=>"000000000",
  54832=>"000000011",
  54833=>"000000000",
  54834=>"001011011",
  54835=>"111111000",
  54836=>"100100000",
  54837=>"001000000",
  54838=>"000000000",
  54839=>"001111111",
  54840=>"000111001",
  54841=>"000000000",
  54842=>"000001000",
  54843=>"110110000",
  54844=>"001101111",
  54845=>"000111111",
  54846=>"000000010",
  54847=>"111111111",
  54848=>"001011111",
  54849=>"111000000",
  54850=>"011111111",
  54851=>"111111111",
  54852=>"111111110",
  54853=>"000000000",
  54854=>"011000000",
  54855=>"111111111",
  54856=>"111111011",
  54857=>"001000001",
  54858=>"000000000",
  54859=>"000000000",
  54860=>"001000000",
  54861=>"101111110",
  54862=>"000000111",
  54863=>"111111111",
  54864=>"000000011",
  54865=>"000000000",
  54866=>"000000000",
  54867=>"000000100",
  54868=>"111111111",
  54869=>"000000000",
  54870=>"000000001",
  54871=>"000000000",
  54872=>"000000111",
  54873=>"000000000",
  54874=>"000000100",
  54875=>"100000100",
  54876=>"000000111",
  54877=>"000000000",
  54878=>"001001001",
  54879=>"000011011",
  54880=>"001000000",
  54881=>"110111111",
  54882=>"010000000",
  54883=>"111100000",
  54884=>"000000000",
  54885=>"101001001",
  54886=>"111111110",
  54887=>"110110111",
  54888=>"000000000",
  54889=>"111111110",
  54890=>"000000001",
  54891=>"111111111",
  54892=>"000011100",
  54893=>"111111110",
  54894=>"110000000",
  54895=>"000000000",
  54896=>"000101110",
  54897=>"001111111",
  54898=>"110000000",
  54899=>"011111111",
  54900=>"111111100",
  54901=>"111010000",
  54902=>"000010000",
  54903=>"001101000",
  54904=>"001001011",
  54905=>"000100111",
  54906=>"100110000",
  54907=>"111111111",
  54908=>"000000000",
  54909=>"000000111",
  54910=>"111000000",
  54911=>"000000000",
  54912=>"111111111",
  54913=>"011111111",
  54914=>"000000000",
  54915=>"000000001",
  54916=>"111101111",
  54917=>"110110110",
  54918=>"100110000",
  54919=>"000011111",
  54920=>"110111111",
  54921=>"111000000",
  54922=>"111111111",
  54923=>"000000000",
  54924=>"011111111",
  54925=>"111111111",
  54926=>"110011011",
  54927=>"000000000",
  54928=>"011011001",
  54929=>"111100100",
  54930=>"011010000",
  54931=>"000000000",
  54932=>"000000000",
  54933=>"000111111",
  54934=>"000000000",
  54935=>"111110000",
  54936=>"000000011",
  54937=>"000111011",
  54938=>"000000000",
  54939=>"011000000",
  54940=>"000100110",
  54941=>"011000001",
  54942=>"000000000",
  54943=>"000001000",
  54944=>"000001011",
  54945=>"010000000",
  54946=>"111111110",
  54947=>"000000000",
  54948=>"000000000",
  54949=>"111101111",
  54950=>"101100101",
  54951=>"110100100",
  54952=>"000001011",
  54953=>"111111111",
  54954=>"111111111",
  54955=>"100001111",
  54956=>"001000000",
  54957=>"000000000",
  54958=>"111011011",
  54959=>"001100000",
  54960=>"011011011",
  54961=>"010000000",
  54962=>"100111111",
  54963=>"000010000",
  54964=>"011000000",
  54965=>"100110000",
  54966=>"000011011",
  54967=>"111110111",
  54968=>"000001011",
  54969=>"000000000",
  54970=>"000000010",
  54971=>"111111100",
  54972=>"111111000",
  54973=>"111111110",
  54974=>"000000000",
  54975=>"100000001",
  54976=>"101100100",
  54977=>"110110010",
  54978=>"000000000",
  54979=>"000100101",
  54980=>"111111111",
  54981=>"000000011",
  54982=>"000111111",
  54983=>"000001111",
  54984=>"100110011",
  54985=>"000001001",
  54986=>"111111111",
  54987=>"110100010",
  54988=>"001101001",
  54989=>"100001111",
  54990=>"111111001",
  54991=>"000000000",
  54992=>"111000000",
  54993=>"111111111",
  54994=>"000000000",
  54995=>"111101111",
  54996=>"000000000",
  54997=>"111111111",
  54998=>"000000000",
  54999=>"000000000",
  55000=>"001011111",
  55001=>"101011000",
  55002=>"000000111",
  55003=>"000000000",
  55004=>"100000000",
  55005=>"111111001",
  55006=>"001011100",
  55007=>"000110111",
  55008=>"000111111",
  55009=>"000000111",
  55010=>"110111111",
  55011=>"000000011",
  55012=>"000000001",
  55013=>"100000001",
  55014=>"110110110",
  55015=>"111111111",
  55016=>"000011000",
  55017=>"000001111",
  55018=>"101000000",
  55019=>"000100101",
  55020=>"111000000",
  55021=>"011011011",
  55022=>"100110001",
  55023=>"011011000",
  55024=>"111111111",
  55025=>"000000111",
  55026=>"100101111",
  55027=>"000000000",
  55028=>"111111111",
  55029=>"000110110",
  55030=>"111111111",
  55031=>"000111111",
  55032=>"000000000",
  55033=>"100101000",
  55034=>"000000111",
  55035=>"111111111",
  55036=>"000000000",
  55037=>"110110110",
  55038=>"100111011",
  55039=>"000000000",
  55040=>"111111111",
  55041=>"000000000",
  55042=>"110110111",
  55043=>"111111000",
  55044=>"000111111",
  55045=>"000000000",
  55046=>"011111111",
  55047=>"000000100",
  55048=>"000000100",
  55049=>"101001000",
  55050=>"111111111",
  55051=>"110110011",
  55052=>"111110010",
  55053=>"110000000",
  55054=>"111111011",
  55055=>"111111111",
  55056=>"011111100",
  55057=>"111111110",
  55058=>"000000101",
  55059=>"001011111",
  55060=>"001000000",
  55061=>"011011100",
  55062=>"011011111",
  55063=>"000000000",
  55064=>"101101011",
  55065=>"000000111",
  55066=>"100111111",
  55067=>"101001100",
  55068=>"100111110",
  55069=>"000010111",
  55070=>"000000000",
  55071=>"010100111",
  55072=>"000100000",
  55073=>"100101000",
  55074=>"000110111",
  55075=>"000000001",
  55076=>"001011011",
  55077=>"011111110",
  55078=>"000111001",
  55079=>"001100100",
  55080=>"000000110",
  55081=>"000000000",
  55082=>"111101111",
  55083=>"111001111",
  55084=>"110110000",
  55085=>"101001001",
  55086=>"000000001",
  55087=>"000000011",
  55088=>"111111011",
  55089=>"111100000",
  55090=>"011111111",
  55091=>"010100110",
  55092=>"000000000",
  55093=>"111111111",
  55094=>"011110111",
  55095=>"111111010",
  55096=>"000000011",
  55097=>"000000010",
  55098=>"111111111",
  55099=>"111110111",
  55100=>"000001001",
  55101=>"110100000",
  55102=>"010110111",
  55103=>"000001001",
  55104=>"111000000",
  55105=>"110110000",
  55106=>"100111111",
  55107=>"000000000",
  55108=>"010111111",
  55109=>"000000000",
  55110=>"000011111",
  55111=>"110111111",
  55112=>"111100111",
  55113=>"111111010",
  55114=>"001000000",
  55115=>"100100110",
  55116=>"111111111",
  55117=>"001011111",
  55118=>"011001001",
  55119=>"100111011",
  55120=>"100110011",
  55121=>"000001001",
  55122=>"000000111",
  55123=>"011011000",
  55124=>"000000100",
  55125=>"011011011",
  55126=>"111011011",
  55127=>"111111111",
  55128=>"111111111",
  55129=>"010111111",
  55130=>"000000001",
  55131=>"011111111",
  55132=>"111111111",
  55133=>"000000000",
  55134=>"000111111",
  55135=>"001001001",
  55136=>"000001000",
  55137=>"100000000",
  55138=>"010001111",
  55139=>"001000000",
  55140=>"111111111",
  55141=>"010000000",
  55142=>"000000111",
  55143=>"111111000",
  55144=>"011001111",
  55145=>"100000000",
  55146=>"000000000",
  55147=>"011000000",
  55148=>"100010000",
  55149=>"000001001",
  55150=>"000000000",
  55151=>"111111011",
  55152=>"110111111",
  55153=>"000000000",
  55154=>"101100000",
  55155=>"100111001",
  55156=>"000000101",
  55157=>"010010011",
  55158=>"111001011",
  55159=>"000000000",
  55160=>"000000000",
  55161=>"111111111",
  55162=>"101101111",
  55163=>"011111111",
  55164=>"000000000",
  55165=>"111111111",
  55166=>"011111111",
  55167=>"000000000",
  55168=>"000000000",
  55169=>"000000110",
  55170=>"000000000",
  55171=>"111000100",
  55172=>"010110000",
  55173=>"000000000",
  55174=>"011001111",
  55175=>"000111111",
  55176=>"000000101",
  55177=>"000011000",
  55178=>"111000000",
  55179=>"111111000",
  55180=>"000000011",
  55181=>"100100000",
  55182=>"000000000",
  55183=>"111111111",
  55184=>"000000000",
  55185=>"000000000",
  55186=>"000000000",
  55187=>"000000000",
  55188=>"000000000",
  55189=>"011000000",
  55190=>"010111111",
  55191=>"000000011",
  55192=>"000000110",
  55193=>"111010000",
  55194=>"111111111",
  55195=>"111111111",
  55196=>"000000000",
  55197=>"111111111",
  55198=>"001000000",
  55199=>"111111111",
  55200=>"000000000",
  55201=>"111111111",
  55202=>"101111111",
  55203=>"000000001",
  55204=>"000100110",
  55205=>"111111111",
  55206=>"000000001",
  55207=>"000000000",
  55208=>"010000000",
  55209=>"011111111",
  55210=>"000100100",
  55211=>"000000000",
  55212=>"001001111",
  55213=>"000000011",
  55214=>"000110111",
  55215=>"111111111",
  55216=>"111011110",
  55217=>"111111111",
  55218=>"000000000",
  55219=>"111111111",
  55220=>"111001101",
  55221=>"100000000",
  55222=>"111101010",
  55223=>"001111111",
  55224=>"111111000",
  55225=>"011011001",
  55226=>"010010110",
  55227=>"110110110",
  55228=>"111111110",
  55229=>"110111010",
  55230=>"100000000",
  55231=>"110111110",
  55232=>"000111001",
  55233=>"011001001",
  55234=>"000000111",
  55235=>"111111111",
  55236=>"011111111",
  55237=>"100010000",
  55238=>"111111111",
  55239=>"111111111",
  55240=>"000000000",
  55241=>"000000000",
  55242=>"000000000",
  55243=>"000000000",
  55244=>"100010000",
  55245=>"000000000",
  55246=>"101111000",
  55247=>"001011011",
  55248=>"100100000",
  55249=>"101000000",
  55250=>"111100110",
  55251=>"010111111",
  55252=>"111111111",
  55253=>"000000001",
  55254=>"011001000",
  55255=>"000000001",
  55256=>"000001011",
  55257=>"000000000",
  55258=>"111000011",
  55259=>"000000000",
  55260=>"000000001",
  55261=>"000000000",
  55262=>"111111110",
  55263=>"000111111",
  55264=>"011000000",
  55265=>"111111111",
  55266=>"111111111",
  55267=>"000100000",
  55268=>"111111111",
  55269=>"000000000",
  55270=>"011001000",
  55271=>"000000000",
  55272=>"000010111",
  55273=>"111111111",
  55274=>"011010111",
  55275=>"000000011",
  55276=>"111000000",
  55277=>"111111000",
  55278=>"000001011",
  55279=>"111111111",
  55280=>"100000111",
  55281=>"111111111",
  55282=>"010010111",
  55283=>"100000000",
  55284=>"000000000",
  55285=>"111111001",
  55286=>"110111111",
  55287=>"001010011",
  55288=>"010000000",
  55289=>"110110110",
  55290=>"010000111",
  55291=>"111100100",
  55292=>"111110000",
  55293=>"111011111",
  55294=>"011010000",
  55295=>"000000000",
  55296=>"000000000",
  55297=>"000000000",
  55298=>"000110111",
  55299=>"111111111",
  55300=>"011111111",
  55301=>"111111111",
  55302=>"111000000",
  55303=>"000111111",
  55304=>"001000000",
  55305=>"101001000",
  55306=>"000101111",
  55307=>"111000000",
  55308=>"110000000",
  55309=>"011111111",
  55310=>"011111011",
  55311=>"011000010",
  55312=>"111101000",
  55313=>"010011111",
  55314=>"011111111",
  55315=>"100111111",
  55316=>"001001000",
  55317=>"111111000",
  55318=>"111111111",
  55319=>"100110100",
  55320=>"010110111",
  55321=>"011011011",
  55322=>"111111110",
  55323=>"000000011",
  55324=>"000000110",
  55325=>"000000101",
  55326=>"010011111",
  55327=>"101100000",
  55328=>"010000000",
  55329=>"000000101",
  55330=>"111111011",
  55331=>"111111111",
  55332=>"100000000",
  55333=>"000000000",
  55334=>"011100000",
  55335=>"001001111",
  55336=>"001001111",
  55337=>"111111000",
  55338=>"000011000",
  55339=>"001111111",
  55340=>"111111111",
  55341=>"111111001",
  55342=>"100111111",
  55343=>"011001000",
  55344=>"111011011",
  55345=>"110010111",
  55346=>"100110000",
  55347=>"010000000",
  55348=>"000001001",
  55349=>"110010010",
  55350=>"000000111",
  55351=>"110110111",
  55352=>"000111100",
  55353=>"000111001",
  55354=>"000000000",
  55355=>"000100110",
  55356=>"111000000",
  55357=>"011111101",
  55358=>"110000011",
  55359=>"111111111",
  55360=>"000011111",
  55361=>"101101111",
  55362=>"000000110",
  55363=>"111000100",
  55364=>"000000000",
  55365=>"000001011",
  55366=>"111000000",
  55367=>"111110000",
  55368=>"100111101",
  55369=>"111000111",
  55370=>"000000000",
  55371=>"100011111",
  55372=>"111111111",
  55373=>"000000001",
  55374=>"001101111",
  55375=>"111111111",
  55376=>"000100111",
  55377=>"101111101",
  55378=>"000011000",
  55379=>"110011011",
  55380=>"111111111",
  55381=>"010011111",
  55382=>"001011101",
  55383=>"111011000",
  55384=>"000111111",
  55385=>"000000110",
  55386=>"000111101",
  55387=>"000000000",
  55388=>"011000011",
  55389=>"000000000",
  55390=>"011000000",
  55391=>"100100111",
  55392=>"001000000",
  55393=>"000101111",
  55394=>"100000000",
  55395=>"001001111",
  55396=>"000001010",
  55397=>"000000101",
  55398=>"000000000",
  55399=>"000000000",
  55400=>"000000000",
  55401=>"111111100",
  55402=>"110100110",
  55403=>"000000000",
  55404=>"000000010",
  55405=>"000111111",
  55406=>"101111111",
  55407=>"000000000",
  55408=>"111111000",
  55409=>"000000111",
  55410=>"010010011",
  55411=>"001000000",
  55412=>"011111110",
  55413=>"000000010",
  55414=>"101111000",
  55415=>"010001001",
  55416=>"001000011",
  55417=>"111111110",
  55418=>"000000111",
  55419=>"000000111",
  55420=>"110000110",
  55421=>"000000000",
  55422=>"000000110",
  55423=>"001111000",
  55424=>"101100000",
  55425=>"011000000",
  55426=>"111100000",
  55427=>"010000111",
  55428=>"001011111",
  55429=>"101100111",
  55430=>"000000000",
  55431=>"111011011",
  55432=>"111001000",
  55433=>"111100000",
  55434=>"011001000",
  55435=>"111111000",
  55436=>"001000011",
  55437=>"000000000",
  55438=>"101111111",
  55439=>"111111111",
  55440=>"000110111",
  55441=>"000001111",
  55442=>"100101100",
  55443=>"001000011",
  55444=>"000110111",
  55445=>"111000010",
  55446=>"000001100",
  55447=>"100000000",
  55448=>"000000100",
  55449=>"111111100",
  55450=>"000000000",
  55451=>"110110011",
  55452=>"111111001",
  55453=>"000100111",
  55454=>"111110111",
  55455=>"011011000",
  55456=>"111000100",
  55457=>"111111111",
  55458=>"111110000",
  55459=>"111110100",
  55460=>"011000000",
  55461=>"001000000",
  55462=>"110111111",
  55463=>"001001110",
  55464=>"010101111",
  55465=>"011000111",
  55466=>"101000000",
  55467=>"000111011",
  55468=>"010110111",
  55469=>"000000101",
  55470=>"111000100",
  55471=>"000001101",
  55472=>"101111111",
  55473=>"110111111",
  55474=>"010011010",
  55475=>"000111111",
  55476=>"111110010",
  55477=>"011001111",
  55478=>"111111111",
  55479=>"111111000",
  55480=>"000000111",
  55481=>"000101111",
  55482=>"111000000",
  55483=>"110000111",
  55484=>"000000000",
  55485=>"111011011",
  55486=>"111111111",
  55487=>"111000110",
  55488=>"111111111",
  55489=>"001111110",
  55490=>"100100000",
  55491=>"000000111",
  55492=>"000000000",
  55493=>"111111000",
  55494=>"111010100",
  55495=>"011010100",
  55496=>"000111011",
  55497=>"011010000",
  55498=>"111000000",
  55499=>"111000000",
  55500=>"001100000",
  55501=>"011011000",
  55502=>"111000000",
  55503=>"010000000",
  55504=>"000000000",
  55505=>"111111111",
  55506=>"000000000",
  55507=>"110111000",
  55508=>"111111000",
  55509=>"110101101",
  55510=>"110111000",
  55511=>"000111111",
  55512=>"000111111",
  55513=>"011101000",
  55514=>"000000000",
  55515=>"011000011",
  55516=>"111110010",
  55517=>"011000000",
  55518=>"111111010",
  55519=>"011111000",
  55520=>"101000000",
  55521=>"101100000",
  55522=>"100101101",
  55523=>"000000111",
  55524=>"111000000",
  55525=>"110110000",
  55526=>"111111000",
  55527=>"111111100",
  55528=>"000001001",
  55529=>"000000100",
  55530=>"111111111",
  55531=>"111101100",
  55532=>"111111111",
  55533=>"111000000",
  55534=>"011001101",
  55535=>"111111000",
  55536=>"000000001",
  55537=>"111111111",
  55538=>"000000111",
  55539=>"111111100",
  55540=>"001011111",
  55541=>"000000000",
  55542=>"010111000",
  55543=>"111010000",
  55544=>"001011111",
  55545=>"000000111",
  55546=>"111111111",
  55547=>"001111111",
  55548=>"110010000",
  55549=>"011111101",
  55550=>"010110110",
  55551=>"001001111",
  55552=>"011001001",
  55553=>"110011000",
  55554=>"000110100",
  55555=>"001101111",
  55556=>"000110111",
  55557=>"101111111",
  55558=>"101101001",
  55559=>"000001111",
  55560=>"111111110",
  55561=>"111111111",
  55562=>"111000000",
  55563=>"001000111",
  55564=>"110110111",
  55565=>"011111111",
  55566=>"011011001",
  55567=>"111010000",
  55568=>"000010111",
  55569=>"111100000",
  55570=>"110000010",
  55571=>"011111000",
  55572=>"111011000",
  55573=>"100000000",
  55574=>"000000111",
  55575=>"111111101",
  55576=>"111111111",
  55577=>"000100100",
  55578=>"110000000",
  55579=>"000111100",
  55580=>"011011111",
  55581=>"000000111",
  55582=>"111110010",
  55583=>"111001001",
  55584=>"100100001",
  55585=>"000100110",
  55586=>"111111000",
  55587=>"111000000",
  55588=>"100010111",
  55589=>"000000000",
  55590=>"001000000",
  55591=>"000000000",
  55592=>"011000000",
  55593=>"011011010",
  55594=>"001100110",
  55595=>"000101110",
  55596=>"100000010",
  55597=>"001011111",
  55598=>"001010010",
  55599=>"011111111",
  55600=>"110111111",
  55601=>"000000010",
  55602=>"000111111",
  55603=>"111001000",
  55604=>"111101010",
  55605=>"000000000",
  55606=>"001000001",
  55607=>"111000000",
  55608=>"000111111",
  55609=>"101000001",
  55610=>"110100000",
  55611=>"111100100",
  55612=>"111110011",
  55613=>"010000000",
  55614=>"010011011",
  55615=>"011001111",
  55616=>"101111000",
  55617=>"001111111",
  55618=>"111001000",
  55619=>"000000110",
  55620=>"111110111",
  55621=>"111001000",
  55622=>"111110111",
  55623=>"111100000",
  55624=>"001111111",
  55625=>"001100110",
  55626=>"010011000",
  55627=>"000111111",
  55628=>"110110000",
  55629=>"111110011",
  55630=>"011000000",
  55631=>"011000000",
  55632=>"110110110",
  55633=>"110000111",
  55634=>"100111111",
  55635=>"000000000",
  55636=>"111111111",
  55637=>"011011011",
  55638=>"000101111",
  55639=>"011000000",
  55640=>"110111111",
  55641=>"100000110",
  55642=>"111101111",
  55643=>"000110111",
  55644=>"101101000",
  55645=>"000000000",
  55646=>"000000000",
  55647=>"000100110",
  55648=>"111111111",
  55649=>"000111111",
  55650=>"000010111",
  55651=>"100101111",
  55652=>"000000110",
  55653=>"000000000",
  55654=>"111000010",
  55655=>"000010000",
  55656=>"000111111",
  55657=>"111111000",
  55658=>"111000100",
  55659=>"001111111",
  55660=>"011011011",
  55661=>"111000101",
  55662=>"000100111",
  55663=>"011011001",
  55664=>"000000111",
  55665=>"000101111",
  55666=>"111000100",
  55667=>"000000000",
  55668=>"000110110",
  55669=>"111111100",
  55670=>"000000100",
  55671=>"000000000",
  55672=>"100000000",
  55673=>"000000111",
  55674=>"000000111",
  55675=>"011000000",
  55676=>"100100111",
  55677=>"001000101",
  55678=>"000000000",
  55679=>"000000000",
  55680=>"110010111",
  55681=>"010110111",
  55682=>"000000101",
  55683=>"000101111",
  55684=>"111111111",
  55685=>"100111111",
  55686=>"100101011",
  55687=>"111111000",
  55688=>"000000000",
  55689=>"111111111",
  55690=>"111111000",
  55691=>"111111101",
  55692=>"101000001",
  55693=>"000010000",
  55694=>"000000111",
  55695=>"000000010",
  55696=>"111111111",
  55697=>"100100011",
  55698=>"110111110",
  55699=>"011011111",
  55700=>"111000001",
  55701=>"011000000",
  55702=>"000000110",
  55703=>"110100000",
  55704=>"001111111",
  55705=>"000010011",
  55706=>"000111111",
  55707=>"001001011",
  55708=>"001000101",
  55709=>"111111111",
  55710=>"010011010",
  55711=>"000101111",
  55712=>"000000000",
  55713=>"100000000",
  55714=>"001001111",
  55715=>"111111000",
  55716=>"001000001",
  55717=>"111001000",
  55718=>"000000000",
  55719=>"101111111",
  55720=>"000111111",
  55721=>"000000111",
  55722=>"110000111",
  55723=>"111101110",
  55724=>"000000000",
  55725=>"111100111",
  55726=>"000111111",
  55727=>"011000000",
  55728=>"100000000",
  55729=>"000000000",
  55730=>"000000000",
  55731=>"111110100",
  55732=>"000101111",
  55733=>"111000100",
  55734=>"110111101",
  55735=>"111111000",
  55736=>"111111110",
  55737=>"111110000",
  55738=>"000000011",
  55739=>"111111111",
  55740=>"111111000",
  55741=>"000111111",
  55742=>"000111111",
  55743=>"010000001",
  55744=>"011000000",
  55745=>"000001000",
  55746=>"111111111",
  55747=>"111001001",
  55748=>"011111101",
  55749=>"111110000",
  55750=>"001100111",
  55751=>"001111111",
  55752=>"000000001",
  55753=>"000000111",
  55754=>"011000000",
  55755=>"000000100",
  55756=>"110110000",
  55757=>"100111110",
  55758=>"000111100",
  55759=>"111000100",
  55760=>"101101101",
  55761=>"011011000",
  55762=>"100000000",
  55763=>"001111111",
  55764=>"010011011",
  55765=>"000000111",
  55766=>"011000001",
  55767=>"000000110",
  55768=>"111011011",
  55769=>"000111111",
  55770=>"011111011",
  55771=>"011111111",
  55772=>"000000111",
  55773=>"000101000",
  55774=>"010000010",
  55775=>"010010000",
  55776=>"101000000",
  55777=>"000000000",
  55778=>"111111100",
  55779=>"000001101",
  55780=>"111111111",
  55781=>"111111111",
  55782=>"001100101",
  55783=>"100100100",
  55784=>"111110110",
  55785=>"100100100",
  55786=>"000011111",
  55787=>"001011111",
  55788=>"000000001",
  55789=>"011000111",
  55790=>"111111011",
  55791=>"000100100",
  55792=>"011011011",
  55793=>"111111111",
  55794=>"111011001",
  55795=>"000101111",
  55796=>"000111110",
  55797=>"111000000",
  55798=>"011000111",
  55799=>"010000000",
  55800=>"101101100",
  55801=>"111010000",
  55802=>"000000000",
  55803=>"000000000",
  55804=>"111111001",
  55805=>"010000000",
  55806=>"111000000",
  55807=>"001011111",
  55808=>"111111111",
  55809=>"111011000",
  55810=>"000000111",
  55811=>"111100011",
  55812=>"111101000",
  55813=>"000000000",
  55814=>"000000000",
  55815=>"000000000",
  55816=>"000000000",
  55817=>"000001101",
  55818=>"011010111",
  55819=>"111111111",
  55820=>"011001000",
  55821=>"011111111",
  55822=>"110110100",
  55823=>"000000000",
  55824=>"111111010",
  55825=>"111000000",
  55826=>"001011100",
  55827=>"000000000",
  55828=>"000000000",
  55829=>"111000101",
  55830=>"000000000",
  55831=>"111111111",
  55832=>"000000000",
  55833=>"111111000",
  55834=>"000000110",
  55835=>"111000000",
  55836=>"000000111",
  55837=>"111111111",
  55838=>"000000000",
  55839=>"111011011",
  55840=>"101111111",
  55841=>"100100110",
  55842=>"001101111",
  55843=>"111011111",
  55844=>"111001000",
  55845=>"010000000",
  55846=>"000000100",
  55847=>"111111010",
  55848=>"001101111",
  55849=>"000000000",
  55850=>"000000000",
  55851=>"000000000",
  55852=>"110000000",
  55853=>"000000111",
  55854=>"000000000",
  55855=>"111111100",
  55856=>"000000100",
  55857=>"111111111",
  55858=>"000000111",
  55859=>"111001111",
  55860=>"000010010",
  55861=>"111110100",
  55862=>"111111111",
  55863=>"000001000",
  55864=>"000000000",
  55865=>"000110111",
  55866=>"001000111",
  55867=>"001001000",
  55868=>"000000100",
  55869=>"000001011",
  55870=>"111101100",
  55871=>"001100111",
  55872=>"001010101",
  55873=>"000001001",
  55874=>"100000100",
  55875=>"111111010",
  55876=>"111111101",
  55877=>"111100000",
  55878=>"000000010",
  55879=>"010010000",
  55880=>"011011011",
  55881=>"101000001",
  55882=>"011011001",
  55883=>"111111111",
  55884=>"000111111",
  55885=>"010010111",
  55886=>"000000000",
  55887=>"000000000",
  55888=>"011111111",
  55889=>"000000000",
  55890=>"111111111",
  55891=>"110110110",
  55892=>"111111111",
  55893=>"111111001",
  55894=>"000000110",
  55895=>"111110110",
  55896=>"111111111",
  55897=>"101000000",
  55898=>"100000000",
  55899=>"000000000",
  55900=>"000000001",
  55901=>"000000111",
  55902=>"111111110",
  55903=>"111111000",
  55904=>"111101111",
  55905=>"111111111",
  55906=>"111111111",
  55907=>"111100000",
  55908=>"000100010",
  55909=>"000000000",
  55910=>"111111111",
  55911=>"111111000",
  55912=>"100000000",
  55913=>"000000000",
  55914=>"111111000",
  55915=>"111111000",
  55916=>"110111111",
  55917=>"111111111",
  55918=>"111111110",
  55919=>"111111000",
  55920=>"111111111",
  55921=>"011001111",
  55922=>"111111111",
  55923=>"111111111",
  55924=>"000000111",
  55925=>"111000000",
  55926=>"110110110",
  55927=>"111111111",
  55928=>"101111111",
  55929=>"111111111",
  55930=>"000000000",
  55931=>"000000000",
  55932=>"000110110",
  55933=>"011000000",
  55934=>"111010000",
  55935=>"011111111",
  55936=>"111111011",
  55937=>"101000100",
  55938=>"010010111",
  55939=>"000000001",
  55940=>"111111111",
  55941=>"111111111",
  55942=>"001001111",
  55943=>"110110110",
  55944=>"000000000",
  55945=>"000000011",
  55946=>"000000000",
  55947=>"011010111",
  55948=>"101111111",
  55949=>"001111111",
  55950=>"011111111",
  55951=>"111010111",
  55952=>"111010000",
  55953=>"011000000",
  55954=>"000000000",
  55955=>"000000111",
  55956=>"111111111",
  55957=>"111111101",
  55958=>"000000101",
  55959=>"000000111",
  55960=>"001000111",
  55961=>"000000000",
  55962=>"111111110",
  55963=>"110100000",
  55964=>"100100010",
  55965=>"000111111",
  55966=>"111111000",
  55967=>"011111111",
  55968=>"000000111",
  55969=>"011111100",
  55970=>"111100100",
  55971=>"000000000",
  55972=>"000000100",
  55973=>"001011111",
  55974=>"000000000",
  55975=>"000011010",
  55976=>"000010110",
  55977=>"001000000",
  55978=>"111100100",
  55979=>"000110000",
  55980=>"000100000",
  55981=>"000110111",
  55982=>"000000111",
  55983=>"011100100",
  55984=>"111111000",
  55985=>"111111011",
  55986=>"000000000",
  55987=>"010100111",
  55988=>"000000000",
  55989=>"010010010",
  55990=>"000000000",
  55991=>"000000000",
  55992=>"011111111",
  55993=>"000111000",
  55994=>"000000000",
  55995=>"000000000",
  55996=>"011011000",
  55997=>"111111111",
  55998=>"111000011",
  55999=>"000101000",
  56000=>"001001000",
  56001=>"000000100",
  56002=>"110111000",
  56003=>"000000000",
  56004=>"111000111",
  56005=>"000000111",
  56006=>"000000000",
  56007=>"000001100",
  56008=>"000000000",
  56009=>"111111111",
  56010=>"000000000",
  56011=>"111111011",
  56012=>"000100110",
  56013=>"000111110",
  56014=>"000000111",
  56015=>"010010010",
  56016=>"000010000",
  56017=>"000000101",
  56018=>"101111111",
  56019=>"001000000",
  56020=>"000000001",
  56021=>"001000000",
  56022=>"000000011",
  56023=>"000111111",
  56024=>"001111000",
  56025=>"000010110",
  56026=>"000000000",
  56027=>"000000000",
  56028=>"110101001",
  56029=>"000000100",
  56030=>"000000000",
  56031=>"000100111",
  56032=>"111111111",
  56033=>"110110110",
  56034=>"000000000",
  56035=>"000010111",
  56036=>"000000000",
  56037=>"000100000",
  56038=>"111111111",
  56039=>"000110111",
  56040=>"000000000",
  56041=>"111111111",
  56042=>"111100000",
  56043=>"001000000",
  56044=>"000000000",
  56045=>"111111111",
  56046=>"000101101",
  56047=>"001000000",
  56048=>"011001000",
  56049=>"000000100",
  56050=>"001000101",
  56051=>"000000000",
  56052=>"101111101",
  56053=>"100100001",
  56054=>"000111111",
  56055=>"100100111",
  56056=>"111111111",
  56057=>"111011000",
  56058=>"000000000",
  56059=>"000000000",
  56060=>"011111110",
  56061=>"111111111",
  56062=>"111111110",
  56063=>"111111111",
  56064=>"000111111",
  56065=>"000000000",
  56066=>"111100100",
  56067=>"000000000",
  56068=>"001100111",
  56069=>"111111000",
  56070=>"000000110",
  56071=>"000000000",
  56072=>"000011000",
  56073=>"000000000",
  56074=>"111111111",
  56075=>"111111111",
  56076=>"000000000",
  56077=>"010111111",
  56078=>"111111110",
  56079=>"110110000",
  56080=>"000000000",
  56081=>"001000001",
  56082=>"000000110",
  56083=>"001011000",
  56084=>"001000000",
  56085=>"011000000",
  56086=>"000000000",
  56087=>"000000111",
  56088=>"000000000",
  56089=>"000000000",
  56090=>"000000000",
  56091=>"011000000",
  56092=>"100000000",
  56093=>"111011000",
  56094=>"000001001",
  56095=>"000000000",
  56096=>"111111110",
  56097=>"000000101",
  56098=>"000111111",
  56099=>"001000111",
  56100=>"000111011",
  56101=>"001000111",
  56102=>"111100100",
  56103=>"111111111",
  56104=>"000000001",
  56105=>"000000111",
  56106=>"001111111",
  56107=>"001110100",
  56108=>"110111110",
  56109=>"000111111",
  56110=>"111111110",
  56111=>"000010011",
  56112=>"111111111",
  56113=>"111111111",
  56114=>"000000000",
  56115=>"110000000",
  56116=>"001000111",
  56117=>"010111111",
  56118=>"111011111",
  56119=>"000110110",
  56120=>"000000111",
  56121=>"100111111",
  56122=>"000000000",
  56123=>"000000001",
  56124=>"000000110",
  56125=>"000000110",
  56126=>"111000000",
  56127=>"000000000",
  56128=>"000000111",
  56129=>"000011000",
  56130=>"001000000",
  56131=>"000000111",
  56132=>"111111111",
  56133=>"101101000",
  56134=>"000000000",
  56135=>"001111111",
  56136=>"000000000",
  56137=>"111101101",
  56138=>"000110111",
  56139=>"000001100",
  56140=>"001010010",
  56141=>"000000000",
  56142=>"011111000",
  56143=>"110110100",
  56144=>"001100100",
  56145=>"000100110",
  56146=>"000110111",
  56147=>"000000001",
  56148=>"111111110",
  56149=>"001000001",
  56150=>"000111111",
  56151=>"000001111",
  56152=>"111111001",
  56153=>"111111111",
  56154=>"000001001",
  56155=>"110011111",
  56156=>"000000111",
  56157=>"111011001",
  56158=>"110111111",
  56159=>"111110111",
  56160=>"010000111",
  56161=>"000000000",
  56162=>"011000000",
  56163=>"111111111",
  56164=>"111101101",
  56165=>"011111000",
  56166=>"101111111",
  56167=>"000000000",
  56168=>"000010000",
  56169=>"111111010",
  56170=>"000000100",
  56171=>"001111111",
  56172=>"110000000",
  56173=>"000000100",
  56174=>"000000000",
  56175=>"000000000",
  56176=>"011001001",
  56177=>"000110000",
  56178=>"000000100",
  56179=>"111011000",
  56180=>"000000101",
  56181=>"000100110",
  56182=>"111111000",
  56183=>"111111111",
  56184=>"000000101",
  56185=>"111111111",
  56186=>"111111111",
  56187=>"000000000",
  56188=>"000000010",
  56189=>"000000000",
  56190=>"110100000",
  56191=>"011111011",
  56192=>"011001100",
  56193=>"111100111",
  56194=>"111111001",
  56195=>"111111100",
  56196=>"000000100",
  56197=>"010111111",
  56198=>"110100000",
  56199=>"100011000",
  56200=>"000000111",
  56201=>"100001000",
  56202=>"111111001",
  56203=>"110011011",
  56204=>"111111111",
  56205=>"000011011",
  56206=>"111011111",
  56207=>"001001111",
  56208=>"000000000",
  56209=>"111111111",
  56210=>"011000000",
  56211=>"000000000",
  56212=>"000000110",
  56213=>"000000000",
  56214=>"101001001",
  56215=>"010100100",
  56216=>"111111111",
  56217=>"000000101",
  56218=>"110110111",
  56219=>"011101000",
  56220=>"111111010",
  56221=>"000000110",
  56222=>"000000000",
  56223=>"000000000",
  56224=>"011111011",
  56225=>"001001000",
  56226=>"011111110",
  56227=>"111111111",
  56228=>"001000111",
  56229=>"111111111",
  56230=>"111101111",
  56231=>"110111111",
  56232=>"000000100",
  56233=>"111111111",
  56234=>"100100000",
  56235=>"011111011",
  56236=>"101001000",
  56237=>"101000100",
  56238=>"111111111",
  56239=>"000000000",
  56240=>"111111111",
  56241=>"000000000",
  56242=>"001000000",
  56243=>"001000000",
  56244=>"111111111",
  56245=>"111111111",
  56246=>"000000111",
  56247=>"111111111",
  56248=>"111111111",
  56249=>"111000000",
  56250=>"111011000",
  56251=>"111111111",
  56252=>"110010100",
  56253=>"001000000",
  56254=>"000011111",
  56255=>"000000110",
  56256=>"000100111",
  56257=>"110000000",
  56258=>"000000111",
  56259=>"000000111",
  56260=>"110000101",
  56261=>"000000000",
  56262=>"010000000",
  56263=>"000000000",
  56264=>"000000001",
  56265=>"100000110",
  56266=>"000000000",
  56267=>"111111111",
  56268=>"010011111",
  56269=>"110000000",
  56270=>"000000111",
  56271=>"100100000",
  56272=>"111110111",
  56273=>"111111011",
  56274=>"111111111",
  56275=>"000000000",
  56276=>"011000000",
  56277=>"000000001",
  56278=>"000000000",
  56279=>"100100100",
  56280=>"000111001",
  56281=>"011011010",
  56282=>"000000000",
  56283=>"001000100",
  56284=>"111111111",
  56285=>"100000000",
  56286=>"000000000",
  56287=>"000000000",
  56288=>"000000111",
  56289=>"000111111",
  56290=>"000000000",
  56291=>"111111111",
  56292=>"111101000",
  56293=>"000000110",
  56294=>"110110111",
  56295=>"100111111",
  56296=>"000000000",
  56297=>"111111111",
  56298=>"000000000",
  56299=>"000001000",
  56300=>"011001111",
  56301=>"001111111",
  56302=>"100111111",
  56303=>"111111111",
  56304=>"000000000",
  56305=>"111111100",
  56306=>"111111111",
  56307=>"000000000",
  56308=>"111111111",
  56309=>"000000000",
  56310=>"111111111",
  56311=>"000100100",
  56312=>"000110111",
  56313=>"100110000",
  56314=>"111111111",
  56315=>"010111100",
  56316=>"000100001",
  56317=>"000000000",
  56318=>"111000001",
  56319=>"111111111",
  56320=>"011111111",
  56321=>"111111111",
  56322=>"101000101",
  56323=>"000000000",
  56324=>"001000100",
  56325=>"000000000",
  56326=>"011011001",
  56327=>"111111111",
  56328=>"000000010",
  56329=>"000000000",
  56330=>"000000001",
  56331=>"001101111",
  56332=>"111110100",
  56333=>"000000000",
  56334=>"101100101",
  56335=>"111111111",
  56336=>"000000000",
  56337=>"000000000",
  56338=>"000111001",
  56339=>"111111000",
  56340=>"100100000",
  56341=>"111110000",
  56342=>"111111011",
  56343=>"001001001",
  56344=>"000000000",
  56345=>"111100100",
  56346=>"111001000",
  56347=>"100000000",
  56348=>"111111111",
  56349=>"110000100",
  56350=>"100000000",
  56351=>"110011011",
  56352=>"000100100",
  56353=>"000000000",
  56354=>"110111110",
  56355=>"110110111",
  56356=>"111111111",
  56357=>"111101101",
  56358=>"000000000",
  56359=>"000000000",
  56360=>"111111111",
  56361=>"000000000",
  56362=>"111111111",
  56363=>"000000000",
  56364=>"000000010",
  56365=>"111111110",
  56366=>"001101111",
  56367=>"110111001",
  56368=>"110110111",
  56369=>"110100111",
  56370=>"000000000",
  56371=>"111100100",
  56372=>"100111000",
  56373=>"111111111",
  56374=>"001000000",
  56375=>"001000000",
  56376=>"000000000",
  56377=>"111000100",
  56378=>"000000000",
  56379=>"111111111",
  56380=>"111111111",
  56381=>"011000010",
  56382=>"110000000",
  56383=>"000001011",
  56384=>"011011011",
  56385=>"110111011",
  56386=>"111111111",
  56387=>"000010111",
  56388=>"111111111",
  56389=>"000000000",
  56390=>"011000010",
  56391=>"111111111",
  56392=>"101111110",
  56393=>"110100111",
  56394=>"000000011",
  56395=>"001000100",
  56396=>"000100100",
  56397=>"000000000",
  56398=>"111111000",
  56399=>"111110000",
  56400=>"000000000",
  56401=>"000000110",
  56402=>"000000000",
  56403=>"111011011",
  56404=>"000000000",
  56405=>"111111001",
  56406=>"001000000",
  56407=>"100000000",
  56408=>"000000001",
  56409=>"000000111",
  56410=>"111100100",
  56411=>"000000000",
  56412=>"111111111",
  56413=>"000000000",
  56414=>"010000000",
  56415=>"100010001",
  56416=>"110110110",
  56417=>"111001111",
  56418=>"111111001",
  56419=>"111111111",
  56420=>"000000010",
  56421=>"111111001",
  56422=>"000000000",
  56423=>"110000000",
  56424=>"000000000",
  56425=>"000000111",
  56426=>"000001111",
  56427=>"111111110",
  56428=>"001000000",
  56429=>"000111111",
  56430=>"111111111",
  56431=>"111111011",
  56432=>"001000111",
  56433=>"000000000",
  56434=>"111111111",
  56435=>"000000110",
  56436=>"111111111",
  56437=>"111111111",
  56438=>"110110000",
  56439=>"001000000",
  56440=>"000000100",
  56441=>"111111111",
  56442=>"000000000",
  56443=>"111111111",
  56444=>"111111111",
  56445=>"111111111",
  56446=>"111111111",
  56447=>"000000011",
  56448=>"000000000",
  56449=>"010000000",
  56450=>"001000111",
  56451=>"111011000",
  56452=>"001100111",
  56453=>"111111111",
  56454=>"111111110",
  56455=>"000000000",
  56456=>"000000000",
  56457=>"101111111",
  56458=>"111111111",
  56459=>"000000000",
  56460=>"111111101",
  56461=>"000000000",
  56462=>"000000000",
  56463=>"000000000",
  56464=>"100000000",
  56465=>"011111010",
  56466=>"001001001",
  56467=>"000000000",
  56468=>"111110111",
  56469=>"000000000",
  56470=>"000000000",
  56471=>"000000000",
  56472=>"111111011",
  56473=>"111111111",
  56474=>"000000000",
  56475=>"000000000",
  56476=>"111110100",
  56477=>"101111111",
  56478=>"111001000",
  56479=>"110000000",
  56480=>"111111110",
  56481=>"111100100",
  56482=>"000000111",
  56483=>"011001000",
  56484=>"011011001",
  56485=>"011000100",
  56486=>"100000000",
  56487=>"011011111",
  56488=>"111111000",
  56489=>"001001001",
  56490=>"000000000",
  56491=>"000000110",
  56492=>"001000000",
  56493=>"110111110",
  56494=>"000000000",
  56495=>"000000001",
  56496=>"000111111",
  56497=>"001011011",
  56498=>"110110010",
  56499=>"100000000",
  56500=>"011000000",
  56501=>"100101101",
  56502=>"000000000",
  56503=>"111111111",
  56504=>"000000111",
  56505=>"111001000",
  56506=>"100100100",
  56507=>"011001101",
  56508=>"000000000",
  56509=>"000000000",
  56510=>"000100101",
  56511=>"000000000",
  56512=>"000000000",
  56513=>"011010111",
  56514=>"000000000",
  56515=>"111111111",
  56516=>"111111111",
  56517=>"111111110",
  56518=>"111010000",
  56519=>"001000000",
  56520=>"110111111",
  56521=>"011010111",
  56522=>"110000001",
  56523=>"110110111",
  56524=>"000000110",
  56525=>"000110110",
  56526=>"111111111",
  56527=>"111000001",
  56528=>"000000000",
  56529=>"110111111",
  56530=>"011011011",
  56531=>"000000000",
  56532=>"000000000",
  56533=>"011001000",
  56534=>"000100110",
  56535=>"111111001",
  56536=>"111001111",
  56537=>"111111111",
  56538=>"111110110",
  56539=>"011011111",
  56540=>"111111010",
  56541=>"011000000",
  56542=>"110111111",
  56543=>"111111111",
  56544=>"000000111",
  56545=>"000111000",
  56546=>"000100111",
  56547=>"000000000",
  56548=>"111111111",
  56549=>"000000110",
  56550=>"000000000",
  56551=>"111111111",
  56552=>"111111011",
  56553=>"000000100",
  56554=>"000000100",
  56555=>"110111100",
  56556=>"111110110",
  56557=>"000010010",
  56558=>"000100111",
  56559=>"000000000",
  56560=>"101101001",
  56561=>"011000000",
  56562=>"000000000",
  56563=>"000000000",
  56564=>"001111111",
  56565=>"000001000",
  56566=>"000111111",
  56567=>"000000111",
  56568=>"111111111",
  56569=>"111111111",
  56570=>"111111111",
  56571=>"111111111",
  56572=>"000000000",
  56573=>"011011011",
  56574=>"000000000",
  56575=>"000000110",
  56576=>"111111000",
  56577=>"111111111",
  56578=>"011110111",
  56579=>"000000000",
  56580=>"000100111",
  56581=>"000001000",
  56582=>"000100000",
  56583=>"111011001",
  56584=>"000000000",
  56585=>"000000000",
  56586=>"111111111",
  56587=>"000000000",
  56588=>"100100100",
  56589=>"000000000",
  56590=>"111111111",
  56591=>"000000000",
  56592=>"111011011",
  56593=>"000000000",
  56594=>"111111011",
  56595=>"011100001",
  56596=>"000000000",
  56597=>"100111111",
  56598=>"000000000",
  56599=>"000000000",
  56600=>"110111111",
  56601=>"000000000",
  56602=>"111001011",
  56603=>"110000100",
  56604=>"011010110",
  56605=>"111010000",
  56606=>"011011011",
  56607=>"111110000",
  56608=>"000100000",
  56609=>"010110111",
  56610=>"111111000",
  56611=>"011111111",
  56612=>"000100110",
  56613=>"000000000",
  56614=>"000000000",
  56615=>"001000000",
  56616=>"010000000",
  56617=>"000000000",
  56618=>"111101101",
  56619=>"000111010",
  56620=>"000111111",
  56621=>"000000000",
  56622=>"100000000",
  56623=>"000000000",
  56624=>"000100100",
  56625=>"000000000",
  56626=>"111111111",
  56627=>"100111000",
  56628=>"111111111",
  56629=>"111111111",
  56630=>"111000011",
  56631=>"111111111",
  56632=>"000000000",
  56633=>"111001100",
  56634=>"111110111",
  56635=>"111111111",
  56636=>"111111111",
  56637=>"000000000",
  56638=>"111111011",
  56639=>"011100000",
  56640=>"001100000",
  56641=>"000000000",
  56642=>"000000000",
  56643=>"111111110",
  56644=>"000000111",
  56645=>"110111111",
  56646=>"010010011",
  56647=>"111111011",
  56648=>"000000000",
  56649=>"010000000",
  56650=>"110110111",
  56651=>"111111101",
  56652=>"111111111",
  56653=>"000110111",
  56654=>"000000111",
  56655=>"000000000",
  56656=>"111011001",
  56657=>"111111111",
  56658=>"111111111",
  56659=>"111001001",
  56660=>"000000000",
  56661=>"011011011",
  56662=>"111000000",
  56663=>"000001001",
  56664=>"111111111",
  56665=>"010110111",
  56666=>"011111111",
  56667=>"000000111",
  56668=>"000000111",
  56669=>"000000000",
  56670=>"000000000",
  56671=>"000001100",
  56672=>"111000111",
  56673=>"000000000",
  56674=>"110100100",
  56675=>"100000111",
  56676=>"110111110",
  56677=>"001000100",
  56678=>"000001111",
  56679=>"011000000",
  56680=>"111111111",
  56681=>"000000101",
  56682=>"111111111",
  56683=>"000000000",
  56684=>"011110110",
  56685=>"000000000",
  56686=>"000000000",
  56687=>"100000100",
  56688=>"111111011",
  56689=>"111111111",
  56690=>"111111101",
  56691=>"110111110",
  56692=>"111001000",
  56693=>"001000111",
  56694=>"000000011",
  56695=>"000110111",
  56696=>"111111111",
  56697=>"110000000",
  56698=>"000000000",
  56699=>"110111011",
  56700=>"001000010",
  56701=>"011010000",
  56702=>"000000000",
  56703=>"111111111",
  56704=>"010110100",
  56705=>"000000000",
  56706=>"000000000",
  56707=>"101111111",
  56708=>"011111111",
  56709=>"000000000",
  56710=>"111111111",
  56711=>"000000000",
  56712=>"110110000",
  56713=>"011001001",
  56714=>"110000000",
  56715=>"000000000",
  56716=>"111111111",
  56717=>"101110110",
  56718=>"000000000",
  56719=>"000000000",
  56720=>"000000000",
  56721=>"111111111",
  56722=>"000000000",
  56723=>"111000000",
  56724=>"001000000",
  56725=>"010011000",
  56726=>"111111111",
  56727=>"111111111",
  56728=>"100110111",
  56729=>"111111111",
  56730=>"111111111",
  56731=>"111110111",
  56732=>"111011000",
  56733=>"111111111",
  56734=>"111111111",
  56735=>"000000000",
  56736=>"001100000",
  56737=>"000000011",
  56738=>"001000000",
  56739=>"000000000",
  56740=>"000000111",
  56741=>"111111110",
  56742=>"100000110",
  56743=>"000000000",
  56744=>"111111111",
  56745=>"110000110",
  56746=>"001101111",
  56747=>"000000100",
  56748=>"000011000",
  56749=>"111011011",
  56750=>"000000110",
  56751=>"001001111",
  56752=>"000000110",
  56753=>"000010111",
  56754=>"110011000",
  56755=>"000000000",
  56756=>"001111111",
  56757=>"111101101",
  56758=>"110110111",
  56759=>"000000010",
  56760=>"000001011",
  56761=>"000110111",
  56762=>"000000111",
  56763=>"111011111",
  56764=>"000010011",
  56765=>"111011011",
  56766=>"111111101",
  56767=>"101111111",
  56768=>"000000000",
  56769=>"000000000",
  56770=>"000000000",
  56771=>"000000000",
  56772=>"111111111",
  56773=>"000000000",
  56774=>"000000000",
  56775=>"110111111",
  56776=>"111000110",
  56777=>"000000000",
  56778=>"000000000",
  56779=>"111111000",
  56780=>"100110100",
  56781=>"111111111",
  56782=>"110111111",
  56783=>"110100000",
  56784=>"000000001",
  56785=>"111100000",
  56786=>"110000000",
  56787=>"111111111",
  56788=>"110110110",
  56789=>"000000000",
  56790=>"000000000",
  56791=>"000000000",
  56792=>"111100111",
  56793=>"000011111",
  56794=>"111111011",
  56795=>"010010111",
  56796=>"011111111",
  56797=>"011111111",
  56798=>"000000000",
  56799=>"011011011",
  56800=>"111011111",
  56801=>"000000000",
  56802=>"001011111",
  56803=>"111111000",
  56804=>"000000001",
  56805=>"001000000",
  56806=>"111111000",
  56807=>"000000000",
  56808=>"101111111",
  56809=>"011001011",
  56810=>"100110000",
  56811=>"000000000",
  56812=>"100101111",
  56813=>"010010110",
  56814=>"000000000",
  56815=>"000000000",
  56816=>"000000101",
  56817=>"010111111",
  56818=>"000000000",
  56819=>"111110111",
  56820=>"110111000",
  56821=>"000010010",
  56822=>"111111000",
  56823=>"000000111",
  56824=>"100000000",
  56825=>"000000100",
  56826=>"000000001",
  56827=>"110100100",
  56828=>"000000000",
  56829=>"111011011",
  56830=>"000000111",
  56831=>"101111111",
  56832=>"000000000",
  56833=>"111001001",
  56834=>"111111111",
  56835=>"111001101",
  56836=>"100111110",
  56837=>"001000100",
  56838=>"111000000",
  56839=>"011111111",
  56840=>"000000000",
  56841=>"000000000",
  56842=>"000111111",
  56843=>"111101101",
  56844=>"000000000",
  56845=>"111010011",
  56846=>"101000000",
  56847=>"001111011",
  56848=>"000000001",
  56849=>"000110100",
  56850=>"000000001",
  56851=>"010011111",
  56852=>"101111111",
  56853=>"111000000",
  56854=>"000010111",
  56855=>"011100000",
  56856=>"000111111",
  56857=>"111111001",
  56858=>"000000000",
  56859=>"111111001",
  56860=>"000000111",
  56861=>"111011001",
  56862=>"100110000",
  56863=>"111111111",
  56864=>"001111111",
  56865=>"000111111",
  56866=>"000000100",
  56867=>"111111001",
  56868=>"011111111",
  56869=>"000000000",
  56870=>"100000000",
  56871=>"111111111",
  56872=>"000100000",
  56873=>"000111111",
  56874=>"001011111",
  56875=>"111111100",
  56876=>"001011000",
  56877=>"000100110",
  56878=>"000000001",
  56879=>"110111000",
  56880=>"111110100",
  56881=>"111111111",
  56882=>"000100000",
  56883=>"000011111",
  56884=>"111111001",
  56885=>"111111100",
  56886=>"111111011",
  56887=>"010111111",
  56888=>"000100110",
  56889=>"010010000",
  56890=>"000000111",
  56891=>"111011111",
  56892=>"101000000",
  56893=>"000000011",
  56894=>"110111110",
  56895=>"000000000",
  56896=>"100000111",
  56897=>"111111010",
  56898=>"000000000",
  56899=>"000000000",
  56900=>"011000000",
  56901=>"001001001",
  56902=>"000000111",
  56903=>"000000000",
  56904=>"111111111",
  56905=>"111000000",
  56906=>"111000000",
  56907=>"000000000",
  56908=>"000000000",
  56909=>"111111100",
  56910=>"111110000",
  56911=>"000000000",
  56912=>"111111111",
  56913=>"111111111",
  56914=>"000000100",
  56915=>"111111101",
  56916=>"111101100",
  56917=>"111000000",
  56918=>"000101111",
  56919=>"011111111",
  56920=>"010010000",
  56921=>"111100000",
  56922=>"000010111",
  56923=>"111011111",
  56924=>"000000000",
  56925=>"000000000",
  56926=>"111010000",
  56927=>"001011011",
  56928=>"000000000",
  56929=>"011000000",
  56930=>"111111000",
  56931=>"000000011",
  56932=>"110000001",
  56933=>"111001001",
  56934=>"111111000",
  56935=>"010000001",
  56936=>"111000000",
  56937=>"111100000",
  56938=>"111000000",
  56939=>"001000000",
  56940=>"111111110",
  56941=>"001000000",
  56942=>"101101111",
  56943=>"111111000",
  56944=>"100100000",
  56945=>"111111111",
  56946=>"001111110",
  56947=>"001000001",
  56948=>"111001001",
  56949=>"000000000",
  56950=>"111111000",
  56951=>"000100000",
  56952=>"000000000",
  56953=>"000111111",
  56954=>"000000000",
  56955=>"111110100",
  56956=>"000110111",
  56957=>"000111111",
  56958=>"000000000",
  56959=>"111111001",
  56960=>"001111001",
  56961=>"001101111",
  56962=>"000000111",
  56963=>"110100111",
  56964=>"000000000",
  56965=>"000000000",
  56966=>"111000011",
  56967=>"111000000",
  56968=>"110000000",
  56969=>"111111111",
  56970=>"100110100",
  56971=>"000110111",
  56972=>"001001111",
  56973=>"111000000",
  56974=>"000000111",
  56975=>"000000000",
  56976=>"000000010",
  56977=>"000000000",
  56978=>"000101100",
  56979=>"000001001",
  56980=>"111111000",
  56981=>"111101100",
  56982=>"000010111",
  56983=>"000000111",
  56984=>"111000000",
  56985=>"111100000",
  56986=>"111001000",
  56987=>"111111111",
  56988=>"001000101",
  56989=>"111111011",
  56990=>"111101101",
  56991=>"000000011",
  56992=>"111001000",
  56993=>"100000011",
  56994=>"101100100",
  56995=>"010111111",
  56996=>"000001001",
  56997=>"111111001",
  56998=>"111110110",
  56999=>"011111000",
  57000=>"111111111",
  57001=>"000111111",
  57002=>"111111111",
  57003=>"111100101",
  57004=>"000000000",
  57005=>"110110110",
  57006=>"111111111",
  57007=>"000110111",
  57008=>"000000000",
  57009=>"111110100",
  57010=>"111111010",
  57011=>"111111110",
  57012=>"111101101",
  57013=>"101111100",
  57014=>"111111111",
  57015=>"111101001",
  57016=>"000000010",
  57017=>"000000110",
  57018=>"000000001",
  57019=>"001000000",
  57020=>"000000111",
  57021=>"000000000",
  57022=>"000110111",
  57023=>"001001000",
  57024=>"000000000",
  57025=>"000000110",
  57026=>"111000000",
  57027=>"111111111",
  57028=>"000001111",
  57029=>"111000111",
  57030=>"111111000",
  57031=>"000101111",
  57032=>"000000111",
  57033=>"100000000",
  57034=>"011001000",
  57035=>"000000000",
  57036=>"010010011",
  57037=>"111110111",
  57038=>"111000001",
  57039=>"000100110",
  57040=>"000000111",
  57041=>"011001010",
  57042=>"011110111",
  57043=>"000000000",
  57044=>"001000000",
  57045=>"111111101",
  57046=>"000000000",
  57047=>"111111111",
  57048=>"000111110",
  57049=>"111110111",
  57050=>"000000000",
  57051=>"111111000",
  57052=>"000001111",
  57053=>"111111111",
  57054=>"111111000",
  57055=>"000000000",
  57056=>"000111111",
  57057=>"110110111",
  57058=>"111111111",
  57059=>"000000010",
  57060=>"000111001",
  57061=>"111110111",
  57062=>"100000001",
  57063=>"100110111",
  57064=>"111111111",
  57065=>"000001111",
  57066=>"111111001",
  57067=>"111111001",
  57068=>"000000000",
  57069=>"000000000",
  57070=>"000000111",
  57071=>"111111111",
  57072=>"000010000",
  57073=>"011111111",
  57074=>"000111111",
  57075=>"001001001",
  57076=>"111110000",
  57077=>"000100110",
  57078=>"011111111",
  57079=>"111111111",
  57080=>"111111000",
  57081=>"000011111",
  57082=>"111111111",
  57083=>"000000010",
  57084=>"111111111",
  57085=>"001100100",
  57086=>"000000000",
  57087=>"111111111",
  57088=>"111110100",
  57089=>"111111000",
  57090=>"111111100",
  57091=>"000111111",
  57092=>"000000000",
  57093=>"110000000",
  57094=>"100101111",
  57095=>"000000111",
  57096=>"000000000",
  57097=>"000000111",
  57098=>"111111111",
  57099=>"110010000",
  57100=>"100100100",
  57101=>"111000000",
  57102=>"111101101",
  57103=>"111111000",
  57104=>"111010000",
  57105=>"000000000",
  57106=>"000000000",
  57107=>"000000100",
  57108=>"111001011",
  57109=>"111111001",
  57110=>"000000000",
  57111=>"000000000",
  57112=>"000000110",
  57113=>"000000000",
  57114=>"111111111",
  57115=>"000000000",
  57116=>"001011001",
  57117=>"110000000",
  57118=>"000000000",
  57119=>"111110111",
  57120=>"000000000",
  57121=>"000000001",
  57122=>"111111111",
  57123=>"000000000",
  57124=>"001111111",
  57125=>"001101111",
  57126=>"100001001",
  57127=>"000010011",
  57128=>"011001111",
  57129=>"111001001",
  57130=>"101111111",
  57131=>"111111111",
  57132=>"000000110",
  57133=>"111000000",
  57134=>"000000110",
  57135=>"111011011",
  57136=>"000101111",
  57137=>"111011001",
  57138=>"111000000",
  57139=>"000000000",
  57140=>"000000000",
  57141=>"000000000",
  57142=>"111111111",
  57143=>"001000000",
  57144=>"010110010",
  57145=>"111111100",
  57146=>"011000000",
  57147=>"111011011",
  57148=>"001001001",
  57149=>"011111111",
  57150=>"010100111",
  57151=>"111111000",
  57152=>"110000000",
  57153=>"111111000",
  57154=>"111111111",
  57155=>"100000111",
  57156=>"101000000",
  57157=>"011010110",
  57158=>"000000000",
  57159=>"000000000",
  57160=>"000000000",
  57161=>"110000111",
  57162=>"111000000",
  57163=>"010111111",
  57164=>"010111111",
  57165=>"001000000",
  57166=>"101100111",
  57167=>"110111110",
  57168=>"001111111",
  57169=>"111111111",
  57170=>"000000000",
  57171=>"000000000",
  57172=>"001001111",
  57173=>"001011011",
  57174=>"000000001",
  57175=>"111000100",
  57176=>"000000000",
  57177=>"000001101",
  57178=>"111111111",
  57179=>"111000001",
  57180=>"000000001",
  57181=>"000000111",
  57182=>"111111111",
  57183=>"011101000",
  57184=>"000000000",
  57185=>"111111000",
  57186=>"001000000",
  57187=>"111111111",
  57188=>"111111000",
  57189=>"000000000",
  57190=>"000000000",
  57191=>"000000111",
  57192=>"001001000",
  57193=>"010001111",
  57194=>"010110000",
  57195=>"100000101",
  57196=>"111000000",
  57197=>"000111110",
  57198=>"111000101",
  57199=>"110110000",
  57200=>"000000011",
  57201=>"000100000",
  57202=>"111111111",
  57203=>"011111011",
  57204=>"000000000",
  57205=>"000000110",
  57206=>"000111111",
  57207=>"111111101",
  57208=>"001111111",
  57209=>"110000000",
  57210=>"111111111",
  57211=>"111000000",
  57212=>"000000000",
  57213=>"111000000",
  57214=>"001000000",
  57215=>"111111111",
  57216=>"111111111",
  57217=>"000000000",
  57218=>"001001001",
  57219=>"111111111",
  57220=>"111111110",
  57221=>"111111111",
  57222=>"111010000",
  57223=>"111111111",
  57224=>"000000000",
  57225=>"100000000",
  57226=>"000001001",
  57227=>"111110111",
  57228=>"000000111",
  57229=>"000111000",
  57230=>"111001001",
  57231=>"111100111",
  57232=>"000000000",
  57233=>"111111111",
  57234=>"100100000",
  57235=>"100100000",
  57236=>"100000000",
  57237=>"010110110",
  57238=>"000000000",
  57239=>"000000000",
  57240=>"111110001",
  57241=>"000000000",
  57242=>"111000000",
  57243=>"101001111",
  57244=>"000000111",
  57245=>"100110110",
  57246=>"110011000",
  57247=>"010010000",
  57248=>"001000100",
  57249=>"001000001",
  57250=>"101001101",
  57251=>"101111000",
  57252=>"101000000",
  57253=>"110111010",
  57254=>"000000000",
  57255=>"000000000",
  57256=>"111010010",
  57257=>"111011111",
  57258=>"111100000",
  57259=>"100000001",
  57260=>"001001101",
  57261=>"111111011",
  57262=>"111111000",
  57263=>"000000100",
  57264=>"111111000",
  57265=>"000011111",
  57266=>"000000000",
  57267=>"111111111",
  57268=>"111111111",
  57269=>"111111111",
  57270=>"000011111",
  57271=>"000000000",
  57272=>"111111111",
  57273=>"000111111",
  57274=>"011001000",
  57275=>"000000001",
  57276=>"000000110",
  57277=>"111111000",
  57278=>"100000000",
  57279=>"000000000",
  57280=>"000110111",
  57281=>"110010000",
  57282=>"111111000",
  57283=>"110000010",
  57284=>"100100000",
  57285=>"100100100",
  57286=>"100000000",
  57287=>"111000000",
  57288=>"111111111",
  57289=>"100000000",
  57290=>"001001001",
  57291=>"111111111",
  57292=>"000000000",
  57293=>"000000000",
  57294=>"000000000",
  57295=>"000010111",
  57296=>"000000000",
  57297=>"000111111",
  57298=>"000011101",
  57299=>"000000000",
  57300=>"110100000",
  57301=>"000101100",
  57302=>"111111111",
  57303=>"110100000",
  57304=>"100101000",
  57305=>"000000000",
  57306=>"011010000",
  57307=>"111100000",
  57308=>"000100000",
  57309=>"111111111",
  57310=>"000000100",
  57311=>"111011111",
  57312=>"000000000",
  57313=>"000000111",
  57314=>"001111110",
  57315=>"111111000",
  57316=>"111111011",
  57317=>"111111111",
  57318=>"111100110",
  57319=>"000101111",
  57320=>"000000101",
  57321=>"111111111",
  57322=>"101000000",
  57323=>"111111000",
  57324=>"111111111",
  57325=>"000000001",
  57326=>"111000000",
  57327=>"000000000",
  57328=>"000110110",
  57329=>"111111101",
  57330=>"001001111",
  57331=>"100110010",
  57332=>"111111111",
  57333=>"000000000",
  57334=>"000010110",
  57335=>"110000000",
  57336=>"111111111",
  57337=>"000000010",
  57338=>"000000000",
  57339=>"000100110",
  57340=>"000110100",
  57341=>"111111111",
  57342=>"000000000",
  57343=>"100110000",
  57344=>"111111111",
  57345=>"000000000",
  57346=>"000000001",
  57347=>"100111111",
  57348=>"010001011",
  57349=>"010000000",
  57350=>"000000011",
  57351=>"100000000",
  57352=>"101000100",
  57353=>"001000000",
  57354=>"111111111",
  57355=>"000110100",
  57356=>"000000100",
  57357=>"111111111",
  57358=>"000000000",
  57359=>"110111000",
  57360=>"000000000",
  57361=>"111111000",
  57362=>"111111111",
  57363=>"111110000",
  57364=>"100100111",
  57365=>"100000000",
  57366=>"000111111",
  57367=>"111110100",
  57368=>"111111001",
  57369=>"111001110",
  57370=>"000000000",
  57371=>"000000000",
  57372=>"010111111",
  57373=>"000000000",
  57374=>"001011011",
  57375=>"000100100",
  57376=>"000000000",
  57377=>"000000000",
  57378=>"000000000",
  57379=>"111111111",
  57380=>"111100101",
  57381=>"111111111",
  57382=>"000000111",
  57383=>"000001000",
  57384=>"110111111",
  57385=>"111111001",
  57386=>"111111111",
  57387=>"000000000",
  57388=>"111110110",
  57389=>"011111111",
  57390=>"111111111",
  57391=>"000000000",
  57392=>"111111111",
  57393=>"111000000",
  57394=>"001011001",
  57395=>"110100100",
  57396=>"010110100",
  57397=>"011111001",
  57398=>"000100111",
  57399=>"110000000",
  57400=>"101100110",
  57401=>"001011111",
  57402=>"111110000",
  57403=>"000000001",
  57404=>"111111111",
  57405=>"111101111",
  57406=>"000000000",
  57407=>"111111111",
  57408=>"001001101",
  57409=>"111101101",
  57410=>"000000101",
  57411=>"111111111",
  57412=>"000000000",
  57413=>"111111111",
  57414=>"100100000",
  57415=>"000000000",
  57416=>"000000001",
  57417=>"000000000",
  57418=>"000000100",
  57419=>"011111111",
  57420=>"100000111",
  57421=>"011011000",
  57422=>"111000000",
  57423=>"000000000",
  57424=>"000000110",
  57425=>"111110111",
  57426=>"110111111",
  57427=>"111111111",
  57428=>"111001001",
  57429=>"000000000",
  57430=>"010000001",
  57431=>"101101111",
  57432=>"000000000",
  57433=>"000001111",
  57434=>"110110010",
  57435=>"010011111",
  57436=>"001111111",
  57437=>"000000000",
  57438=>"000000111",
  57439=>"000001001",
  57440=>"111111111",
  57441=>"000000000",
  57442=>"000000000",
  57443=>"000000010",
  57444=>"101101110",
  57445=>"001000000",
  57446=>"000000000",
  57447=>"111111111",
  57448=>"111110010",
  57449=>"101101101",
  57450=>"000100111",
  57451=>"000010010",
  57452=>"000000000",
  57453=>"111110111",
  57454=>"000011111",
  57455=>"000001000",
  57456=>"000000000",
  57457=>"000001010",
  57458=>"011011000",
  57459=>"110011011",
  57460=>"100001011",
  57461=>"111000100",
  57462=>"111111111",
  57463=>"111111111",
  57464=>"111101111",
  57465=>"000000100",
  57466=>"001001000",
  57467=>"001100101",
  57468=>"010110110",
  57469=>"011001001",
  57470=>"010000000",
  57471=>"000000000",
  57472=>"000000000",
  57473=>"111000000",
  57474=>"000000000",
  57475=>"111111111",
  57476=>"111100000",
  57477=>"000000000",
  57478=>"001000001",
  57479=>"111111110",
  57480=>"110111111",
  57481=>"000000001",
  57482=>"000000000",
  57483=>"000000000",
  57484=>"111110111",
  57485=>"111110000",
  57486=>"000000000",
  57487=>"000000000",
  57488=>"111101000",
  57489=>"111101101",
  57490=>"010111110",
  57491=>"111011000",
  57492=>"111111111",
  57493=>"111101000",
  57494=>"011011111",
  57495=>"010000000",
  57496=>"000111111",
  57497=>"110100100",
  57498=>"000000001",
  57499=>"111000000",
  57500=>"111111111",
  57501=>"110100101",
  57502=>"101101111",
  57503=>"111111111",
  57504=>"010111001",
  57505=>"000000001",
  57506=>"011111111",
  57507=>"001001011",
  57508=>"001001000",
  57509=>"111111111",
  57510=>"000001111",
  57511=>"000010110",
  57512=>"010111111",
  57513=>"111111011",
  57514=>"111111111",
  57515=>"001000001",
  57516=>"100110110",
  57517=>"110001011",
  57518=>"011011001",
  57519=>"011011111",
  57520=>"000000000",
  57521=>"110110101",
  57522=>"111011010",
  57523=>"111001111",
  57524=>"110000100",
  57525=>"000011111",
  57526=>"000000101",
  57527=>"110100000",
  57528=>"000100100",
  57529=>"111011111",
  57530=>"000000000",
  57531=>"010010010",
  57532=>"111011000",
  57533=>"100111111",
  57534=>"000110110",
  57535=>"000000000",
  57536=>"000000000",
  57537=>"000000111",
  57538=>"000000000",
  57539=>"000011000",
  57540=>"111111111",
  57541=>"000000000",
  57542=>"011000100",
  57543=>"000001111",
  57544=>"000000111",
  57545=>"000000000",
  57546=>"000000000",
  57547=>"001000000",
  57548=>"001000000",
  57549=>"101111111",
  57550=>"000011101",
  57551=>"000000000",
  57552=>"000000001",
  57553=>"000000000",
  57554=>"111011111",
  57555=>"000000000",
  57556=>"100110110",
  57557=>"111110000",
  57558=>"000000110",
  57559=>"000000000",
  57560=>"000000001",
  57561=>"111100110",
  57562=>"000000000",
  57563=>"011111111",
  57564=>"000000000",
  57565=>"001011111",
  57566=>"001000111",
  57567=>"000000000",
  57568=>"000000000",
  57569=>"011011010",
  57570=>"000000000",
  57571=>"110000000",
  57572=>"101000001",
  57573=>"110110000",
  57574=>"110110000",
  57575=>"000101111",
  57576=>"100101111",
  57577=>"101101001",
  57578=>"111000000",
  57579=>"000000010",
  57580=>"000000000",
  57581=>"000000000",
  57582=>"000000000",
  57583=>"111010011",
  57584=>"111111111",
  57585=>"000000111",
  57586=>"000011111",
  57587=>"000000000",
  57588=>"110110011",
  57589=>"000010110",
  57590=>"111111111",
  57591=>"111000000",
  57592=>"000000000",
  57593=>"000000001",
  57594=>"000000000",
  57595=>"111111111",
  57596=>"011011111",
  57597=>"000000011",
  57598=>"000000000",
  57599=>"000100110",
  57600=>"000000001",
  57601=>"000011011",
  57602=>"000000000",
  57603=>"000110000",
  57604=>"000000000",
  57605=>"000000110",
  57606=>"111111110",
  57607=>"000000001",
  57608=>"111111111",
  57609=>"110100000",
  57610=>"111111111",
  57611=>"110000010",
  57612=>"000000000",
  57613=>"111111111",
  57614=>"110010000",
  57615=>"111000000",
  57616=>"000000000",
  57617=>"000000000",
  57618=>"000000000",
  57619=>"000000000",
  57620=>"100100001",
  57621=>"111000000",
  57622=>"000000111",
  57623=>"001000000",
  57624=>"111011111",
  57625=>"000100101",
  57626=>"000001111",
  57627=>"111001000",
  57628=>"100110110",
  57629=>"111110000",
  57630=>"000000110",
  57631=>"111111111",
  57632=>"110100111",
  57633=>"000010011",
  57634=>"111111111",
  57635=>"000001111",
  57636=>"100110111",
  57637=>"000000000",
  57638=>"100100000",
  57639=>"011000000",
  57640=>"111111111",
  57641=>"000000000",
  57642=>"111001101",
  57643=>"011000000",
  57644=>"001001001",
  57645=>"001001011",
  57646=>"110000111",
  57647=>"111110000",
  57648=>"011011111",
  57649=>"111111000",
  57650=>"111111111",
  57651=>"111000000",
  57652=>"000000000",
  57653=>"111111111",
  57654=>"000001001",
  57655=>"000000110",
  57656=>"000000000",
  57657=>"001001111",
  57658=>"000001000",
  57659=>"001000110",
  57660=>"000000000",
  57661=>"010110000",
  57662=>"110000000",
  57663=>"111111111",
  57664=>"111010000",
  57665=>"110101111",
  57666=>"001001111",
  57667=>"100100000",
  57668=>"100100000",
  57669=>"000001111",
  57670=>"101101101",
  57671=>"111111111",
  57672=>"110000001",
  57673=>"000000000",
  57674=>"111000000",
  57675=>"000101100",
  57676=>"111001000",
  57677=>"000010000",
  57678=>"000111000",
  57679=>"110001000",
  57680=>"001110101",
  57681=>"000001000",
  57682=>"100110000",
  57683=>"111110000",
  57684=>"010000100",
  57685=>"011011011",
  57686=>"000000100",
  57687=>"110011011",
  57688=>"000000000",
  57689=>"100100111",
  57690=>"001011111",
  57691=>"000111111",
  57692=>"110000000",
  57693=>"000000001",
  57694=>"111011001",
  57695=>"100000000",
  57696=>"111111111",
  57697=>"000000000",
  57698=>"100100110",
  57699=>"111111111",
  57700=>"000110111",
  57701=>"011111001",
  57702=>"000000110",
  57703=>"000000000",
  57704=>"110111111",
  57705=>"111111111",
  57706=>"000000000",
  57707=>"111101111",
  57708=>"111111111",
  57709=>"000000000",
  57710=>"100111111",
  57711=>"000000011",
  57712=>"000000000",
  57713=>"000000010",
  57714=>"000000101",
  57715=>"111001001",
  57716=>"111011000",
  57717=>"000110111",
  57718=>"000000111",
  57719=>"101111000",
  57720=>"000000000",
  57721=>"111011001",
  57722=>"111011001",
  57723=>"111011011",
  57724=>"000000000",
  57725=>"100110110",
  57726=>"000000000",
  57727=>"110111111",
  57728=>"000010010",
  57729=>"000000000",
  57730=>"111111111",
  57731=>"000000001",
  57732=>"111111111",
  57733=>"110111111",
  57734=>"000000000",
  57735=>"010000000",
  57736=>"000110110",
  57737=>"110111100",
  57738=>"000000011",
  57739=>"100000000",
  57740=>"101101111",
  57741=>"111110100",
  57742=>"000000011",
  57743=>"000000000",
  57744=>"000011011",
  57745=>"110110110",
  57746=>"111101111",
  57747=>"110001000",
  57748=>"000000111",
  57749=>"000000000",
  57750=>"000000000",
  57751=>"010011011",
  57752=>"010000000",
  57753=>"111111111",
  57754=>"111111111",
  57755=>"111111111",
  57756=>"001011111",
  57757=>"110000000",
  57758=>"111101001",
  57759=>"110111111",
  57760=>"010010000",
  57761=>"011010010",
  57762=>"000000010",
  57763=>"111011011",
  57764=>"111111111",
  57765=>"111111111",
  57766=>"111111111",
  57767=>"100110111",
  57768=>"110000000",
  57769=>"000000010",
  57770=>"000100100",
  57771=>"011001011",
  57772=>"111111111",
  57773=>"000000100",
  57774=>"000000010",
  57775=>"000000111",
  57776=>"011000000",
  57777=>"000110000",
  57778=>"000000100",
  57779=>"000000000",
  57780=>"000000000",
  57781=>"000000111",
  57782=>"110110111",
  57783=>"001000000",
  57784=>"001111011",
  57785=>"010010000",
  57786=>"001001000",
  57787=>"111111111",
  57788=>"111111100",
  57789=>"100110110",
  57790=>"011000000",
  57791=>"011010010",
  57792=>"000000000",
  57793=>"000000000",
  57794=>"000000000",
  57795=>"010000000",
  57796=>"111111000",
  57797=>"100111111",
  57798=>"000000000",
  57799=>"011000000",
  57800=>"000000111",
  57801=>"100100000",
  57802=>"000000001",
  57803=>"011001111",
  57804=>"111111110",
  57805=>"000000000",
  57806=>"000000000",
  57807=>"001000111",
  57808=>"110111111",
  57809=>"111111011",
  57810=>"111111111",
  57811=>"010010000",
  57812=>"000000000",
  57813=>"110011111",
  57814=>"101100000",
  57815=>"000000011",
  57816=>"000111111",
  57817=>"111000001",
  57818=>"101101001",
  57819=>"000000001",
  57820=>"111111000",
  57821=>"111001000",
  57822=>"111111111",
  57823=>"101111111",
  57824=>"111111110",
  57825=>"111110110",
  57826=>"000011100",
  57827=>"000000000",
  57828=>"000000110",
  57829=>"110111111",
  57830=>"000001111",
  57831=>"000010000",
  57832=>"111100111",
  57833=>"110111111",
  57834=>"110000001",
  57835=>"111111111",
  57836=>"000000000",
  57837=>"001101111",
  57838=>"111111111",
  57839=>"000000000",
  57840=>"011000000",
  57841=>"110110000",
  57842=>"111111111",
  57843=>"111011111",
  57844=>"000000001",
  57845=>"100000000",
  57846=>"000000000",
  57847=>"101111001",
  57848=>"111111100",
  57849=>"110011000",
  57850=>"111111111",
  57851=>"000000000",
  57852=>"111111111",
  57853=>"111111111",
  57854=>"000110111",
  57855=>"010000000",
  57856=>"111111110",
  57857=>"000000100",
  57858=>"111111111",
  57859=>"111111111",
  57860=>"000011111",
  57861=>"111111111",
  57862=>"000000000",
  57863=>"000011111",
  57864=>"000000000",
  57865=>"000000000",
  57866=>"111111111",
  57867=>"110110100",
  57868=>"001011111",
  57869=>"000111111",
  57870=>"111100000",
  57871=>"000110111",
  57872=>"000000110",
  57873=>"000110111",
  57874=>"000000111",
  57875=>"000000111",
  57876=>"111000111",
  57877=>"000000000",
  57878=>"000000100",
  57879=>"100111111",
  57880=>"000000000",
  57881=>"011000011",
  57882=>"110111111",
  57883=>"100000000",
  57884=>"000000000",
  57885=>"000000000",
  57886=>"110011011",
  57887=>"111111100",
  57888=>"000000111",
  57889=>"100100110",
  57890=>"101000000",
  57891=>"101001000",
  57892=>"101111111",
  57893=>"000010111",
  57894=>"001000000",
  57895=>"110110110",
  57896=>"000001111",
  57897=>"111100111",
  57898=>"000000001",
  57899=>"000000000",
  57900=>"100000101",
  57901=>"101111111",
  57902=>"100000000",
  57903=>"111001010",
  57904=>"111111111",
  57905=>"110110111",
  57906=>"000000000",
  57907=>"111111100",
  57908=>"000010111",
  57909=>"000100100",
  57910=>"111111111",
  57911=>"000111111",
  57912=>"101111111",
  57913=>"100000000",
  57914=>"101000000",
  57915=>"011011000",
  57916=>"000000000",
  57917=>"111111011",
  57918=>"011111111",
  57919=>"111101000",
  57920=>"111111101",
  57921=>"000011000",
  57922=>"111111100",
  57923=>"000000111",
  57924=>"111001001",
  57925=>"000000010",
  57926=>"110000001",
  57927=>"000000000",
  57928=>"000110011",
  57929=>"111111111",
  57930=>"111000111",
  57931=>"111001001",
  57932=>"000000000",
  57933=>"110110100",
  57934=>"000000000",
  57935=>"111111111",
  57936=>"000000000",
  57937=>"111111001",
  57938=>"111000000",
  57939=>"111111001",
  57940=>"110110110",
  57941=>"000000111",
  57942=>"111100111",
  57943=>"011000000",
  57944=>"111111001",
  57945=>"111000000",
  57946=>"000000101",
  57947=>"110110000",
  57948=>"101000000",
  57949=>"100000000",
  57950=>"111111111",
  57951=>"000000001",
  57952=>"000111111",
  57953=>"110111111",
  57954=>"101101001",
  57955=>"000000111",
  57956=>"000000000",
  57957=>"010000000",
  57958=>"100001001",
  57959=>"000011011",
  57960=>"000111111",
  57961=>"111111110",
  57962=>"011011111",
  57963=>"111111111",
  57964=>"111111111",
  57965=>"010000000",
  57966=>"111100111",
  57967=>"000000000",
  57968=>"000000111",
  57969=>"000000000",
  57970=>"000000000",
  57971=>"001001011",
  57972=>"111111111",
  57973=>"000111111",
  57974=>"100000000",
  57975=>"111111111",
  57976=>"110100000",
  57977=>"000100110",
  57978=>"000110111",
  57979=>"000000000",
  57980=>"000000010",
  57981=>"000111111",
  57982=>"000001001",
  57983=>"110100000",
  57984=>"011011011",
  57985=>"111111111",
  57986=>"000000000",
  57987=>"111111111",
  57988=>"111111011",
  57989=>"001000000",
  57990=>"110110110",
  57991=>"000000000",
  57992=>"101111011",
  57993=>"000101111",
  57994=>"001000000",
  57995=>"000000000",
  57996=>"111001000",
  57997=>"010011101",
  57998=>"000010000",
  57999=>"111111100",
  58000=>"000111111",
  58001=>"000100000",
  58002=>"111111001",
  58003=>"110111111",
  58004=>"000000001",
  58005=>"111100110",
  58006=>"111111000",
  58007=>"111101000",
  58008=>"000000110",
  58009=>"000000000",
  58010=>"000000000",
  58011=>"000000010",
  58012=>"001000000",
  58013=>"000000000",
  58014=>"000000000",
  58015=>"000011000",
  58016=>"101100000",
  58017=>"001011111",
  58018=>"111111100",
  58019=>"100110111",
  58020=>"000001011",
  58021=>"000100100",
  58022=>"000000111",
  58023=>"011011001",
  58024=>"000100000",
  58025=>"110110110",
  58026=>"001100111",
  58027=>"111110000",
  58028=>"000001111",
  58029=>"101111111",
  58030=>"000000000",
  58031=>"001001100",
  58032=>"111111101",
  58033=>"000011100",
  58034=>"111111111",
  58035=>"000000110",
  58036=>"010010111",
  58037=>"010111111",
  58038=>"110110000",
  58039=>"111111111",
  58040=>"000011001",
  58041=>"111111000",
  58042=>"000100111",
  58043=>"000000000",
  58044=>"100000100",
  58045=>"000000000",
  58046=>"011000101",
  58047=>"110111000",
  58048=>"100000000",
  58049=>"000111111",
  58050=>"001101000",
  58051=>"000000000",
  58052=>"000000000",
  58053=>"000100111",
  58054=>"000000001",
  58055=>"111111111",
  58056=>"000000111",
  58057=>"101111000",
  58058=>"000000000",
  58059=>"000110111",
  58060=>"000000000",
  58061=>"000000100",
  58062=>"111111110",
  58063=>"011011111",
  58064=>"000110111",
  58065=>"000100000",
  58066=>"100000100",
  58067=>"000000000",
  58068=>"000100101",
  58069=>"000000111",
  58070=>"000000000",
  58071=>"111111000",
  58072=>"111111111",
  58073=>"000000000",
  58074=>"110111000",
  58075=>"001000000",
  58076=>"000000000",
  58077=>"000000001",
  58078=>"100101111",
  58079=>"000000010",
  58080=>"001110000",
  58081=>"110111111",
  58082=>"111000000",
  58083=>"101100111",
  58084=>"000000000",
  58085=>"000000000",
  58086=>"001001011",
  58087=>"000000000",
  58088=>"100000111",
  58089=>"111111111",
  58090=>"001000000",
  58091=>"101111111",
  58092=>"000111111",
  58093=>"010000100",
  58094=>"111001000",
  58095=>"111111111",
  58096=>"000001111",
  58097=>"111010000",
  58098=>"000000111",
  58099=>"110111000",
  58100=>"111111111",
  58101=>"110111011",
  58102=>"110111111",
  58103=>"111111111",
  58104=>"111111111",
  58105=>"000000000",
  58106=>"011000110",
  58107=>"000000110",
  58108=>"000000100",
  58109=>"101101100",
  58110=>"111110001",
  58111=>"011011011",
  58112=>"000001001",
  58113=>"010000110",
  58114=>"000000011",
  58115=>"000000000",
  58116=>"111001011",
  58117=>"000000000",
  58118=>"111111101",
  58119=>"000000111",
  58120=>"111111111",
  58121=>"011111111",
  58122=>"001001101",
  58123=>"101011010",
  58124=>"111111000",
  58125=>"000000000",
  58126=>"111101000",
  58127=>"000000000",
  58128=>"000100110",
  58129=>"000110111",
  58130=>"011000000",
  58131=>"110111111",
  58132=>"101111100",
  58133=>"111111111",
  58134=>"000000000",
  58135=>"111111110",
  58136=>"000000000",
  58137=>"111110110",
  58138=>"110111011",
  58139=>"000000000",
  58140=>"110111111",
  58141=>"100111000",
  58142=>"000000000",
  58143=>"000000000",
  58144=>"110111111",
  58145=>"100000111",
  58146=>"110101111",
  58147=>"011111111",
  58148=>"110110010",
  58149=>"001111111",
  58150=>"000000000",
  58151=>"111111000",
  58152=>"100000000",
  58153=>"111110110",
  58154=>"100100001",
  58155=>"111101101",
  58156=>"111111110",
  58157=>"000000000",
  58158=>"000110111",
  58159=>"100001000",
  58160=>"111111110",
  58161=>"000000010",
  58162=>"000000111",
  58163=>"000000000",
  58164=>"000000000",
  58165=>"111100111",
  58166=>"011001000",
  58167=>"001000011",
  58168=>"010010111",
  58169=>"111111111",
  58170=>"111111110",
  58171=>"000011110",
  58172=>"000000000",
  58173=>"110100000",
  58174=>"111111110",
  58175=>"010000000",
  58176=>"111000000",
  58177=>"111111111",
  58178=>"111111111",
  58179=>"111000000",
  58180=>"000000000",
  58181=>"000111111",
  58182=>"111110100",
  58183=>"001001111",
  58184=>"000000111",
  58185=>"111100000",
  58186=>"000000110",
  58187=>"101001001",
  58188=>"000111111",
  58189=>"111111011",
  58190=>"101110111",
  58191=>"010111111",
  58192=>"100000000",
  58193=>"000011111",
  58194=>"111110000",
  58195=>"101000000",
  58196=>"001111111",
  58197=>"001001111",
  58198=>"111001000",
  58199=>"100110111",
  58200=>"000000100",
  58201=>"110110000",
  58202=>"000000110",
  58203=>"110111111",
  58204=>"000000000",
  58205=>"111100111",
  58206=>"110110001",
  58207=>"000000000",
  58208=>"111111111",
  58209=>"000000111",
  58210=>"011111111",
  58211=>"111111001",
  58212=>"000000000",
  58213=>"111111100",
  58214=>"000001111",
  58215=>"001001001",
  58216=>"111111001",
  58217=>"101000000",
  58218=>"111111111",
  58219=>"000000000",
  58220=>"100111111",
  58221=>"111111111",
  58222=>"000000000",
  58223=>"110111011",
  58224=>"000000000",
  58225=>"010100100",
  58226=>"111111110",
  58227=>"000000111",
  58228=>"111111000",
  58229=>"011111001",
  58230=>"000000000",
  58231=>"111111111",
  58232=>"111111011",
  58233=>"000111110",
  58234=>"000000000",
  58235=>"110110000",
  58236=>"111111100",
  58237=>"000100110",
  58238=>"000000111",
  58239=>"000000111",
  58240=>"001001111",
  58241=>"000000000",
  58242=>"000000101",
  58243=>"111110010",
  58244=>"111111110",
  58245=>"110110000",
  58246=>"001111000",
  58247=>"000000000",
  58248=>"110111010",
  58249=>"000000011",
  58250=>"110111111",
  58251=>"111111111",
  58252=>"111111111",
  58253=>"000111111",
  58254=>"010000001",
  58255=>"000000000",
  58256=>"110111111",
  58257=>"000000000",
  58258=>"000000111",
  58259=>"000100000",
  58260=>"000000000",
  58261=>"000000001",
  58262=>"111101101",
  58263=>"111000000",
  58264=>"111111111",
  58265=>"100111111",
  58266=>"101000000",
  58267=>"111111111",
  58268=>"101000000",
  58269=>"000000000",
  58270=>"000000111",
  58271=>"000000000",
  58272=>"000000000",
  58273=>"110000101",
  58274=>"111111110",
  58275=>"111111111",
  58276=>"011110000",
  58277=>"001011011",
  58278=>"000000000",
  58279=>"111111111",
  58280=>"100000000",
  58281=>"110010010",
  58282=>"111110100",
  58283=>"000000000",
  58284=>"011000000",
  58285=>"110100000",
  58286=>"111011011",
  58287=>"101111000",
  58288=>"000011111",
  58289=>"000000000",
  58290=>"111111001",
  58291=>"111111111",
  58292=>"111111011",
  58293=>"100111011",
  58294=>"111111110",
  58295=>"100110111",
  58296=>"100000000",
  58297=>"111111111",
  58298=>"000000111",
  58299=>"000110100",
  58300=>"000000000",
  58301=>"000001000",
  58302=>"111111110",
  58303=>"011001001",
  58304=>"000000111",
  58305=>"000000000",
  58306=>"001111110",
  58307=>"111111000",
  58308=>"001000000",
  58309=>"011000111",
  58310=>"111111111",
  58311=>"000000000",
  58312=>"011110000",
  58313=>"110000000",
  58314=>"111110000",
  58315=>"000011011",
  58316=>"000111111",
  58317=>"000000111",
  58318=>"100000000",
  58319=>"000100100",
  58320=>"110111111",
  58321=>"000011111",
  58322=>"001000000",
  58323=>"000000000",
  58324=>"111111111",
  58325=>"100100100",
  58326=>"111000000",
  58327=>"000100000",
  58328=>"111111111",
  58329=>"110100100",
  58330=>"100110110",
  58331=>"111111000",
  58332=>"101111101",
  58333=>"100000001",
  58334=>"111011011",
  58335=>"111010000",
  58336=>"000110111",
  58337=>"001011001",
  58338=>"000000000",
  58339=>"001111001",
  58340=>"000000000",
  58341=>"000000000",
  58342=>"000001011",
  58343=>"111000100",
  58344=>"001000000",
  58345=>"000000001",
  58346=>"001011011",
  58347=>"111110111",
  58348=>"111111011",
  58349=>"010011111",
  58350=>"111111000",
  58351=>"011011000",
  58352=>"110111111",
  58353=>"111111100",
  58354=>"000100111",
  58355=>"100110111",
  58356=>"111111111",
  58357=>"110110110",
  58358=>"000000111",
  58359=>"000110111",
  58360=>"010111101",
  58361=>"000010111",
  58362=>"011101101",
  58363=>"111111111",
  58364=>"000000100",
  58365=>"000001000",
  58366=>"000110110",
  58367=>"111111110",
  58368=>"111000101",
  58369=>"101000000",
  58370=>"111000000",
  58371=>"111001111",
  58372=>"111111101",
  58373=>"000100000",
  58374=>"111011000",
  58375=>"111111111",
  58376=>"111111111",
  58377=>"000000000",
  58378=>"000000000",
  58379=>"000000001",
  58380=>"000000000",
  58381=>"010011111",
  58382=>"000110111",
  58383=>"111111100",
  58384=>"110110111",
  58385=>"111111101",
  58386=>"111000100",
  58387=>"011111111",
  58388=>"000001011",
  58389=>"111010000",
  58390=>"111000000",
  58391=>"011111111",
  58392=>"000001011",
  58393=>"101011001",
  58394=>"000000000",
  58395=>"000000100",
  58396=>"111111111",
  58397=>"001111000",
  58398=>"111111111",
  58399=>"000111111",
  58400=>"000100111",
  58401=>"101011111",
  58402=>"111111000",
  58403=>"111111111",
  58404=>"000000000",
  58405=>"001000001",
  58406=>"000000000",
  58407=>"000000111",
  58408=>"001111111",
  58409=>"111111000",
  58410=>"000101111",
  58411=>"000000000",
  58412=>"000111111",
  58413=>"111111110",
  58414=>"001111111",
  58415=>"000000110",
  58416=>"111111111",
  58417=>"001001111",
  58418=>"111111011",
  58419=>"111000000",
  58420=>"010000010",
  58421=>"010100000",
  58422=>"000111111",
  58423=>"111111101",
  58424=>"001000000",
  58425=>"111000000",
  58426=>"000000000",
  58427=>"000000100",
  58428=>"111000000",
  58429=>"000000000",
  58430=>"000000100",
  58431=>"001000000",
  58432=>"101001000",
  58433=>"000000011",
  58434=>"111000000",
  58435=>"000000011",
  58436=>"011011101",
  58437=>"111111000",
  58438=>"011010011",
  58439=>"010000000",
  58440=>"000000100",
  58441=>"000000111",
  58442=>"000111111",
  58443=>"111111101",
  58444=>"001100111",
  58445=>"110111111",
  58446=>"001110100",
  58447=>"000010111",
  58448=>"000001111",
  58449=>"000000000",
  58450=>"111101101",
  58451=>"111111111",
  58452=>"000000000",
  58453=>"000000000",
  58454=>"111001000",
  58455=>"000100100",
  58456=>"000100100",
  58457=>"000000000",
  58458=>"000111111",
  58459=>"000110111",
  58460=>"111111000",
  58461=>"111110110",
  58462=>"000100101",
  58463=>"000000000",
  58464=>"111111100",
  58465=>"001000000",
  58466=>"110111110",
  58467=>"111010000",
  58468=>"101000000",
  58469=>"111011001",
  58470=>"000000111",
  58471=>"000000111",
  58472=>"000000111",
  58473=>"111000100",
  58474=>"011111000",
  58475=>"000101110",
  58476=>"011011001",
  58477=>"000100100",
  58478=>"000000011",
  58479=>"000100111",
  58480=>"111100111",
  58481=>"111111001",
  58482=>"100111111",
  58483=>"100100110",
  58484=>"000111110",
  58485=>"100100110",
  58486=>"000001111",
  58487=>"000000101",
  58488=>"000110100",
  58489=>"110101100",
  58490=>"000000011",
  58491=>"000111111",
  58492=>"010010010",
  58493=>"001111100",
  58494=>"000000100",
  58495=>"110111000",
  58496=>"000000000",
  58497=>"101001111",
  58498=>"000011011",
  58499=>"111111111",
  58500=>"000010111",
  58501=>"110000000",
  58502=>"100000100",
  58503=>"111011000",
  58504=>"111000111",
  58505=>"000001000",
  58506=>"001001111",
  58507=>"110000111",
  58508=>"100111000",
  58509=>"000111111",
  58510=>"000000001",
  58511=>"000000010",
  58512=>"110000000",
  58513=>"000111111",
  58514=>"101000000",
  58515=>"111111000",
  58516=>"100000000",
  58517=>"000000111",
  58518=>"110000001",
  58519=>"000000000",
  58520=>"000001101",
  58521=>"000000000",
  58522=>"111111100",
  58523=>"000000111",
  58524=>"001001000",
  58525=>"011111111",
  58526=>"111111111",
  58527=>"100000000",
  58528=>"000000000",
  58529=>"001001001",
  58530=>"001000000",
  58531=>"111111111",
  58532=>"000000000",
  58533=>"011010000",
  58534=>"111111000",
  58535=>"111110110",
  58536=>"001000000",
  58537=>"111111000",
  58538=>"111111011",
  58539=>"111111111",
  58540=>"111111111",
  58541=>"001000000",
  58542=>"111111100",
  58543=>"000000110",
  58544=>"000111111",
  58545=>"000000110",
  58546=>"110110110",
  58547=>"111000000",
  58548=>"000000111",
  58549=>"000000000",
  58550=>"111000000",
  58551=>"000000000",
  58552=>"110111111",
  58553=>"000110111",
  58554=>"000000000",
  58555=>"000000101",
  58556=>"000111111",
  58557=>"110100111",
  58558=>"000000100",
  58559=>"110111111",
  58560=>"111111000",
  58561=>"000000001",
  58562=>"100111111",
  58563=>"111101111",
  58564=>"101100111",
  58565=>"110010000",
  58566=>"111111000",
  58567=>"000000000",
  58568=>"111011001",
  58569=>"001000000",
  58570=>"111101111",
  58571=>"000001001",
  58572=>"000100000",
  58573=>"100011000",
  58574=>"000000000",
  58575=>"000000000",
  58576=>"000000111",
  58577=>"111111111",
  58578=>"111111111",
  58579=>"000000000",
  58580=>"100110001",
  58581=>"111000111",
  58582=>"111111111",
  58583=>"101100000",
  58584=>"111111100",
  58585=>"000000000",
  58586=>"000011001",
  58587=>"000000000",
  58588=>"000100111",
  58589=>"101101111",
  58590=>"000000110",
  58591=>"000000000",
  58592=>"000001011",
  58593=>"000000000",
  58594=>"011111111",
  58595=>"000000000",
  58596=>"000111101",
  58597=>"000000111",
  58598=>"010010111",
  58599=>"000000000",
  58600=>"111111111",
  58601=>"100101111",
  58602=>"111111110",
  58603=>"110000001",
  58604=>"110110010",
  58605=>"110100000",
  58606=>"111000001",
  58607=>"000000000",
  58608=>"110111100",
  58609=>"011111111",
  58610=>"001100111",
  58611=>"000000110",
  58612=>"101111000",
  58613=>"111011000",
  58614=>"111101000",
  58615=>"000111111",
  58616=>"111000000",
  58617=>"000000000",
  58618=>"001000000",
  58619=>"000000000",
  58620=>"000000000",
  58621=>"011001000",
  58622=>"111000000",
  58623=>"000111101",
  58624=>"000000000",
  58625=>"111111000",
  58626=>"111111111",
  58627=>"001111111",
  58628=>"000110101",
  58629=>"111111111",
  58630=>"000000000",
  58631=>"000000001",
  58632=>"111111000",
  58633=>"111111011",
  58634=>"100111111",
  58635=>"011111111",
  58636=>"111110110",
  58637=>"000111111",
  58638=>"000000000",
  58639=>"000110110",
  58640=>"000100111",
  58641=>"000001000",
  58642=>"000100111",
  58643=>"111000000",
  58644=>"110000000",
  58645=>"000000000",
  58646=>"111111110",
  58647=>"000000000",
  58648=>"000000000",
  58649=>"111011100",
  58650=>"111111111",
  58651=>"100100111",
  58652=>"111111111",
  58653=>"000000000",
  58654=>"111111111",
  58655=>"111010011",
  58656=>"111110000",
  58657=>"011111110",
  58658=>"111111101",
  58659=>"100111000",
  58660=>"011000111",
  58661=>"011011011",
  58662=>"100111111",
  58663=>"000100100",
  58664=>"000000000",
  58665=>"000111111",
  58666=>"111111111",
  58667=>"111111100",
  58668=>"000010100",
  58669=>"111110000",
  58670=>"111111111",
  58671=>"001101000",
  58672=>"011111111",
  58673=>"000000000",
  58674=>"100000001",
  58675=>"000100100",
  58676=>"001001011",
  58677=>"111111111",
  58678=>"000010110",
  58679=>"011111100",
  58680=>"000100000",
  58681=>"100000000",
  58682=>"000000111",
  58683=>"011111011",
  58684=>"111101000",
  58685=>"010111000",
  58686=>"101101111",
  58687=>"111111100",
  58688=>"011000000",
  58689=>"111111111",
  58690=>"000000000",
  58691=>"111111000",
  58692=>"111100000",
  58693=>"000101101",
  58694=>"011111111",
  58695=>"100111111",
  58696=>"111111000",
  58697=>"000111000",
  58698=>"111101001",
  58699=>"100100000",
  58700=>"000000000",
  58701=>"001111111",
  58702=>"001000100",
  58703=>"011011001",
  58704=>"000111111",
  58705=>"111101001",
  58706=>"111111111",
  58707=>"111101000",
  58708=>"000110000",
  58709=>"011011001",
  58710=>"111111011",
  58711=>"000000001",
  58712=>"111111111",
  58713=>"110111111",
  58714=>"000000111",
  58715=>"000000000",
  58716=>"111111000",
  58717=>"001011001",
  58718=>"000000000",
  58719=>"100101101",
  58720=>"000001001",
  58721=>"111101000",
  58722=>"100000110",
  58723=>"111111111",
  58724=>"111111110",
  58725=>"111111111",
  58726=>"000000111",
  58727=>"000111000",
  58728=>"111000001",
  58729=>"000111001",
  58730=>"111100000",
  58731=>"000000000",
  58732=>"010011000",
  58733=>"001000101",
  58734=>"111000000",
  58735=>"011001000",
  58736=>"000000110",
  58737=>"110111001",
  58738=>"111111100",
  58739=>"111011001",
  58740=>"001001111",
  58741=>"000111111",
  58742=>"000001111",
  58743=>"000000000",
  58744=>"111010111",
  58745=>"000001111",
  58746=>"111111110",
  58747=>"111111000",
  58748=>"000001111",
  58749=>"000000100",
  58750=>"000000000",
  58751=>"001111111",
  58752=>"111111111",
  58753=>"000000101",
  58754=>"100110000",
  58755=>"000000000",
  58756=>"111000000",
  58757=>"000111000",
  58758=>"000000000",
  58759=>"000100111",
  58760=>"100000101",
  58761=>"000001011",
  58762=>"000111111",
  58763=>"111111111",
  58764=>"000001111",
  58765=>"000000000",
  58766=>"101100101",
  58767=>"000000000",
  58768=>"000000001",
  58769=>"110111111",
  58770=>"000000000",
  58771=>"011001000",
  58772=>"000000000",
  58773=>"111011010",
  58774=>"111111111",
  58775=>"110111000",
  58776=>"100101111",
  58777=>"000111100",
  58778=>"101111111",
  58779=>"111111000",
  58780=>"000000000",
  58781=>"001111000",
  58782=>"010010000",
  58783=>"000000110",
  58784=>"000111111",
  58785=>"111000001",
  58786=>"000000100",
  58787=>"000000000",
  58788=>"000000000",
  58789=>"001001111",
  58790=>"111001011",
  58791=>"111000000",
  58792=>"010111111",
  58793=>"000000000",
  58794=>"000000100",
  58795=>"001011100",
  58796=>"111111000",
  58797=>"101011011",
  58798=>"111000000",
  58799=>"100110111",
  58800=>"111000000",
  58801=>"111111111",
  58802=>"000000000",
  58803=>"000000111",
  58804=>"000000111",
  58805=>"000000000",
  58806=>"100100000",
  58807=>"110111111",
  58808=>"000000111",
  58809=>"000100010",
  58810=>"011000001",
  58811=>"111111000",
  58812=>"000000000",
  58813=>"000000100",
  58814=>"000000000",
  58815=>"000000110",
  58816=>"000000000",
  58817=>"010000011",
  58818=>"011000000",
  58819=>"000000111",
  58820=>"111111111",
  58821=>"111011000",
  58822=>"111011001",
  58823=>"000010010",
  58824=>"000000000",
  58825=>"000000000",
  58826=>"000000100",
  58827=>"000000000",
  58828=>"000000110",
  58829=>"000000000",
  58830=>"000000000",
  58831=>"101000101",
  58832=>"001000000",
  58833=>"111110110",
  58834=>"111111111",
  58835=>"111111011",
  58836=>"000001011",
  58837=>"111111101",
  58838=>"100111111",
  58839=>"011010000",
  58840=>"111011000",
  58841=>"011111111",
  58842=>"000000000",
  58843=>"000000000",
  58844=>"110110100",
  58845=>"100000000",
  58846=>"100110111",
  58847=>"111111110",
  58848=>"111011001",
  58849=>"000001111",
  58850=>"111001000",
  58851=>"000010000",
  58852=>"000000000",
  58853=>"111111111",
  58854=>"101101111",
  58855=>"000110000",
  58856=>"001000000",
  58857=>"000111111",
  58858=>"101100110",
  58859=>"100111111",
  58860=>"000111000",
  58861=>"100111111",
  58862=>"111010000",
  58863=>"001001001",
  58864=>"000000111",
  58865=>"110000101",
  58866=>"001011001",
  58867=>"111011001",
  58868=>"000000110",
  58869=>"110100000",
  58870=>"111111100",
  58871=>"111011000",
  58872=>"000000000",
  58873=>"001001101",
  58874=>"111111000",
  58875=>"100111100",
  58876=>"000000000",
  58877=>"101100111",
  58878=>"000000000",
  58879=>"000001111",
  58880=>"000000000",
  58881=>"000000000",
  58882=>"000000000",
  58883=>"110111111",
  58884=>"111111111",
  58885=>"100100000",
  58886=>"110100111",
  58887=>"000000111",
  58888=>"000000100",
  58889=>"000001011",
  58890=>"111111111",
  58891=>"100111101",
  58892=>"100111111",
  58893=>"111111111",
  58894=>"111011011",
  58895=>"111110100",
  58896=>"000000111",
  58897=>"101101111",
  58898=>"110100111",
  58899=>"111111110",
  58900=>"000000000",
  58901=>"110111111",
  58902=>"110110110",
  58903=>"011111111",
  58904=>"000000000",
  58905=>"100011011",
  58906=>"111111111",
  58907=>"111011000",
  58908=>"000001001",
  58909=>"111111111",
  58910=>"000010011",
  58911=>"011001000",
  58912=>"110000110",
  58913=>"000001000",
  58914=>"000001100",
  58915=>"101100100",
  58916=>"000000001",
  58917=>"000000000",
  58918=>"110100000",
  58919=>"111111111",
  58920=>"111011011",
  58921=>"001000000",
  58922=>"000001000",
  58923=>"000000000",
  58924=>"001001000",
  58925=>"100110100",
  58926=>"000000000",
  58927=>"111110000",
  58928=>"110111110",
  58929=>"111111110",
  58930=>"011001001",
  58931=>"100100100",
  58932=>"111100000",
  58933=>"011010011",
  58934=>"111000000",
  58935=>"000000001",
  58936=>"111111111",
  58937=>"111110010",
  58938=>"111001100",
  58939=>"000011011",
  58940=>"111111000",
  58941=>"111111111",
  58942=>"001000000",
  58943=>"001001111",
  58944=>"111101000",
  58945=>"001001001",
  58946=>"111111111",
  58947=>"011011111",
  58948=>"111001001",
  58949=>"111111110",
  58950=>"111000111",
  58951=>"111000000",
  58952=>"111111111",
  58953=>"000000000",
  58954=>"111100100",
  58955=>"001001000",
  58956=>"111111111",
  58957=>"000000100",
  58958=>"000000000",
  58959=>"000000000",
  58960=>"111111101",
  58961=>"111111111",
  58962=>"010011000",
  58963=>"111111111",
  58964=>"010011110",
  58965=>"000100111",
  58966=>"001000000",
  58967=>"110111111",
  58968=>"000001000",
  58969=>"001001001",
  58970=>"000000000",
  58971=>"000011001",
  58972=>"000000000",
  58973=>"110111111",
  58974=>"000011111",
  58975=>"111111111",
  58976=>"000000000",
  58977=>"011111111",
  58978=>"000110111",
  58979=>"000000000",
  58980=>"001101000",
  58981=>"000000000",
  58982=>"111111111",
  58983=>"110110100",
  58984=>"000000000",
  58985=>"000000000",
  58986=>"000000000",
  58987=>"111111010",
  58988=>"000000000",
  58989=>"000100100",
  58990=>"001011000",
  58991=>"000000001",
  58992=>"100111111",
  58993=>"001011000",
  58994=>"111101000",
  58995=>"010011010",
  58996=>"000000110",
  58997=>"000010111",
  58998=>"000000000",
  58999=>"100000011",
  59000=>"011110111",
  59001=>"111111110",
  59002=>"100110001",
  59003=>"000000000",
  59004=>"100111110",
  59005=>"000000000",
  59006=>"100110111",
  59007=>"110000000",
  59008=>"111111111",
  59009=>"110110000",
  59010=>"111000000",
  59011=>"101111001",
  59012=>"111011011",
  59013=>"001000001",
  59014=>"111111111",
  59015=>"111001001",
  59016=>"111111111",
  59017=>"110111111",
  59018=>"000001000",
  59019=>"000000000",
  59020=>"111111101",
  59021=>"111111111",
  59022=>"000000111",
  59023=>"001000000",
  59024=>"000111111",
  59025=>"000000000",
  59026=>"000000000",
  59027=>"010000000",
  59028=>"000000011",
  59029=>"000001000",
  59030=>"110111111",
  59031=>"000000000",
  59032=>"110100110",
  59033=>"000000000",
  59034=>"111111100",
  59035=>"000000000",
  59036=>"000001011",
  59037=>"110000000",
  59038=>"000100000",
  59039=>"100000111",
  59040=>"000000110",
  59041=>"111111011",
  59042=>"000001000",
  59043=>"111111101",
  59044=>"111111111",
  59045=>"110111111",
  59046=>"000000000",
  59047=>"111111111",
  59048=>"000000000",
  59049=>"000100111",
  59050=>"100111111",
  59051=>"111111000",
  59052=>"101111111",
  59053=>"000001011",
  59054=>"000000111",
  59055=>"111111000",
  59056=>"010000000",
  59057=>"001001001",
  59058=>"111111011",
  59059=>"001001111",
  59060=>"110110100",
  59061=>"000001000",
  59062=>"001001001",
  59063=>"100000100",
  59064=>"111001111",
  59065=>"111111111",
  59066=>"100100100",
  59067=>"100000110",
  59068=>"000000010",
  59069=>"011000110",
  59070=>"111111111",
  59071=>"100111111",
  59072=>"111000000",
  59073=>"111011000",
  59074=>"111111111",
  59075=>"111111111",
  59076=>"111111010",
  59077=>"001111111",
  59078=>"110010011",
  59079=>"000001011",
  59080=>"000000000",
  59081=>"111001111",
  59082=>"111111000",
  59083=>"000000000",
  59084=>"000000000",
  59085=>"110111111",
  59086=>"000000000",
  59087=>"000000000",
  59088=>"000000000",
  59089=>"000000000",
  59090=>"000000000",
  59091=>"000010010",
  59092=>"011111111",
  59093=>"000010000",
  59094=>"000000000",
  59095=>"110000111",
  59096=>"111111100",
  59097=>"000000000",
  59098=>"011001000",
  59099=>"000101111",
  59100=>"100000100",
  59101=>"111111011",
  59102=>"011001000",
  59103=>"000001011",
  59104=>"000000000",
  59105=>"011000000",
  59106=>"000110111",
  59107=>"111000000",
  59108=>"111110000",
  59109=>"001000001",
  59110=>"111111111",
  59111=>"110110111",
  59112=>"011011110",
  59113=>"000001111",
  59114=>"000100111",
  59115=>"000001101",
  59116=>"000000101",
  59117=>"000000000",
  59118=>"000110011",
  59119=>"000110111",
  59120=>"000000000",
  59121=>"000000000",
  59122=>"110110000",
  59123=>"111001000",
  59124=>"000000100",
  59125=>"111111111",
  59126=>"000011011",
  59127=>"011111111",
  59128=>"111111111",
  59129=>"000001011",
  59130=>"001101100",
  59131=>"000000000",
  59132=>"000000000",
  59133=>"000101111",
  59134=>"100111111",
  59135=>"110100000",
  59136=>"000000000",
  59137=>"001001100",
  59138=>"011011011",
  59139=>"000000000",
  59140=>"000000101",
  59141=>"000101011",
  59142=>"000000001",
  59143=>"000111011",
  59144=>"110001100",
  59145=>"111111111",
  59146=>"010011001",
  59147=>"111111101",
  59148=>"000001111",
  59149=>"000101000",
  59150=>"011111011",
  59151=>"100000000",
  59152=>"110111110",
  59153=>"111110101",
  59154=>"111111111",
  59155=>"000100100",
  59156=>"100100000",
  59157=>"000111111",
  59158=>"110100000",
  59159=>"111110111",
  59160=>"000001111",
  59161=>"111111111",
  59162=>"111111111",
  59163=>"000000011",
  59164=>"000000000",
  59165=>"000110111",
  59166=>"100100111",
  59167=>"111100111",
  59168=>"111001001",
  59169=>"000000000",
  59170=>"010011011",
  59171=>"111111111",
  59172=>"111001111",
  59173=>"111110111",
  59174=>"111100111",
  59175=>"000100000",
  59176=>"110111111",
  59177=>"110100100",
  59178=>"110110111",
  59179=>"000100100",
  59180=>"000000111",
  59181=>"111011011",
  59182=>"000001000",
  59183=>"000000000",
  59184=>"000100100",
  59185=>"111011111",
  59186=>"001111111",
  59187=>"000010111",
  59188=>"111100000",
  59189=>"101100100",
  59190=>"100000010",
  59191=>"111011111",
  59192=>"000000000",
  59193=>"011011111",
  59194=>"000011010",
  59195=>"111111111",
  59196=>"000000000",
  59197=>"111110110",
  59198=>"000000110",
  59199=>"100000011",
  59200=>"000000000",
  59201=>"000000000",
  59202=>"000000000",
  59203=>"000000000",
  59204=>"001100100",
  59205=>"000000000",
  59206=>"000000000",
  59207=>"100100100",
  59208=>"000101000",
  59209=>"100000000",
  59210=>"101001111",
  59211=>"000110000",
  59212=>"000000000",
  59213=>"000000000",
  59214=>"111111110",
  59215=>"101101001",
  59216=>"100000100",
  59217=>"001110110",
  59218=>"111111101",
  59219=>"000000100",
  59220=>"111001001",
  59221=>"011111111",
  59222=>"000000000",
  59223=>"111111111",
  59224=>"000000000",
  59225=>"010010000",
  59226=>"111111111",
  59227=>"110111111",
  59228=>"111001000",
  59229=>"111111111",
  59230=>"001001011",
  59231=>"000000000",
  59232=>"000111011",
  59233=>"000100111",
  59234=>"000000011",
  59235=>"011111111",
  59236=>"011001001",
  59237=>"000000001",
  59238=>"111111110",
  59239=>"111111110",
  59240=>"000011000",
  59241=>"001010111",
  59242=>"000000001",
  59243=>"000000000",
  59244=>"100100000",
  59245=>"000100000",
  59246=>"110111111",
  59247=>"000000000",
  59248=>"000000000",
  59249=>"000000100",
  59250=>"111111111",
  59251=>"000000000",
  59252=>"110110110",
  59253=>"000000000",
  59254=>"011001000",
  59255=>"000111000",
  59256=>"000000100",
  59257=>"000000111",
  59258=>"111001000",
  59259=>"000000100",
  59260=>"111100111",
  59261=>"000000000",
  59262=>"110111111",
  59263=>"000000000",
  59264=>"001101100",
  59265=>"000000000",
  59266=>"011111111",
  59267=>"000000000",
  59268=>"000000000",
  59269=>"000111011",
  59270=>"001001111",
  59271=>"000000001",
  59272=>"111111111",
  59273=>"110110010",
  59274=>"000010000",
  59275=>"111111001",
  59276=>"111111101",
  59277=>"000000000",
  59278=>"001001111",
  59279=>"011000000",
  59280=>"000000111",
  59281=>"111111111",
  59282=>"111111011",
  59283=>"000010000",
  59284=>"001111111",
  59285=>"001000000",
  59286=>"111100000",
  59287=>"111000000",
  59288=>"010000000",
  59289=>"000001001",
  59290=>"110110111",
  59291=>"000011110",
  59292=>"011111111",
  59293=>"011011001",
  59294=>"110000000",
  59295=>"111111111",
  59296=>"000000000",
  59297=>"011110110",
  59298=>"001001111",
  59299=>"000000000",
  59300=>"000100111",
  59301=>"000001000",
  59302=>"111111111",
  59303=>"111011011",
  59304=>"111011000",
  59305=>"000000000",
  59306=>"000001111",
  59307=>"000000000",
  59308=>"000110111",
  59309=>"000001001",
  59310=>"100101101",
  59311=>"010001000",
  59312=>"111111111",
  59313=>"111111110",
  59314=>"111111111",
  59315=>"111111111",
  59316=>"001000001",
  59317=>"101101111",
  59318=>"101111000",
  59319=>"000011110",
  59320=>"111111110",
  59321=>"000000000",
  59322=>"011111111",
  59323=>"111000100",
  59324=>"000011111",
  59325=>"000000111",
  59326=>"000000000",
  59327=>"001001000",
  59328=>"000000000",
  59329=>"100111111",
  59330=>"100000000",
  59331=>"000000000",
  59332=>"000000111",
  59333=>"110111011",
  59334=>"111111000",
  59335=>"000100000",
  59336=>"100100100",
  59337=>"111111111",
  59338=>"000000000",
  59339=>"111111111",
  59340=>"111011011",
  59341=>"000000000",
  59342=>"000011001",
  59343=>"011000000",
  59344=>"000000000",
  59345=>"110111111",
  59346=>"100100110",
  59347=>"001000001",
  59348=>"001101100",
  59349=>"111111111",
  59350=>"000000000",
  59351=>"111100111",
  59352=>"111101000",
  59353=>"011011110",
  59354=>"110110000",
  59355=>"100111000",
  59356=>"000000010",
  59357=>"111111011",
  59358=>"111010111",
  59359=>"101111111",
  59360=>"111000011",
  59361=>"000011011",
  59362=>"000000111",
  59363=>"111111001",
  59364=>"000010010",
  59365=>"111111111",
  59366=>"111101111",
  59367=>"000000000",
  59368=>"111111111",
  59369=>"111110111",
  59370=>"111100111",
  59371=>"110011011",
  59372=>"000000000",
  59373=>"110110111",
  59374=>"011111111",
  59375=>"000100111",
  59376=>"000000000",
  59377=>"100000101",
  59378=>"000000001",
  59379=>"000000000",
  59380=>"000101111",
  59381=>"111111111",
  59382=>"110111111",
  59383=>"110110100",
  59384=>"111111111",
  59385=>"000100111",
  59386=>"000000000",
  59387=>"000111011",
  59388=>"000000011",
  59389=>"110100111",
  59390=>"111011000",
  59391=>"000000111",
  59392=>"011011000",
  59393=>"110111101",
  59394=>"111111111",
  59395=>"001000001",
  59396=>"100110111",
  59397=>"111111111",
  59398=>"000010111",
  59399=>"111111111",
  59400=>"101000000",
  59401=>"110110111",
  59402=>"111111110",
  59403=>"000000000",
  59404=>"110110110",
  59405=>"000000001",
  59406=>"100100111",
  59407=>"111111000",
  59408=>"011011011",
  59409=>"000111001",
  59410=>"000000111",
  59411=>"000000110",
  59412=>"000000000",
  59413=>"111111000",
  59414=>"000100100",
  59415=>"000111100",
  59416=>"000000100",
  59417=>"000111111",
  59418=>"111111111",
  59419=>"111111111",
  59420=>"111101100",
  59421=>"000000000",
  59422=>"011011010",
  59423=>"111011000",
  59424=>"111111010",
  59425=>"111010110",
  59426=>"000000100",
  59427=>"011000000",
  59428=>"000000110",
  59429=>"011001000",
  59430=>"000001000",
  59431=>"111000000",
  59432=>"111111111",
  59433=>"110110110",
  59434=>"000000000",
  59435=>"000000010",
  59436=>"000000011",
  59437=>"000111000",
  59438=>"000000001",
  59439=>"010111111",
  59440=>"000000010",
  59441=>"000000101",
  59442=>"111111111",
  59443=>"101111111",
  59444=>"111111101",
  59445=>"111111111",
  59446=>"001000000",
  59447=>"111100100",
  59448=>"111110111",
  59449=>"101111100",
  59450=>"111111111",
  59451=>"111001001",
  59452=>"000000001",
  59453=>"111101100",
  59454=>"111100110",
  59455=>"111101101",
  59456=>"000001111",
  59457=>"000110110",
  59458=>"000000010",
  59459=>"111000000",
  59460=>"111000000",
  59461=>"000000100",
  59462=>"000000000",
  59463=>"000110111",
  59464=>"011111010",
  59465=>"000000000",
  59466=>"000001111",
  59467=>"001000110",
  59468=>"000000000",
  59469=>"110111111",
  59470=>"111100110",
  59471=>"000000011",
  59472=>"110111111",
  59473=>"010111111",
  59474=>"111000000",
  59475=>"011001001",
  59476=>"011111111",
  59477=>"100111111",
  59478=>"111100100",
  59479=>"100111111",
  59480=>"001001001",
  59481=>"101000111",
  59482=>"111110101",
  59483=>"100000000",
  59484=>"000001000",
  59485=>"111001001",
  59486=>"110000000",
  59487=>"111011111",
  59488=>"000000111",
  59489=>"111000000",
  59490=>"110100100",
  59491=>"111111111",
  59492=>"101000000",
  59493=>"000001001",
  59494=>"011001100",
  59495=>"010111111",
  59496=>"010000000",
  59497=>"000000000",
  59498=>"000110110",
  59499=>"011011000",
  59500=>"111111111",
  59501=>"100100000",
  59502=>"111101111",
  59503=>"100111111",
  59504=>"011001011",
  59505=>"111111101",
  59506=>"001111011",
  59507=>"111000011",
  59508=>"110111111",
  59509=>"111100000",
  59510=>"100000000",
  59511=>"010111111",
  59512=>"000000000",
  59513=>"011000000",
  59514=>"001000000",
  59515=>"000100100",
  59516=>"000100111",
  59517=>"000000111",
  59518=>"000000000",
  59519=>"000000000",
  59520=>"011111100",
  59521=>"000000100",
  59522=>"110000110",
  59523=>"000100000",
  59524=>"001001111",
  59525=>"000000000",
  59526=>"000000010",
  59527=>"101101101",
  59528=>"000000000",
  59529=>"000000000",
  59530=>"111011011",
  59531=>"111111000",
  59532=>"000101111",
  59533=>"111000101",
  59534=>"011011001",
  59535=>"000000000",
  59536=>"001000001",
  59537=>"000000000",
  59538=>"011101111",
  59539=>"111111111",
  59540=>"000100111",
  59541=>"010000000",
  59542=>"010111111",
  59543=>"111000000",
  59544=>"000000111",
  59545=>"110111111",
  59546=>"111000000",
  59547=>"001111111",
  59548=>"111111110",
  59549=>"111100110",
  59550=>"111111110",
  59551=>"000100111",
  59552=>"100000000",
  59553=>"111111101",
  59554=>"001001000",
  59555=>"000000000",
  59556=>"111001001",
  59557=>"111111101",
  59558=>"111111111",
  59559=>"001001001",
  59560=>"000110111",
  59561=>"101000000",
  59562=>"000000010",
  59563=>"000001111",
  59564=>"000000000",
  59565=>"011001011",
  59566=>"001000101",
  59567=>"001011101",
  59568=>"000000011",
  59569=>"111011001",
  59570=>"001111000",
  59571=>"111111000",
  59572=>"000011001",
  59573=>"001000001",
  59574=>"000000001",
  59575=>"111111110",
  59576=>"111001111",
  59577=>"000000000",
  59578=>"110111111",
  59579=>"011011111",
  59580=>"111111111",
  59581=>"111111000",
  59582=>"000100000",
  59583=>"000000000",
  59584=>"111001101",
  59585=>"111100100",
  59586=>"111111000",
  59587=>"111111111",
  59588=>"010111111",
  59589=>"001000000",
  59590=>"111110110",
  59591=>"001001000",
  59592=>"010110111",
  59593=>"000000000",
  59594=>"000000000",
  59595=>"000000000",
  59596=>"001000100",
  59597=>"111111111",
  59598=>"111111000",
  59599=>"000111000",
  59600=>"100001111",
  59601=>"110110111",
  59602=>"111111111",
  59603=>"000000000",
  59604=>"000001111",
  59605=>"000000000",
  59606=>"000000000",
  59607=>"000000001",
  59608=>"000100111",
  59609=>"111000000",
  59610=>"111110111",
  59611=>"011011011",
  59612=>"111111101",
  59613=>"000000000",
  59614=>"111111111",
  59615=>"011111100",
  59616=>"000000000",
  59617=>"000110110",
  59618=>"010111011",
  59619=>"000000000",
  59620=>"000000000",
  59621=>"011001111",
  59622=>"110000000",
  59623=>"111111000",
  59624=>"111111000",
  59625=>"000000000",
  59626=>"111111000",
  59627=>"000000100",
  59628=>"000001011",
  59629=>"100000111",
  59630=>"111111111",
  59631=>"000000000",
  59632=>"011111111",
  59633=>"100100111",
  59634=>"000000000",
  59635=>"000000000",
  59636=>"111110110",
  59637=>"110000000",
  59638=>"101000000",
  59639=>"111010000",
  59640=>"000000000",
  59641=>"000010000",
  59642=>"111101101",
  59643=>"111111111",
  59644=>"101111011",
  59645=>"000000011",
  59646=>"000000000",
  59647=>"110110100",
  59648=>"111111100",
  59649=>"111000000",
  59650=>"111111111",
  59651=>"101011011",
  59652=>"111100000",
  59653=>"111101111",
  59654=>"111001111",
  59655=>"111101111",
  59656=>"011100000",
  59657=>"111011000",
  59658=>"000000000",
  59659=>"111111111",
  59660=>"001001000",
  59661=>"010011111",
  59662=>"000000111",
  59663=>"110000000",
  59664=>"000111110",
  59665=>"111100100",
  59666=>"111000111",
  59667=>"111101101",
  59668=>"000000100",
  59669=>"011111111",
  59670=>"001001001",
  59671=>"100000110",
  59672=>"111111100",
  59673=>"000000001",
  59674=>"000000001",
  59675=>"000000000",
  59676=>"111111010",
  59677=>"111111011",
  59678=>"010111111",
  59679=>"111001000",
  59680=>"100000001",
  59681=>"111000000",
  59682=>"110110000",
  59683=>"110001000",
  59684=>"000000000",
  59685=>"000000001",
  59686=>"000011001",
  59687=>"111011011",
  59688=>"101000001",
  59689=>"010111111",
  59690=>"000000000",
  59691=>"000000111",
  59692=>"000000000",
  59693=>"101111001",
  59694=>"111000000",
  59695=>"000000001",
  59696=>"111110110",
  59697=>"100110111",
  59698=>"001111111",
  59699=>"100110111",
  59700=>"100100000",
  59701=>"111111100",
  59702=>"111101000",
  59703=>"000001001",
  59704=>"111110111",
  59705=>"100000001",
  59706=>"000000000",
  59707=>"111111101",
  59708=>"111100100",
  59709=>"000001111",
  59710=>"001101111",
  59711=>"000000010",
  59712=>"111000111",
  59713=>"111111111",
  59714=>"000000110",
  59715=>"001011011",
  59716=>"000101111",
  59717=>"111111110",
  59718=>"010011110",
  59719=>"000000111",
  59720=>"100000000",
  59721=>"011000000",
  59722=>"010001000",
  59723=>"001011011",
  59724=>"100000000",
  59725=>"111010000",
  59726=>"111010011",
  59727=>"000000000",
  59728=>"000000100",
  59729=>"011011111",
  59730=>"111111111",
  59731=>"000100000",
  59732=>"111111110",
  59733=>"001011011",
  59734=>"111111111",
  59735=>"100001001",
  59736=>"011001111",
  59737=>"100000000",
  59738=>"001001111",
  59739=>"111111111",
  59740=>"110000100",
  59741=>"000000000",
  59742=>"011010000",
  59743=>"111111110",
  59744=>"111111000",
  59745=>"111111011",
  59746=>"111111011",
  59747=>"011000000",
  59748=>"000000001",
  59749=>"100100000",
  59750=>"100100110",
  59751=>"011011010",
  59752=>"000000001",
  59753=>"000000000",
  59754=>"001000000",
  59755=>"000000000",
  59756=>"111011000",
  59757=>"000011111",
  59758=>"000010010",
  59759=>"001001101",
  59760=>"111100100",
  59761=>"000000111",
  59762=>"000100111",
  59763=>"100100000",
  59764=>"111111111",
  59765=>"100111111",
  59766=>"111001011",
  59767=>"100000000",
  59768=>"000000000",
  59769=>"100000000",
  59770=>"101100000",
  59771=>"111101011",
  59772=>"111111100",
  59773=>"111110110",
  59774=>"000100110",
  59775=>"000000000",
  59776=>"001001001",
  59777=>"011001100",
  59778=>"100000000",
  59779=>"000000110",
  59780=>"000100111",
  59781=>"111111111",
  59782=>"000000000",
  59783=>"001001001",
  59784=>"100100000",
  59785=>"111111111",
  59786=>"000110010",
  59787=>"010111010",
  59788=>"101000000",
  59789=>"111111000",
  59790=>"111111000",
  59791=>"010011111",
  59792=>"000101000",
  59793=>"011111111",
  59794=>"001001001",
  59795=>"111011001",
  59796=>"001010111",
  59797=>"010000000",
  59798=>"110111010",
  59799=>"011011011",
  59800=>"001000000",
  59801=>"111001000",
  59802=>"111111111",
  59803=>"000101101",
  59804=>"111111000",
  59805=>"001000000",
  59806=>"000000000",
  59807=>"111110110",
  59808=>"100000000",
  59809=>"011011011",
  59810=>"001000101",
  59811=>"100000011",
  59812=>"000000111",
  59813=>"000000111",
  59814=>"000000000",
  59815=>"111111111",
  59816=>"111011001",
  59817=>"000000000",
  59818=>"011001111",
  59819=>"000000110",
  59820=>"111111000",
  59821=>"000100111",
  59822=>"110110011",
  59823=>"101100000",
  59824=>"111100100",
  59825=>"101101111",
  59826=>"000110000",
  59827=>"000000000",
  59828=>"011100100",
  59829=>"000000110",
  59830=>"000000000",
  59831=>"010011111",
  59832=>"000001111",
  59833=>"001001101",
  59834=>"111110110",
  59835=>"000000001",
  59836=>"000000000",
  59837=>"111110111",
  59838=>"011001000",
  59839=>"000001001",
  59840=>"000000101",
  59841=>"000000000",
  59842=>"000000000",
  59843=>"000000000",
  59844=>"111110000",
  59845=>"101000111",
  59846=>"111111110",
  59847=>"111001001",
  59848=>"001000000",
  59849=>"111110110",
  59850=>"000000101",
  59851=>"000000000",
  59852=>"001010011",
  59853=>"011011000",
  59854=>"011111111",
  59855=>"000000110",
  59856=>"000000000",
  59857=>"111100000",
  59858=>"001000000",
  59859=>"001001111",
  59860=>"101011011",
  59861=>"000000110",
  59862=>"110010000",
  59863=>"111111111",
  59864=>"000100111",
  59865=>"011010000",
  59866=>"000100100",
  59867=>"111101001",
  59868=>"000000100",
  59869=>"001001111",
  59870=>"111011000",
  59871=>"000010011",
  59872=>"000000000",
  59873=>"010000111",
  59874=>"000001001",
  59875=>"111100100",
  59876=>"111001001",
  59877=>"111111000",
  59878=>"011011011",
  59879=>"110110000",
  59880=>"111000000",
  59881=>"111111101",
  59882=>"000010011",
  59883=>"000001000",
  59884=>"010111111",
  59885=>"001111111",
  59886=>"100100100",
  59887=>"010110110",
  59888=>"000000101",
  59889=>"000000001",
  59890=>"001000000",
  59891=>"000000011",
  59892=>"111111111",
  59893=>"011011000",
  59894=>"111110000",
  59895=>"100001001",
  59896=>"000000000",
  59897=>"011110110",
  59898=>"100000000",
  59899=>"111111111",
  59900=>"100111111",
  59901=>"000010000",
  59902=>"011100100",
  59903=>"001111111",
  59904=>"100100100",
  59905=>"000000000",
  59906=>"000000000",
  59907=>"000000000",
  59908=>"000000111",
  59909=>"000000000",
  59910=>"000000000",
  59911=>"111101101",
  59912=>"111111111",
  59913=>"000010000",
  59914=>"000000000",
  59915=>"000000000",
  59916=>"000000100",
  59917=>"000000000",
  59918=>"000000000",
  59919=>"000000100",
  59920=>"111111001",
  59921=>"000001111",
  59922=>"000011101",
  59923=>"111011000",
  59924=>"000000000",
  59925=>"000000010",
  59926=>"000000000",
  59927=>"001011001",
  59928=>"000000000",
  59929=>"111111111",
  59930=>"111000000",
  59931=>"011111100",
  59932=>"110110100",
  59933=>"000000000",
  59934=>"000000001",
  59935=>"000110111",
  59936=>"010000111",
  59937=>"111111111",
  59938=>"000100110",
  59939=>"000001001",
  59940=>"111111110",
  59941=>"111111111",
  59942=>"110110011",
  59943=>"000001111",
  59944=>"100000000",
  59945=>"000000000",
  59946=>"000000000",
  59947=>"000000000",
  59948=>"111111011",
  59949=>"100101001",
  59950=>"111111111",
  59951=>"000100111",
  59952=>"000011111",
  59953=>"111111011",
  59954=>"000000011",
  59955=>"100000100",
  59956=>"110111111",
  59957=>"000000000",
  59958=>"000000000",
  59959=>"000000110",
  59960=>"000000000",
  59961=>"000000000",
  59962=>"000000000",
  59963=>"111111011",
  59964=>"100000000",
  59965=>"111110110",
  59966=>"000110110",
  59967=>"000000000",
  59968=>"000000000",
  59969=>"111111111",
  59970=>"000000000",
  59971=>"110111111",
  59972=>"000000000",
  59973=>"000000000",
  59974=>"111000010",
  59975=>"011111111",
  59976=>"001000111",
  59977=>"000000000",
  59978=>"111111111",
  59979=>"000000000",
  59980=>"011111111",
  59981=>"010110111",
  59982=>"010001000",
  59983=>"111110000",
  59984=>"000000000",
  59985=>"000000111",
  59986=>"000000000",
  59987=>"111100000",
  59988=>"001000000",
  59989=>"000001100",
  59990=>"000111111",
  59991=>"111111111",
  59992=>"001100100",
  59993=>"100000001",
  59994=>"000000101",
  59995=>"111100100",
  59996=>"001000110",
  59997=>"100110111",
  59998=>"000000000",
  59999=>"111111111",
  60000=>"111111111",
  60001=>"000000000",
  60002=>"000100000",
  60003=>"000011000",
  60004=>"111111000",
  60005=>"001101111",
  60006=>"000000110",
  60007=>"000001001",
  60008=>"111111111",
  60009=>"111111011",
  60010=>"010000000",
  60011=>"100000000",
  60012=>"000100100",
  60013=>"101111000",
  60014=>"111111111",
  60015=>"111111111",
  60016=>"000111111",
  60017=>"100110111",
  60018=>"111111111",
  60019=>"000000000",
  60020=>"000000000",
  60021=>"111110110",
  60022=>"000000000",
  60023=>"000000000",
  60024=>"000000010",
  60025=>"101111111",
  60026=>"000000000",
  60027=>"000000000",
  60028=>"000000000",
  60029=>"000111100",
  60030=>"011111101",
  60031=>"000010111",
  60032=>"001001000",
  60033=>"000000000",
  60034=>"110111111",
  60035=>"011011111",
  60036=>"111110000",
  60037=>"101000100",
  60038=>"111111110",
  60039=>"111100100",
  60040=>"000001000",
  60041=>"111111111",
  60042=>"001000000",
  60043=>"100100100",
  60044=>"000000000",
  60045=>"000000100",
  60046=>"111011000",
  60047=>"110111111",
  60048=>"000000000",
  60049=>"000001011",
  60050=>"100110111",
  60051=>"111111111",
  60052=>"111111011",
  60053=>"111110100",
  60054=>"111000000",
  60055=>"000000100",
  60056=>"000000000",
  60057=>"110111111",
  60058=>"111000000",
  60059=>"001000000",
  60060=>"011101111",
  60061=>"000000000",
  60062=>"000100100",
  60063=>"111111111",
  60064=>"111111000",
  60065=>"111001000",
  60066=>"000100111",
  60067=>"000001011",
  60068=>"000000000",
  60069=>"011111111",
  60070=>"000110111",
  60071=>"110100110",
  60072=>"111100111",
  60073=>"000000010",
  60074=>"000111111",
  60075=>"000000111",
  60076=>"000001111",
  60077=>"111111111",
  60078=>"111111110",
  60079=>"000111111",
  60080=>"111111111",
  60081=>"110111111",
  60082=>"110111111",
  60083=>"000111111",
  60084=>"111111000",
  60085=>"111111111",
  60086=>"000100100",
  60087=>"000000001",
  60088=>"001000000",
  60089=>"011010000",
  60090=>"000001000",
  60091=>"100000000",
  60092=>"110110111",
  60093=>"111111110",
  60094=>"111111111",
  60095=>"000001101",
  60096=>"111111111",
  60097=>"000000000",
  60098=>"111111111",
  60099=>"000000100",
  60100=>"000000111",
  60101=>"111111000",
  60102=>"011101101",
  60103=>"111111111",
  60104=>"000000000",
  60105=>"111111111",
  60106=>"011000000",
  60107=>"011111111",
  60108=>"111100111",
  60109=>"111100000",
  60110=>"000000000",
  60111=>"110111000",
  60112=>"001001011",
  60113=>"000111111",
  60114=>"000110000",
  60115=>"001001001",
  60116=>"000000000",
  60117=>"000000001",
  60118=>"100000000",
  60119=>"100110110",
  60120=>"000000000",
  60121=>"001100100",
  60122=>"000000000",
  60123=>"100100100",
  60124=>"111111011",
  60125=>"110111110",
  60126=>"000000010",
  60127=>"000001111",
  60128=>"000000000",
  60129=>"110111001",
  60130=>"000000000",
  60131=>"111111100",
  60132=>"111011111",
  60133=>"110110110",
  60134=>"111100000",
  60135=>"000000001",
  60136=>"111111111",
  60137=>"011001111",
  60138=>"011111111",
  60139=>"100111111",
  60140=>"111111000",
  60141=>"000000000",
  60142=>"110010000",
  60143=>"001111111",
  60144=>"011000000",
  60145=>"011011011",
  60146=>"010100100",
  60147=>"000100111",
  60148=>"111111111",
  60149=>"011111111",
  60150=>"111001001",
  60151=>"100100111",
  60152=>"111111111",
  60153=>"111111111",
  60154=>"111111111",
  60155=>"000000000",
  60156=>"000000011",
  60157=>"100100110",
  60158=>"011000000",
  60159=>"001101001",
  60160=>"000000000",
  60161=>"101000000",
  60162=>"000000000",
  60163=>"100110100",
  60164=>"000110100",
  60165=>"000000000",
  60166=>"111111111",
  60167=>"000110111",
  60168=>"000000000",
  60169=>"000000000",
  60170=>"000000000",
  60171=>"000110110",
  60172=>"100000110",
  60173=>"000001001",
  60174=>"111111111",
  60175=>"000100100",
  60176=>"011010000",
  60177=>"000000000",
  60178=>"111101011",
  60179=>"000000000",
  60180=>"000000000",
  60181=>"111101000",
  60182=>"001001001",
  60183=>"111111110",
  60184=>"110010010",
  60185=>"000001011",
  60186=>"000000111",
  60187=>"001100111",
  60188=>"000000111",
  60189=>"000000000",
  60190=>"000011000",
  60191=>"111110100",
  60192=>"000000000",
  60193=>"000000000",
  60194=>"010011010",
  60195=>"111111111",
  60196=>"111101000",
  60197=>"001011111",
  60198=>"110110011",
  60199=>"111101111",
  60200=>"111111111",
  60201=>"000000000",
  60202=>"110110111",
  60203=>"110111110",
  60204=>"001001111",
  60205=>"110011111",
  60206=>"000000100",
  60207=>"000000000",
  60208=>"111111111",
  60209=>"100000100",
  60210=>"111011111",
  60211=>"011111011",
  60212=>"111001000",
  60213=>"111111000",
  60214=>"111111000",
  60215=>"000000100",
  60216=>"100000000",
  60217=>"100000001",
  60218=>"111111111",
  60219=>"110000000",
  60220=>"111111101",
  60221=>"111111101",
  60222=>"011001001",
  60223=>"011011000",
  60224=>"000000110",
  60225=>"111111111",
  60226=>"111111111",
  60227=>"000000000",
  60228=>"100111110",
  60229=>"000000111",
  60230=>"010111111",
  60231=>"001000100",
  60232=>"111011011",
  60233=>"111111111",
  60234=>"000000101",
  60235=>"111111111",
  60236=>"000010000",
  60237=>"010111111",
  60238=>"011001111",
  60239=>"100000000",
  60240=>"100100100",
  60241=>"000110111",
  60242=>"111111111",
  60243=>"100001001",
  60244=>"101000111",
  60245=>"000011011",
  60246=>"000010111",
  60247=>"111111111",
  60248=>"000000000",
  60249=>"111111111",
  60250=>"111111011",
  60251=>"001001011",
  60252=>"000000000",
  60253=>"001011011",
  60254=>"000000000",
  60255=>"101011111",
  60256=>"000000000",
  60257=>"010001000",
  60258=>"100100000",
  60259=>"111111111",
  60260=>"111111000",
  60261=>"100000111",
  60262=>"000000000",
  60263=>"000110111",
  60264=>"111110110",
  60265=>"111111111",
  60266=>"000000110",
  60267=>"110111011",
  60268=>"011000100",
  60269=>"000101100",
  60270=>"000000000",
  60271=>"111111100",
  60272=>"111111111",
  60273=>"111011000",
  60274=>"001111111",
  60275=>"000000110",
  60276=>"111111111",
  60277=>"000000100",
  60278=>"000000100",
  60279=>"000110111",
  60280=>"000000100",
  60281=>"111111110",
  60282=>"111000110",
  60283=>"111000000",
  60284=>"111111111",
  60285=>"000111111",
  60286=>"011001000",
  60287=>"111111111",
  60288=>"110110110",
  60289=>"001001001",
  60290=>"111100100",
  60291=>"011011111",
  60292=>"101111101",
  60293=>"000000001",
  60294=>"101101000",
  60295=>"101001001",
  60296=>"000000000",
  60297=>"011111110",
  60298=>"110100110",
  60299=>"000000011",
  60300=>"100001001",
  60301=>"000110000",
  60302=>"000011101",
  60303=>"000000000",
  60304=>"110011111",
  60305=>"001000001",
  60306=>"000000010",
  60307=>"111111110",
  60308=>"000000000",
  60309=>"011011011",
  60310=>"111111101",
  60311=>"011011001",
  60312=>"011111110",
  60313=>"010110111",
  60314=>"101001101",
  60315=>"001111111",
  60316=>"000000000",
  60317=>"000101111",
  60318=>"000000000",
  60319=>"111111000",
  60320=>"111111111",
  60321=>"011001001",
  60322=>"100100000",
  60323=>"111111111",
  60324=>"100000100",
  60325=>"111111111",
  60326=>"000001101",
  60327=>"111111111",
  60328=>"000001111",
  60329=>"111110110",
  60330=>"000000000",
  60331=>"000000000",
  60332=>"000000000",
  60333=>"111111001",
  60334=>"000000001",
  60335=>"000000000",
  60336=>"001000111",
  60337=>"000000000",
  60338=>"000000000",
  60339=>"110000000",
  60340=>"001011001",
  60341=>"111111111",
  60342=>"111111111",
  60343=>"000000111",
  60344=>"111111010",
  60345=>"111111111",
  60346=>"111111001",
  60347=>"100100000",
  60348=>"111000000",
  60349=>"111111111",
  60350=>"111100110",
  60351=>"111111011",
  60352=>"111110000",
  60353=>"000000111",
  60354=>"000000000",
  60355=>"111100101",
  60356=>"000000000",
  60357=>"100100000",
  60358=>"111111111",
  60359=>"100000000",
  60360=>"001100110",
  60361=>"111111000",
  60362=>"000000110",
  60363=>"000000000",
  60364=>"111000000",
  60365=>"111111010",
  60366=>"000110110",
  60367=>"010000000",
  60368=>"011011010",
  60369=>"100110110",
  60370=>"111111111",
  60371=>"111011000",
  60372=>"100100101",
  60373=>"111111101",
  60374=>"110000100",
  60375=>"001001011",
  60376=>"111000000",
  60377=>"011001001",
  60378=>"001001001",
  60379=>"000111001",
  60380=>"111110110",
  60381=>"001000111",
  60382=>"100110111",
  60383=>"111110100",
  60384=>"111010000",
  60385=>"000000000",
  60386=>"111000000",
  60387=>"100000000",
  60388=>"010111111",
  60389=>"011001001",
  60390=>"111100100",
  60391=>"111011001",
  60392=>"001000000",
  60393=>"111000111",
  60394=>"101100100",
  60395=>"010111000",
  60396=>"110111111",
  60397=>"000110100",
  60398=>"011011111",
  60399=>"000111111",
  60400=>"001001000",
  60401=>"000000000",
  60402=>"111111000",
  60403=>"000110110",
  60404=>"000000000",
  60405=>"000110111",
  60406=>"011011000",
  60407=>"110111111",
  60408=>"100000000",
  60409=>"000010100",
  60410=>"000000000",
  60411=>"000000000",
  60412=>"000110011",
  60413=>"111111111",
  60414=>"001001100",
  60415=>"111011000",
  60416=>"000001011",
  60417=>"000001100",
  60418=>"111000111",
  60419=>"000000000",
  60420=>"111111111",
  60421=>"110100101",
  60422=>"001001111",
  60423=>"111111111",
  60424=>"000000000",
  60425=>"100000000",
  60426=>"000000111",
  60427=>"010111111",
  60428=>"110100101",
  60429=>"000001001",
  60430=>"110100000",
  60431=>"000000000",
  60432=>"110110000",
  60433=>"111111111",
  60434=>"011100100",
  60435=>"000000100",
  60436=>"101101110",
  60437=>"011000010",
  60438=>"101001000",
  60439=>"111111011",
  60440=>"110110110",
  60441=>"001001001",
  60442=>"111000111",
  60443=>"001001000",
  60444=>"000000000",
  60445=>"000110111",
  60446=>"111001001",
  60447=>"111111111",
  60448=>"000000001",
  60449=>"110110010",
  60450=>"110111100",
  60451=>"010000111",
  60452=>"000110110",
  60453=>"000001111",
  60454=>"111111011",
  60455=>"000000000",
  60456=>"001001101",
  60457=>"100101101",
  60458=>"000000010",
  60459=>"000000110",
  60460=>"110000000",
  60461=>"011011000",
  60462=>"000000001",
  60463=>"000111100",
  60464=>"100100101",
  60465=>"000000000",
  60466=>"100111111",
  60467=>"100000010",
  60468=>"000000000",
  60469=>"100011001",
  60470=>"001000100",
  60471=>"000100000",
  60472=>"001111111",
  60473=>"110111111",
  60474=>"000011011",
  60475=>"000000000",
  60476=>"001000001",
  60477=>"111011111",
  60478=>"000000100",
  60479=>"000001111",
  60480=>"010000110",
  60481=>"000001000",
  60482=>"010111111",
  60483=>"110010000",
  60484=>"000100110",
  60485=>"000000101",
  60486=>"111110110",
  60487=>"111100000",
  60488=>"110111011",
  60489=>"000010010",
  60490=>"101101111",
  60491=>"000000111",
  60492=>"000000000",
  60493=>"111111101",
  60494=>"100100000",
  60495=>"101000111",
  60496=>"001001000",
  60497=>"111111111",
  60498=>"110000110",
  60499=>"000000000",
  60500=>"000000000",
  60501=>"101101111",
  60502=>"001011011",
  60503=>"000000000",
  60504=>"100000100",
  60505=>"101000111",
  60506=>"000000100",
  60507=>"111010010",
  60508=>"111111111",
  60509=>"000001111",
  60510=>"001111111",
  60511=>"001111111",
  60512=>"000001101",
  60513=>"000000000",
  60514=>"000001111",
  60515=>"100101000",
  60516=>"111010000",
  60517=>"000000110",
  60518=>"101101001",
  60519=>"000000101",
  60520=>"011111111",
  60521=>"001001001",
  60522=>"000000000",
  60523=>"000000000",
  60524=>"000001111",
  60525=>"000000000",
  60526=>"111111101",
  60527=>"011100110",
  60528=>"001001000",
  60529=>"100001000",
  60530=>"100100101",
  60531=>"000001000",
  60532=>"000111110",
  60533=>"110110110",
  60534=>"001001000",
  60535=>"000110000",
  60536=>"111111110",
  60537=>"010110111",
  60538=>"011000000",
  60539=>"111111111",
  60540=>"110110000",
  60541=>"110110110",
  60542=>"110111111",
  60543=>"111111000",
  60544=>"010000010",
  60545=>"011010000",
  60546=>"001000111",
  60547=>"101000001",
  60548=>"000000000",
  60549=>"111000000",
  60550=>"011010111",
  60551=>"011010010",
  60552=>"000000010",
  60553=>"000000000",
  60554=>"110110110",
  60555=>"101101111",
  60556=>"110110000",
  60557=>"001001111",
  60558=>"101000000",
  60559=>"000110111",
  60560=>"101110100",
  60561=>"101001111",
  60562=>"001011111",
  60563=>"110110110",
  60564=>"000000001",
  60565=>"111110111",
  60566=>"001000100",
  60567=>"111110000",
  60568=>"101001111",
  60569=>"000001111",
  60570=>"011111001",
  60571=>"000010000",
  60572=>"001111111",
  60573=>"000000110",
  60574=>"000000000",
  60575=>"000000100",
  60576=>"000001000",
  60577=>"000110110",
  60578=>"001101001",
  60579=>"011011000",
  60580=>"000000000",
  60581=>"111111000",
  60582=>"011111111",
  60583=>"011111000",
  60584=>"111111011",
  60585=>"001000000",
  60586=>"000111111",
  60587=>"101000000",
  60588=>"000100000",
  60589=>"001001101",
  60590=>"111111111",
  60591=>"000001100",
  60592=>"000000001",
  60593=>"100110110",
  60594=>"111111010",
  60595=>"111111010",
  60596=>"010010110",
  60597=>"111010010",
  60598=>"101111111",
  60599=>"010100000",
  60600=>"111101111",
  60601=>"100000110",
  60602=>"011000010",
  60603=>"110110111",
  60604=>"000000111",
  60605=>"101101100",
  60606=>"000000111",
  60607=>"000001000",
  60608=>"000100000",
  60609=>"111100111",
  60610=>"110110110",
  60611=>"100101111",
  60612=>"000000110",
  60613=>"110100000",
  60614=>"000010110",
  60615=>"010111011",
  60616=>"000001010",
  60617=>"000000111",
  60618=>"101000000",
  60619=>"000000000",
  60620=>"100100100",
  60621=>"010110111",
  60622=>"000111110",
  60623=>"000000100",
  60624=>"001001001",
  60625=>"111110010",
  60626=>"111111000",
  60627=>"110010000",
  60628=>"000100001",
  60629=>"110110111",
  60630=>"000000000",
  60631=>"111111111",
  60632=>"101111111",
  60633=>"111101111",
  60634=>"100000100",
  60635=>"011111111",
  60636=>"001111111",
  60637=>"111111001",
  60638=>"000000001",
  60639=>"000001001",
  60640=>"000000000",
  60641=>"010010000",
  60642=>"111111111",
  60643=>"011111111",
  60644=>"001101001",
  60645=>"110100100",
  60646=>"101111111",
  60647=>"111111111",
  60648=>"111110111",
  60649=>"000001111",
  60650=>"000000110",
  60651=>"000000110",
  60652=>"111100000",
  60653=>"000000000",
  60654=>"000110111",
  60655=>"000110111",
  60656=>"000110111",
  60657=>"001001001",
  60658=>"111011001",
  60659=>"100000100",
  60660=>"110111111",
  60661=>"100110110",
  60662=>"101100100",
  60663=>"000000111",
  60664=>"010000000",
  60665=>"010111111",
  60666=>"101101011",
  60667=>"111111000",
  60668=>"110110001",
  60669=>"001001111",
  60670=>"111000100",
  60671=>"111101001",
  60672=>"101101100",
  60673=>"100000001",
  60674=>"110110000",
  60675=>"110110000",
  60676=>"001111110",
  60677=>"001000100",
  60678=>"111111111",
  60679=>"000000010",
  60680=>"000010111",
  60681=>"000000000",
  60682=>"111111110",
  60683=>"111101111",
  60684=>"111001001",
  60685=>"000000101",
  60686=>"110111000",
  60687=>"111111010",
  60688=>"000000000",
  60689=>"111001001",
  60690=>"001101101",
  60691=>"000101111",
  60692=>"111000000",
  60693=>"000101111",
  60694=>"000010001",
  60695=>"111111101",
  60696=>"111111001",
  60697=>"001000111",
  60698=>"000000101",
  60699=>"010000111",
  60700=>"001011100",
  60701=>"011010111",
  60702=>"001001111",
  60703=>"000001000",
  60704=>"000000001",
  60705=>"111111111",
  60706=>"111111111",
  60707=>"001111001",
  60708=>"100100100",
  60709=>"111001000",
  60710=>"000010001",
  60711=>"000000101",
  60712=>"000000111",
  60713=>"111110000",
  60714=>"000000000",
  60715=>"001101101",
  60716=>"111010000",
  60717=>"001001000",
  60718=>"000000000",
  60719=>"100100000",
  60720=>"001101001",
  60721=>"010000000",
  60722=>"000000111",
  60723=>"100111111",
  60724=>"000000111",
  60725=>"111111011",
  60726=>"000000100",
  60727=>"001000000",
  60728=>"000001000",
  60729=>"000000000",
  60730=>"000000111",
  60731=>"010011001",
  60732=>"111111111",
  60733=>"001001001",
  60734=>"110111111",
  60735=>"000111110",
  60736=>"100100000",
  60737=>"110110000",
  60738=>"110111110",
  60739=>"111111111",
  60740=>"000000010",
  60741=>"110111111",
  60742=>"111111111",
  60743=>"001001111",
  60744=>"000000000",
  60745=>"000110010",
  60746=>"000101101",
  60747=>"011111011",
  60748=>"000000000",
  60749=>"000100111",
  60750=>"101001111",
  60751=>"000000000",
  60752=>"000001000",
  60753=>"011101111",
  60754=>"001000000",
  60755=>"000001101",
  60756=>"001001111",
  60757=>"011011001",
  60758=>"011001111",
  60759=>"101100000",
  60760=>"000111011",
  60761=>"111111111",
  60762=>"000000000",
  60763=>"000100101",
  60764=>"000000011",
  60765=>"000000000",
  60766=>"000100000",
  60767=>"111111111",
  60768=>"000000001",
  60769=>"101101000",
  60770=>"110111101",
  60771=>"000010000",
  60772=>"000111010",
  60773=>"000001000",
  60774=>"000000100",
  60775=>"000000101",
  60776=>"100100111",
  60777=>"001001111",
  60778=>"001001001",
  60779=>"000100101",
  60780=>"111011001",
  60781=>"111011011",
  60782=>"110110010",
  60783=>"000000000",
  60784=>"110110111",
  60785=>"010011000",
  60786=>"001000001",
  60787=>"011111011",
  60788=>"110011001",
  60789=>"010111111",
  60790=>"000001111",
  60791=>"101010111",
  60792=>"001000111",
  60793=>"111111111",
  60794=>"111111010",
  60795=>"000000101",
  60796=>"111001011",
  60797=>"111111111",
  60798=>"000000000",
  60799=>"000000000",
  60800=>"100100110",
  60801=>"001001111",
  60802=>"000001000",
  60803=>"111111111",
  60804=>"111111111",
  60805=>"000010000",
  60806=>"111110111",
  60807=>"101001111",
  60808=>"111111001",
  60809=>"111111010",
  60810=>"100000101",
  60811=>"001100000",
  60812=>"000000111",
  60813=>"110110000",
  60814=>"111111111",
  60815=>"000000110",
  60816=>"000000000",
  60817=>"101111111",
  60818=>"001001111",
  60819=>"111011001",
  60820=>"111000111",
  60821=>"000010000",
  60822=>"011011001",
  60823=>"000000000",
  60824=>"000000110",
  60825=>"010010111",
  60826=>"001001001",
  60827=>"100000000",
  60828=>"001101111",
  60829=>"110111000",
  60830=>"000000000",
  60831=>"001000000",
  60832=>"000000111",
  60833=>"100100000",
  60834=>"110110111",
  60835=>"000000000",
  60836=>"000000001",
  60837=>"000000000",
  60838=>"001001111",
  60839=>"111010000",
  60840=>"111111111",
  60841=>"111000100",
  60842=>"111111111",
  60843=>"001001011",
  60844=>"111001110",
  60845=>"000001111",
  60846=>"000000101",
  60847=>"000000000",
  60848=>"000000111",
  60849=>"000100000",
  60850=>"001000001",
  60851=>"110111111",
  60852=>"000000000",
  60853=>"111011110",
  60854=>"111101111",
  60855=>"111001010",
  60856=>"001000010",
  60857=>"011001001",
  60858=>"001000000",
  60859=>"000000000",
  60860=>"001001111",
  60861=>"111001011",
  60862=>"101001000",
  60863=>"100100000",
  60864=>"111000100",
  60865=>"001000100",
  60866=>"001000000",
  60867=>"000000100",
  60868=>"000000111",
  60869=>"011110111",
  60870=>"001000000",
  60871=>"001001101",
  60872=>"100111111",
  60873=>"000101111",
  60874=>"001001101",
  60875=>"000001001",
  60876=>"111100111",
  60877=>"000001111",
  60878=>"000000000",
  60879=>"000000100",
  60880=>"101000000",
  60881=>"110111000",
  60882=>"001111110",
  60883=>"000001111",
  60884=>"011111111",
  60885=>"111111111",
  60886=>"000001001",
  60887=>"011011101",
  60888=>"001001111",
  60889=>"011011111",
  60890=>"111111000",
  60891=>"000111111",
  60892=>"010111010",
  60893=>"000000000",
  60894=>"111111111",
  60895=>"011000001",
  60896=>"101000000",
  60897=>"111111000",
  60898=>"000000000",
  60899=>"010110000",
  60900=>"110110111",
  60901=>"101101101",
  60902=>"001001111",
  60903=>"000000011",
  60904=>"000000000",
  60905=>"000110111",
  60906=>"001000110",
  60907=>"110111000",
  60908=>"111100100",
  60909=>"001000000",
  60910=>"101000000",
  60911=>"101000111",
  60912=>"001001000",
  60913=>"000000000",
  60914=>"110000111",
  60915=>"000000000",
  60916=>"000011111",
  60917=>"101101000",
  60918=>"110110110",
  60919=>"000000110",
  60920=>"111111111",
  60921=>"001001001",
  60922=>"001101101",
  60923=>"101001100",
  60924=>"111000000",
  60925=>"100110111",
  60926=>"001001011",
  60927=>"111111111",
  60928=>"111111111",
  60929=>"000000000",
  60930=>"000000001",
  60931=>"000000000",
  60932=>"000000000",
  60933=>"100110000",
  60934=>"011000001",
  60935=>"000000001",
  60936=>"000111111",
  60937=>"110111111",
  60938=>"100001001",
  60939=>"101111111",
  60940=>"101000000",
  60941=>"000100000",
  60942=>"110001111",
  60943=>"000000000",
  60944=>"111111111",
  60945=>"111100000",
  60946=>"111111111",
  60947=>"110111111",
  60948=>"111111111",
  60949=>"111000000",
  60950=>"011000000",
  60951=>"111110000",
  60952=>"000000000",
  60953=>"001000000",
  60954=>"000000000",
  60955=>"000100111",
  60956=>"001111111",
  60957=>"111111111",
  60958=>"101100000",
  60959=>"111111000",
  60960=>"111111111",
  60961=>"111111110",
  60962=>"111111111",
  60963=>"100100001",
  60964=>"001000000",
  60965=>"000000000",
  60966=>"111111111",
  60967=>"000000100",
  60968=>"111111000",
  60969=>"111111111",
  60970=>"111000000",
  60971=>"000000000",
  60972=>"000000000",
  60973=>"111111111",
  60974=>"111111111",
  60975=>"111111100",
  60976=>"000101000",
  60977=>"111111000",
  60978=>"111100111",
  60979=>"000000000",
  60980=>"000000000",
  60981=>"111111110",
  60982=>"001000000",
  60983=>"000000000",
  60984=>"000000001",
  60985=>"101000000",
  60986=>"011111001",
  60987=>"111000000",
  60988=>"101100111",
  60989=>"111000000",
  60990=>"111111111",
  60991=>"111111111",
  60992=>"111000000",
  60993=>"000000011",
  60994=>"000000000",
  60995=>"000000100",
  60996=>"100101111",
  60997=>"111111110",
  60998=>"111111011",
  60999=>"110000110",
  61000=>"000000001",
  61001=>"000000001",
  61002=>"111111111",
  61003=>"000000110",
  61004=>"000110110",
  61005=>"111111111",
  61006=>"000000000",
  61007=>"000000111",
  61008=>"110110111",
  61009=>"110100000",
  61010=>"000000110",
  61011=>"000111111",
  61012=>"111111111",
  61013=>"111001000",
  61014=>"100000001",
  61015=>"000000000",
  61016=>"111111100",
  61017=>"111111111",
  61018=>"000000111",
  61019=>"000001110",
  61020=>"000000111",
  61021=>"000000000",
  61022=>"000000111",
  61023=>"001001011",
  61024=>"000000110",
  61025=>"100000000",
  61026=>"100000100",
  61027=>"000000000",
  61028=>"111111000",
  61029=>"001000000",
  61030=>"111111111",
  61031=>"001101110",
  61032=>"111111111",
  61033=>"000000101",
  61034=>"001000000",
  61035=>"011111011",
  61036=>"111111111",
  61037=>"000000000",
  61038=>"111111111",
  61039=>"001001001",
  61040=>"100000000",
  61041=>"111000111",
  61042=>"110010010",
  61043=>"111111111",
  61044=>"000000000",
  61045=>"001000010",
  61046=>"011000001",
  61047=>"111111111",
  61048=>"000000111",
  61049=>"111111000",
  61050=>"111111100",
  61051=>"000000000",
  61052=>"111111111",
  61053=>"001111011",
  61054=>"111111111",
  61055=>"110111111",
  61056=>"001000000",
  61057=>"011111110",
  61058=>"000001111",
  61059=>"110001000",
  61060=>"111111111",
  61061=>"111111111",
  61062=>"111011000",
  61063=>"000000000",
  61064=>"110110000",
  61065=>"000000000",
  61066=>"000000000",
  61067=>"010110111",
  61068=>"111111111",
  61069=>"000000000",
  61070=>"111100000",
  61071=>"111111111",
  61072=>"000000111",
  61073=>"000000000",
  61074=>"101111111",
  61075=>"111111000",
  61076=>"110000000",
  61077=>"001111011",
  61078=>"111111111",
  61079=>"000000000",
  61080=>"000000001",
  61081=>"111111100",
  61082=>"000000000",
  61083=>"011110001",
  61084=>"011000111",
  61085=>"100000000",
  61086=>"000000000",
  61087=>"000000010",
  61088=>"000000000",
  61089=>"110111111",
  61090=>"111111111",
  61091=>"100110110",
  61092=>"000100101",
  61093=>"111010011",
  61094=>"000000001",
  61095=>"111110010",
  61096=>"011011000",
  61097=>"100100110",
  61098=>"011011001",
  61099=>"100111001",
  61100=>"001000111",
  61101=>"001001101",
  61102=>"111111111",
  61103=>"000011111",
  61104=>"000000000",
  61105=>"001101000",
  61106=>"110111110",
  61107=>"111111010",
  61108=>"011111110",
  61109=>"000000000",
  61110=>"111001000",
  61111=>"011111100",
  61112=>"000000000",
  61113=>"111111001",
  61114=>"000000000",
  61115=>"011001001",
  61116=>"000000000",
  61117=>"101111111",
  61118=>"110000000",
  61119=>"000110010",
  61120=>"001111001",
  61121=>"110000001",
  61122=>"000000111",
  61123=>"011011000",
  61124=>"000100001",
  61125=>"000000111",
  61126=>"111111000",
  61127=>"000100010",
  61128=>"001000000",
  61129=>"000000011",
  61130=>"000000111",
  61131=>"001011111",
  61132=>"000000000",
  61133=>"111111011",
  61134=>"011000000",
  61135=>"101100111",
  61136=>"100010000",
  61137=>"000010110",
  61138=>"111001000",
  61139=>"000000111",
  61140=>"110111011",
  61141=>"111110110",
  61142=>"001111111",
  61143=>"000001111",
  61144=>"100000000",
  61145=>"111011101",
  61146=>"111111100",
  61147=>"001001001",
  61148=>"011000000",
  61149=>"000000000",
  61150=>"111111111",
  61151=>"100100111",
  61152=>"110111111",
  61153=>"111111111",
  61154=>"001000000",
  61155=>"011010000",
  61156=>"001111111",
  61157=>"001000110",
  61158=>"111111110",
  61159=>"111111111",
  61160=>"000111111",
  61161=>"000000000",
  61162=>"001101011",
  61163=>"101111111",
  61164=>"000110111",
  61165=>"111111111",
  61166=>"000111111",
  61167=>"000000111",
  61168=>"001000110",
  61169=>"111111111",
  61170=>"001000000",
  61171=>"000000111",
  61172=>"110110111",
  61173=>"111111111",
  61174=>"000000000",
  61175=>"001011001",
  61176=>"111000000",
  61177=>"001011000",
  61178=>"000000000",
  61179=>"000100100",
  61180=>"111011011",
  61181=>"111111111",
  61182=>"111111111",
  61183=>"001000000",
  61184=>"000000000",
  61185=>"100110111",
  61186=>"110100000",
  61187=>"100101111",
  61188=>"000000111",
  61189=>"111111111",
  61190=>"111111111",
  61191=>"000000110",
  61192=>"000000000",
  61193=>"000011011",
  61194=>"000100100",
  61195=>"000000001",
  61196=>"000000110",
  61197=>"110000111",
  61198=>"111000000",
  61199=>"011111111",
  61200=>"001001101",
  61201=>"001001000",
  61202=>"111111111",
  61203=>"000111011",
  61204=>"000111111",
  61205=>"111101101",
  61206=>"001001111",
  61207=>"000001111",
  61208=>"100011000",
  61209=>"000000000",
  61210=>"000000000",
  61211=>"111011011",
  61212=>"000100000",
  61213=>"001111111",
  61214=>"001011011",
  61215=>"000001001",
  61216=>"110111111",
  61217=>"000000001",
  61218=>"000000000",
  61219=>"000000000",
  61220=>"001001001",
  61221=>"000111111",
  61222=>"000000110",
  61223=>"111111000",
  61224=>"001100000",
  61225=>"111111111",
  61226=>"100000001",
  61227=>"011001001",
  61228=>"111111001",
  61229=>"001011000",
  61230=>"111111111",
  61231=>"001000110",
  61232=>"111111111",
  61233=>"000000000",
  61234=>"000000000",
  61235=>"111111100",
  61236=>"111111111",
  61237=>"000100000",
  61238=>"000000000",
  61239=>"111111111",
  61240=>"000000000",
  61241=>"000000111",
  61242=>"111111111",
  61243=>"111111000",
  61244=>"000000001",
  61245=>"111000000",
  61246=>"000000000",
  61247=>"111111111",
  61248=>"000000000",
  61249=>"111111111",
  61250=>"001011110",
  61251=>"000000000",
  61252=>"111111111",
  61253=>"001101111",
  61254=>"111011000",
  61255=>"111110111",
  61256=>"000000000",
  61257=>"000000111",
  61258=>"100000000",
  61259=>"000000000",
  61260=>"000000000",
  61261=>"111001000",
  61262=>"111001001",
  61263=>"111111000",
  61264=>"011001000",
  61265=>"111111100",
  61266=>"011011011",
  61267=>"001011011",
  61268=>"000000000",
  61269=>"001001000",
  61270=>"111111111",
  61271=>"000110110",
  61272=>"111111111",
  61273=>"010111111",
  61274=>"111111111",
  61275=>"110100000",
  61276=>"110000000",
  61277=>"110000011",
  61278=>"110111100",
  61279=>"000000000",
  61280=>"111111111",
  61281=>"111011000",
  61282=>"010010000",
  61283=>"111111010",
  61284=>"111000000",
  61285=>"000001111",
  61286=>"111111000",
  61287=>"101001011",
  61288=>"001001100",
  61289=>"111111110",
  61290=>"111111111",
  61291=>"111111111",
  61292=>"001111111",
  61293=>"111111111",
  61294=>"001011011",
  61295=>"000000000",
  61296=>"111111111",
  61297=>"111111111",
  61298=>"000000000",
  61299=>"010000100",
  61300=>"111100000",
  61301=>"110000001",
  61302=>"110110010",
  61303=>"001111111",
  61304=>"111000000",
  61305=>"000000000",
  61306=>"111000000",
  61307=>"100100110",
  61308=>"111111111",
  61309=>"111111111",
  61310=>"111111111",
  61311=>"101111111",
  61312=>"000000000",
  61313=>"111110110",
  61314=>"111111111",
  61315=>"000000000",
  61316=>"000001001",
  61317=>"010011000",
  61318=>"100110000",
  61319=>"000000111",
  61320=>"111111111",
  61321=>"111111000",
  61322=>"111111111",
  61323=>"001000000",
  61324=>"001001111",
  61325=>"111111110",
  61326=>"111111111",
  61327=>"111111011",
  61328=>"111111110",
  61329=>"000000000",
  61330=>"110111010",
  61331=>"000000100",
  61332=>"110111111",
  61333=>"000000000",
  61334=>"100000000",
  61335=>"111111101",
  61336=>"111001000",
  61337=>"111111111",
  61338=>"111111100",
  61339=>"000000000",
  61340=>"111101110",
  61341=>"111110000",
  61342=>"000000001",
  61343=>"100101111",
  61344=>"011000101",
  61345=>"000000000",
  61346=>"100010000",
  61347=>"000000111",
  61348=>"000000000",
  61349=>"110110111",
  61350=>"000000111",
  61351=>"000111111",
  61352=>"000110011",
  61353=>"001011111",
  61354=>"000000000",
  61355=>"000000000",
  61356=>"000000000",
  61357=>"001100000",
  61358=>"001000000",
  61359=>"000100010",
  61360=>"111100000",
  61361=>"111111111",
  61362=>"111111001",
  61363=>"000000011",
  61364=>"000111111",
  61365=>"001001111",
  61366=>"111111111",
  61367=>"001001000",
  61368=>"111111111",
  61369=>"000011011",
  61370=>"000000000",
  61371=>"111111000",
  61372=>"000000111",
  61373=>"000000000",
  61374=>"111111111",
  61375=>"111001100",
  61376=>"000111000",
  61377=>"000000000",
  61378=>"000000001",
  61379=>"111111111",
  61380=>"100000000",
  61381=>"000000000",
  61382=>"110000000",
  61383=>"000000001",
  61384=>"000001001",
  61385=>"111100000",
  61386=>"100100100",
  61387=>"000010000",
  61388=>"111111111",
  61389=>"111111101",
  61390=>"000000001",
  61391=>"111111110",
  61392=>"110111000",
  61393=>"111111011",
  61394=>"111111111",
  61395=>"011000110",
  61396=>"011111100",
  61397=>"000000000",
  61398=>"110101110",
  61399=>"100000000",
  61400=>"111111111",
  61401=>"110110110",
  61402=>"001101100",
  61403=>"000000000",
  61404=>"011011111",
  61405=>"111011111",
  61406=>"000000001",
  61407=>"000000001",
  61408=>"000000010",
  61409=>"000000110",
  61410=>"111111000",
  61411=>"111001001",
  61412=>"111011000",
  61413=>"111111000",
  61414=>"000001000",
  61415=>"111111111",
  61416=>"111110011",
  61417=>"111111000",
  61418=>"000111100",
  61419=>"000010010",
  61420=>"111011111",
  61421=>"110100100",
  61422=>"111111001",
  61423=>"111111001",
  61424=>"000000110",
  61425=>"000000111",
  61426=>"111111111",
  61427=>"110010000",
  61428=>"111111011",
  61429=>"000000000",
  61430=>"101100111",
  61431=>"001001001",
  61432=>"000100111",
  61433=>"000000000",
  61434=>"000000000",
  61435=>"000010000",
  61436=>"000000101",
  61437=>"101000000",
  61438=>"111111111",
  61439=>"111111111",
  61440=>"011111111",
  61441=>"111111111",
  61442=>"111110110",
  61443=>"000000000",
  61444=>"000001011",
  61445=>"110000000",
  61446=>"000111111",
  61447=>"111101111",
  61448=>"111111110",
  61449=>"001011000",
  61450=>"000001001",
  61451=>"011011111",
  61452=>"011111111",
  61453=>"110011011",
  61454=>"100000100",
  61455=>"000000000",
  61456=>"100000000",
  61457=>"110110111",
  61458=>"011000010",
  61459=>"000000000",
  61460=>"000000000",
  61461=>"111111110",
  61462=>"001011111",
  61463=>"001000001",
  61464=>"110110110",
  61465=>"011111111",
  61466=>"111000000",
  61467=>"111111000",
  61468=>"111111111",
  61469=>"000000111",
  61470=>"111111111",
  61471=>"000100111",
  61472=>"000000000",
  61473=>"100110111",
  61474=>"111011111",
  61475=>"001000000",
  61476=>"110000000",
  61477=>"111111111",
  61478=>"111111111",
  61479=>"000110100",
  61480=>"001000000",
  61481=>"111111111",
  61482=>"000000010",
  61483=>"000000011",
  61484=>"111000000",
  61485=>"101100001",
  61486=>"000010000",
  61487=>"011111100",
  61488=>"110011011",
  61489=>"001011111",
  61490=>"111111111",
  61491=>"111111001",
  61492=>"001001001",
  61493=>"111111111",
  61494=>"000000000",
  61495=>"000111111",
  61496=>"111011111",
  61497=>"000000010",
  61498=>"000000000",
  61499=>"000101000",
  61500=>"111111111",
  61501=>"011110000",
  61502=>"111111111",
  61503=>"100000111",
  61504=>"000000000",
  61505=>"000011111",
  61506=>"000110100",
  61507=>"000000000",
  61508=>"110110110",
  61509=>"000011111",
  61510=>"100111000",
  61511=>"111111111",
  61512=>"001001001",
  61513=>"000111000",
  61514=>"111111111",
  61515=>"110110111",
  61516=>"111111111",
  61517=>"000000000",
  61518=>"000000001",
  61519=>"111111111",
  61520=>"110110010",
  61521=>"000000000",
  61522=>"100110100",
  61523=>"111111111",
  61524=>"000011111",
  61525=>"101001000",
  61526=>"001001111",
  61527=>"000000000",
  61528=>"001000000",
  61529=>"000000110",
  61530=>"110111111",
  61531=>"000000000",
  61532=>"000000000",
  61533=>"111111111",
  61534=>"111111000",
  61535=>"000000010",
  61536=>"000000000",
  61537=>"001001011",
  61538=>"000100000",
  61539=>"111111111",
  61540=>"101001001",
  61541=>"000000000",
  61542=>"010001111",
  61543=>"000000000",
  61544=>"000000000",
  61545=>"000000000",
  61546=>"000010000",
  61547=>"110111111",
  61548=>"111001011",
  61549=>"111011111",
  61550=>"001000010",
  61551=>"111111110",
  61552=>"000000000",
  61553=>"111110110",
  61554=>"001001001",
  61555=>"111111000",
  61556=>"110110110",
  61557=>"111110000",
  61558=>"000000111",
  61559=>"111111011",
  61560=>"000001000",
  61561=>"100100110",
  61562=>"100110111",
  61563=>"111111000",
  61564=>"001111111",
  61565=>"111111011",
  61566=>"111111111",
  61567=>"000001001",
  61568=>"111000000",
  61569=>"000011000",
  61570=>"001001111",
  61571=>"011001000",
  61572=>"110000000",
  61573=>"000000000",
  61574=>"000000000",
  61575=>"011111001",
  61576=>"010000000",
  61577=>"010000000",
  61578=>"000000000",
  61579=>"000000000",
  61580=>"101000000",
  61581=>"000010011",
  61582=>"111100000",
  61583=>"000000111",
  61584=>"101100110",
  61585=>"000000000",
  61586=>"110111101",
  61587=>"100111111",
  61588=>"000000100",
  61589=>"000000000",
  61590=>"111110110",
  61591=>"111111000",
  61592=>"000001001",
  61593=>"000110111",
  61594=>"111111110",
  61595=>"110111110",
  61596=>"111111111",
  61597=>"111011011",
  61598=>"001111111",
  61599=>"111111111",
  61600=>"001111111",
  61601=>"111111110",
  61602=>"011010001",
  61603=>"000110110",
  61604=>"011011011",
  61605=>"111100000",
  61606=>"000100101",
  61607=>"001001001",
  61608=>"111110110",
  61609=>"111111111",
  61610=>"000011011",
  61611=>"111011001",
  61612=>"000001100",
  61613=>"000011011",
  61614=>"111111111",
  61615=>"000000100",
  61616=>"000001111",
  61617=>"111111000",
  61618=>"000101101",
  61619=>"000110111",
  61620=>"011010110",
  61621=>"011111111",
  61622=>"111111111",
  61623=>"000000011",
  61624=>"000001000",
  61625=>"000100110",
  61626=>"011011001",
  61627=>"001011011",
  61628=>"100000101",
  61629=>"000001000",
  61630=>"110111111",
  61631=>"111111000",
  61632=>"111111101",
  61633=>"000100110",
  61634=>"000000000",
  61635=>"111111111",
  61636=>"000000000",
  61637=>"011001000",
  61638=>"000000010",
  61639=>"111111011",
  61640=>"100000000",
  61641=>"111000001",
  61642=>"000000001",
  61643=>"011110000",
  61644=>"000011111",
  61645=>"000101101",
  61646=>"000000000",
  61647=>"111100111",
  61648=>"011000000",
  61649=>"111000000",
  61650=>"000000000",
  61651=>"111000100",
  61652=>"111111111",
  61653=>"001101101",
  61654=>"000000000",
  61655=>"001000000",
  61656=>"111111111",
  61657=>"000000000",
  61658=>"010011011",
  61659=>"111111100",
  61660=>"011000100",
  61661=>"001000000",
  61662=>"111111111",
  61663=>"011001011",
  61664=>"000100101",
  61665=>"110100100",
  61666=>"110111000",
  61667=>"011011000",
  61668=>"111111111",
  61669=>"000000000",
  61670=>"001000100",
  61671=>"111111111",
  61672=>"100000000",
  61673=>"111111111",
  61674=>"110000000",
  61675=>"111101111",
  61676=>"111001001",
  61677=>"111111111",
  61678=>"111100000",
  61679=>"001011111",
  61680=>"000000001",
  61681=>"100100101",
  61682=>"110111111",
  61683=>"011011000",
  61684=>"110111111",
  61685=>"000000000",
  61686=>"111111000",
  61687=>"100111001",
  61688=>"111011001",
  61689=>"000000100",
  61690=>"001000000",
  61691=>"111111111",
  61692=>"011011011",
  61693=>"011000111",
  61694=>"000000110",
  61695=>"110110110",
  61696=>"000000001",
  61697=>"011011000",
  61698=>"111110110",
  61699=>"000000000",
  61700=>"111111110",
  61701=>"000000000",
  61702=>"111000000",
  61703=>"111110000",
  61704=>"000000000",
  61705=>"111111111",
  61706=>"100100000",
  61707=>"010000000",
  61708=>"000000101",
  61709=>"111111101",
  61710=>"101111001",
  61711=>"000000000",
  61712=>"000000011",
  61713=>"111111011",
  61714=>"111111111",
  61715=>"111111001",
  61716=>"001010010",
  61717=>"000101111",
  61718=>"000001000",
  61719=>"000001111",
  61720=>"000000011",
  61721=>"111000000",
  61722=>"100010110",
  61723=>"110110011",
  61724=>"000000100",
  61725=>"110111111",
  61726=>"110111111",
  61727=>"011001011",
  61728=>"011101011",
  61729=>"001111111",
  61730=>"110110000",
  61731=>"000000000",
  61732=>"110110000",
  61733=>"111001001",
  61734=>"111111111",
  61735=>"000111111",
  61736=>"111111011",
  61737=>"000010000",
  61738=>"000001011",
  61739=>"101000000",
  61740=>"000000000",
  61741=>"000001011",
  61742=>"111111000",
  61743=>"001001001",
  61744=>"111111110",
  61745=>"011001001",
  61746=>"000000001",
  61747=>"101001001",
  61748=>"000000000",
  61749=>"000000000",
  61750=>"001000011",
  61751=>"011000000",
  61752=>"001001000",
  61753=>"111000000",
  61754=>"000000000",
  61755=>"111100100",
  61756=>"110111111",
  61757=>"000000000",
  61758=>"000000000",
  61759=>"000001100",
  61760=>"111111000",
  61761=>"000000000",
  61762=>"111111110",
  61763=>"000000000",
  61764=>"011011001",
  61765=>"011000000",
  61766=>"000000111",
  61767=>"001011000",
  61768=>"000000111",
  61769=>"010000100",
  61770=>"100010011",
  61771=>"100000001",
  61772=>"010010010",
  61773=>"010011111",
  61774=>"111001000",
  61775=>"011011001",
  61776=>"001111110",
  61777=>"110111011",
  61778=>"111111111",
  61779=>"111001000",
  61780=>"101111101",
  61781=>"110010111",
  61782=>"000000100",
  61783=>"000000001",
  61784=>"111111111",
  61785=>"000010111",
  61786=>"000000001",
  61787=>"011111111",
  61788=>"111111100",
  61789=>"111111011",
  61790=>"000000000",
  61791=>"001001001",
  61792=>"000000111",
  61793=>"111111111",
  61794=>"111111111",
  61795=>"111111111",
  61796=>"111111111",
  61797=>"000001011",
  61798=>"111111111",
  61799=>"111111011",
  61800=>"001001000",
  61801=>"111011111",
  61802=>"001000000",
  61803=>"111011011",
  61804=>"111111001",
  61805=>"000000001",
  61806=>"110111111",
  61807=>"000000000",
  61808=>"000000000",
  61809=>"000000000",
  61810=>"101110000",
  61811=>"011111011",
  61812=>"000011111",
  61813=>"000000000",
  61814=>"110110111",
  61815=>"000000100",
  61816=>"000010111",
  61817=>"111000000",
  61818=>"010000000",
  61819=>"001001011",
  61820=>"110110110",
  61821=>"111111111",
  61822=>"000000000",
  61823=>"000000000",
  61824=>"000000000",
  61825=>"111011011",
  61826=>"001001000",
  61827=>"111111110",
  61828=>"110111110",
  61829=>"000000000",
  61830=>"000111111",
  61831=>"111111100",
  61832=>"000000100",
  61833=>"000000011",
  61834=>"111111101",
  61835=>"000000000",
  61836=>"111111111",
  61837=>"011100001",
  61838=>"000000011",
  61839=>"000101111",
  61840=>"100000100",
  61841=>"011111111",
  61842=>"111110111",
  61843=>"011111111",
  61844=>"000110111",
  61845=>"000000000",
  61846=>"100101111",
  61847=>"111111111",
  61848=>"000000011",
  61849=>"100110110",
  61850=>"111111000",
  61851=>"011011011",
  61852=>"001001000",
  61853=>"000000001",
  61854=>"000000001",
  61855=>"111111111",
  61856=>"111100100",
  61857=>"100110111",
  61858=>"111110100",
  61859=>"111110100",
  61860=>"001000000",
  61861=>"111111111",
  61862=>"111111110",
  61863=>"111110000",
  61864=>"110110110",
  61865=>"000100100",
  61866=>"000000000",
  61867=>"001001011",
  61868=>"000000000",
  61869=>"000000111",
  61870=>"000000110",
  61871=>"000000000",
  61872=>"000110110",
  61873=>"000000111",
  61874=>"100101001",
  61875=>"111111111",
  61876=>"000000000",
  61877=>"011001000",
  61878=>"000100000",
  61879=>"100000000",
  61880=>"110011000",
  61881=>"100100100",
  61882=>"010000010",
  61883=>"111111111",
  61884=>"111011110",
  61885=>"111100101",
  61886=>"000000000",
  61887=>"001001001",
  61888=>"111011111",
  61889=>"111111000",
  61890=>"000000000",
  61891=>"000011010",
  61892=>"001000100",
  61893=>"001111101",
  61894=>"111111111",
  61895=>"111111111",
  61896=>"000000000",
  61897=>"000000000",
  61898=>"111111100",
  61899=>"000000000",
  61900=>"010011000",
  61901=>"001000111",
  61902=>"000110001",
  61903=>"000110111",
  61904=>"000000101",
  61905=>"000001001",
  61906=>"001000111",
  61907=>"111111011",
  61908=>"000110111",
  61909=>"000000000",
  61910=>"111101000",
  61911=>"011111111",
  61912=>"110000000",
  61913=>"011000010",
  61914=>"011010000",
  61915=>"001111111",
  61916=>"000000011",
  61917=>"011111011",
  61918=>"111111011",
  61919=>"000000001",
  61920=>"000000000",
  61921=>"110111111",
  61922=>"111000000",
  61923=>"111100000",
  61924=>"000000111",
  61925=>"111110100",
  61926=>"000000000",
  61927=>"000000000",
  61928=>"111111011",
  61929=>"111111111",
  61930=>"111111111",
  61931=>"101111011",
  61932=>"110111010",
  61933=>"000101101",
  61934=>"111111111",
  61935=>"000010000",
  61936=>"001101101",
  61937=>"111111111",
  61938=>"111011011",
  61939=>"000000000",
  61940=>"000000011",
  61941=>"000000000",
  61942=>"000000000",
  61943=>"000001001",
  61944=>"111111111",
  61945=>"000011111",
  61946=>"100100000",
  61947=>"100100000",
  61948=>"010011000",
  61949=>"111110010",
  61950=>"000000000",
  61951=>"001001111",
  61952=>"000000010",
  61953=>"000010111",
  61954=>"110111111",
  61955=>"111111111",
  61956=>"100000110",
  61957=>"000000110",
  61958=>"011000000",
  61959=>"100101111",
  61960=>"111111001",
  61961=>"000000011",
  61962=>"000000000",
  61963=>"111111001",
  61964=>"110110100",
  61965=>"001000000",
  61966=>"110111111",
  61967=>"001000000",
  61968=>"011000000",
  61969=>"000011111",
  61970=>"011101101",
  61971=>"111111111",
  61972=>"011000000",
  61973=>"110111111",
  61974=>"000000000",
  61975=>"000111111",
  61976=>"100000110",
  61977=>"000000000",
  61978=>"000000111",
  61979=>"011111111",
  61980=>"000000000",
  61981=>"111111100",
  61982=>"111100000",
  61983=>"111111000",
  61984=>"000000110",
  61985=>"011000000",
  61986=>"111100111",
  61987=>"000000100",
  61988=>"111111010",
  61989=>"000111111",
  61990=>"111111001",
  61991=>"111000111",
  61992=>"101111111",
  61993=>"000010011",
  61994=>"000000111",
  61995=>"111100000",
  61996=>"111111010",
  61997=>"000000011",
  61998=>"100000000",
  61999=>"110111011",
  62000=>"000000101",
  62001=>"000000011",
  62002=>"000001011",
  62003=>"000000000",
  62004=>"100110000",
  62005=>"000111010",
  62006=>"011000000",
  62007=>"110100100",
  62008=>"111011000",
  62009=>"100000000",
  62010=>"000000000",
  62011=>"111111111",
  62012=>"100101101",
  62013=>"111000000",
  62014=>"001001011",
  62015=>"000000000",
  62016=>"111111000",
  62017=>"000011001",
  62018=>"110110110",
  62019=>"111111000",
  62020=>"000100111",
  62021=>"001000110",
  62022=>"111101111",
  62023=>"000001111",
  62024=>"111111110",
  62025=>"101000111",
  62026=>"111111111",
  62027=>"111111111",
  62028=>"111110110",
  62029=>"001000001",
  62030=>"000000000",
  62031=>"000000111",
  62032=>"000000000",
  62033=>"100000001",
  62034=>"000000100",
  62035=>"111000000",
  62036=>"000000000",
  62037=>"000000111",
  62038=>"000100100",
  62039=>"111111111",
  62040=>"110000000",
  62041=>"111000111",
  62042=>"111111000",
  62043=>"111111101",
  62044=>"000111110",
  62045=>"111111111",
  62046=>"111100001",
  62047=>"111110000",
  62048=>"111111100",
  62049=>"000000000",
  62050=>"000011111",
  62051=>"000101111",
  62052=>"110111111",
  62053=>"000000000",
  62054=>"011010111",
  62055=>"111111111",
  62056=>"100100111",
  62057=>"011000110",
  62058=>"111111111",
  62059=>"000000001",
  62060=>"111110100",
  62061=>"101101111",
  62062=>"110100000",
  62063=>"000000000",
  62064=>"001001000",
  62065=>"000000000",
  62066=>"111001001",
  62067=>"000110110",
  62068=>"001000010",
  62069=>"110111111",
  62070=>"011011111",
  62071=>"011011000",
  62072=>"000000100",
  62073=>"001000000",
  62074=>"000011111",
  62075=>"000000111",
  62076=>"111110100",
  62077=>"000000000",
  62078=>"011001111",
  62079=>"001001111",
  62080=>"000111110",
  62081=>"000000111",
  62082=>"111111111",
  62083=>"100000000",
  62084=>"001000100",
  62085=>"100000100",
  62086=>"110110111",
  62087=>"110111010",
  62088=>"111111111",
  62089=>"111000110",
  62090=>"110111000",
  62091=>"111011000",
  62092=>"000001000",
  62093=>"100110111",
  62094=>"100100110",
  62095=>"110000000",
  62096=>"000000111",
  62097=>"111011001",
  62098=>"111111000",
  62099=>"000000100",
  62100=>"111000000",
  62101=>"111001111",
  62102=>"000000111",
  62103=>"111111111",
  62104=>"111111111",
  62105=>"001000110",
  62106=>"001111110",
  62107=>"111111000",
  62108=>"111111111",
  62109=>"001111111",
  62110=>"111111001",
  62111=>"000000111",
  62112=>"000000111",
  62113=>"000000100",
  62114=>"000000111",
  62115=>"111111111",
  62116=>"100110111",
  62117=>"100000101",
  62118=>"111101111",
  62119=>"000100100",
  62120=>"111001000",
  62121=>"000000111",
  62122=>"111111111",
  62123=>"111111111",
  62124=>"111111000",
  62125=>"110110100",
  62126=>"000000110",
  62127=>"111111100",
  62128=>"111011000",
  62129=>"000100100",
  62130=>"111111111",
  62131=>"000000111",
  62132=>"000110111",
  62133=>"111110111",
  62134=>"000110100",
  62135=>"000000001",
  62136=>"000000111",
  62137=>"000000000",
  62138=>"100000111",
  62139=>"100101001",
  62140=>"111000000",
  62141=>"100111000",
  62142=>"111011111",
  62143=>"010011000",
  62144=>"000000000",
  62145=>"110111100",
  62146=>"000000111",
  62147=>"011111111",
  62148=>"111111111",
  62149=>"110110111",
  62150=>"000010010",
  62151=>"001100111",
  62152=>"111111111",
  62153=>"000000111",
  62154=>"100000000",
  62155=>"001001001",
  62156=>"111111100",
  62157=>"000111111",
  62158=>"000100110",
  62159=>"000000000",
  62160=>"000111011",
  62161=>"000000111",
  62162=>"000000111",
  62163=>"011001001",
  62164=>"100000000",
  62165=>"111111000",
  62166=>"000000000",
  62167=>"000000000",
  62168=>"111111111",
  62169=>"000000001",
  62170=>"101000000",
  62171=>"010111111",
  62172=>"100111100",
  62173=>"111110110",
  62174=>"000000011",
  62175=>"000000100",
  62176=>"111111000",
  62177=>"111011000",
  62178=>"111111111",
  62179=>"111110111",
  62180=>"100111110",
  62181=>"111111111",
  62182=>"111111000",
  62183=>"101000111",
  62184=>"111011000",
  62185=>"111111111",
  62186=>"000110111",
  62187=>"111100001",
  62188=>"000110111",
  62189=>"001000111",
  62190=>"010000000",
  62191=>"111111100",
  62192=>"000000001",
  62193=>"000001111",
  62194=>"011011111",
  62195=>"011011011",
  62196=>"000110001",
  62197=>"110111001",
  62198=>"000011011",
  62199=>"111010000",
  62200=>"000000000",
  62201=>"111111111",
  62202=>"100000100",
  62203=>"111111111",
  62204=>"111011001",
  62205=>"110000001",
  62206=>"000111000",
  62207=>"010011011",
  62208=>"000000000",
  62209=>"101001001",
  62210=>"000000000",
  62211=>"000000111",
  62212=>"000111101",
  62213=>"000000000",
  62214=>"011010000",
  62215=>"100101111",
  62216=>"111111100",
  62217=>"000010010",
  62218=>"000000011",
  62219=>"111010000",
  62220=>"000000000",
  62221=>"111101001",
  62222=>"111110111",
  62223=>"000000110",
  62224=>"000100000",
  62225=>"000000100",
  62226=>"111100111",
  62227=>"000000000",
  62228=>"000000010",
  62229=>"001011111",
  62230=>"000000011",
  62231=>"111000111",
  62232=>"010111111",
  62233=>"111111011",
  62234=>"000000000",
  62235=>"000000001",
  62236=>"111111111",
  62237=>"000000000",
  62238=>"000000001",
  62239=>"000000111",
  62240=>"101101100",
  62241=>"000000111",
  62242=>"000000111",
  62243=>"111111110",
  62244=>"110100101",
  62245=>"011111111",
  62246=>"100000000",
  62247=>"000001111",
  62248=>"011111110",
  62249=>"100000000",
  62250=>"110110110",
  62251=>"111101111",
  62252=>"111001000",
  62253=>"111111100",
  62254=>"000111111",
  62255=>"100000000",
  62256=>"011111000",
  62257=>"111011001",
  62258=>"110000000",
  62259=>"000000001",
  62260=>"000000000",
  62261=>"001000001",
  62262=>"000000000",
  62263=>"000000000",
  62264=>"000000000",
  62265=>"000000111",
  62266=>"111100101",
  62267=>"000000000",
  62268=>"000000011",
  62269=>"110111000",
  62270=>"000000000",
  62271=>"111110000",
  62272=>"100000000",
  62273=>"001000001",
  62274=>"111111010",
  62275=>"000000000",
  62276=>"110110111",
  62277=>"011001111",
  62278=>"000000000",
  62279=>"111111000",
  62280=>"000000000",
  62281=>"000000000",
  62282=>"000000100",
  62283=>"100110110",
  62284=>"111111111",
  62285=>"111110000",
  62286=>"111101111",
  62287=>"000110000",
  62288=>"001011111",
  62289=>"000000111",
  62290=>"111111111",
  62291=>"110111111",
  62292=>"000000000",
  62293=>"011011011",
  62294=>"000100100",
  62295=>"111111100",
  62296=>"000000101",
  62297=>"000000111",
  62298=>"111100000",
  62299=>"001000000",
  62300=>"000000111",
  62301=>"000000111",
  62302=>"000000000",
  62303=>"111111111",
  62304=>"011111111",
  62305=>"111111111",
  62306=>"011111110",
  62307=>"111101000",
  62308=>"000011110",
  62309=>"000000110",
  62310=>"000000111",
  62311=>"110110100",
  62312=>"100101001",
  62313=>"001000000",
  62314=>"001000000",
  62315=>"100111111",
  62316=>"000110111",
  62317=>"000010110",
  62318=>"111111111",
  62319=>"111100111",
  62320=>"000000000",
  62321=>"111111011",
  62322=>"111010000",
  62323=>"111111000",
  62324=>"000000100",
  62325=>"000011100",
  62326=>"111111111",
  62327=>"000100110",
  62328=>"111111111",
  62329=>"111011111",
  62330=>"000001011",
  62331=>"000000000",
  62332=>"111001001",
  62333=>"111000000",
  62334=>"000000111",
  62335=>"000000111",
  62336=>"111111110",
  62337=>"111111100",
  62338=>"000000111",
  62339=>"001000111",
  62340=>"001111011",
  62341=>"000010000",
  62342=>"000011111",
  62343=>"000100111",
  62344=>"001001111",
  62345=>"000000000",
  62346=>"111111001",
  62347=>"111000000",
  62348=>"111111111",
  62349=>"100110110",
  62350=>"000101110",
  62351=>"000000000",
  62352=>"001001000",
  62353=>"000100111",
  62354=>"001011000",
  62355=>"100000100",
  62356=>"001111000",
  62357=>"000000010",
  62358=>"000000000",
  62359=>"110001111",
  62360=>"000000000",
  62361=>"111111100",
  62362=>"000001001",
  62363=>"000000011",
  62364=>"111111011",
  62365=>"000111111",
  62366=>"000000111",
  62367=>"101111111",
  62368=>"000000011",
  62369=>"000000000",
  62370=>"100100000",
  62371=>"110000001",
  62372=>"111110000",
  62373=>"001000000",
  62374=>"001001111",
  62375=>"000010110",
  62376=>"001111111",
  62377=>"111111011",
  62378=>"111111011",
  62379=>"111000100",
  62380=>"000000111",
  62381=>"001000000",
  62382=>"000000100",
  62383=>"000101001",
  62384=>"111111111",
  62385=>"000011111",
  62386=>"000000000",
  62387=>"011001000",
  62388=>"111111000",
  62389=>"111000000",
  62390=>"000100100",
  62391=>"000000111",
  62392=>"001000111",
  62393=>"011011111",
  62394=>"000000110",
  62395=>"111111000",
  62396=>"111111111",
  62397=>"000000000",
  62398=>"000000111",
  62399=>"110111000",
  62400=>"111000000",
  62401=>"000000000",
  62402=>"000000001",
  62403=>"000000001",
  62404=>"100111110",
  62405=>"000000000",
  62406=>"000000000",
  62407=>"000000111",
  62408=>"111000010",
  62409=>"000000110",
  62410=>"001000000",
  62411=>"000111110",
  62412=>"111000111",
  62413=>"111111111",
  62414=>"011111000",
  62415=>"111011001",
  62416=>"000000011",
  62417=>"111111010",
  62418=>"000001010",
  62419=>"001000000",
  62420=>"000110111",
  62421=>"111111011",
  62422=>"111111111",
  62423=>"001011011",
  62424=>"100100100",
  62425=>"111111000",
  62426=>"000000000",
  62427=>"000111111",
  62428=>"010011000",
  62429=>"000000110",
  62430=>"001011000",
  62431=>"110000000",
  62432=>"101111000",
  62433=>"011100100",
  62434=>"110000010",
  62435=>"000000111",
  62436=>"100010000",
  62437=>"000000000",
  62438=>"001111001",
  62439=>"111111011",
  62440=>"110000000",
  62441=>"111111111",
  62442=>"011111111",
  62443=>"100100000",
  62444=>"110000110",
  62445=>"000000110",
  62446=>"110111101",
  62447=>"000000000",
  62448=>"000000000",
  62449=>"000111111",
  62450=>"111111011",
  62451=>"000000000",
  62452=>"111011000",
  62453=>"000000011",
  62454=>"100000000",
  62455=>"100100110",
  62456=>"100000000",
  62457=>"000110000",
  62458=>"000000001",
  62459=>"000000000",
  62460=>"000000111",
  62461=>"111111010",
  62462=>"111011100",
  62463=>"111111111",
  62464=>"001000000",
  62465=>"111001111",
  62466=>"111001111",
  62467=>"111000000",
  62468=>"010010001",
  62469=>"111000000",
  62470=>"011011000",
  62471=>"101001111",
  62472=>"111111000",
  62473=>"011011011",
  62474=>"001000001",
  62475=>"100111111",
  62476=>"110111111",
  62477=>"000110111",
  62478=>"111111011",
  62479=>"011011011",
  62480=>"110111111",
  62481=>"111111111",
  62482=>"011111111",
  62483=>"000000000",
  62484=>"000000011",
  62485=>"010010111",
  62486=>"000001111",
  62487=>"110110110",
  62488=>"110110110",
  62489=>"011011000",
  62490=>"000000000",
  62491=>"100101111",
  62492=>"000000101",
  62493=>"000000000",
  62494=>"001001001",
  62495=>"001111111",
  62496=>"010000001",
  62497=>"000000110",
  62498=>"000001000",
  62499=>"111111111",
  62500=>"111000000",
  62501=>"000111111",
  62502=>"100111000",
  62503=>"111111000",
  62504=>"100000000",
  62505=>"000000000",
  62506=>"000000000",
  62507=>"000000000",
  62508=>"000000011",
  62509=>"000000000",
  62510=>"000000000",
  62511=>"000010111",
  62512=>"111001101",
  62513=>"000000000",
  62514=>"000000000",
  62515=>"101000000",
  62516=>"101111111",
  62517=>"000110010",
  62518=>"000000001",
  62519=>"000000001",
  62520=>"101001111",
  62521=>"000111011",
  62522=>"111111111",
  62523=>"110111101",
  62524=>"000000101",
  62525=>"000001101",
  62526=>"111100100",
  62527=>"000000000",
  62528=>"001001101",
  62529=>"100000111",
  62530=>"011000000",
  62531=>"111111111",
  62532=>"000111110",
  62533=>"000000000",
  62534=>"001000010",
  62535=>"100000000",
  62536=>"111001011",
  62537=>"111110111",
  62538=>"010110110",
  62539=>"111111110",
  62540=>"000001001",
  62541=>"000011001",
  62542=>"011000000",
  62543=>"001001111",
  62544=>"000000001",
  62545=>"000111111",
  62546=>"111111000",
  62547=>"111101100",
  62548=>"000000000",
  62549=>"000101000",
  62550=>"111111111",
  62551=>"111111010",
  62552=>"111010000",
  62553=>"111000101",
  62554=>"000010111",
  62555=>"110000000",
  62556=>"000000111",
  62557=>"101101111",
  62558=>"011111010",
  62559=>"000000111",
  62560=>"000111011",
  62561=>"000000011",
  62562=>"111111111",
  62563=>"000000001",
  62564=>"110110000",
  62565=>"100100111",
  62566=>"000000111",
  62567=>"000000000",
  62568=>"000000000",
  62569=>"000000111",
  62570=>"000000000",
  62571=>"111111111",
  62572=>"000000000",
  62573=>"111111010",
  62574=>"001001111",
  62575=>"000011011",
  62576=>"111111111",
  62577=>"000000000",
  62578=>"011011110",
  62579=>"000000111",
  62580=>"111111001",
  62581=>"110111110",
  62582=>"000000111",
  62583=>"001010000",
  62584=>"000000111",
  62585=>"001000001",
  62586=>"000000000",
  62587=>"100110110",
  62588=>"000000011",
  62589=>"001000000",
  62590=>"000000000",
  62591=>"010000000",
  62592=>"011000000",
  62593=>"101100000",
  62594=>"001000000",
  62595=>"111111011",
  62596=>"000101111",
  62597=>"000011000",
  62598=>"111111000",
  62599=>"000000000",
  62600=>"111000000",
  62601=>"111111111",
  62602=>"111111111",
  62603=>"000000000",
  62604=>"100100110",
  62605=>"000000000",
  62606=>"100111000",
  62607=>"010000000",
  62608=>"111111111",
  62609=>"000000000",
  62610=>"000000000",
  62611=>"001111111",
  62612=>"101111111",
  62613=>"110000011",
  62614=>"101000000",
  62615=>"000000111",
  62616=>"101001001",
  62617=>"000100111",
  62618=>"111001010",
  62619=>"000100111",
  62620=>"111000000",
  62621=>"011001111",
  62622=>"001000100",
  62623=>"011011011",
  62624=>"000000000",
  62625=>"011111011",
  62626=>"101000000",
  62627=>"000000000",
  62628=>"100111111",
  62629=>"000101100",
  62630=>"101111110",
  62631=>"111111011",
  62632=>"001001001",
  62633=>"000001111",
  62634=>"111110000",
  62635=>"000000000",
  62636=>"000001010",
  62637=>"100101111",
  62638=>"100111000",
  62639=>"011001111",
  62640=>"111110111",
  62641=>"000011011",
  62642=>"011111010",
  62643=>"000000000",
  62644=>"110011011",
  62645=>"111011011",
  62646=>"001111110",
  62647=>"110111110",
  62648=>"000000111",
  62649=>"110000001",
  62650=>"011011011",
  62651=>"111011000",
  62652=>"100000000",
  62653=>"111111010",
  62654=>"100001001",
  62655=>"001000111",
  62656=>"111111011",
  62657=>"000000000",
  62658=>"000000000",
  62659=>"000001111",
  62660=>"001111111",
  62661=>"011000001",
  62662=>"100100000",
  62663=>"101101111",
  62664=>"000011011",
  62665=>"111111101",
  62666=>"101100101",
  62667=>"000000000",
  62668=>"000111011",
  62669=>"111000000",
  62670=>"111111001",
  62671=>"100000001",
  62672=>"010000101",
  62673=>"111111111",
  62674=>"111111111",
  62675=>"110110000",
  62676=>"000000000",
  62677=>"110111001",
  62678=>"000000000",
  62679=>"111001100",
  62680=>"000000000",
  62681=>"000000000",
  62682=>"101110111",
  62683=>"000111011",
  62684=>"000011011",
  62685=>"000000000",
  62686=>"111111111",
  62687=>"000000000",
  62688=>"011000101",
  62689=>"000000110",
  62690=>"011101000",
  62691=>"100011111",
  62692=>"000000000",
  62693=>"111110000",
  62694=>"001001001",
  62695=>"111111111",
  62696=>"100111010",
  62697=>"011111111",
  62698=>"000000110",
  62699=>"111001000",
  62700=>"111111111",
  62701=>"000000000",
  62702=>"110110010",
  62703=>"000000000",
  62704=>"100100000",
  62705=>"011111111",
  62706=>"011001011",
  62707=>"111000111",
  62708=>"111111111",
  62709=>"001011011",
  62710=>"100111111",
  62711=>"111110001",
  62712=>"111111000",
  62713=>"000000000",
  62714=>"000011000",
  62715=>"111111111",
  62716=>"011111100",
  62717=>"110000000",
  62718=>"111000000",
  62719=>"000000111",
  62720=>"000000000",
  62721=>"111111001",
  62722=>"000000000",
  62723=>"010000000",
  62724=>"111111111",
  62725=>"111111111",
  62726=>"100000100",
  62727=>"000101100",
  62728=>"001000000",
  62729=>"101000000",
  62730=>"000000001",
  62731=>"111111111",
  62732=>"101001001",
  62733=>"111000000",
  62734=>"010111111",
  62735=>"010110000",
  62736=>"001001101",
  62737=>"011111111",
  62738=>"111111001",
  62739=>"000111101",
  62740=>"111111111",
  62741=>"101111111",
  62742=>"100111111",
  62743=>"101111111",
  62744=>"011011000",
  62745=>"011011000",
  62746=>"000000000",
  62747=>"000000000",
  62748=>"100100111",
  62749=>"111000000",
  62750=>"000000001",
  62751=>"000000000",
  62752=>"000000000",
  62753=>"000000000",
  62754=>"111100000",
  62755=>"101101001",
  62756=>"000001001",
  62757=>"111111111",
  62758=>"111111111",
  62759=>"001000000",
  62760=>"000000001",
  62761=>"011111110",
  62762=>"100000001",
  62763=>"111110000",
  62764=>"000001100",
  62765=>"011011000",
  62766=>"111110111",
  62767=>"100000000",
  62768=>"110110111",
  62769=>"000010000",
  62770=>"001101111",
  62771=>"000000100",
  62772=>"000010110",
  62773=>"000000000",
  62774=>"000000000",
  62775=>"001000001",
  62776=>"000000000",
  62777=>"000000000",
  62778=>"101000101",
  62779=>"000000001",
  62780=>"100101111",
  62781=>"000000000",
  62782=>"111101101",
  62783=>"000000000",
  62784=>"111101000",
  62785=>"110111110",
  62786=>"110111010",
  62787=>"111111111",
  62788=>"000110000",
  62789=>"011000000",
  62790=>"111111011",
  62791=>"000000010",
  62792=>"000000000",
  62793=>"000011111",
  62794=>"010111111",
  62795=>"111110111",
  62796=>"000000000",
  62797=>"011001101",
  62798=>"101001001",
  62799=>"110111000",
  62800=>"000000000",
  62801=>"001000000",
  62802=>"111111111",
  62803=>"111101111",
  62804=>"000010111",
  62805=>"001011011",
  62806=>"000000001",
  62807=>"111001001",
  62808=>"000000000",
  62809=>"001000000",
  62810=>"001001101",
  62811=>"100000000",
  62812=>"111111111",
  62813=>"111111111",
  62814=>"011000000",
  62815=>"111111111",
  62816=>"000010110",
  62817=>"111111111",
  62818=>"110111100",
  62819=>"111100111",
  62820=>"110100000",
  62821=>"000000000",
  62822=>"000101101",
  62823=>"001000101",
  62824=>"001001111",
  62825=>"000111111",
  62826=>"100100111",
  62827=>"111111111",
  62828=>"000000000",
  62829=>"111111111",
  62830=>"001000000",
  62831=>"001000000",
  62832=>"010111111",
  62833=>"111000010",
  62834=>"110111011",
  62835=>"111111110",
  62836=>"011011000",
  62837=>"000000000",
  62838=>"111111111",
  62839=>"110000000",
  62840=>"111001000",
  62841=>"110100000",
  62842=>"000000001",
  62843=>"000111111",
  62844=>"000000000",
  62845=>"111110111",
  62846=>"001011111",
  62847=>"001011101",
  62848=>"111111111",
  62849=>"100011011",
  62850=>"000000000",
  62851=>"011000000",
  62852=>"000111111",
  62853=>"111111111",
  62854=>"001001000",
  62855=>"010011011",
  62856=>"001000000",
  62857=>"110000010",
  62858=>"100100111",
  62859=>"000000000",
  62860=>"111111111",
  62861=>"111111111",
  62862=>"001111010",
  62863=>"000000100",
  62864=>"000000000",
  62865=>"111001001",
  62866=>"011010000",
  62867=>"001001100",
  62868=>"111000111",
  62869=>"000000000",
  62870=>"100000001",
  62871=>"000000100",
  62872=>"011111111",
  62873=>"111111001",
  62874=>"001011000",
  62875=>"111111010",
  62876=>"111111111",
  62877=>"111111111",
  62878=>"011011001",
  62879=>"101111111",
  62880=>"111111111",
  62881=>"111111111",
  62882=>"100111110",
  62883=>"000011111",
  62884=>"101101110",
  62885=>"000000000",
  62886=>"111100111",
  62887=>"011010000",
  62888=>"110000000",
  62889=>"000000101",
  62890=>"111111111",
  62891=>"000000001",
  62892=>"000000000",
  62893=>"000001100",
  62894=>"000000111",
  62895=>"000000111",
  62896=>"111111111",
  62897=>"111111111",
  62898=>"000000111",
  62899=>"000001110",
  62900=>"000000001",
  62901=>"000000100",
  62902=>"000000000",
  62903=>"000000000",
  62904=>"000000011",
  62905=>"111111111",
  62906=>"000000000",
  62907=>"011001011",
  62908=>"000000000",
  62909=>"111101101",
  62910=>"011000000",
  62911=>"111111100",
  62912=>"000000000",
  62913=>"111101111",
  62914=>"111111111",
  62915=>"111111111",
  62916=>"000000101",
  62917=>"011111111",
  62918=>"100111110",
  62919=>"100100111",
  62920=>"011001001",
  62921=>"101000000",
  62922=>"001000000",
  62923=>"000000000",
  62924=>"001010000",
  62925=>"000001001",
  62926=>"111101111",
  62927=>"000000000",
  62928=>"011001000",
  62929=>"000000011",
  62930=>"111111101",
  62931=>"111111000",
  62932=>"111111111",
  62933=>"000000001",
  62934=>"000111111",
  62935=>"111111111",
  62936=>"111000001",
  62937=>"011111111",
  62938=>"111000001",
  62939=>"111111000",
  62940=>"000000001",
  62941=>"111001000",
  62942=>"111111110",
  62943=>"000000001",
  62944=>"110111110",
  62945=>"000000000",
  62946=>"100101101",
  62947=>"001001000",
  62948=>"111011011",
  62949=>"100000000",
  62950=>"111111111",
  62951=>"000000000",
  62952=>"101001001",
  62953=>"000010000",
  62954=>"011000000",
  62955=>"110000111",
  62956=>"111111111",
  62957=>"001100100",
  62958=>"100101111",
  62959=>"000000000",
  62960=>"000000001",
  62961=>"000000000",
  62962=>"111111111",
  62963=>"100000100",
  62964=>"100000111",
  62965=>"111111111",
  62966=>"001001000",
  62967=>"000010000",
  62968=>"000000000",
  62969=>"001101001",
  62970=>"001000100",
  62971=>"111111111",
  62972=>"111011000",
  62973=>"111101111",
  62974=>"011011001",
  62975=>"000000000",
  62976=>"111111111",
  62977=>"001111111",
  62978=>"000010000",
  62979=>"111111001",
  62980=>"111000000",
  62981=>"001111111",
  62982=>"111111111",
  62983=>"000010010",
  62984=>"100000000",
  62985=>"111011000",
  62986=>"000000001",
  62987=>"000000101",
  62988=>"111011011",
  62989=>"111111110",
  62990=>"111001000",
  62991=>"110100110",
  62992=>"111111111",
  62993=>"110010000",
  62994=>"011100000",
  62995=>"000000000",
  62996=>"000000101",
  62997=>"111111111",
  62998=>"100101111",
  62999=>"000000000",
  63000=>"010111111",
  63001=>"000000000",
  63002=>"000000000",
  63003=>"100110111",
  63004=>"000000111",
  63005=>"111111100",
  63006=>"001011010",
  63007=>"111111111",
  63008=>"100000111",
  63009=>"111111001",
  63010=>"000111111",
  63011=>"000100111",
  63012=>"011001000",
  63013=>"000011000",
  63014=>"111111000",
  63015=>"111000000",
  63016=>"010010111",
  63017=>"111111111",
  63018=>"111111111",
  63019=>"011011111",
  63020=>"000000000",
  63021=>"111111011",
  63022=>"000011101",
  63023=>"111000000",
  63024=>"111111011",
  63025=>"111111111",
  63026=>"111001000",
  63027=>"101101101",
  63028=>"111110110",
  63029=>"111111010",
  63030=>"011010010",
  63031=>"001001111",
  63032=>"111111110",
  63033=>"111011111",
  63034=>"111111111",
  63035=>"111111111",
  63036=>"000000000",
  63037=>"100100000",
  63038=>"001000111",
  63039=>"111111111",
  63040=>"001101111",
  63041=>"111111111",
  63042=>"000110000",
  63043=>"111100011",
  63044=>"000100000",
  63045=>"000110100",
  63046=>"111111111",
  63047=>"000000000",
  63048=>"100111111",
  63049=>"000010000",
  63050=>"000000001",
  63051=>"011010111",
  63052=>"101111111",
  63053=>"000000000",
  63054=>"111000000",
  63055=>"111101101",
  63056=>"111111111",
  63057=>"111111100",
  63058=>"111011111",
  63059=>"011011111",
  63060=>"000111111",
  63061=>"111111111",
  63062=>"000000001",
  63063=>"011011000",
  63064=>"010011000",
  63065=>"000000000",
  63066=>"111111111",
  63067=>"000000100",
  63068=>"010011111",
  63069=>"101000000",
  63070=>"000100111",
  63071=>"111111110",
  63072=>"111111110",
  63073=>"011111111",
  63074=>"000110000",
  63075=>"111111111",
  63076=>"001111111",
  63077=>"000010011",
  63078=>"000000000",
  63079=>"111111111",
  63080=>"111111011",
  63081=>"010011010",
  63082=>"000000110",
  63083=>"101111111",
  63084=>"001011000",
  63085=>"000000000",
  63086=>"111111001",
  63087=>"111000011",
  63088=>"111111111",
  63089=>"111001100",
  63090=>"000000000",
  63091=>"110111100",
  63092=>"111111111",
  63093=>"000000000",
  63094=>"111111111",
  63095=>"000000000",
  63096=>"000000111",
  63097=>"011011011",
  63098=>"011001001",
  63099=>"000000101",
  63100=>"000100000",
  63101=>"000000000",
  63102=>"000000010",
  63103=>"000000100",
  63104=>"111111111",
  63105=>"110110111",
  63106=>"110000001",
  63107=>"100000100",
  63108=>"100100100",
  63109=>"000000111",
  63110=>"101111111",
  63111=>"000000100",
  63112=>"101000000",
  63113=>"111110001",
  63114=>"110110111",
  63115=>"111111111",
  63116=>"110111111",
  63117=>"111111111",
  63118=>"100000101",
  63119=>"111100001",
  63120=>"110111011",
  63121=>"000000000",
  63122=>"111111111",
  63123=>"000011111",
  63124=>"111111111",
  63125=>"100110110",
  63126=>"111100000",
  63127=>"111111011",
  63128=>"111011111",
  63129=>"110000010",
  63130=>"100000000",
  63131=>"100111111",
  63132=>"100000100",
  63133=>"010011000",
  63134=>"001000010",
  63135=>"000000111",
  63136=>"001000100",
  63137=>"111111111",
  63138=>"000110111",
  63139=>"111111111",
  63140=>"111101111",
  63141=>"101101000",
  63142=>"111111010",
  63143=>"000000000",
  63144=>"111111111",
  63145=>"100000001",
  63146=>"111000001",
  63147=>"111111111",
  63148=>"001101001",
  63149=>"110110111",
  63150=>"111000000",
  63151=>"010111111",
  63152=>"000000000",
  63153=>"100111100",
  63154=>"000010000",
  63155=>"000111000",
  63156=>"101111111",
  63157=>"000001000",
  63158=>"111110000",
  63159=>"000100000",
  63160=>"000000100",
  63161=>"111111111",
  63162=>"011000001",
  63163=>"111101001",
  63164=>"111111011",
  63165=>"111111111",
  63166=>"000000000",
  63167=>"000010111",
  63168=>"000000000",
  63169=>"100000000",
  63170=>"000000000",
  63171=>"000001000",
  63172=>"010000111",
  63173=>"001000010",
  63174=>"111011001",
  63175=>"110000110",
  63176=>"101101111",
  63177=>"000011010",
  63178=>"110110110",
  63179=>"100110111",
  63180=>"011111110",
  63181=>"000000001",
  63182=>"111111111",
  63183=>"111111111",
  63184=>"000000000",
  63185=>"000100100",
  63186=>"000101111",
  63187=>"101111111",
  63188=>"010011001",
  63189=>"000111111",
  63190=>"111011001",
  63191=>"001111111",
  63192=>"111101111",
  63193=>"110100111",
  63194=>"000000000",
  63195=>"010010000",
  63196=>"100100111",
  63197=>"101000000",
  63198=>"000000000",
  63199=>"110010101",
  63200=>"000010000",
  63201=>"000000000",
  63202=>"000000100",
  63203=>"111111111",
  63204=>"011010111",
  63205=>"000000010",
  63206=>"100100000",
  63207=>"000000000",
  63208=>"011011111",
  63209=>"000000000",
  63210=>"000001001",
  63211=>"010111000",
  63212=>"011001000",
  63213=>"111111000",
  63214=>"101111001",
  63215=>"000111111",
  63216=>"111110110",
  63217=>"011011011",
  63218=>"100110110",
  63219=>"110010000",
  63220=>"111111111",
  63221=>"111110110",
  63222=>"000000000",
  63223=>"000110001",
  63224=>"000000000",
  63225=>"111111111",
  63226=>"010000011",
  63227=>"110100111",
  63228=>"001100000",
  63229=>"100111111",
  63230=>"111011000",
  63231=>"000000000",
  63232=>"111111001",
  63233=>"111111111",
  63234=>"001111011",
  63235=>"111111101",
  63236=>"110111111",
  63237=>"110100100",
  63238=>"000000100",
  63239=>"111111111",
  63240=>"000000000",
  63241=>"001101111",
  63242=>"111111111",
  63243=>"000000000",
  63244=>"100000001",
  63245=>"000000001",
  63246=>"111111111",
  63247=>"111100110",
  63248=>"111111100",
  63249=>"111110111",
  63250=>"111110111",
  63251=>"000001111",
  63252=>"111100000",
  63253=>"111111000",
  63254=>"100110111",
  63255=>"110010111",
  63256=>"011011000",
  63257=>"001001001",
  63258=>"111111111",
  63259=>"000101111",
  63260=>"100100111",
  63261=>"111111000",
  63262=>"111111111",
  63263=>"011001111",
  63264=>"111000110",
  63265=>"011011111",
  63266=>"111111111",
  63267=>"100101111",
  63268=>"110100000",
  63269=>"111111111",
  63270=>"001000000",
  63271=>"110000000",
  63272=>"000100100",
  63273=>"000000101",
  63274=>"111011011",
  63275=>"101101111",
  63276=>"111111110",
  63277=>"100100100",
  63278=>"111110111",
  63279=>"101000000",
  63280=>"001001001",
  63281=>"011011111",
  63282=>"011111010",
  63283=>"111100101",
  63284=>"000110110",
  63285=>"110000110",
  63286=>"100001111",
  63287=>"111111111",
  63288=>"010000000",
  63289=>"111111111",
  63290=>"011011111",
  63291=>"111111111",
  63292=>"001101001",
  63293=>"010100000",
  63294=>"000000111",
  63295=>"001000111",
  63296=>"111101111",
  63297=>"111000000",
  63298=>"100000000",
  63299=>"001001111",
  63300=>"000001101",
  63301=>"111111110",
  63302=>"000111000",
  63303=>"001000000",
  63304=>"111111111",
  63305=>"000111111",
  63306=>"000001111",
  63307=>"111111100",
  63308=>"000000001",
  63309=>"111111011",
  63310=>"111000000",
  63311=>"111111011",
  63312=>"001001001",
  63313=>"000000001",
  63314=>"100000000",
  63315=>"000000000",
  63316=>"111111111",
  63317=>"101000000",
  63318=>"100100111",
  63319=>"100110000",
  63320=>"011011111",
  63321=>"000111010",
  63322=>"110111111",
  63323=>"100101110",
  63324=>"111110110",
  63325=>"011010000",
  63326=>"111111111",
  63327=>"111010000",
  63328=>"000001001",
  63329=>"011011010",
  63330=>"100000000",
  63331=>"111111111",
  63332=>"000110111",
  63333=>"111111000",
  63334=>"101111100",
  63335=>"111111111",
  63336=>"100110111",
  63337=>"000000000",
  63338=>"111111111",
  63339=>"011000110",
  63340=>"000000000",
  63341=>"010000000",
  63342=>"000111111",
  63343=>"001001111",
  63344=>"111100111",
  63345=>"000000011",
  63346=>"000000000",
  63347=>"000000110",
  63348=>"000000000",
  63349=>"000000000",
  63350=>"101111111",
  63351=>"000100000",
  63352=>"111111111",
  63353=>"011000000",
  63354=>"011111110",
  63355=>"111111111",
  63356=>"111111101",
  63357=>"011011111",
  63358=>"000000000",
  63359=>"000111111",
  63360=>"111010111",
  63361=>"110111111",
  63362=>"000010001",
  63363=>"100000011",
  63364=>"111111110",
  63365=>"111011011",
  63366=>"010011111",
  63367=>"110011000",
  63368=>"111111111",
  63369=>"000000000",
  63370=>"000000011",
  63371=>"101111111",
  63372=>"111111111",
  63373=>"100110000",
  63374=>"000000011",
  63375=>"111111111",
  63376=>"111111111",
  63377=>"011111111",
  63378=>"111001000",
  63379=>"001011000",
  63380=>"010010000",
  63381=>"000000011",
  63382=>"000000100",
  63383=>"110111110",
  63384=>"111111111",
  63385=>"101001001",
  63386=>"110111000",
  63387=>"011111111",
  63388=>"000000010",
  63389=>"111010110",
  63390=>"111000000",
  63391=>"111111111",
  63392=>"011001111",
  63393=>"000000100",
  63394=>"101001011",
  63395=>"101101001",
  63396=>"111111101",
  63397=>"111000000",
  63398=>"110111111",
  63399=>"011111001",
  63400=>"111111111",
  63401=>"100100110",
  63402=>"111111111",
  63403=>"000000000",
  63404=>"000001000",
  63405=>"000000000",
  63406=>"111001000",
  63407=>"000001000",
  63408=>"111111001",
  63409=>"111111111",
  63410=>"111111011",
  63411=>"000010011",
  63412=>"110111111",
  63413=>"111111111",
  63414=>"000000000",
  63415=>"111111111",
  63416=>"111011111",
  63417=>"111111111",
  63418=>"110110101",
  63419=>"011111111",
  63420=>"111111111",
  63421=>"100100001",
  63422=>"111000000",
  63423=>"110111111",
  63424=>"000000000",
  63425=>"000110010",
  63426=>"111111111",
  63427=>"011111111",
  63428=>"000000111",
  63429=>"011001101",
  63430=>"000000000",
  63431=>"100000000",
  63432=>"111111000",
  63433=>"111000011",
  63434=>"111000101",
  63435=>"111111010",
  63436=>"011000000",
  63437=>"001001000",
  63438=>"111111101",
  63439=>"100000000",
  63440=>"100000000",
  63441=>"111111000",
  63442=>"111001010",
  63443=>"000000000",
  63444=>"100101110",
  63445=>"110110111",
  63446=>"010000000",
  63447=>"111000110",
  63448=>"111100000",
  63449=>"001111111",
  63450=>"111100111",
  63451=>"111101111",
  63452=>"011000100",
  63453=>"000000000",
  63454=>"100110111",
  63455=>"101111011",
  63456=>"110100000",
  63457=>"000000000",
  63458=>"000000111",
  63459=>"111111101",
  63460=>"111011111",
  63461=>"100100000",
  63462=>"111111000",
  63463=>"111111111",
  63464=>"000011010",
  63465=>"111101100",
  63466=>"100101101",
  63467=>"011111111",
  63468=>"111000111",
  63469=>"111111111",
  63470=>"000000000",
  63471=>"011011001",
  63472=>"100111111",
  63473=>"100000111",
  63474=>"111111111",
  63475=>"100100000",
  63476=>"000011111",
  63477=>"111111000",
  63478=>"000000001",
  63479=>"000010001",
  63480=>"101111111",
  63481=>"011111101",
  63482=>"110110110",
  63483=>"111111111",
  63484=>"111111111",
  63485=>"000000011",
  63486=>"000100100",
  63487=>"000000000",
  63488=>"000010111",
  63489=>"111101001",
  63490=>"000001111",
  63491=>"000000000",
  63492=>"110001000",
  63493=>"000000001",
  63494=>"000000000",
  63495=>"111111111",
  63496=>"011111111",
  63497=>"000000000",
  63498=>"010111111",
  63499=>"100100100",
  63500=>"100111011",
  63501=>"000000000",
  63502=>"000000001",
  63503=>"111111111",
  63504=>"000000000",
  63505=>"011000100",
  63506=>"001001001",
  63507=>"000000011",
  63508=>"111111111",
  63509=>"011001000",
  63510=>"111011111",
  63511=>"111111011",
  63512=>"110000000",
  63513=>"110110100",
  63514=>"111111111",
  63515=>"010000101",
  63516=>"010110111",
  63517=>"000000000",
  63518=>"000000000",
  63519=>"110111110",
  63520=>"111111111",
  63521=>"110100100",
  63522=>"111111111",
  63523=>"000000000",
  63524=>"111111111",
  63525=>"000000100",
  63526=>"111000011",
  63527=>"011100100",
  63528=>"110111111",
  63529=>"111111111",
  63530=>"000000000",
  63531=>"011110000",
  63532=>"111111111",
  63533=>"100000000",
  63534=>"111111110",
  63535=>"111100000",
  63536=>"000000000",
  63537=>"000100000",
  63538=>"011110000",
  63539=>"100111111",
  63540=>"111111100",
  63541=>"111111111",
  63542=>"000000000",
  63543=>"100000111",
  63544=>"000001011",
  63545=>"000000000",
  63546=>"111111111",
  63547=>"000000001",
  63548=>"001001000",
  63549=>"011111111",
  63550=>"000000000",
  63551=>"111111111",
  63552=>"000000100",
  63553=>"111111110",
  63554=>"111011011",
  63555=>"111111000",
  63556=>"111111011",
  63557=>"011010000",
  63558=>"111100111",
  63559=>"110000000",
  63560=>"000000000",
  63561=>"000000100",
  63562=>"111111111",
  63563=>"001001111",
  63564=>"000000110",
  63565=>"000000110",
  63566=>"111001000",
  63567=>"111111010",
  63568=>"110000000",
  63569=>"000000000",
  63570=>"000000000",
  63571=>"011011111",
  63572=>"010000100",
  63573=>"000000100",
  63574=>"111111111",
  63575=>"111111000",
  63576=>"111111111",
  63577=>"000000000",
  63578=>"000000111",
  63579=>"110010010",
  63580=>"111111111",
  63581=>"000000000",
  63582=>"111111111",
  63583=>"110111011",
  63584=>"100100000",
  63585=>"000000000",
  63586=>"100100110",
  63587=>"111000000",
  63588=>"011111000",
  63589=>"010000000",
  63590=>"000000000",
  63591=>"011001000",
  63592=>"000000000",
  63593=>"000111111",
  63594=>"001111111",
  63595=>"110100000",
  63596=>"000000000",
  63597=>"000000000",
  63598=>"110000000",
  63599=>"000000110",
  63600=>"000100100",
  63601=>"001111111",
  63602=>"000000000",
  63603=>"000000000",
  63604=>"111111111",
  63605=>"001111111",
  63606=>"000000000",
  63607=>"000100111",
  63608=>"100100000",
  63609=>"111110111",
  63610=>"001000000",
  63611=>"011000101",
  63612=>"100100100",
  63613=>"000000000",
  63614=>"000000000",
  63615=>"100100100",
  63616=>"000000000",
  63617=>"111111111",
  63618=>"111111111",
  63619=>"001101111",
  63620=>"011111111",
  63621=>"111111111",
  63622=>"000000000",
  63623=>"000000100",
  63624=>"111111000",
  63625=>"001000000",
  63626=>"111111111",
  63627=>"000000000",
  63628=>"000000000",
  63629=>"000000000",
  63630=>"111111111",
  63631=>"000010000",
  63632=>"011011110",
  63633=>"000000000",
  63634=>"110110100",
  63635=>"000000000",
  63636=>"000001001",
  63637=>"111011000",
  63638=>"111111111",
  63639=>"111001001",
  63640=>"000000001",
  63641=>"100000000",
  63642=>"110111011",
  63643=>"000000000",
  63644=>"111001111",
  63645=>"001001111",
  63646=>"100000000",
  63647=>"111000000",
  63648=>"111111111",
  63649=>"111001000",
  63650=>"110111111",
  63651=>"000000010",
  63652=>"000100111",
  63653=>"000100110",
  63654=>"100000101",
  63655=>"010110010",
  63656=>"001000000",
  63657=>"000000000",
  63658=>"000000000",
  63659=>"000111111",
  63660=>"111111001",
  63661=>"111111011",
  63662=>"000001001",
  63663=>"110001000",
  63664=>"000000000",
  63665=>"101110100",
  63666=>"111111111",
  63667=>"111111111",
  63668=>"111011010",
  63669=>"000111100",
  63670=>"111101101",
  63671=>"111000000",
  63672=>"111111111",
  63673=>"101111111",
  63674=>"111000000",
  63675=>"000000000",
  63676=>"000000000",
  63677=>"001111111",
  63678=>"001000000",
  63679=>"110111111",
  63680=>"111100000",
  63681=>"000000111",
  63682=>"011001000",
  63683=>"000000111",
  63684=>"000111111",
  63685=>"000000000",
  63686=>"011110111",
  63687=>"000000111",
  63688=>"001000000",
  63689=>"111111111",
  63690=>"001000000",
  63691=>"111111111",
  63692=>"111101111",
  63693=>"111111000",
  63694=>"011111111",
  63695=>"010000000",
  63696=>"100111111",
  63697=>"000000000",
  63698=>"111111101",
  63699=>"000000001",
  63700=>"100100111",
  63701=>"111111110",
  63702=>"000100110",
  63703=>"001000000",
  63704=>"000000100",
  63705=>"100000111",
  63706=>"000000000",
  63707=>"011000000",
  63708=>"111111000",
  63709=>"000000000",
  63710=>"111111111",
  63711=>"000001010",
  63712=>"111111010",
  63713=>"000110111",
  63714=>"111111000",
  63715=>"011111111",
  63716=>"000000000",
  63717=>"111100100",
  63718=>"111111111",
  63719=>"100000000",
  63720=>"000000000",
  63721=>"111111000",
  63722=>"000000011",
  63723=>"011001011",
  63724=>"110110110",
  63725=>"000000000",
  63726=>"111111111",
  63727=>"111111111",
  63728=>"110110100",
  63729=>"111111110",
  63730=>"000000011",
  63731=>"010111111",
  63732=>"111111111",
  63733=>"110110000",
  63734=>"000011111",
  63735=>"000000000",
  63736=>"011000000",
  63737=>"000000000",
  63738=>"000000000",
  63739=>"000000000",
  63740=>"000000000",
  63741=>"000100100",
  63742=>"001000000",
  63743=>"000011000",
  63744=>"111111111",
  63745=>"100100000",
  63746=>"100000000",
  63747=>"000000000",
  63748=>"110110111",
  63749=>"001111111",
  63750=>"000000100",
  63751=>"000000000",
  63752=>"000000001",
  63753=>"100000000",
  63754=>"111101101",
  63755=>"111111111",
  63756=>"111011111",
  63757=>"100000000",
  63758=>"101001111",
  63759=>"000000111",
  63760=>"000000110",
  63761=>"000110111",
  63762=>"110000001",
  63763=>"010000001",
  63764=>"000000001",
  63765=>"000000000",
  63766=>"001001001",
  63767=>"001001101",
  63768=>"111111111",
  63769=>"111111001",
  63770=>"010000000",
  63771=>"111000000",
  63772=>"111111011",
  63773=>"110110111",
  63774=>"000000000",
  63775=>"111111111",
  63776=>"111100100",
  63777=>"111111111",
  63778=>"111111111",
  63779=>"000001111",
  63780=>"000001001",
  63781=>"000000101",
  63782=>"100000000",
  63783=>"001001000",
  63784=>"000000000",
  63785=>"010000001",
  63786=>"111101101",
  63787=>"000000000",
  63788=>"111111111",
  63789=>"110111111",
  63790=>"001011011",
  63791=>"111111000",
  63792=>"000000011",
  63793=>"111111111",
  63794=>"111111111",
  63795=>"010011000",
  63796=>"110111111",
  63797=>"100100100",
  63798=>"001000000",
  63799=>"000000001",
  63800=>"000000100",
  63801=>"000001111",
  63802=>"111000000",
  63803=>"101111111",
  63804=>"000000000",
  63805=>"000000000",
  63806=>"011011000",
  63807=>"101110011",
  63808=>"111111000",
  63809=>"000111001",
  63810=>"111101111",
  63811=>"111111111",
  63812=>"111111110",
  63813=>"000000000",
  63814=>"100000000",
  63815=>"000000000",
  63816=>"000000000",
  63817=>"000001111",
  63818=>"111111111",
  63819=>"000000000",
  63820=>"000000000",
  63821=>"000100111",
  63822=>"111100111",
  63823=>"111111001",
  63824=>"011101000",
  63825=>"000000000",
  63826=>"011000010",
  63827=>"000000001",
  63828=>"000000111",
  63829=>"011011000",
  63830=>"000000000",
  63831=>"000000000",
  63832=>"111111111",
  63833=>"110110111",
  63834=>"111110000",
  63835=>"111110111",
  63836=>"001001011",
  63837=>"000000000",
  63838=>"111111111",
  63839=>"111111111",
  63840=>"010000000",
  63841=>"000000000",
  63842=>"000000110",
  63843=>"000000000",
  63844=>"110011001",
  63845=>"000000000",
  63846=>"111000000",
  63847=>"000000001",
  63848=>"000000000",
  63849=>"110111100",
  63850=>"110101111",
  63851=>"000000000",
  63852=>"110111111",
  63853=>"000000110",
  63854=>"000000000",
  63855=>"000000000",
  63856=>"000000000",
  63857=>"111001000",
  63858=>"000000110",
  63859=>"101111111",
  63860=>"000000000",
  63861=>"000000000",
  63862=>"011011111",
  63863=>"000000010",
  63864=>"001001001",
  63865=>"011011000",
  63866=>"001000100",
  63867=>"011011000",
  63868=>"100110111",
  63869=>"000000100",
  63870=>"000000000",
  63871=>"111111111",
  63872=>"100100111",
  63873=>"100000110",
  63874=>"000000000",
  63875=>"000000111",
  63876=>"000000110",
  63877=>"000111111",
  63878=>"010000111",
  63879=>"001000000",
  63880=>"000000000",
  63881=>"111110000",
  63882=>"111011011",
  63883=>"000000000",
  63884=>"110110111",
  63885=>"111111111",
  63886=>"000000101",
  63887=>"111111111",
  63888=>"000000000",
  63889=>"000000100",
  63890=>"111101000",
  63891=>"100000000",
  63892=>"011000000",
  63893=>"000010000",
  63894=>"111111101",
  63895=>"000000000",
  63896=>"111111100",
  63897=>"111111111",
  63898=>"000000111",
  63899=>"111101111",
  63900=>"111111110",
  63901=>"000100100",
  63902=>"011011001",
  63903=>"000000001",
  63904=>"011111111",
  63905=>"001011011",
  63906=>"110011111",
  63907=>"000000111",
  63908=>"000000001",
  63909=>"111100000",
  63910=>"110010111",
  63911=>"000000001",
  63912=>"000100100",
  63913=>"011110111",
  63914=>"000000110",
  63915=>"000000000",
  63916=>"000000000",
  63917=>"111101111",
  63918=>"000000110",
  63919=>"010111000",
  63920=>"111000000",
  63921=>"110100110",
  63922=>"000000000",
  63923=>"111110100",
  63924=>"111100101",
  63925=>"000001111",
  63926=>"000000000",
  63927=>"000011011",
  63928=>"111111000",
  63929=>"111111111",
  63930=>"000111111",
  63931=>"100000001",
  63932=>"001001000",
  63933=>"100100110",
  63934=>"101000000",
  63935=>"100100100",
  63936=>"000000000",
  63937=>"000000100",
  63938=>"010111000",
  63939=>"111111111",
  63940=>"101001111",
  63941=>"010000100",
  63942=>"001000101",
  63943=>"010110000",
  63944=>"000000101",
  63945=>"000000000",
  63946=>"000000000",
  63947=>"011001000",
  63948=>"000000000",
  63949=>"111000000",
  63950=>"111101111",
  63951=>"110010010",
  63952=>"000000000",
  63953=>"111100010",
  63954=>"110000100",
  63955=>"000011000",
  63956=>"111000000",
  63957=>"111111111",
  63958=>"000001011",
  63959=>"001100100",
  63960=>"111100110",
  63961=>"010000110",
  63962=>"110000000",
  63963=>"001000000",
  63964=>"101001100",
  63965=>"011001101",
  63966=>"111011111",
  63967=>"110010110",
  63968=>"100000100",
  63969=>"111111000",
  63970=>"000100110",
  63971=>"100100100",
  63972=>"000000000",
  63973=>"111111011",
  63974=>"001001011",
  63975=>"010000000",
  63976=>"000000000",
  63977=>"111111111",
  63978=>"111111100",
  63979=>"000000001",
  63980=>"000000000",
  63981=>"111111111",
  63982=>"111111111",
  63983=>"101000000",
  63984=>"000000000",
  63985=>"111011111",
  63986=>"110101101",
  63987=>"000000000",
  63988=>"111111111",
  63989=>"010111110",
  63990=>"111111110",
  63991=>"110110000",
  63992=>"000100100",
  63993=>"101101101",
  63994=>"011111111",
  63995=>"000000001",
  63996=>"000000110",
  63997=>"110000000",
  63998=>"111011101",
  63999=>"111110100",
  64000=>"111100100",
  64001=>"001000000",
  64002=>"111101111",
  64003=>"111111111",
  64004=>"110000000",
  64005=>"000100110",
  64006=>"111000101",
  64007=>"100100111",
  64008=>"000000100",
  64009=>"111111111",
  64010=>"111000000",
  64011=>"010110111",
  64012=>"000000000",
  64013=>"101111111",
  64014=>"010000000",
  64015=>"111111111",
  64016=>"011111000",
  64017=>"000010001",
  64018=>"000000000",
  64019=>"000010010",
  64020=>"111111001",
  64021=>"000000000",
  64022=>"000000000",
  64023=>"011001000",
  64024=>"110100000",
  64025=>"111110111",
  64026=>"100000000",
  64027=>"000000100",
  64028=>"111111000",
  64029=>"111111001",
  64030=>"110100000",
  64031=>"000001011",
  64032=>"000110000",
  64033=>"100000000",
  64034=>"001000000",
  64035=>"111111111",
  64036=>"000000111",
  64037=>"111110111",
  64038=>"000100111",
  64039=>"100100000",
  64040=>"111111000",
  64041=>"001101100",
  64042=>"000100000",
  64043=>"000000000",
  64044=>"000000000",
  64045=>"111111111",
  64046=>"111111001",
  64047=>"111111111",
  64048=>"000000000",
  64049=>"001011010",
  64050=>"111111001",
  64051=>"000000000",
  64052=>"011011001",
  64053=>"001001001",
  64054=>"000000100",
  64055=>"100111111",
  64056=>"000100000",
  64057=>"000110111",
  64058=>"111111000",
  64059=>"111111111",
  64060=>"100000110",
  64061=>"000000100",
  64062=>"111111111",
  64063=>"000000000",
  64064=>"011011011",
  64065=>"010010010",
  64066=>"111000000",
  64067=>"110110111",
  64068=>"001000000",
  64069=>"110110111",
  64070=>"000000000",
  64071=>"111111001",
  64072=>"011111111",
  64073=>"111000111",
  64074=>"000000000",
  64075=>"001000001",
  64076=>"000111010",
  64077=>"111111111",
  64078=>"000100000",
  64079=>"111111111",
  64080=>"001001011",
  64081=>"110000000",
  64082=>"000000111",
  64083=>"101000111",
  64084=>"000000100",
  64085=>"111011100",
  64086=>"101101000",
  64087=>"000000100",
  64088=>"111111000",
  64089=>"000000000",
  64090=>"100010000",
  64091=>"110111110",
  64092=>"111000000",
  64093=>"101100001",
  64094=>"111111110",
  64095=>"111011001",
  64096=>"111111110",
  64097=>"000000011",
  64098=>"000000000",
  64099=>"111111111",
  64100=>"000000001",
  64101=>"000001001",
  64102=>"000110111",
  64103=>"001111000",
  64104=>"111010000",
  64105=>"111111100",
  64106=>"110110100",
  64107=>"110110000",
  64108=>"001100000",
  64109=>"111101111",
  64110=>"111111111",
  64111=>"111111111",
  64112=>"000000000",
  64113=>"000110010",
  64114=>"000000000",
  64115=>"111001000",
  64116=>"000000000",
  64117=>"111011011",
  64118=>"000000010",
  64119=>"000111111",
  64120=>"000000001",
  64121=>"111111111",
  64122=>"001001001",
  64123=>"000111000",
  64124=>"100110110",
  64125=>"000000000",
  64126=>"001000100",
  64127=>"000000000",
  64128=>"100111111",
  64129=>"011111111",
  64130=>"111111110",
  64131=>"000000000",
  64132=>"100000001",
  64133=>"000000000",
  64134=>"000000000",
  64135=>"111000000",
  64136=>"000000000",
  64137=>"000000000",
  64138=>"111111111",
  64139=>"000100000",
  64140=>"110111101",
  64141=>"000000000",
  64142=>"111111000",
  64143=>"000000000",
  64144=>"111111111",
  64145=>"110000000",
  64146=>"000000011",
  64147=>"111011111",
  64148=>"110010000",
  64149=>"111111100",
  64150=>"001000000",
  64151=>"111111111",
  64152=>"000000110",
  64153=>"111111111",
  64154=>"000000100",
  64155=>"011001000",
  64156=>"111111011",
  64157=>"111111111",
  64158=>"111000000",
  64159=>"000000000",
  64160=>"000010000",
  64161=>"111111111",
  64162=>"000000000",
  64163=>"100000000",
  64164=>"011111111",
  64165=>"100111111",
  64166=>"000001111",
  64167=>"011011000",
  64168=>"111111111",
  64169=>"000000000",
  64170=>"000000100",
  64171=>"001001111",
  64172=>"111111100",
  64173=>"001000000",
  64174=>"000000000",
  64175=>"000001001",
  64176=>"111111111",
  64177=>"100111111",
  64178=>"000010000",
  64179=>"110101100",
  64180=>"101100000",
  64181=>"111111111",
  64182=>"111111111",
  64183=>"100000000",
  64184=>"111000000",
  64185=>"111111111",
  64186=>"100100100",
  64187=>"000110110",
  64188=>"100100000",
  64189=>"111111111",
  64190=>"000100111",
  64191=>"000011011",
  64192=>"111111111",
  64193=>"001001111",
  64194=>"111111000",
  64195=>"000000000",
  64196=>"000000111",
  64197=>"001101111",
  64198=>"000001001",
  64199=>"000010010",
  64200=>"111110000",
  64201=>"000000000",
  64202=>"000000010",
  64203=>"111100111",
  64204=>"000000111",
  64205=>"000111111",
  64206=>"100000100",
  64207=>"111100000",
  64208=>"111111101",
  64209=>"111111111",
  64210=>"111111100",
  64211=>"111111111",
  64212=>"001000001",
  64213=>"001010000",
  64214=>"000000111",
  64215=>"000000000",
  64216=>"111011000",
  64217=>"111111111",
  64218=>"111011011",
  64219=>"010010000",
  64220=>"111111111",
  64221=>"010000011",
  64222=>"000000000",
  64223=>"110111100",
  64224=>"010010010",
  64225=>"011110000",
  64226=>"000000111",
  64227=>"000000111",
  64228=>"000101111",
  64229=>"111111111",
  64230=>"111111111",
  64231=>"110100000",
  64232=>"000000000",
  64233=>"111111111",
  64234=>"111111011",
  64235=>"001111111",
  64236=>"111111111",
  64237=>"000011111",
  64238=>"000100111",
  64239=>"010111111",
  64240=>"100000001",
  64241=>"000001111",
  64242=>"000110110",
  64243=>"110000000",
  64244=>"100111100",
  64245=>"111011011",
  64246=>"010000000",
  64247=>"000000000",
  64248=>"001001001",
  64249=>"001001011",
  64250=>"000000000",
  64251=>"000100101",
  64252=>"011110100",
  64253=>"000000000",
  64254=>"111110000",
  64255=>"111111001",
  64256=>"100000000",
  64257=>"011011011",
  64258=>"110000111",
  64259=>"111111111",
  64260=>"110111111",
  64261=>"101101111",
  64262=>"111111111",
  64263=>"100100000",
  64264=>"001010000",
  64265=>"000000000",
  64266=>"101000100",
  64267=>"100100000",
  64268=>"100100111",
  64269=>"000110000",
  64270=>"101011111",
  64271=>"100111111",
  64272=>"000000111",
  64273=>"000000000",
  64274=>"111000000",
  64275=>"001100000",
  64276=>"000111000",
  64277=>"000001001",
  64278=>"000110000",
  64279=>"111111101",
  64280=>"110000000",
  64281=>"111111111",
  64282=>"000000000",
  64283=>"000111111",
  64284=>"111111111",
  64285=>"111111110",
  64286=>"000000000",
  64287=>"000000000",
  64288=>"111111111",
  64289=>"111111000",
  64290=>"000000000",
  64291=>"101111111",
  64292=>"000100100",
  64293=>"011010000",
  64294=>"110111011",
  64295=>"111001111",
  64296=>"000111111",
  64297=>"000000000",
  64298=>"000000000",
  64299=>"111111001",
  64300=>"111111111",
  64301=>"100100101",
  64302=>"111111000",
  64303=>"111111111",
  64304=>"100101111",
  64305=>"101000000",
  64306=>"001111111",
  64307=>"111110000",
  64308=>"000000111",
  64309=>"111011001",
  64310=>"000110010",
  64311=>"000000000",
  64312=>"011000000",
  64313=>"001000000",
  64314=>"001111111",
  64315=>"001110000",
  64316=>"111111111",
  64317=>"000000000",
  64318=>"111111111",
  64319=>"111111111",
  64320=>"001001000",
  64321=>"001001011",
  64322=>"001111111",
  64323=>"111111111",
  64324=>"111111111",
  64325=>"010010000",
  64326=>"001100111",
  64327=>"100100000",
  64328=>"000000111",
  64329=>"000010111",
  64330=>"000000000",
  64331=>"000001001",
  64332=>"111011111",
  64333=>"010000000",
  64334=>"111111100",
  64335=>"000110111",
  64336=>"001111111",
  64337=>"000000100",
  64338=>"110000000",
  64339=>"000111111",
  64340=>"101101000",
  64341=>"001001011",
  64342=>"111111111",
  64343=>"000100100",
  64344=>"000101111",
  64345=>"111111011",
  64346=>"111010000",
  64347=>"010010000",
  64348=>"000000000",
  64349=>"111111111",
  64350=>"100100000",
  64351=>"001000000",
  64352=>"000001111",
  64353=>"111110000",
  64354=>"000000000",
  64355=>"000000101",
  64356=>"111111110",
  64357=>"011000010",
  64358=>"111111010",
  64359=>"111111111",
  64360=>"000100000",
  64361=>"001001000",
  64362=>"001011000",
  64363=>"000000001",
  64364=>"000001000",
  64365=>"111111111",
  64366=>"111111010",
  64367=>"000000000",
  64368=>"000000011",
  64369=>"000000101",
  64370=>"000000000",
  64371=>"100110110",
  64372=>"000000110",
  64373=>"111111111",
  64374=>"000000000",
  64375=>"000000000",
  64376=>"001111111",
  64377=>"111111000",
  64378=>"000100000",
  64379=>"000001111",
  64380=>"111111011",
  64381=>"111111001",
  64382=>"110100000",
  64383=>"111111111",
  64384=>"000000000",
  64385=>"011000011",
  64386=>"011111111",
  64387=>"000000000",
  64388=>"000000111",
  64389=>"111111111",
  64390=>"000000011",
  64391=>"110111111",
  64392=>"111001000",
  64393=>"001000000",
  64394=>"000000000",
  64395=>"000000111",
  64396=>"111111111",
  64397=>"110111111",
  64398=>"101001111",
  64399=>"111000100",
  64400=>"000000000",
  64401=>"111111111",
  64402=>"110010100",
  64403=>"100110111",
  64404=>"000000000",
  64405=>"000110111",
  64406=>"100000000",
  64407=>"000000000",
  64408=>"011001000",
  64409=>"000000000",
  64410=>"111010111",
  64411=>"000000000",
  64412=>"000010111",
  64413=>"000111111",
  64414=>"100000001",
  64415=>"011111111",
  64416=>"111111111",
  64417=>"110110111",
  64418=>"000001001",
  64419=>"010000000",
  64420=>"000000000",
  64421=>"111111111",
  64422=>"100000000",
  64423=>"111111010",
  64424=>"110010110",
  64425=>"000000100",
  64426=>"111111100",
  64427=>"000000000",
  64428=>"000000000",
  64429=>"000000100",
  64430=>"000011011",
  64431=>"100110000",
  64432=>"111111111",
  64433=>"000100110",
  64434=>"111111111",
  64435=>"000000000",
  64436=>"100101111",
  64437=>"000000100",
  64438=>"000000000",
  64439=>"110000000",
  64440=>"111111111",
  64441=>"101001000",
  64442=>"000000000",
  64443=>"111111110",
  64444=>"000111111",
  64445=>"111101001",
  64446=>"111111111",
  64447=>"001000000",
  64448=>"000000000",
  64449=>"000000000",
  64450=>"000000010",
  64451=>"111101000",
  64452=>"011111101",
  64453=>"000000011",
  64454=>"110001111",
  64455=>"000000000",
  64456=>"111000000",
  64457=>"111111111",
  64458=>"000100110",
  64459=>"111111000",
  64460=>"011111000",
  64461=>"001000000",
  64462=>"000000000",
  64463=>"111111111",
  64464=>"000111111",
  64465=>"100001000",
  64466=>"111111010",
  64467=>"011000000",
  64468=>"000000000",
  64469=>"110110000",
  64470=>"000000000",
  64471=>"110110100",
  64472=>"000000000",
  64473=>"000111111",
  64474=>"001111111",
  64475=>"110011000",
  64476=>"011111100",
  64477=>"000000000",
  64478=>"111111111",
  64479=>"001000100",
  64480=>"111111000",
  64481=>"111011011",
  64482=>"000000110",
  64483=>"100100000",
  64484=>"111000001",
  64485=>"111111101",
  64486=>"000000000",
  64487=>"000000000",
  64488=>"110110111",
  64489=>"000000110",
  64490=>"100000000",
  64491=>"001001111",
  64492=>"000000000",
  64493=>"000000000",
  64494=>"111010000",
  64495=>"000111111",
  64496=>"111111111",
  64497=>"110111111",
  64498=>"000000000",
  64499=>"000000000",
  64500=>"111111111",
  64501=>"100101111",
  64502=>"000110100",
  64503=>"110111111",
  64504=>"111111011",
  64505=>"000010100",
  64506=>"000000000",
  64507=>"000110100",
  64508=>"000000001",
  64509=>"000000000",
  64510=>"000000000",
  64511=>"000000000",
  64512=>"110111111",
  64513=>"111111111",
  64514=>"111111111",
  64515=>"000000000",
  64516=>"011011011",
  64517=>"000000111",
  64518=>"011001011",
  64519=>"111101111",
  64520=>"000000001",
  64521=>"000000000",
  64522=>"001001000",
  64523=>"000110111",
  64524=>"110110110",
  64525=>"000100101",
  64526=>"000110000",
  64527=>"000000000",
  64528=>"110011001",
  64529=>"000110111",
  64530=>"001001000",
  64531=>"000000000",
  64532=>"111111111",
  64533=>"000000000",
  64534=>"111100000",
  64535=>"011000110",
  64536=>"001000001",
  64537=>"011100110",
  64538=>"001111100",
  64539=>"010000110",
  64540=>"111111110",
  64541=>"000100100",
  64542=>"001001001",
  64543=>"000011111",
  64544=>"111111111",
  64545=>"111111000",
  64546=>"100110011",
  64547=>"111111111",
  64548=>"001000000",
  64549=>"000000000",
  64550=>"000000000",
  64551=>"000000000",
  64552=>"111000000",
  64553=>"111111111",
  64554=>"111111111",
  64555=>"000000000",
  64556=>"000000100",
  64557=>"000111111",
  64558=>"111111111",
  64559=>"111111110",
  64560=>"000000001",
  64561=>"101100111",
  64562=>"111111111",
  64563=>"000100100",
  64564=>"111111111",
  64565=>"110110100",
  64566=>"111001011",
  64567=>"000000000",
  64568=>"111111111",
  64569=>"110100000",
  64570=>"101100111",
  64571=>"111110111",
  64572=>"111111111",
  64573=>"011001011",
  64574=>"111111111",
  64575=>"000000000",
  64576=>"111110110",
  64577=>"000000111",
  64578=>"000111110",
  64579=>"000111111",
  64580=>"000010011",
  64581=>"001001110",
  64582=>"011000000",
  64583=>"000000000",
  64584=>"001001000",
  64585=>"110000000",
  64586=>"000000000",
  64587=>"000000000",
  64588=>"111100110",
  64589=>"000000111",
  64590=>"001000000",
  64591=>"000000110",
  64592=>"111111111",
  64593=>"111000000",
  64594=>"101100100",
  64595=>"000101111",
  64596=>"000000000",
  64597=>"000000000",
  64598=>"101100000",
  64599=>"111111111",
  64600=>"000000001",
  64601=>"000000110",
  64602=>"101000000",
  64603=>"110110110",
  64604=>"001000001",
  64605=>"111111011",
  64606=>"000101111",
  64607=>"000000000",
  64608=>"100000000",
  64609=>"100101000",
  64610=>"111111011",
  64611=>"000000000",
  64612=>"000000000",
  64613=>"010000111",
  64614=>"100110111",
  64615=>"000001001",
  64616=>"111111111",
  64617=>"000000111",
  64618=>"000000000",
  64619=>"111111011",
  64620=>"011111111",
  64621=>"000000000",
  64622=>"111111111",
  64623=>"111111101",
  64624=>"011000110",
  64625=>"100111111",
  64626=>"010000000",
  64627=>"000000001",
  64628=>"111100000",
  64629=>"000000110",
  64630=>"111111111",
  64631=>"001001000",
  64632=>"010110111",
  64633=>"111111111",
  64634=>"000000000",
  64635=>"111111111",
  64636=>"000000000",
  64637=>"111001000",
  64638=>"000000000",
  64639=>"000000000",
  64640=>"111111111",
  64641=>"111110100",
  64642=>"110000000",
  64643=>"001000000",
  64644=>"100100111",
  64645=>"000000000",
  64646=>"001000110",
  64647=>"000000000",
  64648=>"111111001",
  64649=>"001000110",
  64650=>"000110110",
  64651=>"011111111",
  64652=>"000010000",
  64653=>"000000000",
  64654=>"011111111",
  64655=>"111111101",
  64656=>"111111011",
  64657=>"100110111",
  64658=>"111000101",
  64659=>"111110000",
  64660=>"101111111",
  64661=>"111111111",
  64662=>"111111111",
  64663=>"000000000",
  64664=>"110111111",
  64665=>"111111000",
  64666=>"011011011",
  64667=>"111111111",
  64668=>"111111111",
  64669=>"111111001",
  64670=>"000000000",
  64671=>"111011001",
  64672=>"111111111",
  64673=>"000100100",
  64674=>"101111100",
  64675=>"000000000",
  64676=>"000000000",
  64677=>"000000110",
  64678=>"000000001",
  64679=>"000000001",
  64680=>"011001111",
  64681=>"100101111",
  64682=>"000000000",
  64683=>"111110110",
  64684=>"111000000",
  64685=>"110110100",
  64686=>"111111111",
  64687=>"101100100",
  64688=>"000000000",
  64689=>"011011111",
  64690=>"000011001",
  64691=>"000010110",
  64692=>"100100000",
  64693=>"111111010",
  64694=>"000000000",
  64695=>"111111111",
  64696=>"011010000",
  64697=>"110000010",
  64698=>"000000000",
  64699=>"000000111",
  64700=>"000000100",
  64701=>"111111111",
  64702=>"011000000",
  64703=>"000000000",
  64704=>"111100110",
  64705=>"001001001",
  64706=>"011000000",
  64707=>"111000000",
  64708=>"101111100",
  64709=>"111111111",
  64710=>"111111111",
  64711=>"000011000",
  64712=>"000000000",
  64713=>"111111111",
  64714=>"111110110",
  64715=>"000000000",
  64716=>"111111111",
  64717=>"111001000",
  64718=>"011111111",
  64719=>"111111111",
  64720=>"001111000",
  64721=>"100000000",
  64722=>"011111111",
  64723=>"000000001",
  64724=>"011100000",
  64725=>"001101111",
  64726=>"111111111",
  64727=>"001001111",
  64728=>"110111111",
  64729=>"110000000",
  64730=>"000000000",
  64731=>"000000000",
  64732=>"111111111",
  64733=>"001000000",
  64734=>"000000000",
  64735=>"111111111",
  64736=>"001001111",
  64737=>"000000111",
  64738=>"111100000",
  64739=>"011011011",
  64740=>"111111110",
  64741=>"001101101",
  64742=>"000000000",
  64743=>"001111111",
  64744=>"100100111",
  64745=>"000000100",
  64746=>"111111111",
  64747=>"001101111",
  64748=>"010010000",
  64749=>"100000110",
  64750=>"000000101",
  64751=>"111010000",
  64752=>"000110000",
  64753=>"100000000",
  64754=>"111111111",
  64755=>"000000000",
  64756=>"111111111",
  64757=>"010110010",
  64758=>"110000000",
  64759=>"000011000",
  64760=>"010000000",
  64761=>"111111111",
  64762=>"001111000",
  64763=>"001011000",
  64764=>"101100000",
  64765=>"111110000",
  64766=>"000000000",
  64767=>"111101000",
  64768=>"010010010",
  64769=>"111011011",
  64770=>"000001001",
  64771=>"111011101",
  64772=>"100100111",
  64773=>"000000001",
  64774=>"000000000",
  64775=>"111110000",
  64776=>"111111111",
  64777=>"111110110",
  64778=>"111111111",
  64779=>"111111111",
  64780=>"000000000",
  64781=>"000110110",
  64782=>"100011111",
  64783=>"001011111",
  64784=>"110000000",
  64785=>"011111000",
  64786=>"100111000",
  64787=>"111111111",
  64788=>"111011000",
  64789=>"000000000",
  64790=>"111111011",
  64791=>"111111011",
  64792=>"000000000",
  64793=>"000000000",
  64794=>"001000000",
  64795=>"111111111",
  64796=>"100110110",
  64797=>"000000111",
  64798=>"111111111",
  64799=>"100111111",
  64800=>"000000010",
  64801=>"000001011",
  64802=>"100100111",
  64803=>"000000111",
  64804=>"111111111",
  64805=>"111111000",
  64806=>"011111111",
  64807=>"000000000",
  64808=>"111111111",
  64809=>"000000111",
  64810=>"110111111",
  64811=>"000000000",
  64812=>"000000111",
  64813=>"000100111",
  64814=>"111111111",
  64815=>"000000000",
  64816=>"111111111",
  64817=>"011111111",
  64818=>"111111110",
  64819=>"100111101",
  64820=>"111111011",
  64821=>"011011011",
  64822=>"000100111",
  64823=>"100100000",
  64824=>"000000100",
  64825=>"000000000",
  64826=>"000000000",
  64827=>"111111111",
  64828=>"111111111",
  64829=>"111111000",
  64830=>"100000000",
  64831=>"110110111",
  64832=>"111111111",
  64833=>"111111111",
  64834=>"101111111",
  64835=>"111110111",
  64836=>"000000000",
  64837=>"111111111",
  64838=>"111111111",
  64839=>"000000000",
  64840=>"000000000",
  64841=>"011111111",
  64842=>"110110111",
  64843=>"100100000",
  64844=>"011111011",
  64845=>"111111111",
  64846=>"111100000",
  64847=>"110100100",
  64848=>"011001001",
  64849=>"111011010",
  64850=>"111111001",
  64851=>"000000000",
  64852=>"000000000",
  64853=>"010011111",
  64854=>"000000000",
  64855=>"111100000",
  64856=>"111111111",
  64857=>"100111101",
  64858=>"111111000",
  64859=>"000000000",
  64860=>"111111111",
  64861=>"110111111",
  64862=>"110000000",
  64863=>"011111111",
  64864=>"000100100",
  64865=>"000000000",
  64866=>"010000000",
  64867=>"000000000",
  64868=>"111111110",
  64869=>"111111111",
  64870=>"000101001",
  64871=>"110110110",
  64872=>"111111000",
  64873=>"000010000",
  64874=>"111111111",
  64875=>"111111110",
  64876=>"011001001",
  64877=>"000001000",
  64878=>"001000000",
  64879=>"111001000",
  64880=>"000000000",
  64881=>"111111111",
  64882=>"010000000",
  64883=>"000000000",
  64884=>"100000000",
  64885=>"101111111",
  64886=>"101001000",
  64887=>"110100100",
  64888=>"111111111",
  64889=>"001001000",
  64890=>"000000000",
  64891=>"000000000",
  64892=>"000100000",
  64893=>"001000001",
  64894=>"111111111",
  64895=>"111111111",
  64896=>"111111011",
  64897=>"000000001",
  64898=>"000000001",
  64899=>"100100111",
  64900=>"111111011",
  64901=>"000000000",
  64902=>"011011111",
  64903=>"010011101",
  64904=>"000111111",
  64905=>"111111011",
  64906=>"110111111",
  64907=>"000000000",
  64908=>"000000100",
  64909=>"110110000",
  64910=>"000101111",
  64911=>"111111111",
  64912=>"000100011",
  64913=>"111111111",
  64914=>"111111000",
  64915=>"111111111",
  64916=>"000000000",
  64917=>"000000111",
  64918=>"111110000",
  64919=>"011011000",
  64920=>"000000000",
  64921=>"110110000",
  64922=>"000111111",
  64923=>"000101111",
  64924=>"000000000",
  64925=>"101111111",
  64926=>"011001000",
  64927=>"011111111",
  64928=>"110111111",
  64929=>"001001001",
  64930=>"101101111",
  64931=>"111111100",
  64932=>"000000000",
  64933=>"000000000",
  64934=>"101000100",
  64935=>"000110110",
  64936=>"111111111",
  64937=>"000000101",
  64938=>"000000000",
  64939=>"000000000",
  64940=>"001000000",
  64941=>"111111111",
  64942=>"000001000",
  64943=>"010111111",
  64944=>"111111110",
  64945=>"101000000",
  64946=>"111011011",
  64947=>"000000010",
  64948=>"000101101",
  64949=>"101111111",
  64950=>"111111100",
  64951=>"111101001",
  64952=>"111111111",
  64953=>"111001000",
  64954=>"011000001",
  64955=>"111111111",
  64956=>"011111111",
  64957=>"111000100",
  64958=>"000000000",
  64959=>"110000000",
  64960=>"000000010",
  64961=>"111111000",
  64962=>"000000000",
  64963=>"111111111",
  64964=>"011000001",
  64965=>"001000000",
  64966=>"001111111",
  64967=>"101000000",
  64968=>"001000000",
  64969=>"110111110",
  64970=>"000000100",
  64971=>"000000000",
  64972=>"000000000",
  64973=>"111111111",
  64974=>"000000000",
  64975=>"111101100",
  64976=>"000000100",
  64977=>"111110111",
  64978=>"000000000",
  64979=>"111111111",
  64980=>"111110111",
  64981=>"011111111",
  64982=>"111111111",
  64983=>"100100100",
  64984=>"000000100",
  64985=>"111111010",
  64986=>"111111111",
  64987=>"111000000",
  64988=>"111111000",
  64989=>"000000000",
  64990=>"111011001",
  64991=>"111000000",
  64992=>"111111100",
  64993=>"010001011",
  64994=>"010111111",
  64995=>"011000000",
  64996=>"000000000",
  64997=>"111111011",
  64998=>"000000010",
  64999=>"000101101",
  65000=>"000100000",
  65001=>"001111010",
  65002=>"011011000",
  65003=>"111110100",
  65004=>"001000111",
  65005=>"111111011",
  65006=>"011011011",
  65007=>"000000000",
  65008=>"000000000",
  65009=>"111010000",
  65010=>"111111111",
  65011=>"111111111",
  65012=>"000110000",
  65013=>"000000110",
  65014=>"011000000",
  65015=>"000000000",
  65016=>"111111111",
  65017=>"011001001",
  65018=>"110100111",
  65019=>"101101000",
  65020=>"111111111",
  65021=>"110110001",
  65022=>"111111110",
  65023=>"000000000",
  65024=>"000000000",
  65025=>"001111111",
  65026=>"000000000",
  65027=>"000110000",
  65028=>"000001111",
  65029=>"111011001",
  65030=>"001000000",
  65031=>"000000000",
  65032=>"110111111",
  65033=>"000111111",
  65034=>"011010001",
  65035=>"000000000",
  65036=>"100110110",
  65037=>"111110000",
  65038=>"101001101",
  65039=>"000000000",
  65040=>"111000000",
  65041=>"000011001",
  65042=>"110110000",
  65043=>"000010110",
  65044=>"000000000",
  65045=>"001111111",
  65046=>"011111111",
  65047=>"011011000",
  65048=>"001001001",
  65049=>"001001001",
  65050=>"011000000",
  65051=>"011111101",
  65052=>"001000000",
  65053=>"000000010",
  65054=>"011011010",
  65055=>"101101110",
  65056=>"111011111",
  65057=>"110000000",
  65058=>"111111100",
  65059=>"000000000",
  65060=>"100000000",
  65061=>"000100000",
  65062=>"100000000",
  65063=>"000101101",
  65064=>"111111101",
  65065=>"000000101",
  65066=>"001000000",
  65067=>"000000000",
  65068=>"111111000",
  65069=>"111011000",
  65070=>"001000000",
  65071=>"000000000",
  65072=>"000010111",
  65073=>"000000000",
  65074=>"100110100",
  65075=>"111010000",
  65076=>"000000000",
  65077=>"110111011",
  65078=>"000000111",
  65079=>"000000111",
  65080=>"111111111",
  65081=>"111011111",
  65082=>"000000001",
  65083=>"100000000",
  65084=>"011000111",
  65085=>"111111111",
  65086=>"111110100",
  65087=>"100111111",
  65088=>"001001001",
  65089=>"011111000",
  65090=>"111111111",
  65091=>"111000000",
  65092=>"111111111",
  65093=>"000001111",
  65094=>"111000000",
  65095=>"111001011",
  65096=>"100001001",
  65097=>"000000000",
  65098=>"111111111",
  65099=>"000000010",
  65100=>"111111111",
  65101=>"001101111",
  65102=>"000000000",
  65103=>"001000011",
  65104=>"100111000",
  65105=>"111010000",
  65106=>"101010001",
  65107=>"001001001",
  65108=>"000000000",
  65109=>"111111111",
  65110=>"000101111",
  65111=>"011001101",
  65112=>"001111111",
  65113=>"111000111",
  65114=>"111101111",
  65115=>"110110111",
  65116=>"100000101",
  65117=>"100101111",
  65118=>"000010111",
  65119=>"111010001",
  65120=>"000000000",
  65121=>"111110110",
  65122=>"101101101",
  65123=>"111101100",
  65124=>"000000000",
  65125=>"000000111",
  65126=>"111111001",
  65127=>"111111111",
  65128=>"111000000",
  65129=>"111100000",
  65130=>"111111111",
  65131=>"111111000",
  65132=>"011011011",
  65133=>"100000000",
  65134=>"111111110",
  65135=>"000101111",
  65136=>"111111000",
  65137=>"100000000",
  65138=>"001001001",
  65139=>"111101101",
  65140=>"000001000",
  65141=>"000001111",
  65142=>"000000000",
  65143=>"100000000",
  65144=>"000000000",
  65145=>"100000000",
  65146=>"001001000",
  65147=>"000000000",
  65148=>"101001011",
  65149=>"000101111",
  65150=>"111011000",
  65151=>"000111111",
  65152=>"000000000",
  65153=>"100000000",
  65154=>"000111111",
  65155=>"100000000",
  65156=>"000000111",
  65157=>"000000111",
  65158=>"111101000",
  65159=>"000000000",
  65160=>"111111011",
  65161=>"111111000",
  65162=>"000000000",
  65163=>"111111011",
  65164=>"000111111",
  65165=>"111111110",
  65166=>"000000000",
  65167=>"000000000",
  65168=>"000001000",
  65169=>"001101101",
  65170=>"101100101",
  65171=>"001001000",
  65172=>"111111000",
  65173=>"101010010",
  65174=>"111111111",
  65175=>"011011011",
  65176=>"000000001",
  65177=>"000100000",
  65178=>"111000000",
  65179=>"111111110",
  65180=>"100110111",
  65181=>"000000001",
  65182=>"111101111",
  65183=>"000000000",
  65184=>"111111111",
  65185=>"111101000",
  65186=>"000000111",
  65187=>"111111110",
  65188=>"111111001",
  65189=>"111000000",
  65190=>"111111111",
  65191=>"111111101",
  65192=>"001000001",
  65193=>"100000110",
  65194=>"111111111",
  65195=>"111111111",
  65196=>"101000001",
  65197=>"111001000",
  65198=>"111010000",
  65199=>"101111000",
  65200=>"111011000",
  65201=>"000000000",
  65202=>"100101100",
  65203=>"011101111",
  65204=>"000000000",
  65205=>"111001110",
  65206=>"111111111",
  65207=>"000000000",
  65208=>"111111000",
  65209=>"100111111",
  65210=>"101101111",
  65211=>"011011111",
  65212=>"000000000",
  65213=>"000100000",
  65214=>"111000000",
  65215=>"011111111",
  65216=>"011011110",
  65217=>"000000111",
  65218=>"011001001",
  65219=>"000111111",
  65220=>"000000000",
  65221=>"111111111",
  65222=>"111111000",
  65223=>"111111111",
  65224=>"110110111",
  65225=>"001000110",
  65226=>"111111111",
  65227=>"000000111",
  65228=>"111111000",
  65229=>"000111111",
  65230=>"011000000",
  65231=>"001000100",
  65232=>"000000111",
  65233=>"101111111",
  65234=>"111111000",
  65235=>"011000000",
  65236=>"000000000",
  65237=>"110100111",
  65238=>"000110111",
  65239=>"000000000",
  65240=>"111111011",
  65241=>"101000111",
  65242=>"011111111",
  65243=>"011000000",
  65244=>"001000001",
  65245=>"111100000",
  65246=>"011100100",
  65247=>"000000001",
  65248=>"110000000",
  65249=>"000001101",
  65250=>"111111111",
  65251=>"001000000",
  65252=>"000110111",
  65253=>"111110110",
  65254=>"111111110",
  65255=>"111110100",
  65256=>"000001001",
  65257=>"000000001",
  65258=>"001000111",
  65259=>"111011111",
  65260=>"000000000",
  65261=>"000000111",
  65262=>"111111000",
  65263=>"100111111",
  65264=>"000110110",
  65265=>"111111111",
  65266=>"111001000",
  65267=>"111000111",
  65268=>"001111111",
  65269=>"011000001",
  65270=>"111111000",
  65271=>"111000001",
  65272=>"001111000",
  65273=>"111111111",
  65274=>"111001111",
  65275=>"000010011",
  65276=>"100000011",
  65277=>"111110110",
  65278=>"111000000",
  65279=>"100000000",
  65280=>"001000000",
  65281=>"011011111",
  65282=>"010011111",
  65283=>"111111100",
  65284=>"001011000",
  65285=>"011011111",
  65286=>"000000000",
  65287=>"001111111",
  65288=>"111111111",
  65289=>"111110100",
  65290=>"111100000",
  65291=>"000000000",
  65292=>"100000000",
  65293=>"111000000",
  65294=>"111110110",
  65295=>"111010000",
  65296=>"111100000",
  65297=>"011001001",
  65298=>"011000000",
  65299=>"110110110",
  65300=>"111111011",
  65301=>"100100101",
  65302=>"111011001",
  65303=>"101101000",
  65304=>"100110010",
  65305=>"111111111",
  65306=>"000101101",
  65307=>"000000111",
  65308=>"011100100",
  65309=>"000111111",
  65310=>"111111011",
  65311=>"111001111",
  65312=>"111111011",
  65313=>"111000000",
  65314=>"000000000",
  65315=>"101001011",
  65316=>"000000000",
  65317=>"111111111",
  65318=>"111111111",
  65319=>"111100100",
  65320=>"000000000",
  65321=>"000100100",
  65322=>"000100110",
  65323=>"001000000",
  65324=>"111110111",
  65325=>"000110100",
  65326=>"111110111",
  65327=>"000000101",
  65328=>"101100000",
  65329=>"011111111",
  65330=>"001000000",
  65331=>"000000111",
  65332=>"100101011",
  65333=>"100100000",
  65334=>"111111000",
  65335=>"111110100",
  65336=>"111111001",
  65337=>"111000000",
  65338=>"111110100",
  65339=>"000000111",
  65340=>"000000111",
  65341=>"101100000",
  65342=>"101111111",
  65343=>"011111110",
  65344=>"001111000",
  65345=>"000000100",
  65346=>"111111111",
  65347=>"000010111",
  65348=>"001001000",
  65349=>"111111000",
  65350=>"000000000",
  65351=>"111111000",
  65352=>"111000000",
  65353=>"111111111",
  65354=>"111111011",
  65355=>"000100100",
  65356=>"111111000",
  65357=>"001111111",
  65358=>"111100111",
  65359=>"000011111",
  65360=>"000111011",
  65361=>"100100100",
  65362=>"000000111",
  65363=>"111111111",
  65364=>"010111111",
  65365=>"010110111",
  65366=>"111011001",
  65367=>"101111000",
  65368=>"111011010",
  65369=>"111111011",
  65370=>"000111001",
  65371=>"101000000",
  65372=>"111110110",
  65373=>"000001001",
  65374=>"000000000",
  65375=>"001001111",
  65376=>"000111001",
  65377=>"000000001",
  65378=>"110111111",
  65379=>"000001001",
  65380=>"001000000",
  65381=>"111001001",
  65382=>"001111111",
  65383=>"000111011",
  65384=>"000000000",
  65385=>"000010111",
  65386=>"011111111",
  65387=>"111001000",
  65388=>"101001001",
  65389=>"000000000",
  65390=>"000000000",
  65391=>"111111001",
  65392=>"111000100",
  65393=>"000111110",
  65394=>"000000101",
  65395=>"000000010",
  65396=>"000101111",
  65397=>"000000000",
  65398=>"000000000",
  65399=>"111111111",
  65400=>"000000000",
  65401=>"001101111",
  65402=>"110111111",
  65403=>"000000000",
  65404=>"100000000",
  65405=>"111011111",
  65406=>"000000000",
  65407=>"000000000",
  65408=>"111111001",
  65409=>"111000000",
  65410=>"000101101",
  65411=>"000000000",
  65412=>"010000000",
  65413=>"000110110",
  65414=>"000000000",
  65415=>"000011011",
  65416=>"000000000",
  65417=>"111111111",
  65418=>"100000000",
  65419=>"111111111",
  65420=>"111001000",
  65421=>"101001111",
  65422=>"000000110",
  65423=>"000000111",
  65424=>"100100111",
  65425=>"000000000",
  65426=>"100000010",
  65427=>"111101111",
  65428=>"111111110",
  65429=>"010011000",
  65430=>"100000000",
  65431=>"001000111",
  65432=>"000000011",
  65433=>"000000000",
  65434=>"111110111",
  65435=>"111111111",
  65436=>"111101001",
  65437=>"001000000",
  65438=>"000001101",
  65439=>"000000000",
  65440=>"100111111",
  65441=>"010110000",
  65442=>"100000110",
  65443=>"111011000",
  65444=>"000011111",
  65445=>"111111100",
  65446=>"111111110",
  65447=>"000000000",
  65448=>"000000000",
  65449=>"111111001",
  65450=>"111000000",
  65451=>"011001011",
  65452=>"000001111",
  65453=>"111011111",
  65454=>"111000001",
  65455=>"111001001",
  65456=>"111101000",
  65457=>"111000000",
  65458=>"000000101",
  65459=>"111101111",
  65460=>"000000111",
  65461=>"011001111",
  65462=>"011111010",
  65463=>"001000000",
  65464=>"000110010",
  65465=>"111010110",
  65466=>"000001101",
  65467=>"000110111",
  65468=>"001000111",
  65469=>"111111111",
  65470=>"001000000",
  65471=>"111011000",
  65472=>"111111101",
  65473=>"001000000",
  65474=>"111000000",
  65475=>"000000011",
  65476=>"101111111",
  65477=>"111110000",
  65478=>"001010000",
  65479=>"111001000",
  65480=>"111100111",
  65481=>"110100110",
  65482=>"101101000",
  65483=>"111000000",
  65484=>"111111000",
  65485=>"111111000",
  65486=>"000000000",
  65487=>"111110000",
  65488=>"000000011",
  65489=>"101001000",
  65490=>"000000000",
  65491=>"000000000",
  65492=>"100100110",
  65493=>"101100100",
  65494=>"111111111",
  65495=>"011011011",
  65496=>"000000000",
  65497=>"000000111",
  65498=>"100100111",
  65499=>"111111110",
  65500=>"001111000",
  65501=>"111101100",
  65502=>"100100111",
  65503=>"000011011",
  65504=>"111001000",
  65505=>"110111111",
  65506=>"000000111",
  65507=>"101011111",
  65508=>"111111001",
  65509=>"111110000",
  65510=>"111000000",
  65511=>"101111111",
  65512=>"000000101",
  65513=>"111000000",
  65514=>"010010000",
  65515=>"000000001",
  65516=>"100101111",
  65517=>"111111000",
  65518=>"000000000",
  65519=>"010011111",
  65520=>"000000000",
  65521=>"000000000",
  65522=>"111001011",
  65523=>"111011111",
  65524=>"001000000",
  65525=>"110110000",
  65526=>"100110111",
  65527=>"000000000",
  65528=>"000001111",
  65529=>"110100000",
  65530=>"011011000",
  65531=>"111000000",
  65532=>"110000000",
  65533=>"101011111",
  65534=>"111000001",
  65535=>"110000000");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;