LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L5_2_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    address : IN unsigned(6 DOWNTO 0));
END L5_2_BNROM;

ARCHITECTURE RTL OF L5_2_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 127) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  --Contenido bias || scale
  (0=>"1111110011011010"&"0001100000101011",
  1=>"0000001111000111"&"0001011010011001",
  2=>"0000001001010011"&"0001001111100000",
  3=>"0000000010000111"&"0001101001000101",
  4=>"1111110110010011"&"0001010100011110",
  5=>"1111111100110011"&"0001010111001010",
  6=>"1111011101100111"&"0001101110011100",
  7=>"1111010010000111"&"0001100001011011",
  8=>"1111111110001010"&"0001100000101101",
  9=>"1111100110011001"&"0001011001111010",
  10=>"1111110101111100"&"0001001110100110",
  11=>"1111101010001110"&"0001101000111010",
  12=>"0000010110000010"&"0001001100000101",
  13=>"1111001111001111"&"0001101011100000",
  14=>"1111011110100111"&"0001010111100011",
  15=>"1101010011111000"&"0001110001110111",
  16=>"0000010011011111"&"0001101011011010",
  17=>"1111110110011011"&"0001010110111101",
  18=>"1111101100111101"&"0001011000010111",
  19=>"1111001000111010"&"0001100011001111",
  20=>"1111011001001011"&"0001101100100100",
  21=>"0000010111001111"&"0001001010101010",
  22=>"0000011111010010"&"0001000011101000",
  23=>"1111110101010011"&"0001100001001100",
  24=>"1111110111101010"&"0001010010001001",
  25=>"0000000001000001"&"0001110110010100",
  26=>"0000011011001101"&"0000111011010111",
  27=>"1111101000000011"&"0001011100110101",
  28=>"1111111011101101"&"0001011001101010",
  29=>"1111010000110000"&"0001011001011100",
  30=>"1111110101001001"&"0001011010110000",
  31=>"1110011011100111"&"0001010101111101",
  32=>"1111101101011001"&"0001111010010000",
  33=>"0000001001101000"&"0001010000111101",
  34=>"0000001000101000"&"0001001010100101",
  35=>"1111001110011001"&"0001111110010100",
  36=>"0000010100010110"&"0001011100101101",
  37=>"0000000101101000"&"0001010011010011",
  38=>"1111111001001101"&"0001110010111100",
  39=>"0000001100111101"&"0001010001100111",
  40=>"1111111100111100"&"0001011000100010",
  41=>"0000000100101000"&"0001101011010001",
  42=>"0000001000111101"&"0001010010100001",
  43=>"1110111000111101"&"0001010001000000",
  44=>"1111110110001101"&"0010001101110100",
  45=>"0000000110001100"&"0001100010101101",
  46=>"0000010011100111"&"0001010010101110",
  47=>"0000011110101010"&"0001001011110100",
  48=>"1111011111010001"&"0010001111001100",
  49=>"1111101111100010"&"0001101110011010",
  50=>"1111100100011100"&"0001010010100010",
  51=>"1111101011111101"&"0001100010111001",
  52=>"0000000101100110"&"0001011101011110",
  53=>"1111010111110101"&"0001011100110001",
  54=>"1111011100100110"&"0001101110111101",
  55=>"0000001011001101"&"0001101011101100",
  56=>"1111011101000000"&"0001101011011001",
  57=>"1111100001011001"&"0001101101111001",
  58=>"1111110000000100"&"0001100010000001",
  59=>"0000001100011110"&"0001100000000001",
  60=>"0000000001001000"&"0001100011110011",
  61=>"0000011101000000"&"0001011011100010",
  62=>"1111110110110001"&"0001110100000110",
  63=>"1111101001001011"&"0001010001100111",
  64=>"1111110000011110"&"0001000101000010",
  65=>"1111001001011110"&"0000111101101001",
  66=>"1111100000100010"&"0001101110000011",
  67=>"1111111001000110"&"0001111000100000",
  68=>"0000011000100111"&"0001010101101100",
  69=>"1111011111000111"&"0001111100001110",
  70=>"0000001111111011"&"0001001101110011",
  71=>"1111111110101101"&"0001011100111010",
  72=>"1111001011111101"&"0010000011100111",
  73=>"0000001010100011"&"0001100001101100",
  74=>"1111111101100110"&"0001101001110001",
  75=>"0000011111001100"&"0001001000000100",
  76=>"1111100110000011"&"0001001001010101",
  77=>"1111010011101000"&"0001101101110110",
  78=>"1111001110011101"&"0001010011111101",
  79=>"1111111000101101"&"0001011001100001",
  80=>"0000100111100100"&"0000111111001110",
  81=>"0000010111011110"&"0001011011110101",
  82=>"0000000001010001"&"0001011101001001",
  83=>"0000001110111110"&"0001010010110100",
  84=>"0000001010110000"&"0001000110010011",
  85=>"1111111100100110"&"0001100011101100",
  86=>"0000100110001110"&"0000111011001101",
  87=>"1111111001001111"&"0001100011010000",
  88=>"0000100011001000"&"0000110000101100",
  89=>"0000001010110000"&"0001001100111111",
  90=>"1111000110100001"&"0010011001110100",
  91=>"1111111111100111"&"0001001000010101",
  92=>"0000001111110000"&"0001010110111011",
  93=>"0000001111001000"&"0001101010110000",
  94=>"1111101111100001"&"0001011001111001",
  95=>"1111111110001000"&"0001010101100000",
  96=>"1111110011101111"&"0001001111000111",
  97=>"0000011111100011"&"0001010101011011",
  98=>"0000101101111101"&"0001001001110100",
  99=>"0000010111101010"&"0001100101001101",
  100=>"1110111110100011"&"0001010000000100",
  101=>"0000011111000010"&"0001000111110110",
  102=>"1111111011110110"&"0001001000111110",
  103=>"0000000000111111"&"0001010010011011",
  104=>"1111101000001111"&"0001011000111100",
  105=>"1111110110110111"&"0001100110111101",
  106=>"1111110000100101"&"0001001110100100",
  107=>"0000000100001011"&"0001100110100100",
  108=>"0000100111100101"&"0001000101001100",
  109=>"0000000111111000"&"0001100101001011",
  110=>"0000001101000110"&"0001011110011111",
  111=>"1110111000011110"&"0001100110011110",
  112=>"0000001001010011"&"0001000010010010",
  113=>"1111100001011011"&"0001110100101001",
  114=>"0000001100011011"&"0001011011011101",
  115=>"1111111010011000"&"0001001101101110",
  116=>"1111110101001111"&"0001100011010001",
  117=>"0000101111110011"&"0001001000001000",
  118=>"1110100110111001"&"0001100110011111",
  119=>"1111010000110011"&"0001011001100110",
  120=>"0000010100110110"&"0000111100001110",
  121=>"1111111001010111"&"0001010110001110",
  122=>"0000000001001110"&"0000111100011010",
  123=>"0000010011010100"&"0001100011011101",
  124=>"1111111001000110"&"0001000000110111",
  125=>"1111110111010000"&"0001000011110000",
  126=>"1111110101111111"&"0001011110110101",
  127=>"1111100000011100"&"0001001110001101");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;