LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L6_2_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(6)-1 DOWNTO 0));
END L6_2_WROM;

ARCHITECTURE RTL OF L6_2_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"111001011",
  1=>"001101011",
  2=>"000000100",
  3=>"000010111",
  4=>"100000001",
  5=>"111010000",
  6=>"000101011",
  7=>"010000111",
  8=>"000000111",
  9=>"111000000",
  10=>"010000000",
  11=>"000010101",
  12=>"111111111",
  13=>"011000101",
  14=>"100001001",
  15=>"101000000",
  16=>"000000100",
  17=>"111110000",
  18=>"000010000",
  19=>"111000111",
  20=>"111011111",
  21=>"000100010",
  22=>"000010000",
  23=>"011001011",
  24=>"111000000",
  25=>"001101000",
  26=>"000000000",
  27=>"000011000",
  28=>"011000100",
  29=>"100100111",
  30=>"111001100",
  31=>"000101111",
  32=>"000010000",
  33=>"011111111",
  34=>"000010110",
  35=>"010000000",
  36=>"110011111",
  37=>"110110111",
  38=>"000011111",
  39=>"000111111",
  40=>"111111111",
  41=>"111111111",
  42=>"000000000",
  43=>"000110110",
  44=>"011111111",
  45=>"111110011",
  46=>"111101000",
  47=>"000001111",
  48=>"000000000",
  49=>"110000000",
  50=>"000000100",
  51=>"101000000",
  52=>"100000000",
  53=>"111111101",
  54=>"000000000",
  55=>"000000001",
  56=>"111101001",
  57=>"001110110",
  58=>"000010110",
  59=>"111111001",
  60=>"100000111",
  61=>"010111011",
  62=>"000000000",
  63=>"011010110",
  64=>"000000000",
  65=>"111110000",
  66=>"111111111",
  67=>"011001011",
  68=>"100111111",
  69=>"111110010",
  70=>"000000000",
  71=>"010000001",
  72=>"111011110",
  73=>"010000100",
  74=>"010010000",
  75=>"100000000",
  76=>"000000011",
  77=>"110110100",
  78=>"011001100",
  79=>"111111110",
  80=>"000110111",
  81=>"010011000",
  82=>"011101111",
  83=>"011101011",
  84=>"000000010",
  85=>"100110111",
  86=>"001001101",
  87=>"000000000",
  88=>"111111010",
  89=>"111111111",
  90=>"100100111",
  91=>"001100111",
  92=>"000100100",
  93=>"011001001",
  94=>"011111000",
  95=>"100100100",
  96=>"000010111",
  97=>"000010111",
  98=>"111000111",
  99=>"000000010",
  100=>"111111000",
  101=>"000010011",
  102=>"000000111",
  103=>"101100000",
  104=>"011100000",
  105=>"010000110",
  106=>"000000000",
  107=>"111111100",
  108=>"010110101",
  109=>"100011000",
  110=>"000001010",
  111=>"111111001",
  112=>"100100111",
  113=>"000000111",
  114=>"000000000",
  115=>"011111011",
  116=>"111000000",
  117=>"101000000",
  118=>"000010111",
  119=>"011011111",
  120=>"000001111",
  121=>"111100010",
  122=>"001001111",
  123=>"110101100",
  124=>"000000000",
  125=>"110100100",
  126=>"000011110",
  127=>"000000100",
  128=>"111111110",
  129=>"111000100",
  130=>"000010111",
  131=>"101101010",
  132=>"000000010",
  133=>"101101011",
  134=>"011011011",
  135=>"001001100",
  136=>"100001101",
  137=>"001101101",
  138=>"000011000",
  139=>"011011000",
  140=>"000010101",
  141=>"110111100",
  142=>"110011000",
  143=>"000000000",
  144=>"100000100",
  145=>"001000101",
  146=>"101101111",
  147=>"101100000",
  148=>"000001001",
  149=>"000010001",
  150=>"010001000",
  151=>"011011111",
  152=>"010010000",
  153=>"000010011",
  154=>"101000110",
  155=>"000000000",
  156=>"000000000",
  157=>"110110000",
  158=>"001001001",
  159=>"000001000",
  160=>"011000100",
  161=>"101000000",
  162=>"111111111",
  163=>"011001100",
  164=>"010000000",
  165=>"100100110",
  166=>"010110001",
  167=>"010101000",
  168=>"000111000",
  169=>"000000111",
  170=>"010010001",
  171=>"111010000",
  172=>"100110001",
  173=>"111111111",
  174=>"100001000",
  175=>"011111111",
  176=>"011001010",
  177=>"101001011",
  178=>"110010000",
  179=>"010010000",
  180=>"001101110",
  181=>"111110100",
  182=>"000111111",
  183=>"010111000",
  184=>"011100111",
  185=>"100101001",
  186=>"111011000",
  187=>"111000000",
  188=>"111111111",
  189=>"000111011",
  190=>"011011011",
  191=>"000000011",
  192=>"000000000",
  193=>"010111000",
  194=>"000000111",
  195=>"100100111",
  196=>"000011010",
  197=>"011010001",
  198=>"000000100",
  199=>"010111011",
  200=>"000000111",
  201=>"000010010",
  202=>"111111110",
  203=>"001000001",
  204=>"100000101",
  205=>"000000010",
  206=>"001010111",
  207=>"010011000",
  208=>"000011111",
  209=>"110110111",
  210=>"100001010",
  211=>"111101111",
  212=>"000000001",
  213=>"000000100",
  214=>"111111001",
  215=>"000111010",
  216=>"001101111",
  217=>"001000011",
  218=>"111111111",
  219=>"000101010",
  220=>"000000101",
  221=>"010011011",
  222=>"100111111",
  223=>"111101101",
  224=>"100010111",
  225=>"000001001",
  226=>"111111111",
  227=>"100000000",
  228=>"111111111",
  229=>"000000101",
  230=>"010000110",
  231=>"001000000",
  232=>"000010111",
  233=>"100100000",
  234=>"110100000",
  235=>"000000010",
  236=>"011111111",
  237=>"000000110",
  238=>"010000000",
  239=>"000000001",
  240=>"000000111",
  241=>"000001000",
  242=>"111111101",
  243=>"111111111",
  244=>"110100010",
  245=>"000000000",
  246=>"101000000",
  247=>"000000000",
  248=>"000000000",
  249=>"111111010",
  250=>"000000000",
  251=>"000000111",
  252=>"111111100",
  253=>"000000100",
  254=>"000000100",
  255=>"010101000",
  256=>"000000000",
  257=>"110001011",
  258=>"001001001",
  259=>"100111111",
  260=>"101100101",
  261=>"101101111",
  262=>"110010010",
  263=>"100110100",
  264=>"101000111",
  265=>"011011011",
  266=>"111111111",
  267=>"011001011",
  268=>"011011001",
  269=>"000000001",
  270=>"010011100",
  271=>"001000000",
  272=>"001001001",
  273=>"110000111",
  274=>"101100100",
  275=>"000011010",
  276=>"000100100",
  277=>"011011011",
  278=>"011011011",
  279=>"000101101",
  280=>"000000100",
  281=>"100101110",
  282=>"001100000",
  283=>"011011011",
  284=>"010100011",
  285=>"011010000",
  286=>"011011001",
  287=>"001000100",
  288=>"010011000",
  289=>"100100101",
  290=>"010001000",
  291=>"000010011",
  292=>"100100101",
  293=>"100100000",
  294=>"111100100",
  295=>"110100111",
  296=>"100100110",
  297=>"100100110",
  298=>"101001101",
  299=>"011010001",
  300=>"111111100",
  301=>"011001101",
  302=>"010100110",
  303=>"111110110",
  304=>"111001011",
  305=>"101100100",
  306=>"001001011",
  307=>"011101111",
  308=>"111100000",
  309=>"101100101",
  310=>"111010001",
  311=>"000000000",
  312=>"110000100",
  313=>"111000110",
  314=>"000011111",
  315=>"011000111",
  316=>"000010100",
  317=>"100100100",
  318=>"010011011",
  319=>"100101101",
  320=>"111111111",
  321=>"110100100",
  322=>"101100010",
  323=>"011011011",
  324=>"100100000",
  325=>"011000000",
  326=>"001001000",
  327=>"110111110",
  328=>"000011001",
  329=>"101101101",
  330=>"110011000",
  331=>"100100101",
  332=>"111101111",
  333=>"100100100",
  334=>"100100100",
  335=>"101100011",
  336=>"100100100",
  337=>"100000111",
  338=>"100000101",
  339=>"011001000",
  340=>"100110111",
  341=>"111101111",
  342=>"110100101",
  343=>"011011011",
  344=>"100100100",
  345=>"100100000",
  346=>"100100100",
  347=>"000100000",
  348=>"011111111",
  349=>"000000011",
  350=>"011011011",
  351=>"111011000",
  352=>"011011011",
  353=>"101011011",
  354=>"010011111",
  355=>"100110000",
  356=>"000011000",
  357=>"101100001",
  358=>"111111000",
  359=>"000000010",
  360=>"010111111",
  361=>"000001100",
  362=>"110111111",
  363=>"100001011",
  364=>"100101111",
  365=>"000101101",
  366=>"011000001",
  367=>"010100011",
  368=>"111111111",
  369=>"011001010",
  370=>"011101011",
  371=>"110110011",
  372=>"000001111",
  373=>"000000010",
  374=>"111111001",
  375=>"111111010",
  376=>"011010011",
  377=>"100100100",
  378=>"111110110",
  379=>"001011000",
  380=>"100000111",
  381=>"000000110",
  382=>"000011001",
  383=>"111111101",
  384=>"101000000",
  385=>"000000011",
  386=>"011011011",
  387=>"000110110",
  388=>"101111101",
  389=>"111111001",
  390=>"100101110",
  391=>"100100100",
  392=>"100100000",
  393=>"011000100",
  394=>"001011011",
  395=>"011000110",
  396=>"011011001",
  397=>"111111000",
  398=>"111111010",
  399=>"000000111",
  400=>"110110100",
  401=>"101001011",
  402=>"000001111",
  403=>"101111100",
  404=>"100101101",
  405=>"011011011",
  406=>"101100100",
  407=>"001001000",
  408=>"110100110",
  409=>"001111011",
  410=>"001011011",
  411=>"010011010",
  412=>"100010000",
  413=>"010110110",
  414=>"100001100",
  415=>"110110111",
  416=>"000011000",
  417=>"111011011",
  418=>"000000001",
  419=>"000111100",
  420=>"101011110",
  421=>"111110111",
  422=>"100010000",
  423=>"100100000",
  424=>"011000011",
  425=>"011011011",
  426=>"011011011",
  427=>"010000110",
  428=>"000000101",
  429=>"100110110",
  430=>"111101111",
  431=>"000111100",
  432=>"111011001",
  433=>"000110110",
  434=>"101000000",
  435=>"111111111",
  436=>"000000001",
  437=>"001000001",
  438=>"000000000",
  439=>"100100000",
  440=>"011011011",
  441=>"001010111",
  442=>"001001100",
  443=>"101101100",
  444=>"010000000",
  445=>"101100110",
  446=>"001001001",
  447=>"011011011",
  448=>"111111110",
  449=>"110110101",
  450=>"000001111",
  451=>"000100100",
  452=>"011011011",
  453=>"110100000",
  454=>"111101001",
  455=>"000011000",
  456=>"100000101",
  457=>"000111110",
  458=>"101101000",
  459=>"011111100",
  460=>"011010010",
  461=>"111111010",
  462=>"100100100",
  463=>"000011011",
  464=>"100100111",
  465=>"100100100",
  466=>"111001101",
  467=>"100100000",
  468=>"110100100",
  469=>"110101000",
  470=>"101111111",
  471=>"000000111",
  472=>"011011001",
  473=>"100010000",
  474=>"111011101",
  475=>"100100101",
  476=>"101100111",
  477=>"001010010",
  478=>"100000100",
  479=>"011011111",
  480=>"011011001",
  481=>"100100100",
  482=>"011011011",
  483=>"100110101",
  484=>"010011011",
  485=>"011011011",
  486=>"001000101",
  487=>"100110111",
  488=>"000000000",
  489=>"010111001",
  490=>"111101111",
  491=>"001110011",
  492=>"011011011",
  493=>"000101111",
  494=>"000000000",
  495=>"001011011",
  496=>"011001001",
  497=>"000110110",
  498=>"011010010",
  499=>"110111111",
  500=>"101001101",
  501=>"000110101",
  502=>"000010000",
  503=>"000011011",
  504=>"011011011",
  505=>"000000000",
  506=>"110010110",
  507=>"000010100",
  508=>"100100100",
  509=>"001000000",
  510=>"110100100",
  511=>"111111111",
  512=>"011101111",
  513=>"111100100",
  514=>"010010111",
  515=>"101111111",
  516=>"000000111",
  517=>"001111111",
  518=>"101111000",
  519=>"111111000",
  520=>"001000100",
  521=>"000111000",
  522=>"100001001",
  523=>"000011000",
  524=>"000110001",
  525=>"000000000",
  526=>"000110111",
  527=>"000100101",
  528=>"100101100",
  529=>"111111100",
  530=>"110100110",
  531=>"111000000",
  532=>"010000000",
  533=>"101000000",
  534=>"001100000",
  535=>"111010010",
  536=>"101101101",
  537=>"000110101",
  538=>"000000010",
  539=>"010111010",
  540=>"010111000",
  541=>"000000001",
  542=>"000010010",
  543=>"001000000",
  544=>"010111110",
  545=>"101111000",
  546=>"111111110",
  547=>"000000000",
  548=>"000000000",
  549=>"110110100",
  550=>"000000000",
  551=>"000101110",
  552=>"011101111",
  553=>"101000000",
  554=>"000000000",
  555=>"010101111",
  556=>"000011011",
  557=>"000001011",
  558=>"111010111",
  559=>"000000000",
  560=>"000100110",
  561=>"001001000",
  562=>"010000100",
  563=>"101011011",
  564=>"111111110",
  565=>"011110000",
  566=>"011000000",
  567=>"111100100",
  568=>"111111000",
  569=>"111101001",
  570=>"111010000",
  571=>"111111110",
  572=>"100110100",
  573=>"000111111",
  574=>"000010011",
  575=>"110010100",
  576=>"110110000",
  577=>"111010000",
  578=>"000000101",
  579=>"111001001",
  580=>"000000000",
  581=>"101000101",
  582=>"000000110",
  583=>"001100010",
  584=>"001000000",
  585=>"010111010",
  586=>"100000000",
  587=>"111010100",
  588=>"111100000",
  589=>"000000110",
  590=>"010011011",
  591=>"000011010",
  592=>"111000101",
  593=>"111111000",
  594=>"000111011",
  595=>"010111110",
  596=>"010010000",
  597=>"001000000",
  598=>"000110011",
  599=>"010111111",
  600=>"111111111",
  601=>"110111000",
  602=>"111111011",
  603=>"100110000",
  604=>"111111010",
  605=>"010011110",
  606=>"111101111",
  607=>"010100110",
  608=>"101100111",
  609=>"100101101",
  610=>"010111111",
  611=>"111111111",
  612=>"000111011",
  613=>"101111100",
  614=>"110111010",
  615=>"001000101",
  616=>"101111011",
  617=>"111111000",
  618=>"111111101",
  619=>"000010111",
  620=>"000000000",
  621=>"000000000",
  622=>"100111111",
  623=>"111111000",
  624=>"110110100",
  625=>"100111111",
  626=>"011000000",
  627=>"010010110",
  628=>"111111011",
  629=>"001000100",
  630=>"000111111",
  631=>"000100101",
  632=>"111111010",
  633=>"010000000",
  634=>"001000100",
  635=>"010101111",
  636=>"000100110",
  637=>"000010011",
  638=>"000000111",
  639=>"110111110",
  640=>"000111111",
  641=>"010110010",
  642=>"010111111",
  643=>"111111000",
  644=>"000100001",
  645=>"011011000",
  646=>"011011001",
  647=>"000100010",
  648=>"001111111",
  649=>"110000010",
  650=>"010011011",
  651=>"001101010",
  652=>"000000101",
  653=>"110111111",
  654=>"111101111",
  655=>"000000110",
  656=>"010000000",
  657=>"111101000",
  658=>"000101100",
  659=>"111000111",
  660=>"011011111",
  661=>"101111000",
  662=>"110111000",
  663=>"111110100",
  664=>"111111101",
  665=>"111000000",
  666=>"000110000",
  667=>"011111111",
  668=>"001000000",
  669=>"010111101",
  670=>"000101000",
  671=>"000110111",
  672=>"000110011",
  673=>"111111111",
  674=>"010000010",
  675=>"100000000",
  676=>"000000111",
  677=>"110011010",
  678=>"011001010",
  679=>"000110000",
  680=>"001101111",
  681=>"011101101",
  682=>"010000000",
  683=>"000111011",
  684=>"101111111",
  685=>"111111111",
  686=>"010110000",
  687=>"101001101",
  688=>"111011001",
  689=>"001101101",
  690=>"000111000",
  691=>"111111000",
  692=>"000111011",
  693=>"111111010",
  694=>"101111101",
  695=>"011111111",
  696=>"001001001",
  697=>"000100110",
  698=>"111000010",
  699=>"000111111",
  700=>"000010111",
  701=>"010111111",
  702=>"011100101",
  703=>"111100000",
  704=>"111101010",
  705=>"111000000",
  706=>"000100110",
  707=>"000011011",
  708=>"000011000",
  709=>"111011111",
  710=>"001111110",
  711=>"110111000",
  712=>"000101001",
  713=>"110100100",
  714=>"001101110",
  715=>"111100110",
  716=>"000000000",
  717=>"000000011",
  718=>"110010010",
  719=>"110101001",
  720=>"111111010",
  721=>"110011011",
  722=>"111011011",
  723=>"000000010",
  724=>"000011111",
  725=>"110001111",
  726=>"000010010",
  727=>"011001000",
  728=>"111111111",
  729=>"000001011",
  730=>"101011101",
  731=>"110010000",
  732=>"100110111",
  733=>"111101100",
  734=>"111100000",
  735=>"000000000",
  736=>"100111111",
  737=>"000111111",
  738=>"111000000",
  739=>"011111111",
  740=>"010010010",
  741=>"000000111",
  742=>"010111000",
  743=>"110010101",
  744=>"101101111",
  745=>"000100010",
  746=>"001001011",
  747=>"101111111",
  748=>"001001000",
  749=>"101000000",
  750=>"010110010",
  751=>"100011011",
  752=>"111000111",
  753=>"111100111",
  754=>"000111111",
  755=>"010010000",
  756=>"000000111",
  757=>"101000101",
  758=>"000001000",
  759=>"010000000",
  760=>"000000000",
  761=>"101001010",
  762=>"101100111",
  763=>"000111111",
  764=>"111001000",
  765=>"011000101",
  766=>"001110100",
  767=>"000010000",
  768=>"000011111",
  769=>"000000000",
  770=>"000000100",
  771=>"110111010",
  772=>"000000000",
  773=>"000010000",
  774=>"110000001",
  775=>"111110011",
  776=>"000111111",
  777=>"000000000",
  778=>"011001000",
  779=>"000000000",
  780=>"000000000",
  781=>"000111111",
  782=>"000011011",
  783=>"000000000",
  784=>"101111001",
  785=>"110000011",
  786=>"111000000",
  787=>"111111000",
  788=>"101010000",
  789=>"010011010",
  790=>"000000010",
  791=>"111111011",
  792=>"010010000",
  793=>"000110011",
  794=>"000111000",
  795=>"101111111",
  796=>"000001000",
  797=>"111000000",
  798=>"111011111",
  799=>"111000000",
  800=>"000111111",
  801=>"010010000",
  802=>"111001000",
  803=>"000011111",
  804=>"111101110",
  805=>"001110110",
  806=>"000111110",
  807=>"000110110",
  808=>"000010111",
  809=>"000111111",
  810=>"000000000",
  811=>"000010000",
  812=>"011001000",
  813=>"111000111",
  814=>"111111100",
  815=>"000001101",
  816=>"000000111",
  817=>"000011001",
  818=>"000111100",
  819=>"000000001",
  820=>"001000000",
  821=>"010000101",
  822=>"100100001",
  823=>"001101000",
  824=>"001000010",
  825=>"111000001",
  826=>"110101111",
  827=>"111101011",
  828=>"011000001",
  829=>"010111000",
  830=>"001000000",
  831=>"010111111",
  832=>"000110101",
  833=>"101101101",
  834=>"110111111",
  835=>"000110110",
  836=>"110000000",
  837=>"011001000",
  838=>"011100110",
  839=>"111001000",
  840=>"111100100",
  841=>"111111111",
  842=>"010100101",
  843=>"111101100",
  844=>"010000100",
  845=>"001001101",
  846=>"000100100",
  847=>"111101001",
  848=>"101101101",
  849=>"010011000",
  850=>"111111111",
  851=>"111001000",
  852=>"101000101",
  853=>"010100111",
  854=>"111011001",
  855=>"000111111",
  856=>"001111111",
  857=>"011101001",
  858=>"111100100",
  859=>"111111100",
  860=>"101010010",
  861=>"110001001",
  862=>"111000001",
  863=>"000011111",
  864=>"000010110",
  865=>"110000110",
  866=>"000000001",
  867=>"111100110",
  868=>"010111100",
  869=>"110111101",
  870=>"111111110",
  871=>"000001010",
  872=>"101100110",
  873=>"010111111",
  874=>"111111000",
  875=>"111111101",
  876=>"111111111",
  877=>"111100110",
  878=>"001101000",
  879=>"000000000",
  880=>"000110111",
  881=>"010011010",
  882=>"000001100",
  883=>"111000000",
  884=>"111001000",
  885=>"111001111",
  886=>"000001110",
  887=>"000111111",
  888=>"000001010",
  889=>"000111101",
  890=>"101000100",
  891=>"111101001",
  892=>"001010110",
  893=>"111101000",
  894=>"110110000",
  895=>"000000101",
  896=>"101000111",
  897=>"010100100",
  898=>"111111110",
  899=>"111101111",
  900=>"000100110",
  901=>"111111111",
  902=>"100111011",
  903=>"000010011",
  904=>"000001011",
  905=>"101101000",
  906=>"010000010",
  907=>"101101000",
  908=>"000000000",
  909=>"010110110",
  910=>"010000000",
  911=>"001101000",
  912=>"011001011",
  913=>"000100101",
  914=>"001101000",
  915=>"100011101",
  916=>"000110010",
  917=>"000011111",
  918=>"000000101",
  919=>"010110111",
  920=>"000000000",
  921=>"010000111",
  922=>"100000111",
  923=>"111100000",
  924=>"111010010",
  925=>"110011011",
  926=>"100000000",
  927=>"111101101",
  928=>"111000100",
  929=>"010000110",
  930=>"000111111",
  931=>"000011111",
  932=>"111111101",
  933=>"011001111",
  934=>"111001010",
  935=>"000101000",
  936=>"000100000",
  937=>"000111111",
  938=>"101111111",
  939=>"000000000",
  940=>"111101001",
  941=>"000111111",
  942=>"011001000",
  943=>"111111111",
  944=>"100101000",
  945=>"111110001",
  946=>"111000001",
  947=>"010110110",
  948=>"110000100",
  949=>"101000000",
  950=>"000000111",
  951=>"000010111",
  952=>"110000010",
  953=>"000110101",
  954=>"000000010",
  955=>"000010111",
  956=>"110010111",
  957=>"010111111",
  958=>"001011111",
  959=>"000000101",
  960=>"111000111",
  961=>"111011000",
  962=>"000001111",
  963=>"000110111",
  964=>"101000011",
  965=>"011000001",
  966=>"011000011",
  967=>"001000000",
  968=>"111111000",
  969=>"111100000",
  970=>"000001011",
  971=>"110100001",
  972=>"000011111",
  973=>"100010011",
  974=>"101000000",
  975=>"000111000",
  976=>"000010110",
  977=>"001000010",
  978=>"000010000",
  979=>"111000010",
  980=>"000111111",
  981=>"111000011",
  982=>"000000001",
  983=>"000111010",
  984=>"111100000",
  985=>"001000100",
  986=>"110001101",
  987=>"111000010",
  988=>"100001001",
  989=>"000000111",
  990=>"110100111",
  991=>"011111000",
  992=>"111000100",
  993=>"000000001",
  994=>"000111111",
  995=>"110111111",
  996=>"000010111",
  997=>"000000111",
  998=>"001111111",
  999=>"111111101",
  1000=>"010111110",
  1001=>"010111111",
  1002=>"110100000",
  1003=>"101000000",
  1004=>"000000111",
  1005=>"000110111",
  1006=>"000010000",
  1007=>"101000010",
  1008=>"111000000",
  1009=>"100000100",
  1010=>"101111110",
  1011=>"010001000",
  1012=>"000100111",
  1013=>"111000000",
  1014=>"000000110",
  1015=>"111100001",
  1016=>"101000000",
  1017=>"111000010",
  1018=>"111111111",
  1019=>"000000000",
  1020=>"001000000",
  1021=>"111011011",
  1022=>"110101111",
  1023=>"111110000",
  1024=>"010001000",
  1025=>"000111111",
  1026=>"000000000",
  1027=>"000000111",
  1028=>"110110110",
  1029=>"110111110",
  1030=>"101111100",
  1031=>"000001111",
  1032=>"000000000",
  1033=>"101101011",
  1034=>"010011100",
  1035=>"101000101",
  1036=>"111111100",
  1037=>"100000011",
  1038=>"011100011",
  1039=>"110000000",
  1040=>"000000111",
  1041=>"110010000",
  1042=>"111000101",
  1043=>"111101000",
  1044=>"000000011",
  1045=>"111111100",
  1046=>"011110100",
  1047=>"000001010",
  1048=>"111000000",
  1049=>"111111111",
  1050=>"000001000",
  1051=>"000000001",
  1052=>"000000110",
  1053=>"001101010",
  1054=>"111100000",
  1055=>"100111001",
  1056=>"110111111",
  1057=>"111111011",
  1058=>"000010001",
  1059=>"010010000",
  1060=>"000001100",
  1061=>"111111111",
  1062=>"111100000",
  1063=>"000110000",
  1064=>"100011111",
  1065=>"101101010",
  1066=>"000000011",
  1067=>"010101111",
  1068=>"001001011",
  1069=>"111110110",
  1070=>"101111111",
  1071=>"000000111",
  1072=>"110001101",
  1073=>"110110110",
  1074=>"000010001",
  1075=>"010010000",
  1076=>"000001100",
  1077=>"010000000",
  1078=>"110110100",
  1079=>"000000110",
  1080=>"010101001",
  1081=>"000000000",
  1082=>"011100000",
  1083=>"011010011",
  1084=>"011011110",
  1085=>"111111010",
  1086=>"000000000",
  1087=>"110110110",
  1088=>"010101111",
  1089=>"101111100",
  1090=>"110111010",
  1091=>"011001111",
  1092=>"000110110",
  1093=>"000110110",
  1094=>"010000000",
  1095=>"011000000",
  1096=>"001000110",
  1097=>"111010111",
  1098=>"101100111",
  1099=>"111000000",
  1100=>"000011001",
  1101=>"110110010",
  1102=>"111111111",
  1103=>"100110110",
  1104=>"110010000",
  1105=>"111000010",
  1106=>"111000010",
  1107=>"000000000",
  1108=>"101001111",
  1109=>"011010110",
  1110=>"010011001",
  1111=>"111001111",
  1112=>"000000100",
  1113=>"100100001",
  1114=>"001101101",
  1115=>"100000000",
  1116=>"111100100",
  1117=>"000001000",
  1118=>"001100011",
  1119=>"100101001",
  1120=>"101010000",
  1121=>"000001111",
  1122=>"100010010",
  1123=>"000000100",
  1124=>"001001000",
  1125=>"110000000",
  1126=>"111011111",
  1127=>"010001000",
  1128=>"111010111",
  1129=>"000000000",
  1130=>"000010101",
  1131=>"001011111",
  1132=>"100001101",
  1133=>"010111111",
  1134=>"110010000",
  1135=>"000000110",
  1136=>"001000000",
  1137=>"000111111",
  1138=>"111011100",
  1139=>"111110011",
  1140=>"101110111",
  1141=>"000000000",
  1142=>"000111101",
  1143=>"000000000",
  1144=>"101101100",
  1145=>"000010000",
  1146=>"000110111",
  1147=>"111000001",
  1148=>"011100111",
  1149=>"100000000",
  1150=>"101001111",
  1151=>"001000101",
  1152=>"001001110",
  1153=>"010000111",
  1154=>"100000010",
  1155=>"010101111",
  1156=>"101101110",
  1157=>"000000000",
  1158=>"100011111",
  1159=>"110100111",
  1160=>"000101001",
  1161=>"100000010",
  1162=>"001101101",
  1163=>"111100101",
  1164=>"001001001",
  1165=>"111111001",
  1166=>"000000000",
  1167=>"001000000",
  1168=>"011001100",
  1169=>"100101001",
  1170=>"010001001",
  1171=>"101001100",
  1172=>"100010011",
  1173=>"000110100",
  1174=>"111010010",
  1175=>"000001111",
  1176=>"110110000",
  1177=>"101100101",
  1178=>"101101111",
  1179=>"000000000",
  1180=>"101000100",
  1181=>"111010111",
  1182=>"010000000",
  1183=>"111011111",
  1184=>"000111110",
  1185=>"000000110",
  1186=>"000011001",
  1187=>"101000111",
  1188=>"001000000",
  1189=>"001011010",
  1190=>"110110000",
  1191=>"000000000",
  1192=>"110011000",
  1193=>"000000000",
  1194=>"101101010",
  1195=>"110010000",
  1196=>"011111101",
  1197=>"110110000",
  1198=>"100001010",
  1199=>"110010000",
  1200=>"101000111",
  1201=>"010001000",
  1202=>"000001101",
  1203=>"001100000",
  1204=>"101101100",
  1205=>"001100111",
  1206=>"111111111",
  1207=>"010111111",
  1208=>"100011011",
  1209=>"110010110",
  1210=>"111000000",
  1211=>"001000111",
  1212=>"111110010",
  1213=>"100010111",
  1214=>"011000011",
  1215=>"110100000",
  1216=>"111001111",
  1217=>"101111111",
  1218=>"000111110",
  1219=>"001100110",
  1220=>"000010000",
  1221=>"100100011",
  1222=>"110100110",
  1223=>"111111111",
  1224=>"001110111",
  1225=>"000101000",
  1226=>"000111111",
  1227=>"010111111",
  1228=>"111101101",
  1229=>"110011011",
  1230=>"000010111",
  1231=>"111111111",
  1232=>"000001001",
  1233=>"000000110",
  1234=>"111001111",
  1235=>"000111111",
  1236=>"111011101",
  1237=>"000000011",
  1238=>"001000000",
  1239=>"100000001",
  1240=>"111101110",
  1241=>"001000100",
  1242=>"100000001",
  1243=>"000000000",
  1244=>"010011001",
  1245=>"000101101",
  1246=>"111111000",
  1247=>"110010001",
  1248=>"111110000",
  1249=>"000010000",
  1250=>"001000001",
  1251=>"111111000",
  1252=>"101000100",
  1253=>"111111001",
  1254=>"011001101",
  1255=>"001011010",
  1256=>"000110111",
  1257=>"110110100",
  1258=>"000000011",
  1259=>"001111110",
  1260=>"000000111",
  1261=>"111101100",
  1262=>"000000000",
  1263=>"110110000",
  1264=>"010100000",
  1265=>"011011010",
  1266=>"001000000",
  1267=>"001001001",
  1268=>"011010000",
  1269=>"000000101",
  1270=>"010010010",
  1271=>"000000001",
  1272=>"000000111",
  1273=>"101001000",
  1274=>"001101111",
  1275=>"001001000",
  1276=>"110110000",
  1277=>"011011101",
  1278=>"011010000",
  1279=>"000000000",
  1280=>"100100100",
  1281=>"101000110",
  1282=>"000000101",
  1283=>"101000000",
  1284=>"111101011",
  1285=>"101101000",
  1286=>"000000010",
  1287=>"110111111",
  1288=>"010000000",
  1289=>"000000000",
  1290=>"001110000",
  1291=>"000101100",
  1292=>"011000100",
  1293=>"111111000",
  1294=>"011000000",
  1295=>"111100100",
  1296=>"111000001",
  1297=>"100000000",
  1298=>"100101110",
  1299=>"110111011",
  1300=>"000101101",
  1301=>"000111111",
  1302=>"111011111",
  1303=>"000110111",
  1304=>"000000101",
  1305=>"010111101",
  1306=>"000000000",
  1307=>"000000000",
  1308=>"100000011",
  1309=>"100010000",
  1310=>"000001000",
  1311=>"001111010",
  1312=>"101000101",
  1313=>"111111111",
  1314=>"111101111",
  1315=>"111110111",
  1316=>"111000000",
  1317=>"000011100",
  1318=>"000010000",
  1319=>"111111000",
  1320=>"010111111",
  1321=>"000001000",
  1322=>"101101000",
  1323=>"011111010",
  1324=>"000100111",
  1325=>"111010100",
  1326=>"101110000",
  1327=>"101111110",
  1328=>"101011101",
  1329=>"111000000",
  1330=>"000111111",
  1331=>"000100000",
  1332=>"000010011",
  1333=>"111111111",
  1334=>"001011110",
  1335=>"111010000",
  1336=>"111100111",
  1337=>"000101000",
  1338=>"000100010",
  1339=>"011000111",
  1340=>"001011111",
  1341=>"010111010",
  1342=>"000000000",
  1343=>"001100000",
  1344=>"100000111",
  1345=>"000100000",
  1346=>"111110010",
  1347=>"110100000",
  1348=>"000000000",
  1349=>"000101001",
  1350=>"100101100",
  1351=>"101100010",
  1352=>"111111110",
  1353=>"101101111",
  1354=>"001010010",
  1355=>"000000000",
  1356=>"010000100",
  1357=>"100100100",
  1358=>"011000000",
  1359=>"001000001",
  1360=>"010010000",
  1361=>"111010111",
  1362=>"001000101",
  1363=>"000000000",
  1364=>"000000111",
  1365=>"011010110",
  1366=>"011000000",
  1367=>"101100000",
  1368=>"000000010",
  1369=>"110000000",
  1370=>"000011011",
  1371=>"100000010",
  1372=>"011000001",
  1373=>"001001111",
  1374=>"100101101",
  1375=>"011001001",
  1376=>"111000000",
  1377=>"111110010",
  1378=>"000000000",
  1379=>"000110110",
  1380=>"110000001",
  1381=>"100000000",
  1382=>"111100101",
  1383=>"100000100",
  1384=>"101111010",
  1385=>"111111111",
  1386=>"101101111",
  1387=>"111000000",
  1388=>"100010100",
  1389=>"100011000",
  1390=>"010000000",
  1391=>"000101111",
  1392=>"111000000",
  1393=>"100101101",
  1394=>"000111111",
  1395=>"111000000",
  1396=>"101001000",
  1397=>"000000000",
  1398=>"001001000",
  1399=>"010000000",
  1400=>"001000000",
  1401=>"000100000",
  1402=>"101100001",
  1403=>"000000001",
  1404=>"101100111",
  1405=>"001001001",
  1406=>"011111111",
  1407=>"000001010",
  1408=>"110101101",
  1409=>"000111011",
  1410=>"000000111",
  1411=>"101001100",
  1412=>"000000101",
  1413=>"101111010",
  1414=>"000110000",
  1415=>"011001000",
  1416=>"111000100",
  1417=>"000110010",
  1418=>"000000000",
  1419=>"010000000",
  1420=>"101000100",
  1421=>"101101000",
  1422=>"111010100",
  1423=>"010000000",
  1424=>"110101001",
  1425=>"000001000",
  1426=>"000000000",
  1427=>"000100111",
  1428=>"101100000",
  1429=>"101000101",
  1430=>"111111011",
  1431=>"000101100",
  1432=>"100000000",
  1433=>"000110010",
  1434=>"000011111",
  1435=>"111000001",
  1436=>"011000000",
  1437=>"101111111",
  1438=>"101111111",
  1439=>"010101101",
  1440=>"111111111",
  1441=>"000010011",
  1442=>"011111011",
  1443=>"111111011",
  1444=>"001101000",
  1445=>"011000000",
  1446=>"111101000",
  1447=>"111111111",
  1448=>"110110000",
  1449=>"010011000",
  1450=>"110111111",
  1451=>"101100010",
  1452=>"011000000",
  1453=>"110100100",
  1454=>"001111110",
  1455=>"011101101",
  1456=>"100000101",
  1457=>"111011011",
  1458=>"001111111",
  1459=>"100100111",
  1460=>"101001011",
  1461=>"100100111",
  1462=>"001001111",
  1463=>"111001000",
  1464=>"010111110",
  1465=>"111010000",
  1466=>"010111111",
  1467=>"011010000",
  1468=>"101011011",
  1469=>"111111111",
  1470=>"000100100",
  1471=>"011011000",
  1472=>"000000101",
  1473=>"101100001",
  1474=>"111111000",
  1475=>"110000001",
  1476=>"000000000",
  1477=>"001101000",
  1478=>"110100000",
  1479=>"101010010",
  1480=>"111010111",
  1481=>"111001000",
  1482=>"111010011",
  1483=>"101101000",
  1484=>"111100000",
  1485=>"011011110",
  1486=>"000000000",
  1487=>"001000000",
  1488=>"000001001",
  1489=>"111011000",
  1490=>"011001010",
  1491=>"111101000",
  1492=>"111101111",
  1493=>"110111111",
  1494=>"010011000",
  1495=>"001001000",
  1496=>"000000000",
  1497=>"101111111",
  1498=>"011001100",
  1499=>"001101001",
  1500=>"110101110",
  1501=>"111111000",
  1502=>"001000110",
  1503=>"000000000",
  1504=>"111000000",
  1505=>"000001010",
  1506=>"000101111",
  1507=>"010001000",
  1508=>"000000001",
  1509=>"001101101",
  1510=>"000000000",
  1511=>"000101011",
  1512=>"111000111",
  1513=>"101111111",
  1514=>"000010000",
  1515=>"001000000",
  1516=>"111111001",
  1517=>"111111010",
  1518=>"010000010",
  1519=>"001101100",
  1520=>"100000000",
  1521=>"100100000",
  1522=>"101101100",
  1523=>"011100110",
  1524=>"001001001",
  1525=>"001111010",
  1526=>"010010000",
  1527=>"111101011",
  1528=>"000000111",
  1529=>"000111111",
  1530=>"100101011",
  1531=>"101010000",
  1532=>"111111111",
  1533=>"011111101",
  1534=>"000001111",
  1535=>"100000000",
  1536=>"001000001",
  1537=>"100000100",
  1538=>"101101111",
  1539=>"110010110",
  1540=>"110100100",
  1541=>"100001000",
  1542=>"111011010",
  1543=>"111111010",
  1544=>"000000000",
  1545=>"010010000",
  1546=>"001001011",
  1547=>"101101101",
  1548=>"110000001",
  1549=>"110011000",
  1550=>"100100010",
  1551=>"010110011",
  1552=>"011000000",
  1553=>"010010000",
  1554=>"010100101",
  1555=>"111011000",
  1556=>"010111001",
  1557=>"100100101",
  1558=>"101101101",
  1559=>"101101110",
  1560=>"010010010",
  1561=>"110100001",
  1562=>"110110111",
  1563=>"101100000",
  1564=>"011011000",
  1565=>"001001001",
  1566=>"110010000",
  1567=>"111011010",
  1568=>"001101111",
  1569=>"010000111",
  1570=>"110111111",
  1571=>"000000000",
  1572=>"011011111",
  1573=>"100100000",
  1574=>"000000000",
  1575=>"111111111",
  1576=>"010111011",
  1577=>"100111110",
  1578=>"100000000",
  1579=>"111111111",
  1580=>"100010010",
  1581=>"100101001",
  1582=>"000000011",
  1583=>"100000010",
  1584=>"000010010",
  1585=>"101101101",
  1586=>"111000000",
  1587=>"111100100",
  1588=>"000000100",
  1589=>"111101000",
  1590=>"000100100",
  1591=>"111011110",
  1592=>"101101101",
  1593=>"111100110",
  1594=>"000000101",
  1595=>"111111010",
  1596=>"110110100",
  1597=>"111111111",
  1598=>"000100101",
  1599=>"101101100",
  1600=>"000010010",
  1601=>"010100010",
  1602=>"101111111",
  1603=>"111001001",
  1604=>"010010000",
  1605=>"010000000",
  1606=>"100000000",
  1607=>"011110110",
  1608=>"001100110",
  1609=>"111010010",
  1610=>"000001001",
  1611=>"111000000",
  1612=>"110000000",
  1613=>"011110110",
  1614=>"111111000",
  1615=>"101111011",
  1616=>"100100000",
  1617=>"111111111",
  1618=>"011001100",
  1619=>"000001111",
  1620=>"110100110",
  1621=>"111101111",
  1622=>"000100100",
  1623=>"100100101",
  1624=>"101000000",
  1625=>"011100001",
  1626=>"010000010",
  1627=>"000000101",
  1628=>"010111010",
  1629=>"010001101",
  1630=>"100000000",
  1631=>"100000100",
  1632=>"000110000",
  1633=>"001001000",
  1634=>"111101101",
  1635=>"000110110",
  1636=>"001000100",
  1637=>"000000000",
  1638=>"111101111",
  1639=>"110101111",
  1640=>"111110110",
  1641=>"000010110",
  1642=>"000000000",
  1643=>"111001001",
  1644=>"000000011",
  1645=>"111111110",
  1646=>"000000111",
  1647=>"000000001",
  1648=>"001100000",
  1649=>"100101101",
  1650=>"000001001",
  1651=>"101011001",
  1652=>"010011010",
  1653=>"000000000",
  1654=>"000010000",
  1655=>"101011000",
  1656=>"000000101",
  1657=>"111111000",
  1658=>"100101111",
  1659=>"000001111",
  1660=>"100000111",
  1661=>"001010100",
  1662=>"101100110",
  1663=>"001101001",
  1664=>"101000010",
  1665=>"111011010",
  1666=>"010111000",
  1667=>"001111011",
  1668=>"001000110",
  1669=>"110100000",
  1670=>"001001001",
  1671=>"100101011",
  1672=>"100110100",
  1673=>"000000000",
  1674=>"000110000",
  1675=>"000000001",
  1676=>"110110101",
  1677=>"111111000",
  1678=>"111111111",
  1679=>"001000000",
  1680=>"000100111",
  1681=>"111100100",
  1682=>"010000011",
  1683=>"110010110",
  1684=>"001011010",
  1685=>"101100111",
  1686=>"000010000",
  1687=>"110000111",
  1688=>"010010110",
  1689=>"110111111",
  1690=>"000000000",
  1691=>"011111111",
  1692=>"000000010",
  1693=>"111001111",
  1694=>"010011000",
  1695=>"000000000",
  1696=>"000000011",
  1697=>"010100011",
  1698=>"000101011",
  1699=>"010110010",
  1700=>"001111011",
  1701=>"000000100",
  1702=>"010110001",
  1703=>"100000000",
  1704=>"110010000",
  1705=>"110111100",
  1706=>"000000000",
  1707=>"000011010",
  1708=>"111101101",
  1709=>"000101111",
  1710=>"111110110",
  1711=>"000110000",
  1712=>"101000101",
  1713=>"001000110",
  1714=>"111101111",
  1715=>"000001000",
  1716=>"011111110",
  1717=>"000010011",
  1718=>"010011010",
  1719=>"101100001",
  1720=>"111001001",
  1721=>"000000110",
  1722=>"000010010",
  1723=>"000010110",
  1724=>"101001011",
  1725=>"111111111",
  1726=>"000000000",
  1727=>"001000100",
  1728=>"101000100",
  1729=>"000000010",
  1730=>"000000000",
  1731=>"101100000",
  1732=>"100010011",
  1733=>"100100011",
  1734=>"000000011",
  1735=>"000000000",
  1736=>"100111100",
  1737=>"001000000",
  1738=>"000100010",
  1739=>"000000000",
  1740=>"010100000",
  1741=>"111010110",
  1742=>"000100110",
  1743=>"110110100",
  1744=>"111001010",
  1745=>"101000011",
  1746=>"111100000",
  1747=>"000011111",
  1748=>"111000001",
  1749=>"101101111",
  1750=>"101111111",
  1751=>"010000010",
  1752=>"101000101",
  1753=>"000001100",
  1754=>"000111110",
  1755=>"111100000",
  1756=>"111111101",
  1757=>"000111111",
  1758=>"111000111",
  1759=>"000000000",
  1760=>"111101101",
  1761=>"101000000",
  1762=>"111011000",
  1763=>"011011111",
  1764=>"000000000",
  1765=>"111100000",
  1766=>"000000000",
  1767=>"010010110",
  1768=>"001111010",
  1769=>"000010000",
  1770=>"111100111",
  1771=>"000000111",
  1772=>"000000000",
  1773=>"111111110",
  1774=>"111111000",
  1775=>"000010010",
  1776=>"111101100",
  1777=>"011101111",
  1778=>"000000101",
  1779=>"111110000",
  1780=>"000001100",
  1781=>"101100111",
  1782=>"000000000",
  1783=>"101111001",
  1784=>"000000000",
  1785=>"001010111",
  1786=>"011001011",
  1787=>"011111111",
  1788=>"000000101",
  1789=>"101111101",
  1790=>"001011001",
  1791=>"011111111",
  1792=>"001001011",
  1793=>"000000000",
  1794=>"101100000",
  1795=>"110111111",
  1796=>"101100101",
  1797=>"111101000",
  1798=>"000111010",
  1799=>"110111010",
  1800=>"000000101",
  1801=>"111101000",
  1802=>"111100000",
  1803=>"000000111",
  1804=>"111100101",
  1805=>"000000111",
  1806=>"000100110",
  1807=>"010010010",
  1808=>"111101001",
  1809=>"010010000",
  1810=>"101111010",
  1811=>"000001010",
  1812=>"100000000",
  1813=>"001000000",
  1814=>"111110000",
  1815=>"001111111",
  1816=>"101101101",
  1817=>"000000000",
  1818=>"000011111",
  1819=>"000000111",
  1820=>"000011001",
  1821=>"110111011",
  1822=>"111100101",
  1823=>"000010010",
  1824=>"011010101",
  1825=>"000111101",
  1826=>"110111010",
  1827=>"001010111",
  1828=>"100101011",
  1829=>"000000000",
  1830=>"010111000",
  1831=>"000000000",
  1832=>"001111111",
  1833=>"010111111",
  1834=>"000000100",
  1835=>"110110010",
  1836=>"000110000",
  1837=>"111110000",
  1838=>"010011001",
  1839=>"000000001",
  1840=>"000101101",
  1841=>"100001011",
  1842=>"111111111",
  1843=>"000111111",
  1844=>"101011111",
  1845=>"111010100",
  1846=>"010000000",
  1847=>"100100011",
  1848=>"010011101",
  1849=>"101000000",
  1850=>"000010111",
  1851=>"010010011",
  1852=>"001000010",
  1853=>"101111111",
  1854=>"101101000",
  1855=>"001000001",
  1856=>"111101010",
  1857=>"010000101",
  1858=>"111111110",
  1859=>"011001100",
  1860=>"111000010",
  1861=>"000000101",
  1862=>"110111110",
  1863=>"111110111",
  1864=>"111111100",
  1865=>"000010101",
  1866=>"111001001",
  1867=>"000110111",
  1868=>"011111000",
  1869=>"000000110",
  1870=>"001000111",
  1871=>"000010111",
  1872=>"000111111",
  1873=>"010111010",
  1874=>"000011111",
  1875=>"001001001",
  1876=>"000000111",
  1877=>"011011000",
  1878=>"001111111",
  1879=>"111101101",
  1880=>"100010110",
  1881=>"000010010",
  1882=>"000011011",
  1883=>"000000011",
  1884=>"000010000",
  1885=>"100111111",
  1886=>"111111001",
  1887=>"100100110",
  1888=>"101001000",
  1889=>"110110010",
  1890=>"111101100",
  1891=>"000110110",
  1892=>"000001111",
  1893=>"000011011",
  1894=>"000000111",
  1895=>"111000000",
  1896=>"000010010",
  1897=>"111101101",
  1898=>"000101100",
  1899=>"011111010",
  1900=>"000010010",
  1901=>"000101000",
  1902=>"101111101",
  1903=>"000111111",
  1904=>"000000110",
  1905=>"000100101",
  1906=>"000001001",
  1907=>"111001000",
  1908=>"111011000",
  1909=>"000001111",
  1910=>"000000000",
  1911=>"111101101",
  1912=>"010010000",
  1913=>"000010010",
  1914=>"101111111",
  1915=>"000000000",
  1916=>"000010010",
  1917=>"000100110",
  1918=>"000011010",
  1919=>"101001010",
  1920=>"000001001",
  1921=>"110111100",
  1922=>"011000111",
  1923=>"000001000",
  1924=>"100101111",
  1925=>"111111100",
  1926=>"100000100",
  1927=>"100001111",
  1928=>"001101110",
  1929=>"111000110",
  1930=>"111111000",
  1931=>"111000000",
  1932=>"111101111",
  1933=>"111000000",
  1934=>"000010011",
  1935=>"100000000",
  1936=>"000111111",
  1937=>"101000010",
  1938=>"001000000",
  1939=>"101111111",
  1940=>"000001011",
  1941=>"111101101",
  1942=>"111110000",
  1943=>"000100111",
  1944=>"010011010",
  1945=>"101001000",
  1946=>"001101111",
  1947=>"010111101",
  1948=>"000111111",
  1949=>"000000101",
  1950=>"111011111",
  1951=>"101101000",
  1952=>"101011001",
  1953=>"010111111",
  1954=>"000110010",
  1955=>"000000010",
  1956=>"001011100",
  1957=>"000100100",
  1958=>"000001000",
  1959=>"000000111",
  1960=>"000000101",
  1961=>"010000010",
  1962=>"010111111",
  1963=>"000111110",
  1964=>"010110111",
  1965=>"111101100",
  1966=>"100111110",
  1967=>"000011111",
  1968=>"000110111",
  1969=>"000111011",
  1970=>"010000110",
  1971=>"001101001",
  1972=>"000000000",
  1973=>"000001011",
  1974=>"011100001",
  1975=>"000110111",
  1976=>"000000000",
  1977=>"001001011",
  1978=>"010111000",
  1979=>"000010000",
  1980=>"010010011",
  1981=>"111001111",
  1982=>"110101101",
  1983=>"011111111",
  1984=>"111111100",
  1985=>"110110011",
  1986=>"111111101",
  1987=>"101001111",
  1988=>"100000010",
  1989=>"111111101",
  1990=>"001111011",
  1991=>"111101000",
  1992=>"111001111",
  1993=>"111011111",
  1994=>"101000110",
  1995=>"101000010",
  1996=>"000000111",
  1997=>"100010010",
  1998=>"100111111",
  1999=>"000000100",
  2000=>"111101000",
  2001=>"000101110",
  2002=>"100000111",
  2003=>"010010000",
  2004=>"101101111",
  2005=>"001111010",
  2006=>"000010001",
  2007=>"010110111",
  2008=>"000010011",
  2009=>"000000010",
  2010=>"011111110",
  2011=>"111101101",
  2012=>"111011010",
  2013=>"101101111",
  2014=>"010000010",
  2015=>"110110111",
  2016=>"101000001",
  2017=>"111111101",
  2018=>"111111100",
  2019=>"110011011",
  2020=>"100000100",
  2021=>"010010000",
  2022=>"000000110",
  2023=>"000110110",
  2024=>"010111111",
  2025=>"000011000",
  2026=>"011101001",
  2027=>"000101110",
  2028=>"111101001",
  2029=>"111111011",
  2030=>"110111000",
  2031=>"000000100",
  2032=>"001000011",
  2033=>"100010001",
  2034=>"001111111",
  2035=>"000110000",
  2036=>"000010110",
  2037=>"101100111",
  2038=>"111000100",
  2039=>"000100100",
  2040=>"000101111",
  2041=>"100111111",
  2042=>"100111100",
  2043=>"101111001",
  2044=>"100010111",
  2045=>"000010000",
  2046=>"110000111",
  2047=>"000011011",
  2048=>"000100001",
  2049=>"111111000",
  2050=>"000000100",
  2051=>"000000000",
  2052=>"011111111",
  2053=>"101000101",
  2054=>"110101101",
  2055=>"000111010",
  2056=>"000000010",
  2057=>"101101101",
  2058=>"100000001",
  2059=>"000010110",
  2060=>"100000000",
  2061=>"000101000",
  2062=>"001011001",
  2063=>"000010001",
  2064=>"000010111",
  2065=>"111101111",
  2066=>"000100000",
  2067=>"011100000",
  2068=>"111111111",
  2069=>"110100000",
  2070=>"111011011",
  2071=>"111000111",
  2072=>"010101000",
  2073=>"101110010",
  2074=>"011001000",
  2075=>"000000000",
  2076=>"111111110",
  2077=>"100100001",
  2078=>"111000100",
  2079=>"000100000",
  2080=>"000101100",
  2081=>"111100000",
  2082=>"000100010",
  2083=>"000010010",
  2084=>"111001011",
  2085=>"111011000",
  2086=>"000000000",
  2087=>"001000110",
  2088=>"010111011",
  2089=>"100110010",
  2090=>"000000000",
  2091=>"100011010",
  2092=>"010101110",
  2093=>"111101000",
  2094=>"101101101",
  2095=>"111101010",
  2096=>"111000100",
  2097=>"111111111",
  2098=>"101111010",
  2099=>"100000111",
  2100=>"110100001",
  2101=>"010111010",
  2102=>"110000001",
  2103=>"000001111",
  2104=>"010010011",
  2105=>"010000101",
  2106=>"101101000",
  2107=>"000000100",
  2108=>"110010100",
  2109=>"110101000",
  2110=>"101100000",
  2111=>"011001000",
  2112=>"000011011",
  2113=>"111010100",
  2114=>"111111000",
  2115=>"110000001",
  2116=>"010000111",
  2117=>"001011011",
  2118=>"101001101",
  2119=>"111001001",
  2120=>"111001100",
  2121=>"100000101",
  2122=>"010000000",
  2123=>"101000001",
  2124=>"111101100",
  2125=>"111110110",
  2126=>"110111111",
  2127=>"010010010",
  2128=>"000000000",
  2129=>"111000000",
  2130=>"001101111",
  2131=>"011000111",
  2132=>"100111101",
  2133=>"110100000",
  2134=>"000000110",
  2135=>"111000000",
  2136=>"101101001",
  2137=>"111000100",
  2138=>"100110000",
  2139=>"010011100",
  2140=>"111010110",
  2141=>"001001000",
  2142=>"100111010",
  2143=>"000001100",
  2144=>"011111111",
  2145=>"111000000",
  2146=>"111000000",
  2147=>"000111010",
  2148=>"000110000",
  2149=>"100011011",
  2150=>"111111101",
  2151=>"000111001",
  2152=>"000000111",
  2153=>"101100101",
  2154=>"100000111",
  2155=>"000000000",
  2156=>"010110011",
  2157=>"000010000",
  2158=>"111100101",
  2159=>"011001100",
  2160=>"110110011",
  2161=>"000000101",
  2162=>"001000100",
  2163=>"000001000",
  2164=>"100000000",
  2165=>"101101101",
  2166=>"101101100",
  2167=>"111110100",
  2168=>"101001000",
  2169=>"010000100",
  2170=>"001111111",
  2171=>"101101111",
  2172=>"000111010",
  2173=>"110100100",
  2174=>"011000000",
  2175=>"010000100",
  2176=>"010010000",
  2177=>"101000000",
  2178=>"111111110",
  2179=>"000000100",
  2180=>"000011101",
  2181=>"101111001",
  2182=>"111010000",
  2183=>"000001001",
  2184=>"110001010",
  2185=>"000000001",
  2186=>"000101000",
  2187=>"000111000",
  2188=>"000010110",
  2189=>"100000111",
  2190=>"110000011",
  2191=>"100000001",
  2192=>"001011111",
  2193=>"110100010",
  2194=>"001000000",
  2195=>"000011011",
  2196=>"000000010",
  2197=>"101000000",
  2198=>"111101111",
  2199=>"000011011",
  2200=>"111110111",
  2201=>"101001000",
  2202=>"111000111",
  2203=>"101100101",
  2204=>"111000100",
  2205=>"111100000",
  2206=>"111000011",
  2207=>"111101000",
  2208=>"011011001",
  2209=>"011000010",
  2210=>"010001001",
  2211=>"000101100",
  2212=>"010000110",
  2213=>"000110100",
  2214=>"100110000",
  2215=>"010001000",
  2216=>"111111101",
  2217=>"000000111",
  2218=>"011100000",
  2219=>"011000000",
  2220=>"000101101",
  2221=>"111000000",
  2222=>"110001001",
  2223=>"111111111",
  2224=>"101111010",
  2225=>"000001100",
  2226=>"110001010",
  2227=>"001100100",
  2228=>"000001001",
  2229=>"000100000",
  2230=>"000011111",
  2231=>"010011010",
  2232=>"011011000",
  2233=>"000000000",
  2234=>"100100000",
  2235=>"111101101",
  2236=>"000101101",
  2237=>"111111111",
  2238=>"111100010",
  2239=>"000010001",
  2240=>"111100101",
  2241=>"111101101",
  2242=>"101000000",
  2243=>"101110111",
  2244=>"000000000",
  2245=>"110110001",
  2246=>"000000110",
  2247=>"000000111",
  2248=>"000000101",
  2249=>"000111010",
  2250=>"000111111",
  2251=>"000011001",
  2252=>"000000010",
  2253=>"000111111",
  2254=>"000111000",
  2255=>"000111110",
  2256=>"100100000",
  2257=>"000110111",
  2258=>"000010000",
  2259=>"000000101",
  2260=>"111000010",
  2261=>"000001000",
  2262=>"111000100",
  2263=>"000000111",
  2264=>"000000010",
  2265=>"000011011",
  2266=>"110110110",
  2267=>"001000000",
  2268=>"111110010",
  2269=>"100111000",
  2270=>"100011111",
  2271=>"001000101",
  2272=>"000000000",
  2273=>"111100100",
  2274=>"000010110",
  2275=>"100000011",
  2276=>"101000101",
  2277=>"111101111",
  2278=>"111101111",
  2279=>"011111110",
  2280=>"111111111",
  2281=>"100111001",
  2282=>"011100100",
  2283=>"000000110",
  2284=>"010111000",
  2285=>"010010101",
  2286=>"000000000",
  2287=>"011110110",
  2288=>"000001111",
  2289=>"011011100",
  2290=>"000010001",
  2291=>"110101101",
  2292=>"110001110",
  2293=>"001101000",
  2294=>"000000101",
  2295=>"101100101",
  2296=>"000000010",
  2297=>"001101011",
  2298=>"111001101",
  2299=>"000000001",
  2300=>"110001111",
  2301=>"001000000",
  2302=>"110011111",
  2303=>"111101101",
  2304=>"000110111",
  2305=>"000000000",
  2306=>"101111111",
  2307=>"000111000",
  2308=>"000100001",
  2309=>"000111110",
  2310=>"000000010",
  2311=>"111000100",
  2312=>"110111001",
  2313=>"010111011",
  2314=>"111111011",
  2315=>"111011000",
  2316=>"111111111",
  2317=>"000110110",
  2318=>"111111111",
  2319=>"001111111",
  2320=>"111111001",
  2321=>"111100000",
  2322=>"111111110",
  2323=>"000000001",
  2324=>"000000111",
  2325=>"000000000",
  2326=>"000000000",
  2327=>"110111011",
  2328=>"111111011",
  2329=>"101001001",
  2330=>"000000000",
  2331=>"101111111",
  2332=>"111111111",
  2333=>"111111101",
  2334=>"111111111",
  2335=>"111000011",
  2336=>"111110111",
  2337=>"000010000",
  2338=>"111111111",
  2339=>"110111010",
  2340=>"000000000",
  2341=>"001011011",
  2342=>"110111111",
  2343=>"000111111",
  2344=>"000000101",
  2345=>"000000111",
  2346=>"101111000",
  2347=>"100000101",
  2348=>"100000100",
  2349=>"001101001",
  2350=>"000111001",
  2351=>"111000000",
  2352=>"011111000",
  2353=>"001000110",
  2354=>"001000011",
  2355=>"000000101",
  2356=>"100110111",
  2357=>"001000111",
  2358=>"111110000",
  2359=>"000000000",
  2360=>"111000101",
  2361=>"111111111",
  2362=>"000000111",
  2363=>"110101011",
  2364=>"010110111",
  2365=>"011010010",
  2366=>"000000000",
  2367=>"111011011",
  2368=>"001101001",
  2369=>"110111111",
  2370=>"000000001",
  2371=>"100111011",
  2372=>"000000001",
  2373=>"111101101",
  2374=>"000001111",
  2375=>"101001000",
  2376=>"011011111",
  2377=>"111111111",
  2378=>"111001111",
  2379=>"111111010",
  2380=>"110000000",
  2381=>"001000011",
  2382=>"000000000",
  2383=>"001000101",
  2384=>"011111001",
  2385=>"111010000",
  2386=>"000101100",
  2387=>"110100010",
  2388=>"111000010",
  2389=>"010011011",
  2390=>"000001001",
  2391=>"111111111",
  2392=>"000000100",
  2393=>"000000000",
  2394=>"000000000",
  2395=>"111010000",
  2396=>"111111000",
  2397=>"010110010",
  2398=>"100111111",
  2399=>"011111110",
  2400=>"000000000",
  2401=>"111110010",
  2402=>"000010000",
  2403=>"100000000",
  2404=>"111000011",
  2405=>"100100010",
  2406=>"111111111",
  2407=>"111111111",
  2408=>"001000000",
  2409=>"100111111",
  2410=>"001101000",
  2411=>"111111101",
  2412=>"000001001",
  2413=>"010010010",
  2414=>"001111000",
  2415=>"000000111",
  2416=>"011000011",
  2417=>"000000000",
  2418=>"110111001",
  2419=>"111110111",
  2420=>"000000110",
  2421=>"101000000",
  2422=>"000000001",
  2423=>"000000001",
  2424=>"000101000",
  2425=>"000111111",
  2426=>"101101001",
  2427=>"000010010",
  2428=>"001001011",
  2429=>"011011010",
  2430=>"001111001",
  2431=>"111111111",
  2432=>"000101101",
  2433=>"011011111",
  2434=>"111111000",
  2435=>"110010000",
  2436=>"000000000",
  2437=>"111111111",
  2438=>"110010111",
  2439=>"001000111",
  2440=>"111001110",
  2441=>"000000000",
  2442=>"010111111",
  2443=>"000101010",
  2444=>"000111111",
  2445=>"000001000",
  2446=>"111111111",
  2447=>"100000000",
  2448=>"010000001",
  2449=>"101101111",
  2450=>"110100000",
  2451=>"000000000",
  2452=>"001011111",
  2453=>"111111101",
  2454=>"000111111",
  2455=>"110010000",
  2456=>"000000000",
  2457=>"000100000",
  2458=>"111111000",
  2459=>"010111000",
  2460=>"101011010",
  2461=>"000000000",
  2462=>"100000010",
  2463=>"110110010",
  2464=>"000100111",
  2465=>"111101000",
  2466=>"000000111",
  2467=>"111111010",
  2468=>"101001100",
  2469=>"000000000",
  2470=>"101111111",
  2471=>"110111111",
  2472=>"001101000",
  2473=>"000000001",
  2474=>"001000000",
  2475=>"110111000",
  2476=>"000000000",
  2477=>"100000000",
  2478=>"010011001",
  2479=>"001000000",
  2480=>"111101111",
  2481=>"110000111",
  2482=>"100111111",
  2483=>"100100000",
  2484=>"111111111",
  2485=>"011011011",
  2486=>"000100000",
  2487=>"101101111",
  2488=>"100011111",
  2489=>"100001101",
  2490=>"111111100",
  2491=>"111111010",
  2492=>"000000110",
  2493=>"000111111",
  2494=>"011100100",
  2495=>"001000000",
  2496=>"010111111",
  2497=>"111011000",
  2498=>"101111101",
  2499=>"101000010",
  2500=>"001001010",
  2501=>"001001011",
  2502=>"111101000",
  2503=>"111111111",
  2504=>"110001111",
  2505=>"111010110",
  2506=>"010111000",
  2507=>"101101111",
  2508=>"111111010",
  2509=>"101100100",
  2510=>"000000000",
  2511=>"000010000",
  2512=>"110110010",
  2513=>"010010011",
  2514=>"100101001",
  2515=>"000101111",
  2516=>"111111000",
  2517=>"101011100",
  2518=>"010111111",
  2519=>"110000000",
  2520=>"001000111",
  2521=>"000100001",
  2522=>"011001000",
  2523=>"000111111",
  2524=>"001000001",
  2525=>"111110101",
  2526=>"000000000",
  2527=>"001101000",
  2528=>"000000000",
  2529=>"111010101",
  2530=>"001000101",
  2531=>"100000000",
  2532=>"000110010",
  2533=>"001001111",
  2534=>"110110010",
  2535=>"000010100",
  2536=>"000111000",
  2537=>"100000000",
  2538=>"111111110",
  2539=>"111111111",
  2540=>"101101111",
  2541=>"001000101",
  2542=>"110111111",
  2543=>"010111110",
  2544=>"111110110",
  2545=>"100100101",
  2546=>"101111111",
  2547=>"010010001",
  2548=>"110101110",
  2549=>"100100101",
  2550=>"110000000",
  2551=>"111001111",
  2552=>"111001011",
  2553=>"101000010",
  2554=>"110111111",
  2555=>"010111111",
  2556=>"011011000",
  2557=>"000110111",
  2558=>"000000000",
  2559=>"111000000",
  2560=>"011011000",
  2561=>"001000000",
  2562=>"000000001",
  2563=>"101110110",
  2564=>"100111011",
  2565=>"110100000",
  2566=>"111010011",
  2567=>"000010010",
  2568=>"001111100",
  2569=>"001000110",
  2570=>"101000000",
  2571=>"111000000",
  2572=>"010111000",
  2573=>"000001000",
  2574=>"100011011",
  2575=>"110100111",
  2576=>"111110111",
  2577=>"000000000",
  2578=>"000000000",
  2579=>"000000010",
  2580=>"111001001",
  2581=>"000101101",
  2582=>"000101101",
  2583=>"000000110",
  2584=>"100111110",
  2585=>"000110111",
  2586=>"000101000",
  2587=>"111101000",
  2588=>"000000000",
  2589=>"001000111",
  2590=>"110000110",
  2591=>"000001000",
  2592=>"100000011",
  2593=>"010111010",
  2594=>"101000001",
  2595=>"000010000",
  2596=>"110111001",
  2597=>"111111101",
  2598=>"111000111",
  2599=>"011110000",
  2600=>"111111111",
  2601=>"111010010",
  2602=>"000010010",
  2603=>"111011111",
  2604=>"011001011",
  2605=>"000101010",
  2606=>"011000101",
  2607=>"000000110",
  2608=>"000001010",
  2609=>"101011011",
  2610=>"000000000",
  2611=>"101000111",
  2612=>"111000001",
  2613=>"111111000",
  2614=>"100100001",
  2615=>"000000001",
  2616=>"100000100",
  2617=>"111001000",
  2618=>"011100010",
  2619=>"011001000",
  2620=>"110110000",
  2621=>"001101000",
  2622=>"000000000",
  2623=>"011010000",
  2624=>"111111000",
  2625=>"111101101",
  2626=>"110111010",
  2627=>"001100000",
  2628=>"000000110",
  2629=>"111000101",
  2630=>"011001001",
  2631=>"011111111",
  2632=>"000000000",
  2633=>"110010010",
  2634=>"111000101",
  2635=>"000110000",
  2636=>"010000000",
  2637=>"000100100",
  2638=>"001101100",
  2639=>"111111111",
  2640=>"000001000",
  2641=>"111111001",
  2642=>"000001000",
  2643=>"001000000",
  2644=>"110000101",
  2645=>"000000001",
  2646=>"000101100",
  2647=>"000000000",
  2648=>"110100001",
  2649=>"111111011",
  2650=>"010100000",
  2651=>"110111000",
  2652=>"111011000",
  2653=>"001001011",
  2654=>"111111111",
  2655=>"001101001",
  2656=>"101000000",
  2657=>"111111010",
  2658=>"101000111",
  2659=>"000011000",
  2660=>"000111000",
  2661=>"111100100",
  2662=>"111111000",
  2663=>"111111101",
  2664=>"000000000",
  2665=>"111111000",
  2666=>"111110110",
  2667=>"111111111",
  2668=>"000000111",
  2669=>"000001010",
  2670=>"111110100",
  2671=>"000001001",
  2672=>"111001000",
  2673=>"010110111",
  2674=>"001000100",
  2675=>"101010111",
  2676=>"001011000",
  2677=>"100100000",
  2678=>"000110110",
  2679=>"111010001",
  2680=>"101111101",
  2681=>"110101000",
  2682=>"000000000",
  2683=>"001101111",
  2684=>"000110110",
  2685=>"100100001",
  2686=>"101111110",
  2687=>"000000000",
  2688=>"111111000",
  2689=>"111000001",
  2690=>"010000000",
  2691=>"111111111",
  2692=>"000101000",
  2693=>"001000000",
  2694=>"011101010",
  2695=>"011011000",
  2696=>"000101000",
  2697=>"001110001",
  2698=>"111111011",
  2699=>"010010111",
  2700=>"001000101",
  2701=>"001001111",
  2702=>"001000000",
  2703=>"011000001",
  2704=>"011001101",
  2705=>"111000000",
  2706=>"000000101",
  2707=>"001000100",
  2708=>"000110111",
  2709=>"000000111",
  2710=>"010111101",
  2711=>"110000001",
  2712=>"111111000",
  2713=>"111001110",
  2714=>"000000000",
  2715=>"101000000",
  2716=>"000000010",
  2717=>"000000001",
  2718=>"110001000",
  2719=>"001000011",
  2720=>"000000001",
  2721=>"111111011",
  2722=>"001010010",
  2723=>"111111000",
  2724=>"000000001",
  2725=>"110110000",
  2726=>"001001101",
  2727=>"111110111",
  2728=>"000000011",
  2729=>"111010111",
  2730=>"111111111",
  2731=>"000000000",
  2732=>"011000100",
  2733=>"111111000",
  2734=>"100000001",
  2735=>"000101011",
  2736=>"010000010",
  2737=>"000000000",
  2738=>"010001111",
  2739=>"001100100",
  2740=>"100101010",
  2741=>"000000011",
  2742=>"010110011",
  2743=>"111110111",
  2744=>"011011100",
  2745=>"000111110",
  2746=>"111101010",
  2747=>"001001111",
  2748=>"110110000",
  2749=>"001001001",
  2750=>"101110000",
  2751=>"001001101",
  2752=>"110101000",
  2753=>"010010000",
  2754=>"111000000",
  2755=>"101011000",
  2756=>"011010010",
  2757=>"001001111",
  2758=>"000100111",
  2759=>"110110000",
  2760=>"111110010",
  2761=>"001001001",
  2762=>"110111100",
  2763=>"110110111",
  2764=>"110010000",
  2765=>"000011011",
  2766=>"010000000",
  2767=>"111111101",
  2768=>"000000010",
  2769=>"011100010",
  2770=>"111111010",
  2771=>"110110010",
  2772=>"000000001",
  2773=>"101000000",
  2774=>"111111000",
  2775=>"001101010",
  2776=>"000001001",
  2777=>"011000000",
  2778=>"110100001",
  2779=>"000000111",
  2780=>"001100011",
  2781=>"011011111",
  2782=>"010100101",
  2783=>"000010111",
  2784=>"110111001",
  2785=>"000010001",
  2786=>"000001000",
  2787=>"011111011",
  2788=>"001001001",
  2789=>"000010011",
  2790=>"110110100",
  2791=>"011000100",
  2792=>"111101000",
  2793=>"000000000",
  2794=>"001100000",
  2795=>"001111111",
  2796=>"000110110",
  2797=>"101001001",
  2798=>"000000000",
  2799=>"000001011",
  2800=>"101001111",
  2801=>"100100111",
  2802=>"000000010",
  2803=>"001110110",
  2804=>"110101001",
  2805=>"000000000",
  2806=>"000010000",
  2807=>"110000110",
  2808=>"000000101",
  2809=>"010011110",
  2810=>"111111101",
  2811=>"110111111",
  2812=>"111100001",
  2813=>"001000010",
  2814=>"111111000",
  2815=>"111110010",
  2816=>"011011011",
  2817=>"000001000",
  2818=>"101000000",
  2819=>"001001101",
  2820=>"111100100",
  2821=>"111000000",
  2822=>"000111100",
  2823=>"001000011",
  2824=>"000111011",
  2825=>"001001111",
  2826=>"000000001",
  2827=>"000110000",
  2828=>"000010010",
  2829=>"010011100",
  2830=>"000100111",
  2831=>"000010110",
  2832=>"000000000",
  2833=>"101000111",
  2834=>"111010000",
  2835=>"111000000",
  2836=>"101101111",
  2837=>"111101000",
  2838=>"100100000",
  2839=>"000101111",
  2840=>"000000000",
  2841=>"001111110",
  2842=>"000001000",
  2843=>"111001111",
  2844=>"001001111",
  2845=>"100001000",
  2846=>"110100000",
  2847=>"100000110",
  2848=>"011001000",
  2849=>"001101111",
  2850=>"000111000",
  2851=>"000000000",
  2852=>"100110110",
  2853=>"110000110",
  2854=>"101000000",
  2855=>"000110000",
  2856=>"000010010",
  2857=>"001001001",
  2858=>"000000000",
  2859=>"111101111",
  2860=>"011111111",
  2861=>"000111111",
  2862=>"111111100",
  2863=>"001101000",
  2864=>"110101000",
  2865=>"001001010",
  2866=>"111111000",
  2867=>"101000000",
  2868=>"001000000",
  2869=>"111110111",
  2870=>"110000001",
  2871=>"101011110",
  2872=>"111101111",
  2873=>"101001101",
  2874=>"111111000",
  2875=>"000001011",
  2876=>"100000101",
  2877=>"010111010",
  2878=>"001000000",
  2879=>"000000010",
  2880=>"001010110",
  2881=>"110000011",
  2882=>"000000111",
  2883=>"001001001",
  2884=>"110010110",
  2885=>"001001000",
  2886=>"001000000",
  2887=>"010010010",
  2888=>"010111111",
  2889=>"111001000",
  2890=>"101000101",
  2891=>"111000101",
  2892=>"000010010",
  2893=>"011111110",
  2894=>"000110110",
  2895=>"100111110",
  2896=>"100000011",
  2897=>"010111000",
  2898=>"010111000",
  2899=>"011011001",
  2900=>"000000001",
  2901=>"000100100",
  2902=>"010011011",
  2903=>"101000001",
  2904=>"110111110",
  2905=>"001001000",
  2906=>"100101011",
  2907=>"000011010",
  2908=>"001000010",
  2909=>"100001001",
  2910=>"111111011",
  2911=>"000000010",
  2912=>"010000000",
  2913=>"110101101",
  2914=>"110000101",
  2915=>"001001000",
  2916=>"001100111",
  2917=>"111000101",
  2918=>"011001101",
  2919=>"111011000",
  2920=>"100110000",
  2921=>"000100000",
  2922=>"110001101",
  2923=>"101111000",
  2924=>"111001001",
  2925=>"101011001",
  2926=>"000000110",
  2927=>"001101101",
  2928=>"111111111",
  2929=>"001000000",
  2930=>"001000100",
  2931=>"000010000",
  2932=>"000100010",
  2933=>"101001000",
  2934=>"001000110",
  2935=>"110110100",
  2936=>"110001101",
  2937=>"011011111",
  2938=>"001111110",
  2939=>"000111111",
  2940=>"001001000",
  2941=>"010100101",
  2942=>"011000100",
  2943=>"101000001",
  2944=>"000110111",
  2945=>"111000000",
  2946=>"111001001",
  2947=>"000110110",
  2948=>"100011000",
  2949=>"111111111",
  2950=>"011100110",
  2951=>"000100001",
  2952=>"101111110",
  2953=>"100000000",
  2954=>"101100100",
  2955=>"110010000",
  2956=>"001001111",
  2957=>"000110010",
  2958=>"011001000",
  2959=>"001000110",
  2960=>"100100110",
  2961=>"101110110",
  2962=>"101000011",
  2963=>"111101000",
  2964=>"001110000",
  2965=>"111000001",
  2966=>"101111111",
  2967=>"000010000",
  2968=>"001000100",
  2969=>"101110100",
  2970=>"000010000",
  2971=>"000000101",
  2972=>"101001001",
  2973=>"111111011",
  2974=>"011001111",
  2975=>"010000010",
  2976=>"000011111",
  2977=>"001000100",
  2978=>"111001001",
  2979=>"010101001",
  2980=>"010111000",
  2981=>"000110110",
  2982=>"000110000",
  2983=>"000000000",
  2984=>"110010011",
  2985=>"110111101",
  2986=>"110111000",
  2987=>"101000111",
  2988=>"000010010",
  2989=>"111001001",
  2990=>"011001110",
  2991=>"000110010",
  2992=>"100000000",
  2993=>"100011010",
  2994=>"010001110",
  2995=>"001000000",
  2996=>"100011010",
  2997=>"000000101",
  2998=>"000011011",
  2999=>"011110100",
  3000=>"011000001",
  3001=>"000111110",
  3002=>"111000111",
  3003=>"010000001",
  3004=>"100110001",
  3005=>"000110110",
  3006=>"011011011",
  3007=>"111110010",
  3008=>"101000000",
  3009=>"001000000",
  3010=>"001101111",
  3011=>"000100110",
  3012=>"111000000",
  3013=>"000011011",
  3014=>"000100100",
  3015=>"000101111",
  3016=>"111101000",
  3017=>"000010100",
  3018=>"111001000",
  3019=>"111010010",
  3020=>"111000100",
  3021=>"000000000",
  3022=>"101000100",
  3023=>"010111000",
  3024=>"010110000",
  3025=>"011011110",
  3026=>"101010010",
  3027=>"000010111",
  3028=>"000011111",
  3029=>"001100110",
  3030=>"001001101",
  3031=>"000001111",
  3032=>"110010000",
  3033=>"000000000",
  3034=>"001111110",
  3035=>"101001001",
  3036=>"000001001",
  3037=>"110110101",
  3038=>"111110110",
  3039=>"001110100",
  3040=>"110000110",
  3041=>"101001000",
  3042=>"010011110",
  3043=>"011101111",
  3044=>"111000000",
  3045=>"010001011",
  3046=>"010111111",
  3047=>"111001111",
  3048=>"111000000",
  3049=>"111110001",
  3050=>"101000000",
  3051=>"000000000",
  3052=>"000001010",
  3053=>"010110010",
  3054=>"100000000",
  3055=>"000111001",
  3056=>"010010010",
  3057=>"000001110",
  3058=>"110111101",
  3059=>"000110010",
  3060=>"100111110",
  3061=>"111000000",
  3062=>"000000000",
  3063=>"001000000",
  3064=>"001000111",
  3065=>"100010101",
  3066=>"000101110",
  3067=>"000111111",
  3068=>"110000011",
  3069=>"111101000",
  3070=>"100110001",
  3071=>"111010001",
  3072=>"011011010",
  3073=>"110110110",
  3074=>"110110010",
  3075=>"110010010",
  3076=>"110111010",
  3077=>"100111110",
  3078=>"000000111",
  3079=>"010110010",
  3080=>"100000000",
  3081=>"100100110",
  3082=>"110011010",
  3083=>"111100100",
  3084=>"110010010",
  3085=>"101000000",
  3086=>"000100110",
  3087=>"000010110",
  3088=>"110110000",
  3089=>"111101101",
  3090=>"001011001",
  3091=>"100100110",
  3092=>"101000000",
  3093=>"000010100",
  3094=>"110100110",
  3095=>"001011011",
  3096=>"000101111",
  3097=>"000110000",
  3098=>"111101001",
  3099=>"110110110",
  3100=>"101111111",
  3101=>"100010110",
  3102=>"100011110",
  3103=>"010000010",
  3104=>"111011010",
  3105=>"010011011",
  3106=>"011101001",
  3107=>"000111010",
  3108=>"110100110",
  3109=>"011001011",
  3110=>"110110110",
  3111=>"000000100",
  3112=>"001111111",
  3113=>"001000101",
  3114=>"110110110",
  3115=>"110010010",
  3116=>"011111111",
  3117=>"000110110",
  3118=>"000000010",
  3119=>"111111110",
  3120=>"110000000",
  3121=>"000000010",
  3122=>"001011011",
  3123=>"110110110",
  3124=>"011011000",
  3125=>"110000000",
  3126=>"110110011",
  3127=>"110110100",
  3128=>"010010100",
  3129=>"111001011",
  3130=>"001101001",
  3131=>"110110010",
  3132=>"110010100",
  3133=>"011011011",
  3134=>"100000100",
  3135=>"100000000",
  3136=>"110110110",
  3137=>"111111111",
  3138=>"111000000",
  3139=>"110110110",
  3140=>"111011000",
  3141=>"011001000",
  3142=>"100000110",
  3143=>"001000111",
  3144=>"110010100",
  3145=>"011101111",
  3146=>"100110110",
  3147=>"110100010",
  3148=>"001001001",
  3149=>"001000101",
  3150=>"000111111",
  3151=>"011010011",
  3152=>"110111111",
  3153=>"000000000",
  3154=>"110010111",
  3155=>"110110100",
  3156=>"100110010",
  3157=>"000100100",
  3158=>"100100100",
  3159=>"000111111",
  3160=>"101101000",
  3161=>"001111111",
  3162=>"110110011",
  3163=>"110110000",
  3164=>"110100100",
  3165=>"100100100",
  3166=>"110110110",
  3167=>"100011110",
  3168=>"110110110",
  3169=>"110110000",
  3170=>"110110110",
  3171=>"011100110",
  3172=>"110110111",
  3173=>"001111110",
  3174=>"000001000",
  3175=>"100000100",
  3176=>"000010010",
  3177=>"000000100",
  3178=>"000111000",
  3179=>"100010101",
  3180=>"111011010",
  3181=>"001001001",
  3182=>"111000110",
  3183=>"110111110",
  3184=>"110100000",
  3185=>"110010000",
  3186=>"110110110",
  3187=>"000000110",
  3188=>"011010100",
  3189=>"100100100",
  3190=>"111110011",
  3191=>"110110000",
  3192=>"100100000",
  3193=>"111001000",
  3194=>"000001010",
  3195=>"011101111",
  3196=>"100110000",
  3197=>"001001000",
  3198=>"101101001",
  3199=>"100100111",
  3200=>"110110000",
  3201=>"000100110",
  3202=>"110110000",
  3203=>"110011111",
  3204=>"000000010",
  3205=>"111010111",
  3206=>"000010100",
  3207=>"110100100",
  3208=>"111111111",
  3209=>"110000010",
  3210=>"100100110",
  3211=>"000001001",
  3212=>"001000011",
  3213=>"011110011",
  3214=>"111100111",
  3215=>"100100110",
  3216=>"110000000",
  3217=>"011111110",
  3218=>"000000111",
  3219=>"110000000",
  3220=>"100110110",
  3221=>"010110110",
  3222=>"010011010",
  3223=>"101000100",
  3224=>"010110110",
  3225=>"111000001",
  3226=>"000010000",
  3227=>"100110010",
  3228=>"110000000",
  3229=>"100111000",
  3230=>"001010101",
  3231=>"001011111",
  3232=>"110110100",
  3233=>"110110001",
  3234=>"000000000",
  3235=>"111111110",
  3236=>"100011111",
  3237=>"110110010",
  3238=>"011001001",
  3239=>"000001001",
  3240=>"110110110",
  3241=>"110100000",
  3242=>"011010011",
  3243=>"111000110",
  3244=>"101001001",
  3245=>"000000100",
  3246=>"110011010",
  3247=>"000000000",
  3248=>"000011111",
  3249=>"100100010",
  3250=>"000001001",
  3251=>"110010000",
  3252=>"001001111",
  3253=>"111110111",
  3254=>"000010101",
  3255=>"000011111",
  3256=>"110110100",
  3257=>"011011011",
  3258=>"010010000",
  3259=>"100110000",
  3260=>"101000100",
  3261=>"011011011",
  3262=>"000000000",
  3263=>"100000110",
  3264=>"100010000",
  3265=>"110110010",
  3266=>"000011011",
  3267=>"001011111",
  3268=>"111101101",
  3269=>"100110100",
  3270=>"110010110",
  3271=>"011011011",
  3272=>"000101101",
  3273=>"111110010",
  3274=>"110010100",
  3275=>"100100110",
  3276=>"100100100",
  3277=>"110000111",
  3278=>"100111111",
  3279=>"011011011",
  3280=>"011111011",
  3281=>"100000000",
  3282=>"110000100",
  3283=>"010010010",
  3284=>"000011011",
  3285=>"111111000",
  3286=>"110010110",
  3287=>"011110111",
  3288=>"110110100",
  3289=>"100100110",
  3290=>"011100101",
  3291=>"001101101",
  3292=>"110110000",
  3293=>"001000001",
  3294=>"000100100",
  3295=>"110110110",
  3296=>"000000000",
  3297=>"000000010",
  3298=>"000011111",
  3299=>"110110000",
  3300=>"110110110",
  3301=>"111111010",
  3302=>"110010110",
  3303=>"000010111",
  3304=>"001000000",
  3305=>"111011000",
  3306=>"011011011",
  3307=>"111111111",
  3308=>"100110110",
  3309=>"110010010",
  3310=>"011011011",
  3311=>"000100111",
  3312=>"111000100",
  3313=>"011001111",
  3314=>"100100110",
  3315=>"100100100",
  3316=>"111101111",
  3317=>"110000000",
  3318=>"000000110",
  3319=>"100100101",
  3320=>"100110110",
  3321=>"011000000",
  3322=>"000000001",
  3323=>"000111111",
  3324=>"000111111",
  3325=>"010011110",
  3326=>"000010111",
  3327=>"111110111",
  3328=>"001000111",
  3329=>"110010100",
  3330=>"100000111",
  3331=>"010110100",
  3332=>"000100110",
  3333=>"110101011",
  3334=>"111111011",
  3335=>"111111111",
  3336=>"101000010",
  3337=>"101000010",
  3338=>"010011000",
  3339=>"000101101",
  3340=>"001101000",
  3341=>"101101111",
  3342=>"100100110",
  3343=>"111100000",
  3344=>"111101000",
  3345=>"101000000",
  3346=>"100000000",
  3347=>"100010000",
  3348=>"110110001",
  3349=>"101000111",
  3350=>"111011000",
  3351=>"011000000",
  3352=>"000100100",
  3353=>"101001011",
  3354=>"101101111",
  3355=>"101101101",
  3356=>"101101101",
  3357=>"111010111",
  3358=>"000111111",
  3359=>"101000111",
  3360=>"000000000",
  3361=>"000000000",
  3362=>"011010011",
  3363=>"000011000",
  3364=>"101001001",
  3365=>"001001011",
  3366=>"000110111",
  3367=>"011011000",
  3368=>"011010010",
  3369=>"010100111",
  3370=>"110000110",
  3371=>"010010000",
  3372=>"010000010",
  3373=>"000111111",
  3374=>"000100110",
  3375=>"100000001",
  3376=>"000000000",
  3377=>"001111101",
  3378=>"000000000",
  3379=>"101101101",
  3380=>"010010001",
  3381=>"111000101",
  3382=>"111110100",
  3383=>"100000010",
  3384=>"000000001",
  3385=>"000000111",
  3386=>"101111110",
  3387=>"111000000",
  3388=>"100001001",
  3389=>"111111000",
  3390=>"000000000",
  3391=>"100110100",
  3392=>"000000000",
  3393=>"000101100",
  3394=>"001000000",
  3395=>"011011001",
  3396=>"001101010",
  3397=>"111000000",
  3398=>"000010110",
  3399=>"111000011",
  3400=>"111001101",
  3401=>"111111011",
  3402=>"000001011",
  3403=>"000101111",
  3404=>"000100111",
  3405=>"100100000",
  3406=>"000001011",
  3407=>"110000111",
  3408=>"000000010",
  3409=>"000100000",
  3410=>"111111111",
  3411=>"111001000",
  3412=>"000000111",
  3413=>"110011001",
  3414=>"000100101",
  3415=>"000000000",
  3416=>"001110111",
  3417=>"001011110",
  3418=>"000000111",
  3419=>"001001111",
  3420=>"000000110",
  3421=>"001111111",
  3422=>"101111001",
  3423=>"110110110",
  3424=>"100101101",
  3425=>"010110010",
  3426=>"000000111",
  3427=>"011011000",
  3428=>"000111110",
  3429=>"111100011",
  3430=>"111111100",
  3431=>"101000010",
  3432=>"000100111",
  3433=>"011101100",
  3434=>"101010111",
  3435=>"011101111",
  3436=>"000110101",
  3437=>"000000010",
  3438=>"101000011",
  3439=>"100010011",
  3440=>"000100100",
  3441=>"000000000",
  3442=>"110111001",
  3443=>"000101111",
  3444=>"000000000",
  3445=>"001001101",
  3446=>"101000000",
  3447=>"110010100",
  3448=>"011000101",
  3449=>"111110101",
  3450=>"000110001",
  3451=>"111000101",
  3452=>"010111001",
  3453=>"100000000",
  3454=>"111111000",
  3455=>"010010011",
  3456=>"101000000",
  3457=>"100100010",
  3458=>"001011111",
  3459=>"111010010",
  3460=>"000111111",
  3461=>"011010001",
  3462=>"100110100",
  3463=>"000000010",
  3464=>"001011000",
  3465=>"000010010",
  3466=>"101111110",
  3467=>"010000000",
  3468=>"110000000",
  3469=>"110000100",
  3470=>"101001000",
  3471=>"100000000",
  3472=>"100000111",
  3473=>"111000000",
  3474=>"111000000",
  3475=>"000111011",
  3476=>"111010010",
  3477=>"100000000",
  3478=>"101110111",
  3479=>"101110111",
  3480=>"111111000",
  3481=>"010000111",
  3482=>"101100111",
  3483=>"110000000",
  3484=>"000000011",
  3485=>"101101110",
  3486=>"010101101",
  3487=>"000011000",
  3488=>"011110110",
  3489=>"111110000",
  3490=>"011010010",
  3491=>"101111000",
  3492=>"000010110",
  3493=>"000100111",
  3494=>"110101101",
  3495=>"000000111",
  3496=>"000100110",
  3497=>"000101101",
  3498=>"100000001",
  3499=>"000000000",
  3500=>"000111111",
  3501=>"001111010",
  3502=>"010011010",
  3503=>"111111010",
  3504=>"001110000",
  3505=>"001001011",
  3506=>"100110001",
  3507=>"111011011",
  3508=>"111100000",
  3509=>"111001100",
  3510=>"111000110",
  3511=>"000100101",
  3512=>"101100110",
  3513=>"000000100",
  3514=>"101110111",
  3515=>"101111001",
  3516=>"010111111",
  3517=>"111000000",
  3518=>"001001101",
  3519=>"010000000",
  3520=>"101101101",
  3521=>"101000000",
  3522=>"111101100",
  3523=>"000000100",
  3524=>"000000000",
  3525=>"111111011",
  3526=>"000111011",
  3527=>"000000001",
  3528=>"010000110",
  3529=>"000100000",
  3530=>"111011011",
  3531=>"010000101",
  3532=>"100100011",
  3533=>"000110100",
  3534=>"110101000",
  3535=>"000000100",
  3536=>"000110111",
  3537=>"001001011",
  3538=>"100111111",
  3539=>"011111111",
  3540=>"001001010",
  3541=>"101101000",
  3542=>"000101111",
  3543=>"000000000",
  3544=>"011111000",
  3545=>"101111110",
  3546=>"110101111",
  3547=>"000000100",
  3548=>"111111000",
  3549=>"000010111",
  3550=>"000001100",
  3551=>"001000111",
  3552=>"001000000",
  3553=>"000100100",
  3554=>"111111111",
  3555=>"000110110",
  3556=>"001000000",
  3557=>"111111001",
  3558=>"000010110",
  3559=>"111110110",
  3560=>"100111000",
  3561=>"000001100",
  3562=>"010110001",
  3563=>"101101111",
  3564=>"110010000",
  3565=>"001110111",
  3566=>"000010010",
  3567=>"101110111",
  3568=>"000100000",
  3569=>"011100100",
  3570=>"000110010",
  3571=>"110110010",
  3572=>"100101011",
  3573=>"000000111",
  3574=>"001000110",
  3575=>"010010010",
  3576=>"000000000",
  3577=>"100100000",
  3578=>"111111010",
  3579=>"010101000",
  3580=>"101100111",
  3581=>"011011101",
  3582=>"000111110",
  3583=>"000000111",
  3584=>"110101011",
  3585=>"111110000",
  3586=>"000000000",
  3587=>"111000110",
  3588=>"111000000",
  3589=>"111100000",
  3590=>"111000101",
  3591=>"000111111",
  3592=>"000101010",
  3593=>"010010001",
  3594=>"100100000",
  3595=>"011000000",
  3596=>"000011111",
  3597=>"110100010",
  3598=>"111111111",
  3599=>"111000011",
  3600=>"101101101",
  3601=>"100000100",
  3602=>"000000100",
  3603=>"111000000",
  3604=>"101000111",
  3605=>"000001000",
  3606=>"101001001",
  3607=>"001110010",
  3608=>"000101011",
  3609=>"100010010",
  3610=>"111111100",
  3611=>"111101101",
  3612=>"101100010",
  3613=>"001000111",
  3614=>"011010000",
  3615=>"111101000",
  3616=>"000111011",
  3617=>"000000001",
  3618=>"000111111",
  3619=>"000010010",
  3620=>"000010110",
  3621=>"010110000",
  3622=>"101111011",
  3623=>"001110111",
  3624=>"000000111",
  3625=>"111101101",
  3626=>"111000000",
  3627=>"010001010",
  3628=>"111011111",
  3629=>"111001111",
  3630=>"011000000",
  3631=>"000011000",
  3632=>"000010001",
  3633=>"011100110",
  3634=>"000111000",
  3635=>"010001111",
  3636=>"000000001",
  3637=>"010000100",
  3638=>"010000000",
  3639=>"000111000",
  3640=>"100010000",
  3641=>"100000000",
  3642=>"000100000",
  3643=>"000000010",
  3644=>"000000000",
  3645=>"001111010",
  3646=>"000000000",
  3647=>"111011000",
  3648=>"111111111",
  3649=>"111110000",
  3650=>"010010000",
  3651=>"101110100",
  3652=>"110000010",
  3653=>"101010000",
  3654=>"010110100",
  3655=>"111110111",
  3656=>"011101011",
  3657=>"000111011",
  3658=>"111101101",
  3659=>"111010100",
  3660=>"111011010",
  3661=>"110110110",
  3662=>"011001001",
  3663=>"111100111",
  3664=>"101000000",
  3665=>"111111111",
  3666=>"001101111",
  3667=>"010001001",
  3668=>"010000100",
  3669=>"111100100",
  3670=>"000111011",
  3671=>"111010111",
  3672=>"011111001",
  3673=>"011010000",
  3674=>"101111101",
  3675=>"001011011",
  3676=>"110010010",
  3677=>"110001000",
  3678=>"111101101",
  3679=>"000101000",
  3680=>"111011001",
  3681=>"101000000",
  3682=>"000000001",
  3683=>"100011011",
  3684=>"110110010",
  3685=>"110111101",
  3686=>"010111110",
  3687=>"010111010",
  3688=>"000010111",
  3689=>"001000000",
  3690=>"000010101",
  3691=>"111111111",
  3692=>"001111110",
  3693=>"111101101",
  3694=>"000011011",
  3695=>"111111101",
  3696=>"111101001",
  3697=>"010000000",
  3698=>"111000000",
  3699=>"000111110",
  3700=>"000000000",
  3701=>"101000000",
  3702=>"011111111",
  3703=>"010000000",
  3704=>"101001001",
  3705=>"010110111",
  3706=>"101000000",
  3707=>"000000101",
  3708=>"100100100",
  3709=>"000100100",
  3710=>"011001001",
  3711=>"101100111",
  3712=>"000010010",
  3713=>"011111001",
  3714=>"000000010",
  3715=>"010000000",
  3716=>"110101101",
  3717=>"111110000",
  3718=>"110011100",
  3719=>"000000010",
  3720=>"110000110",
  3721=>"001000000",
  3722=>"111101111",
  3723=>"000010111",
  3724=>"111101101",
  3725=>"000101111",
  3726=>"110111111",
  3727=>"100000000",
  3728=>"100101101",
  3729=>"101111110",
  3730=>"111111001",
  3731=>"110011111",
  3732=>"000100011",
  3733=>"111100000",
  3734=>"011111111",
  3735=>"111101100",
  3736=>"011111010",
  3737=>"011000000",
  3738=>"000010010",
  3739=>"111000000",
  3740=>"000110111",
  3741=>"000101101",
  3742=>"010010100",
  3743=>"000010010",
  3744=>"000110001",
  3745=>"100000010",
  3746=>"010110010",
  3747=>"000111111",
  3748=>"111100100",
  3749=>"000110110",
  3750=>"000110110",
  3751=>"010010000",
  3752=>"101000000",
  3753=>"100111000",
  3754=>"010100000",
  3755=>"101100000",
  3756=>"000011010",
  3757=>"111000001",
  3758=>"110010001",
  3759=>"100100000",
  3760=>"011000000",
  3761=>"001001001",
  3762=>"111000011",
  3763=>"010100101",
  3764=>"010001001",
  3765=>"011011010",
  3766=>"000011001",
  3767=>"010011110",
  3768=>"001001000",
  3769=>"001101110",
  3770=>"111010010",
  3771=>"111010011",
  3772=>"010111111",
  3773=>"111111010",
  3774=>"111111110",
  3775=>"000000000",
  3776=>"101000001",
  3777=>"000000111",
  3778=>"001010011",
  3779=>"011011011",
  3780=>"000000011",
  3781=>"011100101",
  3782=>"111111110",
  3783=>"000010010",
  3784=>"011001000",
  3785=>"111010111",
  3786=>"000111111",
  3787=>"010000000",
  3788=>"111000100",
  3789=>"000111100",
  3790=>"010010000",
  3791=>"111101101",
  3792=>"000111111",
  3793=>"110011010",
  3794=>"001000000",
  3795=>"111101111",
  3796=>"000010010",
  3797=>"110100110",
  3798=>"000100000",
  3799=>"111101000",
  3800=>"010110100",
  3801=>"100101000",
  3802=>"110001000",
  3803=>"011000101",
  3804=>"111111001",
  3805=>"010101101",
  3806=>"000010010",
  3807=>"101101000",
  3808=>"101000110",
  3809=>"010100101",
  3810=>"110111111",
  3811=>"010000010",
  3812=>"110000101",
  3813=>"111111100",
  3814=>"011100000",
  3815=>"111110100",
  3816=>"111100111",
  3817=>"001000100",
  3818=>"101000000",
  3819=>"000111110",
  3820=>"111101001",
  3821=>"010000000",
  3822=>"000000001",
  3823=>"000000111",
  3824=>"011100000",
  3825=>"111001110",
  3826=>"010110100",
  3827=>"110100000",
  3828=>"010011011",
  3829=>"101101101",
  3830=>"001000000",
  3831=>"000000100",
  3832=>"111111010",
  3833=>"101111010",
  3834=>"010000000",
  3835=>"001101111",
  3836=>"100000011",
  3837=>"011000000",
  3838=>"000001011",
  3839=>"000010110",
  3840=>"101100010",
  3841=>"011111011",
  3842=>"100110010",
  3843=>"111111000",
  3844=>"000000110",
  3845=>"111001111",
  3846=>"111100111",
  3847=>"000111101",
  3848=>"000010110",
  3849=>"000000111",
  3850=>"111001100",
  3851=>"000101110",
  3852=>"000000000",
  3853=>"000010111",
  3854=>"000000000",
  3855=>"111111010",
  3856=>"110000011",
  3857=>"111000000",
  3858=>"100010111",
  3859=>"000111100",
  3860=>"111100100",
  3861=>"000001111",
  3862=>"011110010",
  3863=>"011111000",
  3864=>"100100101",
  3865=>"000011110",
  3866=>"010011011",
  3867=>"000010011",
  3868=>"011100010",
  3869=>"000000011",
  3870=>"000001000",
  3871=>"010110110",
  3872=>"111111000",
  3873=>"011111000",
  3874=>"111110101",
  3875=>"111111101",
  3876=>"110100110",
  3877=>"011011000",
  3878=>"000100010",
  3879=>"000111010",
  3880=>"000100010",
  3881=>"011101111",
  3882=>"000000101",
  3883=>"000010111",
  3884=>"000000000",
  3885=>"000110111",
  3886=>"111111110",
  3887=>"111000101",
  3888=>"000000010",
  3889=>"101111110",
  3890=>"111111011",
  3891=>"111101100",
  3892=>"111101111",
  3893=>"111000000",
  3894=>"000000011",
  3895=>"000100100",
  3896=>"000000010",
  3897=>"000000100",
  3898=>"110000100",
  3899=>"011011101",
  3900=>"111000000",
  3901=>"001111111",
  3902=>"110000000",
  3903=>"000011011",
  3904=>"111111000",
  3905=>"101111001",
  3906=>"111111011",
  3907=>"001100000",
  3908=>"011111011",
  3909=>"101111100",
  3910=>"000111110",
  3911=>"111111111",
  3912=>"100010000",
  3913=>"100101000",
  3914=>"010010010",
  3915=>"111000000",
  3916=>"111111000",
  3917=>"011111111",
  3918=>"000011001",
  3919=>"000000000",
  3920=>"000000000",
  3921=>"011111110",
  3922=>"111101100",
  3923=>"110110100",
  3924=>"000010111",
  3925=>"000000100",
  3926=>"000100111",
  3927=>"101000001",
  3928=>"110111110",
  3929=>"111111000",
  3930=>"010010001",
  3931=>"111111010",
  3932=>"000010010",
  3933=>"111110010",
  3934=>"000000001",
  3935=>"100000001",
  3936=>"110100000",
  3937=>"111011000",
  3938=>"000100111",
  3939=>"001001000",
  3940=>"010011011",
  3941=>"011111011",
  3942=>"000000000",
  3943=>"111011010",
  3944=>"111111111",
  3945=>"000000111",
  3946=>"000000111",
  3947=>"001010000",
  3948=>"000000000",
  3949=>"010111000",
  3950=>"000000100",
  3951=>"111000000",
  3952=>"100111110",
  3953=>"110001001",
  3954=>"101000110",
  3955=>"111011111",
  3956=>"100111111",
  3957=>"011011001",
  3958=>"000001000",
  3959=>"000000100",
  3960=>"111110111",
  3961=>"011011000",
  3962=>"111101111",
  3963=>"110110100",
  3964=>"000001100",
  3965=>"010011011",
  3966=>"101111111",
  3967=>"000010011",
  3968=>"101000101",
  3969=>"111010001",
  3970=>"000111011",
  3971=>"111111100",
  3972=>"011100000",
  3973=>"000000000",
  3974=>"110110000",
  3975=>"100100000",
  3976=>"001111011",
  3977=>"110100100",
  3978=>"100000000",
  3979=>"000111111",
  3980=>"000000111",
  3981=>"111100000",
  3982=>"000000000",
  3983=>"011000000",
  3984=>"111100111",
  3985=>"101000100",
  3986=>"000000111",
  3987=>"000010000",
  3988=>"010101000",
  3989=>"111000000",
  3990=>"111001000",
  3991=>"000000000",
  3992=>"000000000",
  3993=>"011000011",
  3994=>"011111111",
  3995=>"111000100",
  3996=>"111101111",
  3997=>"011111111",
  3998=>"000111111",
  3999=>"100000000",
  4000=>"111111000",
  4001=>"111011000",
  4002=>"000001111",
  4003=>"011111000",
  4004=>"100000110",
  4005=>"111011011",
  4006=>"011010010",
  4007=>"000100000",
  4008=>"011011101",
  4009=>"000111101",
  4010=>"011000101",
  4011=>"111000100",
  4012=>"101101111",
  4013=>"111111101",
  4014=>"111001000",
  4015=>"000000000",
  4016=>"101001111",
  4017=>"000110000",
  4018=>"011011010",
  4019=>"111011001",
  4020=>"111111110",
  4021=>"111000010",
  4022=>"100111011",
  4023=>"000100111",
  4024=>"011000010",
  4025=>"001001100",
  4026=>"000000001",
  4027=>"001111111",
  4028=>"110000001",
  4029=>"010111111",
  4030=>"000111100",
  4031=>"000000111",
  4032=>"111111000",
  4033=>"000000101",
  4034=>"010001000",
  4035=>"111111011",
  4036=>"000000001",
  4037=>"011111011",
  4038=>"111111100",
  4039=>"111000101",
  4040=>"111111101",
  4041=>"000111111",
  4042=>"101111111",
  4043=>"000000011",
  4044=>"100100110",
  4045=>"110110000",
  4046=>"111111111",
  4047=>"111010100",
  4048=>"000111111",
  4049=>"100000000",
  4050=>"101101101",
  4051=>"100101100",
  4052=>"001100101",
  4053=>"010011011",
  4054=>"111100000",
  4055=>"110100100",
  4056=>"100000111",
  4057=>"000111100",
  4058=>"111111000",
  4059=>"111011000",
  4060=>"000000011",
  4061=>"100011000",
  4062=>"010000000",
  4063=>"100111111",
  4064=>"000111110",
  4065=>"001000000",
  4066=>"111000001",
  4067=>"000001000",
  4068=>"101000000",
  4069=>"010000000",
  4070=>"111111111",
  4071=>"110110000",
  4072=>"100111110",
  4073=>"000010111",
  4074=>"100000001",
  4075=>"001000000",
  4076=>"111001001",
  4077=>"000001111",
  4078=>"010000110",
  4079=>"011000100",
  4080=>"111000101",
  4081=>"111110111",
  4082=>"000100011",
  4083=>"111111011",
  4084=>"001011001",
  4085=>"000000111",
  4086=>"001001000",
  4087=>"011000000",
  4088=>"110111111",
  4089=>"111111111",
  4090=>"001000000",
  4091=>"111101101",
  4092=>"111011000",
  4093=>"000000111",
  4094=>"000110011",
  4095=>"011111010",
  4096=>"001001010",
  4097=>"111110010",
  4098=>"010000011",
  4099=>"001110110",
  4100=>"100011001",
  4101=>"000011111",
  4102=>"011110101",
  4103=>"010000000",
  4104=>"111110000",
  4105=>"111111000",
  4106=>"100100100",
  4107=>"000000111",
  4108=>"010000000",
  4109=>"000000011",
  4110=>"011001010",
  4111=>"001000000",
  4112=>"111111111",
  4113=>"010111001",
  4114=>"000000000",
  4115=>"111000011",
  4116=>"110110100",
  4117=>"011000000",
  4118=>"011000001",
  4119=>"001000011",
  4120=>"010010110",
  4121=>"111111111",
  4122=>"100111111",
  4123=>"111111011",
  4124=>"111111100",
  4125=>"010100000",
  4126=>"000111011",
  4127=>"101101111",
  4128=>"111100001",
  4129=>"010110111",
  4130=>"111001011",
  4131=>"010111010",
  4132=>"001001000",
  4133=>"100100000",
  4134=>"000011110",
  4135=>"101111000",
  4136=>"110100000",
  4137=>"000110100",
  4138=>"111001001",
  4139=>"100000000",
  4140=>"101001111",
  4141=>"110111010",
  4142=>"001110111",
  4143=>"101000000",
  4144=>"111111000",
  4145=>"101101001",
  4146=>"010001000",
  4147=>"111011101",
  4148=>"101000000",
  4149=>"101111011",
  4150=>"100100001",
  4151=>"000111000",
  4152=>"001000101",
  4153=>"000100111",
  4154=>"100100111",
  4155=>"100001001",
  4156=>"011101000",
  4157=>"101101011",
  4158=>"010000000",
  4159=>"100000000",
  4160=>"011110010",
  4161=>"100101010",
  4162=>"010111100",
  4163=>"000100100",
  4164=>"000000111",
  4165=>"001000000",
  4166=>"110111101",
  4167=>"010000111",
  4168=>"001000000",
  4169=>"111110100",
  4170=>"010010010",
  4171=>"000000000",
  4172=>"000111101",
  4173=>"101101111",
  4174=>"001101100",
  4175=>"111010111",
  4176=>"101111111",
  4177=>"000000111",
  4178=>"001111010",
  4179=>"111000000",
  4180=>"101111111",
  4181=>"000100100",
  4182=>"111101100",
  4183=>"110011000",
  4184=>"111001101",
  4185=>"100101001",
  4186=>"100111001",
  4187=>"100100000",
  4188=>"010111101",
  4189=>"001100001",
  4190=>"010111111",
  4191=>"001001001",
  4192=>"100010011",
  4193=>"010010110",
  4194=>"110111001",
  4195=>"111111110",
  4196=>"100000100",
  4197=>"001001101",
  4198=>"111111111",
  4199=>"111111000",
  4200=>"010101001",
  4201=>"000111111",
  4202=>"111101000",
  4203=>"101100101",
  4204=>"000101111",
  4205=>"011110010",
  4206=>"111111011",
  4207=>"111101101",
  4208=>"100000100",
  4209=>"000111111",
  4210=>"000001001",
  4211=>"000000010",
  4212=>"111001100",
  4213=>"000000010",
  4214=>"000010110",
  4215=>"111111000",
  4216=>"010101010",
  4217=>"110110111",
  4218=>"011000000",
  4219=>"001000101",
  4220=>"000000001",
  4221=>"100000000",
  4222=>"111000000",
  4223=>"000010111",
  4224=>"111010000",
  4225=>"000111000",
  4226=>"111100000",
  4227=>"111000101",
  4228=>"110111000",
  4229=>"101110110",
  4230=>"001001000",
  4231=>"010000001",
  4232=>"001000000",
  4233=>"010000110",
  4234=>"000011111",
  4235=>"000010101",
  4236=>"111100010",
  4237=>"011001001",
  4238=>"111111101",
  4239=>"001010000",
  4240=>"101100011",
  4241=>"010000010",
  4242=>"101000000",
  4243=>"011010011",
  4244=>"011011111",
  4245=>"111110111",
  4246=>"101101101",
  4247=>"000000000",
  4248=>"111011101",
  4249=>"100111110",
  4250=>"011011000",
  4251=>"010011110",
  4252=>"000011100",
  4253=>"110111111",
  4254=>"101100110",
  4255=>"111000111",
  4256=>"100000100",
  4257=>"010000000",
  4258=>"101001000",
  4259=>"111111111",
  4260=>"110110111",
  4261=>"000000000",
  4262=>"000010000",
  4263=>"000000010",
  4264=>"111111111",
  4265=>"010010111",
  4266=>"101000000",
  4267=>"000010111",
  4268=>"000000111",
  4269=>"000111101",
  4270=>"100100100",
  4271=>"110111111",
  4272=>"010100001",
  4273=>"000011000",
  4274=>"000001111",
  4275=>"000100100",
  4276=>"101100101",
  4277=>"011100001",
  4278=>"010100000",
  4279=>"010011111",
  4280=>"100001000",
  4281=>"110100100",
  4282=>"110011001",
  4283=>"111101111",
  4284=>"111000010",
  4285=>"011111001",
  4286=>"001001100",
  4287=>"010101000",
  4288=>"001101101",
  4289=>"000000100",
  4290=>"000001110",
  4291=>"101000001",
  4292=>"111000101",
  4293=>"100010001",
  4294=>"101001101",
  4295=>"010011000",
  4296=>"001001111",
  4297=>"110111010",
  4298=>"000000010",
  4299=>"000001101",
  4300=>"111101000",
  4301=>"100000000",
  4302=>"000001000",
  4303=>"000101110",
  4304=>"110101100",
  4305=>"001000000",
  4306=>"010111101",
  4307=>"100100110",
  4308=>"011111101",
  4309=>"000111000",
  4310=>"000001101",
  4311=>"100101111",
  4312=>"101000000",
  4313=>"010010000",
  4314=>"100000000",
  4315=>"010000110",
  4316=>"001001011",
  4317=>"111010000",
  4318=>"001111000",
  4319=>"100101111",
  4320=>"110111100",
  4321=>"011011011",
  4322=>"010100101",
  4323=>"110110111",
  4324=>"111001110",
  4325=>"111101101",
  4326=>"000001011",
  4327=>"001011001",
  4328=>"010111111",
  4329=>"111111010",
  4330=>"001001001",
  4331=>"111111111",
  4332=>"010110011",
  4333=>"100110110",
  4334=>"000000001",
  4335=>"111001001",
  4336=>"001000010",
  4337=>"110101000",
  4338=>"010010111",
  4339=>"000001100",
  4340=>"100100001",
  4341=>"011111111",
  4342=>"001111000",
  4343=>"001111101",
  4344=>"000000000",
  4345=>"100111111",
  4346=>"111111011",
  4347=>"101000111",
  4348=>"101101101",
  4349=>"010000101",
  4350=>"001000000",
  4351=>"000010101",
  4352=>"011001010",
  4353=>"000000000",
  4354=>"001000101",
  4355=>"110000000",
  4356=>"111111111",
  4357=>"101101111",
  4358=>"110010010",
  4359=>"000110000",
  4360=>"111110000",
  4361=>"101001101",
  4362=>"100101100",
  4363=>"011011010",
  4364=>"000000111",
  4365=>"010111010",
  4366=>"111011001",
  4367=>"000111111",
  4368=>"111111011",
  4369=>"111001000",
  4370=>"000000111",
  4371=>"100000000",
  4372=>"101101111",
  4373=>"001111001",
  4374=>"001101101",
  4375=>"000111111",
  4376=>"101100110",
  4377=>"110000000",
  4378=>"111110001",
  4379=>"000000000",
  4380=>"000000110",
  4381=>"110110111",
  4382=>"111101000",
  4383=>"000000000",
  4384=>"111100000",
  4385=>"001111111",
  4386=>"110001000",
  4387=>"111000001",
  4388=>"011011000",
  4389=>"110100000",
  4390=>"101101111",
  4391=>"110000111",
  4392=>"000101000",
  4393=>"100110000",
  4394=>"000100111",
  4395=>"000001111",
  4396=>"111111111",
  4397=>"111100111",
  4398=>"111010000",
  4399=>"100100010",
  4400=>"101001100",
  4401=>"001111010",
  4402=>"001111110",
  4403=>"101001000",
  4404=>"010000111",
  4405=>"000001100",
  4406=>"000111111",
  4407=>"010110110",
  4408=>"000101000",
  4409=>"000000011",
  4410=>"110100000",
  4411=>"001000000",
  4412=>"100111100",
  4413=>"111000010",
  4414=>"110000000",
  4415=>"001000000",
  4416=>"101000110",
  4417=>"111001000",
  4418=>"111011000",
  4419=>"100100000",
  4420=>"000000011",
  4421=>"010000000",
  4422=>"111111001",
  4423=>"101011000",
  4424=>"011111111",
  4425=>"000000000",
  4426=>"000000010",
  4427=>"010111000",
  4428=>"111000000",
  4429=>"011011010",
  4430=>"100100100",
  4431=>"101101111",
  4432=>"111000000",
  4433=>"000010010",
  4434=>"111101000",
  4435=>"101001001",
  4436=>"000000111",
  4437=>"000011111",
  4438=>"110110100",
  4439=>"001000000",
  4440=>"000110100",
  4441=>"001000011",
  4442=>"100000111",
  4443=>"111111111",
  4444=>"111001101",
  4445=>"011011000",
  4446=>"010110111",
  4447=>"011001000",
  4448=>"111111000",
  4449=>"000000000",
  4450=>"101000000",
  4451=>"100110110",
  4452=>"101000000",
  4453=>"010111111",
  4454=>"000010000",
  4455=>"111000110",
  4456=>"000111111",
  4457=>"101111110",
  4458=>"010000111",
  4459=>"111000100",
  4460=>"000110110",
  4461=>"000000100",
  4462=>"000010111",
  4463=>"100111111",
  4464=>"100101000",
  4465=>"011111110",
  4466=>"011100111",
  4467=>"111111000",
  4468=>"111111111",
  4469=>"001000000",
  4470=>"010000101",
  4471=>"110000101",
  4472=>"100000110",
  4473=>"110000000",
  4474=>"001001111",
  4475=>"000000101",
  4476=>"100011001",
  4477=>"100100000",
  4478=>"000111111",
  4479=>"000000001",
  4480=>"101000001",
  4481=>"101010110",
  4482=>"000000111",
  4483=>"010000111",
  4484=>"111000000",
  4485=>"010100101",
  4486=>"001100110",
  4487=>"110000100",
  4488=>"001000000",
  4489=>"000001000",
  4490=>"101100101",
  4491=>"010000000",
  4492=>"000110100",
  4493=>"111111000",
  4494=>"001000101",
  4495=>"110000001",
  4496=>"110110000",
  4497=>"111111111",
  4498=>"000110000",
  4499=>"101101000",
  4500=>"110100000",
  4501=>"101001101",
  4502=>"111010000",
  4503=>"011011011",
  4504=>"001101000",
  4505=>"000011010",
  4506=>"000111010",
  4507=>"101100000",
  4508=>"101010010",
  4509=>"000000000",
  4510=>"111110111",
  4511=>"101100101",
  4512=>"000110111",
  4513=>"101001010",
  4514=>"000101110",
  4515=>"111000011",
  4516=>"001011111",
  4517=>"110001000",
  4518=>"111110110",
  4519=>"110110000",
  4520=>"110101111",
  4521=>"111110000",
  4522=>"001000000",
  4523=>"111000000",
  4524=>"111000000",
  4525=>"000000001",
  4526=>"100110100",
  4527=>"011000000",
  4528=>"000110110",
  4529=>"001011011",
  4530=>"000000000",
  4531=>"000000100",
  4532=>"110110000",
  4533=>"111111101",
  4534=>"010000000",
  4535=>"011011101",
  4536=>"011011000",
  4537=>"011001000",
  4538=>"111100010",
  4539=>"111111100",
  4540=>"000010010",
  4541=>"111111011",
  4542=>"110110000",
  4543=>"011111000",
  4544=>"100001111",
  4545=>"000101111",
  4546=>"101111110",
  4547=>"001011000",
  4548=>"000000111",
  4549=>"011000100",
  4550=>"010000000",
  4551=>"101001000",
  4552=>"111000000",
  4553=>"000000001",
  4554=>"011001101",
  4555=>"101001110",
  4556=>"100000000",
  4557=>"011110100",
  4558=>"000011111",
  4559=>"001000111",
  4560=>"000000111",
  4561=>"110110000",
  4562=>"111000000",
  4563=>"110010111",
  4564=>"010000000",
  4565=>"100110100",
  4566=>"111110100",
  4567=>"110000111",
  4568=>"000111111",
  4569=>"110000010",
  4570=>"100000101",
  4571=>"000000111",
  4572=>"101101111",
  4573=>"000110110",
  4574=>"111101110",
  4575=>"000110111",
  4576=>"000000001",
  4577=>"101000000",
  4578=>"000000111",
  4579=>"111111000",
  4580=>"100011011",
  4581=>"010110000",
  4582=>"010110110",
  4583=>"011111000",
  4584=>"000000111",
  4585=>"010011001",
  4586=>"001101001",
  4587=>"000010001",
  4588=>"110110011",
  4589=>"110000000",
  4590=>"000000000",
  4591=>"010100001",
  4592=>"000000000",
  4593=>"101001111",
  4594=>"010011000",
  4595=>"110100111",
  4596=>"110001010",
  4597=>"001000101",
  4598=>"010000000",
  4599=>"010001110",
  4600=>"000110111",
  4601=>"111111111",
  4602=>"001000111",
  4603=>"110011001",
  4604=>"111111001",
  4605=>"000000111",
  4606=>"100100000",
  4607=>"111000110",
  4608=>"000000000",
  4609=>"111111111",
  4610=>"010111101",
  4611=>"111111111",
  4612=>"000100111",
  4613=>"110000000",
  4614=>"101111110",
  4615=>"011111111",
  4616=>"011111010",
  4617=>"000001000",
  4618=>"110000000",
  4619=>"000000001",
  4620=>"011011000",
  4621=>"101101000",
  4622=>"000000000",
  4623=>"000000100",
  4624=>"111111111",
  4625=>"000001101",
  4626=>"000000110",
  4627=>"000000010",
  4628=>"000000000",
  4629=>"011110100",
  4630=>"111111111",
  4631=>"111111111",
  4632=>"000000111",
  4633=>"110101001",
  4634=>"000000000",
  4635=>"000111111",
  4636=>"000110010",
  4637=>"111111001",
  4638=>"110010011",
  4639=>"111111111",
  4640=>"000000000",
  4641=>"111011101",
  4642=>"000001000",
  4643=>"001010110",
  4644=>"000000111",
  4645=>"100101010",
  4646=>"011001001",
  4647=>"001100010",
  4648=>"010000101",
  4649=>"000000000",
  4650=>"101000100",
  4651=>"111111111",
  4652=>"110010011",
  4653=>"001000110",
  4654=>"001011111",
  4655=>"110111011",
  4656=>"000000000",
  4657=>"001011001",
  4658=>"000000000",
  4659=>"111100000",
  4660=>"000000000",
  4661=>"010111101",
  4662=>"111110100",
  4663=>"000000010",
  4664=>"000000000",
  4665=>"000000000",
  4666=>"010000000",
  4667=>"100111110",
  4668=>"000000001",
  4669=>"111111111",
  4670=>"010000000",
  4671=>"000000010",
  4672=>"000000100",
  4673=>"000111101",
  4674=>"110010000",
  4675=>"111111101",
  4676=>"000000000",
  4677=>"000000000",
  4678=>"101000100",
  4679=>"101001111",
  4680=>"000000000",
  4681=>"000001001",
  4682=>"000110000",
  4683=>"000100111",
  4684=>"000000100",
  4685=>"000000001",
  4686=>"110110010",
  4687=>"111111111",
  4688=>"010111111",
  4689=>"111111111",
  4690=>"000000111",
  4691=>"001001001",
  4692=>"111110000",
  4693=>"011000001",
  4694=>"100010110",
  4695=>"000000000",
  4696=>"111001101",
  4697=>"001100111",
  4698=>"011110010",
  4699=>"001011100",
  4700=>"000000000",
  4701=>"001000100",
  4702=>"001111111",
  4703=>"111110000",
  4704=>"000001011",
  4705=>"110000000",
  4706=>"000111000",
  4707=>"111111111",
  4708=>"000010010",
  4709=>"000000011",
  4710=>"100010000",
  4711=>"000000000",
  4712=>"010000000",
  4713=>"000000000",
  4714=>"000011011",
  4715=>"000000000",
  4716=>"000001000",
  4717=>"000000000",
  4718=>"110000000",
  4719=>"000110101",
  4720=>"000110011",
  4721=>"000010010",
  4722=>"111011011",
  4723=>"001000001",
  4724=>"000000000",
  4725=>"000000000",
  4726=>"101000000",
  4727=>"000000000",
  4728=>"111111111",
  4729=>"000100111",
  4730=>"000000000",
  4731=>"000001010",
  4732=>"010000011",
  4733=>"100100000",
  4734=>"111111110",
  4735=>"000000000",
  4736=>"101010110",
  4737=>"111011011",
  4738=>"000110010",
  4739=>"111110111",
  4740=>"001010111",
  4741=>"111111111",
  4742=>"000110100",
  4743=>"000000000",
  4744=>"001000000",
  4745=>"000111111",
  4746=>"000000000",
  4747=>"000000011",
  4748=>"111111111",
  4749=>"110111101",
  4750=>"000000110",
  4751=>"000000000",
  4752=>"110110110",
  4753=>"111001111",
  4754=>"000000110",
  4755=>"111111001",
  4756=>"000000000",
  4757=>"001000000",
  4758=>"101001001",
  4759=>"110000000",
  4760=>"010111011",
  4761=>"000010101",
  4762=>"010111010",
  4763=>"011111011",
  4764=>"000000000",
  4765=>"010010110",
  4766=>"000010000",
  4767=>"101111011",
  4768=>"111000001",
  4769=>"111110111",
  4770=>"111111000",
  4771=>"100111111",
  4772=>"010001101",
  4773=>"100010010",
  4774=>"111010011",
  4775=>"110101010",
  4776=>"111111111",
  4777=>"010001001",
  4778=>"111111111",
  4779=>"000000100",
  4780=>"111101111",
  4781=>"000000000",
  4782=>"110110100",
  4783=>"010001111",
  4784=>"111111101",
  4785=>"111001001",
  4786=>"000100010",
  4787=>"000000011",
  4788=>"011111000",
  4789=>"000010111",
  4790=>"001011111",
  4791=>"100101111",
  4792=>"000000110",
  4793=>"011000001",
  4794=>"000000010",
  4795=>"010000111",
  4796=>"100100000",
  4797=>"101101111",
  4798=>"000011000",
  4799=>"111101011",
  4800=>"110111110",
  4801=>"000000011",
  4802=>"000000000",
  4803=>"001011001",
  4804=>"000000000",
  4805=>"001001000",
  4806=>"000000100",
  4807=>"000000011",
  4808=>"111000000",
  4809=>"001001110",
  4810=>"000000000",
  4811=>"010110001",
  4812=>"110101011",
  4813=>"110110110",
  4814=>"111011111",
  4815=>"001101111",
  4816=>"100111100",
  4817=>"111011100",
  4818=>"000000000",
  4819=>"000000001",
  4820=>"111111111",
  4821=>"110110111",
  4822=>"000010100",
  4823=>"000011000",
  4824=>"111111110",
  4825=>"000001011",
  4826=>"011001111",
  4827=>"011001001",
  4828=>"110110111",
  4829=>"111001001",
  4830=>"010000001",
  4831=>"000000000",
  4832=>"010101000",
  4833=>"101000011",
  4834=>"111110111",
  4835=>"000110111",
  4836=>"000101000",
  4837=>"110000111",
  4838=>"001000000",
  4839=>"110110111",
  4840=>"000000011",
  4841=>"001001000",
  4842=>"001001001",
  4843=>"001000001",
  4844=>"000000000",
  4845=>"111111111",
  4846=>"101110000",
  4847=>"010111010",
  4848=>"111101100",
  4849=>"000000000",
  4850=>"101000011",
  4851=>"100111010",
  4852=>"000001010",
  4853=>"111111111",
  4854=>"000000000",
  4855=>"111111111",
  4856=>"010110000",
  4857=>"100111111",
  4858=>"011111111",
  4859=>"010010000",
  4860=>"000000000",
  4861=>"010110000",
  4862=>"000010110",
  4863=>"000110111",
  4864=>"111001111",
  4865=>"000000011",
  4866=>"000101111",
  4867=>"001010000",
  4868=>"111111111",
  4869=>"000000101",
  4870=>"000100000",
  4871=>"011000100",
  4872=>"000110111",
  4873=>"001111111",
  4874=>"111101101",
  4875=>"110001000",
  4876=>"000000111",
  4877=>"000100000",
  4878=>"111001011",
  4879=>"111000111",
  4880=>"011000100",
  4881=>"100101101",
  4882=>"000000000",
  4883=>"000001000",
  4884=>"011010001",
  4885=>"000000110",
  4886=>"001001011",
  4887=>"111111000",
  4888=>"101000000",
  4889=>"111001010",
  4890=>"011011011",
  4891=>"000111111",
  4892=>"000101000",
  4893=>"111000001",
  4894=>"000000001",
  4895=>"111000000",
  4896=>"111111010",
  4897=>"111011000",
  4898=>"011011000",
  4899=>"000010110",
  4900=>"100000001",
  4901=>"110100000",
  4902=>"111100000",
  4903=>"010111010",
  4904=>"111000000",
  4905=>"010000110",
  4906=>"111101000",
  4907=>"000100001",
  4908=>"001001001",
  4909=>"101000000",
  4910=>"110000000",
  4911=>"001111011",
  4912=>"000000110",
  4913=>"011100100",
  4914=>"000000111",
  4915=>"111100000",
  4916=>"111111110",
  4917=>"111011111",
  4918=>"100111111",
  4919=>"101111111",
  4920=>"100001101",
  4921=>"000101111",
  4922=>"000111000",
  4923=>"111010010",
  4924=>"000000000",
  4925=>"111011000",
  4926=>"000000000",
  4927=>"110011000",
  4928=>"000100010",
  4929=>"010000101",
  4930=>"110000100",
  4931=>"000100111",
  4932=>"000000000",
  4933=>"111000001",
  4934=>"000110000",
  4935=>"101100111",
  4936=>"110100001",
  4937=>"000000000",
  4938=>"000111111",
  4939=>"111000000",
  4940=>"000000000",
  4941=>"100110110",
  4942=>"111111001",
  4943=>"111010000",
  4944=>"101101111",
  4945=>"000011011",
  4946=>"001001111",
  4947=>"011010000",
  4948=>"000000000",
  4949=>"010110111",
  4950=>"111001000",
  4951=>"000000001",
  4952=>"000100000",
  4953=>"011010000",
  4954=>"110100100",
  4955=>"111010000",
  4956=>"000000000",
  4957=>"001000000",
  4958=>"100110111",
  4959=>"110001111",
  4960=>"000111111",
  4961=>"000000011",
  4962=>"100111111",
  4963=>"101001001",
  4964=>"010100100",
  4965=>"111100001",
  4966=>"101000000",
  4967=>"111010001",
  4968=>"111111000",
  4969=>"111010000",
  4970=>"010110111",
  4971=>"010000111",
  4972=>"111110010",
  4973=>"111011001",
  4974=>"001010000",
  4975=>"011000000",
  4976=>"100100101",
  4977=>"111000000",
  4978=>"001110011",
  4979=>"101000011",
  4980=>"010000000",
  4981=>"000000000",
  4982=>"000000000",
  4983=>"111011111",
  4984=>"000111000",
  4985=>"111111111",
  4986=>"101111111",
  4987=>"101111111",
  4988=>"110010010",
  4989=>"010001000",
  4990=>"010010000",
  4991=>"100100111",
  4992=>"011000000",
  4993=>"111000111",
  4994=>"000000000",
  4995=>"111111111",
  4996=>"010101100",
  4997=>"011001101",
  4998=>"001001100",
  4999=>"011010100",
  5000=>"001001111",
  5001=>"001001101",
  5002=>"111110001",
  5003=>"010011111",
  5004=>"000000000",
  5005=>"111111011",
  5006=>"000111111",
  5007=>"110111111",
  5008=>"111100001",
  5009=>"101000000",
  5010=>"010000000",
  5011=>"010101111",
  5012=>"011010010",
  5013=>"010010101",
  5014=>"101101111",
  5015=>"011001011",
  5016=>"011011000",
  5017=>"011010101",
  5018=>"000000111",
  5019=>"111111000",
  5020=>"000000000",
  5021=>"000000110",
  5022=>"000000101",
  5023=>"000001111",
  5024=>"001101001",
  5025=>"000000000",
  5026=>"000000101",
  5027=>"100111110",
  5028=>"110101011",
  5029=>"110001000",
  5030=>"111000000",
  5031=>"011111000",
  5032=>"000011111",
  5033=>"010110010",
  5034=>"100001101",
  5035=>"000100011",
  5036=>"111111111",
  5037=>"000111010",
  5038=>"000000001",
  5039=>"011000111",
  5040=>"111011111",
  5041=>"000001001",
  5042=>"111111000",
  5043=>"010000001",
  5044=>"011000100",
  5045=>"000011100",
  5046=>"010001010",
  5047=>"111000000",
  5048=>"000000001",
  5049=>"110110000",
  5050=>"011000000",
  5051=>"000111111",
  5052=>"011000000",
  5053=>"000000111",
  5054=>"001011011",
  5055=>"000000000",
  5056=>"011000000",
  5057=>"111000000",
  5058=>"000100100",
  5059=>"111110110",
  5060=>"000011000",
  5061=>"011001011",
  5062=>"011011000",
  5063=>"101111111",
  5064=>"010000000",
  5065=>"000001111",
  5066=>"000111110",
  5067=>"111111111",
  5068=>"010000000",
  5069=>"011110010",
  5070=>"110101001",
  5071=>"011000000",
  5072=>"011000000",
  5073=>"011101111",
  5074=>"111010000",
  5075=>"011111000",
  5076=>"010000000",
  5077=>"100100110",
  5078=>"001001111",
  5079=>"011010000",
  5080=>"111000000",
  5081=>"111101100",
  5082=>"110110100",
  5083=>"000111111",
  5084=>"000000110",
  5085=>"001000111",
  5086=>"111100000",
  5087=>"111011010",
  5088=>"111011000",
  5089=>"000100111",
  5090=>"111010001",
  5091=>"110101111",
  5092=>"010000000",
  5093=>"001000111",
  5094=>"000101111",
  5095=>"000011011",
  5096=>"000100111",
  5097=>"100111111",
  5098=>"101001001",
  5099=>"000000011",
  5100=>"000111111",
  5101=>"000000111",
  5102=>"000000000",
  5103=>"000000000",
  5104=>"000000000",
  5105=>"111000101",
  5106=>"011111111",
  5107=>"110100000",
  5108=>"000000100",
  5109=>"000001001",
  5110=>"100001010",
  5111=>"111010000",
  5112=>"111111001",
  5113=>"111001000",
  5114=>"001001111",
  5115=>"111010001",
  5116=>"011111010",
  5117=>"111111100",
  5118=>"000101111",
  5119=>"100000001",
  5120=>"000000000",
  5121=>"001100000",
  5122=>"111011000",
  5123=>"011100110",
  5124=>"001011011",
  5125=>"000000011",
  5126=>"111111000",
  5127=>"011111111",
  5128=>"101101111",
  5129=>"000101100",
  5130=>"001001111",
  5131=>"111000010",
  5132=>"111010000",
  5133=>"010000001",
  5134=>"001011001",
  5135=>"001111111",
  5136=>"111111111",
  5137=>"010000001",
  5138=>"000000001",
  5139=>"101110000",
  5140=>"000111011",
  5141=>"000100110",
  5142=>"010001000",
  5143=>"000001000",
  5144=>"111100000",
  5145=>"000000000",
  5146=>"101111000",
  5147=>"111000000",
  5148=>"000000100",
  5149=>"101111111",
  5150=>"001000000",
  5151=>"111111010",
  5152=>"000100111",
  5153=>"111100111",
  5154=>"100111111",
  5155=>"000111010",
  5156=>"001101000",
  5157=>"000000001",
  5158=>"110000111",
  5159=>"110000000",
  5160=>"010111101",
  5161=>"001111110",
  5162=>"100000000",
  5163=>"101000001",
  5164=>"011001000",
  5165=>"111101011",
  5166=>"000000001",
  5167=>"000000111",
  5168=>"000000010",
  5169=>"011101111",
  5170=>"000011111",
  5171=>"000000000",
  5172=>"010010000",
  5173=>"000010010",
  5174=>"110110100",
  5175=>"000111111",
  5176=>"000000000",
  5177=>"000000000",
  5178=>"010110111",
  5179=>"001101100",
  5180=>"110001101",
  5181=>"111111111",
  5182=>"111000000",
  5183=>"100111110",
  5184=>"111101000",
  5185=>"111011011",
  5186=>"100111011",
  5187=>"000100110",
  5188=>"111100100",
  5189=>"010011010",
  5190=>"101111110",
  5191=>"011000011",
  5192=>"111111111",
  5193=>"111110000",
  5194=>"111011111",
  5195=>"101100010",
  5196=>"000001001",
  5197=>"011001001",
  5198=>"100110110",
  5199=>"111111011",
  5200=>"111000000",
  5201=>"000100111",
  5202=>"000000000",
  5203=>"101100000",
  5204=>"011000000",
  5205=>"011001111",
  5206=>"011101100",
  5207=>"011010000",
  5208=>"010000000",
  5209=>"001000010",
  5210=>"110110000",
  5211=>"100100100",
  5212=>"001000000",
  5213=>"001001011",
  5214=>"000011000",
  5215=>"011001011",
  5216=>"000111000",
  5217=>"111110000",
  5218=>"111010000",
  5219=>"011011111",
  5220=>"100100000",
  5221=>"000001111",
  5222=>"110111111",
  5223=>"000111111",
  5224=>"000000000",
  5225=>"010000101",
  5226=>"110111111",
  5227=>"000101111",
  5228=>"101100100",
  5229=>"000010111",
  5230=>"100111000",
  5231=>"000000111",
  5232=>"100111011",
  5233=>"000000110",
  5234=>"001010001",
  5235=>"000010000",
  5236=>"000101111",
  5237=>"000000000",
  5238=>"110000000",
  5239=>"111111111",
  5240=>"011011111",
  5241=>"101100000",
  5242=>"101000000",
  5243=>"000001001",
  5244=>"110100001",
  5245=>"100001000",
  5246=>"000111010",
  5247=>"111010000",
  5248=>"000000000",
  5249=>"000000010",
  5250=>"111111111",
  5251=>"111101111",
  5252=>"101101001",
  5253=>"000000000",
  5254=>"001001011",
  5255=>"111011000",
  5256=>"001001110",
  5257=>"000100100",
  5258=>"000110011",
  5259=>"010000000",
  5260=>"000000000",
  5261=>"000000000",
  5262=>"101100100",
  5263=>"000010000",
  5264=>"100110101",
  5265=>"010000000",
  5266=>"010111010",
  5267=>"011000100",
  5268=>"100001000",
  5269=>"000001111",
  5270=>"110101111",
  5271=>"000001011",
  5272=>"110000111",
  5273=>"010000111",
  5274=>"010111111",
  5275=>"000001111",
  5276=>"000001010",
  5277=>"000000111",
  5278=>"000100111",
  5279=>"111000000",
  5280=>"110111101",
  5281=>"000000111",
  5282=>"111000000",
  5283=>"111111111",
  5284=>"000000111",
  5285=>"011011000",
  5286=>"100110110",
  5287=>"100101111",
  5288=>"001000000",
  5289=>"001101111",
  5290=>"110110111",
  5291=>"111110001",
  5292=>"000000000",
  5293=>"111111000",
  5294=>"000001001",
  5295=>"111111001",
  5296=>"000000000",
  5297=>"001000001",
  5298=>"000000111",
  5299=>"110110100",
  5300=>"110100001",
  5301=>"000000000",
  5302=>"010010000",
  5303=>"000000000",
  5304=>"001000101",
  5305=>"011001000",
  5306=>"011010111",
  5307=>"000111111",
  5308=>"000010110",
  5309=>"000000111",
  5310=>"001011011",
  5311=>"000010111",
  5312=>"101000000",
  5313=>"101101001",
  5314=>"000111011",
  5315=>"101100000",
  5316=>"000000101",
  5317=>"000001001",
  5318=>"001111111",
  5319=>"010001111",
  5320=>"101111010",
  5321=>"111111000",
  5322=>"000000000",
  5323=>"101111010",
  5324=>"000000011",
  5325=>"001100100",
  5326=>"000000000",
  5327=>"001111100",
  5328=>"111111010",
  5329=>"101100110",
  5330=>"111111000",
  5331=>"000001000",
  5332=>"111011000",
  5333=>"000000101",
  5334=>"011010111",
  5335=>"000111111",
  5336=>"000000000",
  5337=>"100111111",
  5338=>"001101101",
  5339=>"011000000",
  5340=>"110100001",
  5341=>"110111111",
  5342=>"010010000",
  5343=>"000000001",
  5344=>"111111010",
  5345=>"000000101",
  5346=>"111011000",
  5347=>"100100100",
  5348=>"100000111",
  5349=>"111010110",
  5350=>"111111001",
  5351=>"101001111",
  5352=>"111000111",
  5353=>"010001000",
  5354=>"100100111",
  5355=>"011111111",
  5356=>"101110000",
  5357=>"000010000",
  5358=>"110000000",
  5359=>"010000011",
  5360=>"010000010",
  5361=>"001101100",
  5362=>"101100011",
  5363=>"100001001",
  5364=>"111101000",
  5365=>"100000000",
  5366=>"010010111",
  5367=>"000000101",
  5368=>"111010111",
  5369=>"000111111",
  5370=>"101111111",
  5371=>"111100000",
  5372=>"000101011",
  5373=>"111010000",
  5374=>"110100101",
  5375=>"000110011",
  5376=>"110000000",
  5377=>"000000000",
  5378=>"111001111",
  5379=>"001000011",
  5380=>"101111011",
  5381=>"110110000",
  5382=>"000111111",
  5383=>"000010111",
  5384=>"101001000",
  5385=>"000000111",
  5386=>"001100110",
  5387=>"110110100",
  5388=>"111010000",
  5389=>"110110000",
  5390=>"110000011",
  5391=>"000001101",
  5392=>"101111111",
  5393=>"000000111",
  5394=>"111010010",
  5395=>"000000111",
  5396=>"001111111",
  5397=>"110000111",
  5398=>"000110000",
  5399=>"000000010",
  5400=>"111001001",
  5401=>"000101111",
  5402=>"000011010",
  5403=>"111000110",
  5404=>"000000100",
  5405=>"001111001",
  5406=>"000011111",
  5407=>"101001001",
  5408=>"111000010",
  5409=>"111110000",
  5410=>"110110011",
  5411=>"110000000",
  5412=>"110111001",
  5413=>"000000000",
  5414=>"101000000",
  5415=>"110000001",
  5416=>"111001000",
  5417=>"110110101",
  5418=>"000101101",
  5419=>"011111000",
  5420=>"000111111",
  5421=>"001111010",
  5422=>"000110111",
  5423=>"000111000",
  5424=>"000111111",
  5425=>"111011000",
  5426=>"111110100",
  5427=>"000111111",
  5428=>"000101111",
  5429=>"100000111",
  5430=>"000001011",
  5431=>"000000000",
  5432=>"000111000",
  5433=>"000001111",
  5434=>"000000001",
  5435=>"000000000",
  5436=>"011001000",
  5437=>"001000101",
  5438=>"100000001",
  5439=>"011011001",
  5440=>"101110111",
  5441=>"110011010",
  5442=>"000000000",
  5443=>"011100110",
  5444=>"110110000",
  5445=>"000000001",
  5446=>"000001110",
  5447=>"101001101",
  5448=>"011000010",
  5449=>"000111111",
  5450=>"000111111",
  5451=>"000101001",
  5452=>"011000000",
  5453=>"110110000",
  5454=>"110110100",
  5455=>"100110111",
  5456=>"101001000",
  5457=>"111111010",
  5458=>"000111111",
  5459=>"101101100",
  5460=>"000101111",
  5461=>"000110100",
  5462=>"011011001",
  5463=>"000101111",
  5464=>"010101001",
  5465=>"011001000",
  5466=>"000100000",
  5467=>"011100100",
  5468=>"000001011",
  5469=>"010001001",
  5470=>"101111010",
  5471=>"100011010",
  5472=>"111100000",
  5473=>"011110111",
  5474=>"111001000",
  5475=>"000001011",
  5476=>"100100000",
  5477=>"000000011",
  5478=>"000000111",
  5479=>"001111110",
  5480=>"110000001",
  5481=>"000000111",
  5482=>"111110000",
  5483=>"000001111",
  5484=>"100111100",
  5485=>"000001111",
  5486=>"000000001",
  5487=>"000000000",
  5488=>"110110000",
  5489=>"010110100",
  5490=>"000100110",
  5491=>"000010111",
  5492=>"111111111",
  5493=>"000000101",
  5494=>"100000000",
  5495=>"110110011",
  5496=>"001000111",
  5497=>"000000110",
  5498=>"111010001",
  5499=>"111111000",
  5500=>"111110110",
  5501=>"000011000",
  5502=>"001000000",
  5503=>"010000000",
  5504=>"100100110",
  5505=>"101000000",
  5506=>"000010010",
  5507=>"101111111",
  5508=>"001111111",
  5509=>"001000000",
  5510=>"000000101",
  5511=>"101100011",
  5512=>"011000000",
  5513=>"010110111",
  5514=>"000110111",
  5515=>"001001111",
  5516=>"110000000",
  5517=>"100000001",
  5518=>"000110111",
  5519=>"000001111",
  5520=>"000100001",
  5521=>"100101100",
  5522=>"010000000",
  5523=>"001001111",
  5524=>"100111111",
  5525=>"001111000",
  5526=>"101000101",
  5527=>"111111100",
  5528=>"101101111",
  5529=>"001001100",
  5530=>"011000000",
  5531=>"001001010",
  5532=>"000111110",
  5533=>"111100000",
  5534=>"000111111",
  5535=>"000111100",
  5536=>"011011000",
  5537=>"000111111",
  5538=>"111010000",
  5539=>"001111111",
  5540=>"000000010",
  5541=>"110111111",
  5542=>"000001111",
  5543=>"101111111",
  5544=>"000111111",
  5545=>"110110100",
  5546=>"111010000",
  5547=>"111111000",
  5548=>"111011000",
  5549=>"110000000",
  5550=>"011001001",
  5551=>"010001111",
  5552=>"111111001",
  5553=>"111110110",
  5554=>"001111000",
  5555=>"111010000",
  5556=>"001001101",
  5557=>"001111111",
  5558=>"111111010",
  5559=>"000010100",
  5560=>"100000000",
  5561=>"101111111",
  5562=>"000110111",
  5563=>"000111111",
  5564=>"000001110",
  5565=>"111111101",
  5566=>"111100000",
  5567=>"000011111",
  5568=>"001001111",
  5569=>"111101111",
  5570=>"011000111",
  5571=>"000001000",
  5572=>"110000000",
  5573=>"111110111",
  5574=>"000101011",
  5575=>"111000000",
  5576=>"110101110",
  5577=>"111110000",
  5578=>"111110000",
  5579=>"110100011",
  5580=>"000101101",
  5581=>"111100001",
  5582=>"100111101",
  5583=>"111111011",
  5584=>"000011101",
  5585=>"110111001",
  5586=>"000000100",
  5587=>"110000101",
  5588=>"111001111",
  5589=>"000010000",
  5590=>"111111000",
  5591=>"001111111",
  5592=>"000001111",
  5593=>"000000000",
  5594=>"110100001",
  5595=>"000000111",
  5596=>"001111101",
  5597=>"001111000",
  5598=>"000101101",
  5599=>"010100111",
  5600=>"000000110",
  5601=>"110111111",
  5602=>"000000001",
  5603=>"111010000",
  5604=>"000000010",
  5605=>"001111110",
  5606=>"111111000",
  5607=>"000000001",
  5608=>"111000000",
  5609=>"000000001",
  5610=>"000001011",
  5611=>"100000001",
  5612=>"110110000",
  5613=>"111111100",
  5614=>"110000000",
  5615=>"110110000",
  5616=>"010000001",
  5617=>"100111011",
  5618=>"000010001",
  5619=>"110011011",
  5620=>"011000000",
  5621=>"000011111",
  5622=>"000000111",
  5623=>"111111000",
  5624=>"111111000",
  5625=>"111111000",
  5626=>"000110110",
  5627=>"000011111",
  5628=>"000101111",
  5629=>"000110000",
  5630=>"011100100",
  5631=>"000101111",
  5632=>"101000000",
  5633=>"010010011",
  5634=>"100001000",
  5635=>"110111111",
  5636=>"000000000",
  5637=>"100100101",
  5638=>"011011011",
  5639=>"001001001",
  5640=>"001100110",
  5641=>"000100000",
  5642=>"001100000",
  5643=>"001000001",
  5644=>"100110110",
  5645=>"110100100",
  5646=>"100100000",
  5647=>"000111101",
  5648=>"111001100",
  5649=>"011011001",
  5650=>"100011001",
  5651=>"011011011",
  5652=>"100100000",
  5653=>"001001011",
  5654=>"011101001",
  5655=>"000110111",
  5656=>"001100000",
  5657=>"111011110",
  5658=>"011011011",
  5659=>"001000000",
  5660=>"011110110",
  5661=>"100100110",
  5662=>"011010000",
  5663=>"110010010",
  5664=>"100101100",
  5665=>"000011111",
  5666=>"100000011",
  5667=>"100100011",
  5668=>"111111111",
  5669=>"011101101",
  5670=>"011011011",
  5671=>"100111111",
  5672=>"010000110",
  5673=>"110111101",
  5674=>"011111001",
  5675=>"111001011",
  5676=>"000001100",
  5677=>"111101011",
  5678=>"001100000",
  5679=>"000100010",
  5680=>"100001110",
  5681=>"000000000",
  5682=>"100001101",
  5683=>"100000001",
  5684=>"000000000",
  5685=>"011001001",
  5686=>"011011001",
  5687=>"001001001",
  5688=>"001001111",
  5689=>"010100101",
  5690=>"100100100",
  5691=>"000100010",
  5692=>"010100100",
  5693=>"100110110",
  5694=>"010000100",
  5695=>"000111001",
  5696=>"001001111",
  5697=>"011110100",
  5698=>"101111001",
  5699=>"010001000",
  5700=>"010110110",
  5701=>"000000000",
  5702=>"001011001",
  5703=>"111101010",
  5704=>"100101110",
  5705=>"010010110",
  5706=>"000000000",
  5707=>"001000000",
  5708=>"011011001",
  5709=>"000000000",
  5710=>"111111111",
  5711=>"100100011",
  5712=>"011011010",
  5713=>"011100110",
  5714=>"000000000",
  5715=>"000000010",
  5716=>"001000010",
  5717=>"111101110",
  5718=>"111110110",
  5719=>"101001100",
  5720=>"111110110",
  5721=>"001001000",
  5722=>"101001101",
  5723=>"100001011",
  5724=>"100100100",
  5725=>"000000000",
  5726=>"111011101",
  5727=>"001011011",
  5728=>"000011000",
  5729=>"010110010",
  5730=>"100001100",
  5731=>"001111111",
  5732=>"110110110",
  5733=>"101111111",
  5734=>"100000010",
  5735=>"100000100",
  5736=>"100111011",
  5737=>"111100100",
  5738=>"011001001",
  5739=>"000011111",
  5740=>"110100110",
  5741=>"100100100",
  5742=>"001100111",
  5743=>"001100100",
  5744=>"000000000",
  5745=>"000000101",
  5746=>"011001010",
  5747=>"111011001",
  5748=>"011000011",
  5749=>"001000000",
  5750=>"001011011",
  5751=>"011011001",
  5752=>"100011001",
  5753=>"110110110",
  5754=>"001011001",
  5755=>"100100110",
  5756=>"111000100",
  5757=>"111100100",
  5758=>"110001100",
  5759=>"000000110",
  5760=>"100000100",
  5761=>"100110000",
  5762=>"001000000",
  5763=>"100100100",
  5764=>"010000000",
  5765=>"000001110",
  5766=>"001000000",
  5767=>"001001000",
  5768=>"111111111",
  5769=>"011010110",
  5770=>"111110110",
  5771=>"001001100",
  5772=>"000001100",
  5773=>"001001101",
  5774=>"010000001",
  5775=>"101000100",
  5776=>"111110011",
  5777=>"010000011",
  5778=>"000000000",
  5779=>"011010011",
  5780=>"011011000",
  5781=>"000001000",
  5782=>"111111111",
  5783=>"001000011",
  5784=>"001000000",
  5785=>"000010010",
  5786=>"011100110",
  5787=>"100100010",
  5788=>"000001010",
  5789=>"011101100",
  5790=>"001111011",
  5791=>"001001001",
  5792=>"100000100",
  5793=>"110100111",
  5794=>"100011111",
  5795=>"111100100",
  5796=>"011111100",
  5797=>"000000100",
  5798=>"000011011",
  5799=>"000100010",
  5800=>"001001001",
  5801=>"010010011",
  5802=>"110100100",
  5803=>"011010001",
  5804=>"000101010",
  5805=>"011011000",
  5806=>"110100101",
  5807=>"000001001",
  5808=>"110101110",
  5809=>"101100100",
  5810=>"100100110",
  5811=>"100000100",
  5812=>"111100111",
  5813=>"000000001",
  5814=>"111110100",
  5815=>"000011101",
  5816=>"100011011",
  5817=>"000000000",
  5818=>"011000001",
  5819=>"101000001",
  5820=>"100011100",
  5821=>"111011111",
  5822=>"000001000",
  5823=>"100011011",
  5824=>"001000001",
  5825=>"011011001",
  5826=>"001001011",
  5827=>"000111101",
  5828=>"000100100",
  5829=>"111100111",
  5830=>"000110110",
  5831=>"111101100",
  5832=>"101100100",
  5833=>"011011010",
  5834=>"100110110",
  5835=>"001001001",
  5836=>"011001010",
  5837=>"011010011",
  5838=>"001000100",
  5839=>"001110000",
  5840=>"011011011",
  5841=>"111101111",
  5842=>"011011010",
  5843=>"001011011",
  5844=>"011011011",
  5845=>"000100100",
  5846=>"000000000",
  5847=>"100000000",
  5848=>"110111011",
  5849=>"110011011",
  5850=>"101101111",
  5851=>"101100100",
  5852=>"111100110",
  5853=>"100110010",
  5854=>"011000010",
  5855=>"111001000",
  5856=>"001000010",
  5857=>"100001101",
  5858=>"001011001",
  5859=>"100110111",
  5860=>"100000010",
  5861=>"000100110",
  5862=>"001011011",
  5863=>"100000100",
  5864=>"000011001",
  5865=>"100001011",
  5866=>"111000000",
  5867=>"100110100",
  5868=>"001011010",
  5869=>"000001111",
  5870=>"000100000",
  5871=>"000100110",
  5872=>"010110110",
  5873=>"000100101",
  5874=>"011111000",
  5875=>"100110100",
  5876=>"111111101",
  5877=>"101000001",
  5878=>"000001011",
  5879=>"011011011",
  5880=>"000000111",
  5881=>"000111011",
  5882=>"110100100",
  5883=>"101000010",
  5884=>"001001000",
  5885=>"110100110",
  5886=>"111111101",
  5887=>"011111001",
  5888=>"111011001",
  5889=>"011100000",
  5890=>"001110100",
  5891=>"010101000",
  5892=>"111111110",
  5893=>"111111110",
  5894=>"000111000",
  5895=>"011101000",
  5896=>"110000000",
  5897=>"000000011",
  5898=>"001010011",
  5899=>"101111011",
  5900=>"100100000",
  5901=>"101110011",
  5902=>"011001011",
  5903=>"111100010",
  5904=>"000011101",
  5905=>"000000110",
  5906=>"111000000",
  5907=>"000000011",
  5908=>"001100000",
  5909=>"011100100",
  5910=>"111001100",
  5911=>"000100101",
  5912=>"001110000",
  5913=>"010000111",
  5914=>"110010001",
  5915=>"011011000",
  5916=>"111111111",
  5917=>"100000000",
  5918=>"001000101",
  5919=>"101101011",
  5920=>"111000000",
  5921=>"000001101",
  5922=>"000111000",
  5923=>"111101000",
  5924=>"100100100",
  5925=>"110111111",
  5926=>"000000000",
  5927=>"000100010",
  5928=>"010111111",
  5929=>"110111111",
  5930=>"000000010",
  5931=>"111010010",
  5932=>"111101011",
  5933=>"000000101",
  5934=>"001101011",
  5935=>"001001000",
  5936=>"000011101",
  5937=>"111101111",
  5938=>"000000000",
  5939=>"000010100",
  5940=>"101111010",
  5941=>"011000000",
  5942=>"110100100",
  5943=>"111100000",
  5944=>"010111000",
  5945=>"010110010",
  5946=>"111100000",
  5947=>"010110100",
  5948=>"100000010",
  5949=>"011101101",
  5950=>"000000000",
  5951=>"111111110",
  5952=>"000000000",
  5953=>"111111111",
  5954=>"100100110",
  5955=>"110110001",
  5956=>"111111100",
  5957=>"111001110",
  5958=>"100000000",
  5959=>"110100001",
  5960=>"000111001",
  5961=>"010011000",
  5962=>"010000000",
  5963=>"001111101",
  5964=>"000111111",
  5965=>"100111011",
  5966=>"110110110",
  5967=>"111111001",
  5968=>"001001010",
  5969=>"001010111",
  5970=>"111110010",
  5971=>"001001001",
  5972=>"111000000",
  5973=>"000000010",
  5974=>"000101011",
  5975=>"011001111",
  5976=>"100000001",
  5977=>"111101111",
  5978=>"111110111",
  5979=>"000011111",
  5980=>"100010010",
  5981=>"001001001",
  5982=>"010010111",
  5983=>"001011000",
  5984=>"110000000",
  5985=>"000000000",
  5986=>"111111111",
  5987=>"100101001",
  5988=>"100111111",
  5989=>"001011001",
  5990=>"110010010",
  5991=>"000000000",
  5992=>"110000000",
  5993=>"010010010",
  5994=>"000110011",
  5995=>"111111000",
  5996=>"000111111",
  5997=>"000011100",
  5998=>"100001000",
  5999=>"111111010",
  6000=>"111101001",
  6001=>"111111000",
  6002=>"001000100",
  6003=>"000101111",
  6004=>"000101111",
  6005=>"101000000",
  6006=>"000000000",
  6007=>"111110110",
  6008=>"011000000",
  6009=>"011010111",
  6010=>"101000000",
  6011=>"010000000",
  6012=>"110000000",
  6013=>"100100100",
  6014=>"010010111",
  6015=>"000110000",
  6016=>"011111100",
  6017=>"010001111",
  6018=>"001111111",
  6019=>"010111010",
  6020=>"000000110",
  6021=>"110110000",
  6022=>"011111111",
  6023=>"000001010",
  6024=>"100100100",
  6025=>"010110010",
  6026=>"010011101",
  6027=>"111000100",
  6028=>"000000010",
  6029=>"001111010",
  6030=>"000101101",
  6031=>"000001000",
  6032=>"100101100",
  6033=>"111111111",
  6034=>"010011001",
  6035=>"111000000",
  6036=>"000000000",
  6037=>"000000000",
  6038=>"111111100",
  6039=>"001011010",
  6040=>"101111011",
  6041=>"000101111",
  6042=>"111101101",
  6043=>"000100100",
  6044=>"110111101",
  6045=>"111101101",
  6046=>"010011001",
  6047=>"111001101",
  6048=>"111010101",
  6049=>"000100000",
  6050=>"010000000",
  6051=>"011101000",
  6052=>"111110100",
  6053=>"000000010",
  6054=>"100100001",
  6055=>"111111010",
  6056=>"000000111",
  6057=>"000000000",
  6058=>"000100100",
  6059=>"111010111",
  6060=>"000110011",
  6061=>"100000100",
  6062=>"110010001",
  6063=>"111000011",
  6064=>"111111111",
  6065=>"001001001",
  6066=>"000111111",
  6067=>"100100110",
  6068=>"000100100",
  6069=>"111111010",
  6070=>"000000011",
  6071=>"111010110",
  6072=>"001000000",
  6073=>"000000000",
  6074=>"111001010",
  6075=>"111101111",
  6076=>"110101011",
  6077=>"111111110",
  6078=>"001000000",
  6079=>"000110010",
  6080=>"001101000",
  6081=>"000010111",
  6082=>"000000111",
  6083=>"011111001",
  6084=>"000010000",
  6085=>"000001000",
  6086=>"010000010",
  6087=>"010110000",
  6088=>"000101111",
  6089=>"001000111",
  6090=>"011111011",
  6091=>"111001101",
  6092=>"000000001",
  6093=>"011000000",
  6094=>"000000000",
  6095=>"101100000",
  6096=>"000010010",
  6097=>"100111101",
  6098=>"100000000",
  6099=>"111111110",
  6100=>"110101000",
  6101=>"100100000",
  6102=>"111000000",
  6103=>"110110010",
  6104=>"101100000",
  6105=>"100000000",
  6106=>"010110101",
  6107=>"000000010",
  6108=>"001000000",
  6109=>"111101000",
  6110=>"000101100",
  6111=>"000001000",
  6112=>"000000011",
  6113=>"000000000",
  6114=>"000000000",
  6115=>"011101010",
  6116=>"010000111",
  6117=>"111111101",
  6118=>"010011101",
  6119=>"110011000",
  6120=>"000010110",
  6121=>"000000000",
  6122=>"110110111",
  6123=>"111111110",
  6124=>"000000000",
  6125=>"111110010",
  6126=>"001000100",
  6127=>"010010111",
  6128=>"100110001",
  6129=>"000000000",
  6130=>"111110010",
  6131=>"000001011",
  6132=>"110110110",
  6133=>"000111111",
  6134=>"000000010",
  6135=>"101000111",
  6136=>"000000000",
  6137=>"000001000",
  6138=>"001001111",
  6139=>"000000000",
  6140=>"110101011",
  6141=>"111111101",
  6142=>"011111000",
  6143=>"000100100",
  6144=>"101110111",
  6145=>"110011110",
  6146=>"100100100",
  6147=>"000001111",
  6148=>"001111011",
  6149=>"100100101",
  6150=>"011001000",
  6151=>"101011001",
  6152=>"000100100",
  6153=>"100100100",
  6154=>"011011110",
  6155=>"000011011",
  6156=>"000011011",
  6157=>"000011111",
  6158=>"101110110",
  6159=>"111000011",
  6160=>"110000000",
  6161=>"101000100",
  6162=>"101101011",
  6163=>"111111000",
  6164=>"111101110",
  6165=>"111100010",
  6166=>"100101110",
  6167=>"111111100",
  6168=>"000100100",
  6169=>"101111111",
  6170=>"010100110",
  6171=>"000000100",
  6172=>"101100111",
  6173=>"000001011",
  6174=>"000100101",
  6175=>"000000001",
  6176=>"111100000",
  6177=>"111111010",
  6178=>"001101111",
  6179=>"000000000",
  6180=>"111110101",
  6181=>"000011011",
  6182=>"001011000",
  6183=>"100000000",
  6184=>"111110110",
  6185=>"010111101",
  6186=>"110111111",
  6187=>"001000000",
  6188=>"111111011",
  6189=>"011011111",
  6190=>"111011000",
  6191=>"000000011",
  6192=>"011100100",
  6193=>"111001001",
  6194=>"101101000",
  6195=>"000000000",
  6196=>"001111111",
  6197=>"111011011",
  6198=>"010000000",
  6199=>"010111001",
  6200=>"111000000",
  6201=>"110000100",
  6202=>"011101011",
  6203=>"100100100",
  6204=>"001001000",
  6205=>"110010010",
  6206=>"100100100",
  6207=>"000010000",
  6208=>"111000001",
  6209=>"000100010",
  6210=>"100110111",
  6211=>"111100011",
  6212=>"100100000",
  6213=>"010000000",
  6214=>"001011111",
  6215=>"111100111",
  6216=>"101011001",
  6217=>"011100101",
  6218=>"111000110",
  6219=>"111000000",
  6220=>"101100100",
  6221=>"101011001",
  6222=>"110110111",
  6223=>"110011111",
  6224=>"000000100",
  6225=>"111111111",
  6226=>"110010111",
  6227=>"000000001",
  6228=>"000011001",
  6229=>"011000010",
  6230=>"100110001",
  6231=>"100100000",
  6232=>"110010111",
  6233=>"000000001",
  6234=>"000100001",
  6235=>"100000100",
  6236=>"111100111",
  6237=>"001000001",
  6238=>"011011011",
  6239=>"110110000",
  6240=>"010000001",
  6241=>"000001001",
  6242=>"100100100",
  6243=>"100110111",
  6244=>"111000001",
  6245=>"000001000",
  6246=>"011011011",
  6247=>"000001001",
  6248=>"000000000",
  6249=>"100101011",
  6250=>"000111011",
  6251=>"110111111",
  6252=>"000100000",
  6253=>"101011001",
  6254=>"111100100",
  6255=>"100100000",
  6256=>"100000000",
  6257=>"100000010",
  6258=>"001000100",
  6259=>"000011110",
  6260=>"000000001",
  6261=>"100100101",
  6262=>"010010011",
  6263=>"000000100",
  6264=>"000100110",
  6265=>"010100000",
  6266=>"100100000",
  6267=>"101111001",
  6268=>"011101000",
  6269=>"000001000",
  6270=>"000000000",
  6271=>"000000100",
  6272=>"011100001",
  6273=>"111110110",
  6274=>"000000101",
  6275=>"100111111",
  6276=>"011001000",
  6277=>"111100111",
  6278=>"110110100",
  6279=>"111000000",
  6280=>"111111111",
  6281=>"111010100",
  6282=>"000001000",
  6283=>"000100000",
  6284=>"011000001",
  6285=>"111101111",
  6286=>"000100011",
  6287=>"111100000",
  6288=>"100110101",
  6289=>"000101111",
  6290=>"011000000",
  6291=>"010111000",
  6292=>"110101000",
  6293=>"100100100",
  6294=>"000010111",
  6295=>"001101110",
  6296=>"100100100",
  6297=>"100011000",
  6298=>"000000110",
  6299=>"100100000",
  6300=>"111010011",
  6301=>"100100000",
  6302=>"000000011",
  6303=>"000100111",
  6304=>"100011001",
  6305=>"000000100",
  6306=>"000011000",
  6307=>"100101111",
  6308=>"000100111",
  6309=>"011100111",
  6310=>"000001100",
  6311=>"001100000",
  6312=>"111111110",
  6313=>"011010011",
  6314=>"000100111",
  6315=>"111000100",
  6316=>"101111111",
  6317=>"100100100",
  6318=>"000000110",
  6319=>"011011000",
  6320=>"000110100",
  6321=>"111110000",
  6322=>"000100111",
  6323=>"100000000",
  6324=>"010001101",
  6325=>"110111111",
  6326=>"000100100",
  6327=>"000000000",
  6328=>"110100000",
  6329=>"001001100",
  6330=>"010000000",
  6331=>"111111111",
  6332=>"110001001",
  6333=>"111110100",
  6334=>"000100100",
  6335=>"000000011",
  6336=>"110000000",
  6337=>"010100100",
  6338=>"010011011",
  6339=>"000000001",
  6340=>"001000001",
  6341=>"001101111",
  6342=>"001110111",
  6343=>"011100100",
  6344=>"111111010",
  6345=>"010000000",
  6346=>"010011110",
  6347=>"110111111",
  6348=>"000100000",
  6349=>"011010000",
  6350=>"100100101",
  6351=>"111000011",
  6352=>"100111111",
  6353=>"000011011",
  6354=>"110100000",
  6355=>"100110001",
  6356=>"100100100",
  6357=>"100000000",
  6358=>"000000000",
  6359=>"000111010",
  6360=>"010011011",
  6361=>"000001011",
  6362=>"111001111",
  6363=>"101100100",
  6364=>"111111010",
  6365=>"100000011",
  6366=>"000000011",
  6367=>"101101100",
  6368=>"000000100",
  6369=>"001100100",
  6370=>"000011011",
  6371=>"011001000",
  6372=>"010000000",
  6373=>"000010010",
  6374=>"111100000",
  6375=>"110110111",
  6376=>"111100100",
  6377=>"111011000",
  6378=>"100001000",
  6379=>"100100100",
  6380=>"000010000",
  6381=>"011010001",
  6382=>"010000000",
  6383=>"000100111",
  6384=>"000000000",
  6385=>"110110111",
  6386=>"100000100",
  6387=>"100100011",
  6388=>"011000100",
  6389=>"100101100",
  6390=>"000000101",
  6391=>"111000000",
  6392=>"000000000",
  6393=>"111011011",
  6394=>"111110111",
  6395=>"101111111",
  6396=>"111111111",
  6397=>"000111111",
  6398=>"111111111",
  6399=>"011000000",
  6400=>"000000001",
  6401=>"000000111",
  6402=>"111000000",
  6403=>"010001111",
  6404=>"110000111",
  6405=>"000000000",
  6406=>"000010110",
  6407=>"001001111",
  6408=>"111100101",
  6409=>"000010000",
  6410=>"001011011",
  6411=>"000000000",
  6412=>"101000001",
  6413=>"000000101",
  6414=>"100000110",
  6415=>"110100100",
  6416=>"101111001",
  6417=>"000010000",
  6418=>"000100000",
  6419=>"000000111",
  6420=>"111111100",
  6421=>"111000000",
  6422=>"010111101",
  6423=>"111000111",
  6424=>"000000000",
  6425=>"001111001",
  6426=>"000000100",
  6427=>"111111000",
  6428=>"000000110",
  6429=>"010000111",
  6430=>"111111100",
  6431=>"101000000",
  6432=>"000000111",
  6433=>"000101111",
  6434=>"101111101",
  6435=>"100100111",
  6436=>"000000011",
  6437=>"011011000",
  6438=>"000000000",
  6439=>"000101101",
  6440=>"100011101",
  6441=>"100010001",
  6442=>"000010000",
  6443=>"010001000",
  6444=>"000111111",
  6445=>"111111111",
  6446=>"000011010",
  6447=>"111111010",
  6448=>"000000111",
  6449=>"111001000",
  6450=>"111111000",
  6451=>"111111111",
  6452=>"001010000",
  6453=>"110010111",
  6454=>"000111110",
  6455=>"101001001",
  6456=>"110111110",
  6457=>"111001011",
  6458=>"011111110",
  6459=>"110001100",
  6460=>"001001011",
  6461=>"111110111",
  6462=>"000000000",
  6463=>"011100101",
  6464=>"111001000",
  6465=>"101111000",
  6466=>"111111111",
  6467=>"011110010",
  6468=>"000000000",
  6469=>"111110000",
  6470=>"110000111",
  6471=>"111111000",
  6472=>"010110111",
  6473=>"110111010",
  6474=>"000101101",
  6475=>"111100000",
  6476=>"101110000",
  6477=>"111000100",
  6478=>"110000000",
  6479=>"111001111",
  6480=>"000000000",
  6481=>"111110111",
  6482=>"000000110",
  6483=>"001100110",
  6484=>"000000110",
  6485=>"001001100",
  6486=>"110011100",
  6487=>"000000001",
  6488=>"001111000",
  6489=>"111110011",
  6490=>"011000000",
  6491=>"000100100",
  6492=>"000000000",
  6493=>"110000001",
  6494=>"111111111",
  6495=>"101111110",
  6496=>"001101111",
  6497=>"111001000",
  6498=>"000010011",
  6499=>"110000000",
  6500=>"111001000",
  6501=>"111111001",
  6502=>"000111100",
  6503=>"111000000",
  6504=>"001000110",
  6505=>"111111000",
  6506=>"101111000",
  6507=>"110000111",
  6508=>"010010111",
  6509=>"001010111",
  6510=>"111000000",
  6511=>"001111110",
  6512=>"111011111",
  6513=>"000010000",
  6514=>"000111011",
  6515=>"000000000",
  6516=>"101110010",
  6517=>"110000000",
  6518=>"101110111",
  6519=>"001100001",
  6520=>"101111011",
  6521=>"101111000",
  6522=>"100000011",
  6523=>"111100000",
  6524=>"001101010",
  6525=>"000100000",
  6526=>"000000010",
  6527=>"110000000",
  6528=>"000101111",
  6529=>"010011011",
  6530=>"000000101",
  6531=>"010001101",
  6532=>"000000111",
  6533=>"111111010",
  6534=>"000110010",
  6535=>"000100000",
  6536=>"010000000",
  6537=>"111000000",
  6538=>"111000100",
  6539=>"101100000",
  6540=>"000000000",
  6541=>"101000101",
  6542=>"010000000",
  6543=>"011000000",
  6544=>"111111111",
  6545=>"111101000",
  6546=>"010000000",
  6547=>"101100000",
  6548=>"000001111",
  6549=>"000111101",
  6550=>"111010000",
  6551=>"000000011",
  6552=>"000110111",
  6553=>"001000111",
  6554=>"111000000",
  6555=>"111000010",
  6556=>"111100100",
  6557=>"111000011",
  6558=>"101111111",
  6559=>"111000000",
  6560=>"001100011",
  6561=>"111111000",
  6562=>"000101101",
  6563=>"001000101",
  6564=>"001011000",
  6565=>"010111111",
  6566=>"000111110",
  6567=>"000111111",
  6568=>"000000110",
  6569=>"000111111",
  6570=>"110000000",
  6571=>"011010000",
  6572=>"111001100",
  6573=>"001001000",
  6574=>"111000000",
  6575=>"001000111",
  6576=>"111111001",
  6577=>"000000000",
  6578=>"000000011",
  6579=>"000001100",
  6580=>"111100111",
  6581=>"111110000",
  6582=>"011000101",
  6583=>"011101101",
  6584=>"000000101",
  6585=>"000000111",
  6586=>"000000000",
  6587=>"000101001",
  6588=>"000000000",
  6589=>"110111111",
  6590=>"110001000",
  6591=>"011110000",
  6592=>"111000000",
  6593=>"111000000",
  6594=>"111111111",
  6595=>"111101110",
  6596=>"111111000",
  6597=>"111100000",
  6598=>"010110111",
  6599=>"111010001",
  6600=>"011100001",
  6601=>"101000111",
  6602=>"000000000",
  6603=>"100000001",
  6604=>"111100000",
  6605=>"000101010",
  6606=>"111111101",
  6607=>"000111111",
  6608=>"100000000",
  6609=>"110000001",
  6610=>"100100100",
  6611=>"110111111",
  6612=>"101000001",
  6613=>"011100000",
  6614=>"001111111",
  6615=>"111001111",
  6616=>"001101110",
  6617=>"000011011",
  6618=>"011001110",
  6619=>"000000000",
  6620=>"010111101",
  6621=>"000001100",
  6622=>"000000000",
  6623=>"001111110",
  6624=>"111111001",
  6625=>"111000000",
  6626=>"111000000",
  6627=>"111000010",
  6628=>"000001000",
  6629=>"000010111",
  6630=>"000000111",
  6631=>"111000000",
  6632=>"111101010",
  6633=>"000000110",
  6634=>"100110010",
  6635=>"010000101",
  6636=>"011100101",
  6637=>"101100000",
  6638=>"010000000",
  6639=>"111000000",
  6640=>"000000000",
  6641=>"111001010",
  6642=>"000111110",
  6643=>"110111110",
  6644=>"001000000",
  6645=>"010000000",
  6646=>"111000000",
  6647=>"111101001",
  6648=>"000111101",
  6649=>"100000110",
  6650=>"111000111",
  6651=>"110001101",
  6652=>"111010111",
  6653=>"000010000",
  6654=>"110001001",
  6655=>"100100000",
  6656=>"010110000",
  6657=>"100000011",
  6658=>"101000000",
  6659=>"000111111",
  6660=>"100111111",
  6661=>"000000000",
  6662=>"100000000",
  6663=>"000001111",
  6664=>"101000000",
  6665=>"000010000",
  6666=>"011110110",
  6667=>"111111111",
  6668=>"100000000",
  6669=>"000001000",
  6670=>"111101011",
  6671=>"000000000",
  6672=>"110111000",
  6673=>"011111011",
  6674=>"111011101",
  6675=>"010010110",
  6676=>"111111111",
  6677=>"100010100",
  6678=>"110000000",
  6679=>"110010111",
  6680=>"000111000",
  6681=>"110111111",
  6682=>"101111111",
  6683=>"000001000",
  6684=>"111101001",
  6685=>"111001111",
  6686=>"111011000",
  6687=>"010010000",
  6688=>"000000000",
  6689=>"000010001",
  6690=>"101011000",
  6691=>"011001000",
  6692=>"000100110",
  6693=>"001010010",
  6694=>"110111100",
  6695=>"000000111",
  6696=>"110111111",
  6697=>"111111111",
  6698=>"001100000",
  6699=>"111100000",
  6700=>"100011011",
  6701=>"111110111",
  6702=>"101100101",
  6703=>"011101001",
  6704=>"111001100",
  6705=>"000001001",
  6706=>"000101110",
  6707=>"111010000",
  6708=>"110110111",
  6709=>"101100110",
  6710=>"011011110",
  6711=>"000000000",
  6712=>"010000000",
  6713=>"000000000",
  6714=>"101000101",
  6715=>"000111001",
  6716=>"010011001",
  6717=>"011111110",
  6718=>"000000000",
  6719=>"100110111",
  6720=>"110111100",
  6721=>"000011111",
  6722=>"101000000",
  6723=>"100110111",
  6724=>"111000000",
  6725=>"101000000",
  6726=>"111000101",
  6727=>"111111001",
  6728=>"110110111",
  6729=>"000110110",
  6730=>"001000000",
  6731=>"011110010",
  6732=>"000010010",
  6733=>"010011001",
  6734=>"000100110",
  6735=>"010101000",
  6736=>"111111111",
  6737=>"010010000",
  6738=>"001100101",
  6739=>"111001000",
  6740=>"110000000",
  6741=>"010001111",
  6742=>"100011000",
  6743=>"000111100",
  6744=>"111110110",
  6745=>"001001001",
  6746=>"001000111",
  6747=>"111111111",
  6748=>"000000000",
  6749=>"000001001",
  6750=>"111111010",
  6751=>"001011110",
  6752=>"100000010",
  6753=>"110110011",
  6754=>"101000100",
  6755=>"110100000",
  6756=>"011111101",
  6757=>"011001001",
  6758=>"110110110",
  6759=>"111111100",
  6760=>"010010111",
  6761=>"000000000",
  6762=>"110111100",
  6763=>"111101110",
  6764=>"101111111",
  6765=>"000110011",
  6766=>"111101101",
  6767=>"111111111",
  6768=>"000100100",
  6769=>"000000001",
  6770=>"110110010",
  6771=>"000110010",
  6772=>"010010000",
  6773=>"000000000",
  6774=>"000011010",
  6775=>"101000000",
  6776=>"100000000",
  6777=>"110100010",
  6778=>"011010011",
  6779=>"011111010",
  6780=>"110111011",
  6781=>"111100000",
  6782=>"010000000",
  6783=>"111001001",
  6784=>"001000011",
  6785=>"111101100",
  6786=>"111000010",
  6787=>"011100101",
  6788=>"111111101",
  6789=>"111101010",
  6790=>"000010010",
  6791=>"000110110",
  6792=>"101001011",
  6793=>"000010110",
  6794=>"010011000",
  6795=>"111111010",
  6796=>"000110010",
  6797=>"111000010",
  6798=>"000001011",
  6799=>"000000000",
  6800=>"100111110",
  6801=>"010110101",
  6802=>"000111111",
  6803=>"110111110",
  6804=>"001111100",
  6805=>"001000101",
  6806=>"111111010",
  6807=>"100100011",
  6808=>"111111111",
  6809=>"110111111",
  6810=>"000100111",
  6811=>"111101000",
  6812=>"110101000",
  6813=>"000000000",
  6814=>"001111111",
  6815=>"110100100",
  6816=>"001101101",
  6817=>"111000000",
  6818=>"001101111",
  6819=>"010001111",
  6820=>"110111100",
  6821=>"100011010",
  6822=>"111110110",
  6823=>"001001000",
  6824=>"001100111",
  6825=>"000000111",
  6826=>"000000111",
  6827=>"111000000",
  6828=>"111011010",
  6829=>"100000100",
  6830=>"111110110",
  6831=>"011010100",
  6832=>"101000000",
  6833=>"010111011",
  6834=>"011100111",
  6835=>"011100100",
  6836=>"100101111",
  6837=>"111110001",
  6838=>"000010011",
  6839=>"000000010",
  6840=>"010010111",
  6841=>"000111111",
  6842=>"010110011",
  6843=>"000111110",
  6844=>"110011011",
  6845=>"111111111",
  6846=>"101100100",
  6847=>"010000000",
  6848=>"111000000",
  6849=>"010000010",
  6850=>"111111111",
  6851=>"100110100",
  6852=>"111001000",
  6853=>"111110110",
  6854=>"100110100",
  6855=>"010111010",
  6856=>"010001010",
  6857=>"100000000",
  6858=>"110000111",
  6859=>"000100111",
  6860=>"010111011",
  6861=>"011111110",
  6862=>"111111111",
  6863=>"000000000",
  6864=>"100110000",
  6865=>"000110110",
  6866=>"000010001",
  6867=>"000000010",
  6868=>"000000100",
  6869=>"010100100",
  6870=>"000010000",
  6871=>"000010110",
  6872=>"110111111",
  6873=>"010010000",
  6874=>"101100100",
  6875=>"010110110",
  6876=>"111100101",
  6877=>"101001011",
  6878=>"010111110",
  6879=>"000000000",
  6880=>"101001000",
  6881=>"111000000",
  6882=>"101100100",
  6883=>"000100100",
  6884=>"000000000",
  6885=>"111000101",
  6886=>"111000000",
  6887=>"100101110",
  6888=>"010000000",
  6889=>"000000000",
  6890=>"110011011",
  6891=>"011111111",
  6892=>"100000000",
  6893=>"000000000",
  6894=>"000001111",
  6895=>"110100000",
  6896=>"110111101",
  6897=>"111011001",
  6898=>"000001000",
  6899=>"111101110",
  6900=>"001110100",
  6901=>"000001111",
  6902=>"100000010",
  6903=>"111000111",
  6904=>"111111111",
  6905=>"111000111",
  6906=>"010000001",
  6907=>"000011010",
  6908=>"000000000",
  6909=>"101000000",
  6910=>"010111111",
  6911=>"100000000",
  6912=>"101110010",
  6913=>"000111111",
  6914=>"010000110",
  6915=>"000111111",
  6916=>"101011000",
  6917=>"000001000",
  6918=>"000010000",
  6919=>"101111010",
  6920=>"100000000",
  6921=>"010000110",
  6922=>"000001000",
  6923=>"111000000",
  6924=>"111111000",
  6925=>"000111111",
  6926=>"011010000",
  6927=>"000000100",
  6928=>"000001000",
  6929=>"000000101",
  6930=>"011011000",
  6931=>"000000010",
  6932=>"101101111",
  6933=>"010111111",
  6934=>"011111111",
  6935=>"111110110",
  6936=>"011101001",
  6937=>"000000101",
  6938=>"000000101",
  6939=>"111100000",
  6940=>"111000011",
  6941=>"001000001",
  6942=>"010110001",
  6943=>"000011111",
  6944=>"111101111",
  6945=>"000101001",
  6946=>"111101000",
  6947=>"101111000",
  6948=>"001001011",
  6949=>"011001000",
  6950=>"011011000",
  6951=>"001000000",
  6952=>"000011111",
  6953=>"111111001",
  6954=>"000000111",
  6955=>"000000111",
  6956=>"111001001",
  6957=>"111000010",
  6958=>"100000100",
  6959=>"000010000",
  6960=>"000110111",
  6961=>"110000000",
  6962=>"101110111",
  6963=>"101000011",
  6964=>"111000000",
  6965=>"100100000",
  6966=>"110000011",
  6967=>"111100000",
  6968=>"111101000",
  6969=>"101001000",
  6970=>"001101111",
  6971=>"111010010",
  6972=>"111001000",
  6973=>"010111011",
  6974=>"000001100",
  6975=>"100110011",
  6976=>"001000000",
  6977=>"100000000",
  6978=>"110111000",
  6979=>"001000000",
  6980=>"100111001",
  6981=>"000000100",
  6982=>"000000111",
  6983=>"000001000",
  6984=>"101101000",
  6985=>"000001000",
  6986=>"000010001",
  6987=>"000101111",
  6988=>"111000000",
  6989=>"000000000",
  6990=>"001011000",
  6991=>"111101000",
  6992=>"010010000",
  6993=>"011001010",
  6994=>"010000001",
  6995=>"000000000",
  6996=>"000011010",
  6997=>"110000100",
  6998=>"000011110",
  6999=>"000010011",
  7000=>"101111111",
  7001=>"010100100",
  7002=>"000100111",
  7003=>"110110000",
  7004=>"000000000",
  7005=>"000101111",
  7006=>"111110000",
  7007=>"010010000",
  7008=>"111011000",
  7009=>"000110111",
  7010=>"000000111",
  7011=>"111001001",
  7012=>"101111000",
  7013=>"110000000",
  7014=>"111000000",
  7015=>"111111111",
  7016=>"100110000",
  7017=>"000100000",
  7018=>"111111000",
  7019=>"000010000",
  7020=>"011111111",
  7021=>"000101111",
  7022=>"111111000",
  7023=>"011111110",
  7024=>"011011011",
  7025=>"001111111",
  7026=>"011000010",
  7027=>"111110010",
  7028=>"111101000",
  7029=>"000000000",
  7030=>"010111001",
  7031=>"111010000",
  7032=>"111100101",
  7033=>"110010011",
  7034=>"100000000",
  7035=>"000000000",
  7036=>"111011100",
  7037=>"000001001",
  7038=>"110001111",
  7039=>"000001111",
  7040=>"000010001",
  7041=>"000000000",
  7042=>"000000100",
  7043=>"000101000",
  7044=>"101101000",
  7045=>"111111010",
  7046=>"110110100",
  7047=>"110100100",
  7048=>"010000111",
  7049=>"000000101",
  7050=>"100010111",
  7051=>"000110000",
  7052=>"000000111",
  7053=>"010010101",
  7054=>"000110110",
  7055=>"000000000",
  7056=>"111000000",
  7057=>"111000000",
  7058=>"101001110",
  7059=>"000000110",
  7060=>"100100100",
  7061=>"000000100",
  7062=>"011010000",
  7063=>"101111011",
  7064=>"010010000",
  7065=>"000011111",
  7066=>"000010111",
  7067=>"111000000",
  7068=>"100000111",
  7069=>"111111011",
  7070=>"100011111",
  7071=>"000000000",
  7072=>"010111101",
  7073=>"101011111",
  7074=>"000010011",
  7075=>"011001000",
  7076=>"000000000",
  7077=>"011001000",
  7078=>"111010000",
  7079=>"000000011",
  7080=>"100000100",
  7081=>"110011111",
  7082=>"011101111",
  7083=>"001000000",
  7084=>"001101101",
  7085=>"000010110",
  7086=>"101011111",
  7087=>"111111000",
  7088=>"100100000",
  7089=>"001001111",
  7090=>"000000101",
  7091=>"010110100",
  7092=>"110100000",
  7093=>"001101101",
  7094=>"000100100",
  7095=>"111010111",
  7096=>"111000000",
  7097=>"101101001",
  7098=>"111010010",
  7099=>"011000011",
  7100=>"111001010",
  7101=>"111111111",
  7102=>"000001110",
  7103=>"010111111",
  7104=>"000100101",
  7105=>"000000000",
  7106=>"111111000",
  7107=>"110011111",
  7108=>"101101111",
  7109=>"000101100",
  7110=>"000101111",
  7111=>"101100111",
  7112=>"001100000",
  7113=>"111001000",
  7114=>"000010001",
  7115=>"010000000",
  7116=>"011011000",
  7117=>"111111000",
  7118=>"000000000",
  7119=>"000000111",
  7120=>"110111000",
  7121=>"011111100",
  7122=>"101101100",
  7123=>"010000000",
  7124=>"111101000",
  7125=>"000110111",
  7126=>"111011010",
  7127=>"000100111",
  7128=>"111010000",
  7129=>"111101000",
  7130=>"010111110",
  7131=>"001000111",
  7132=>"011011110",
  7133=>"000010011",
  7134=>"111100011",
  7135=>"000001000",
  7136=>"000000100",
  7137=>"000110111",
  7138=>"111101000",
  7139=>"100111011",
  7140=>"110000010",
  7141=>"010010000",
  7142=>"011001000",
  7143=>"101101111",
  7144=>"111111000",
  7145=>"011001111",
  7146=>"001000100",
  7147=>"111101101",
  7148=>"001111000",
  7149=>"001001000",
  7150=>"010010010",
  7151=>"011000001",
  7152=>"101100011",
  7153=>"110111110",
  7154=>"011110100",
  7155=>"000001100",
  7156=>"110101001",
  7157=>"000000000",
  7158=>"011111000",
  7159=>"111110000",
  7160=>"000100000",
  7161=>"111111011",
  7162=>"101111111",
  7163=>"111000000",
  7164=>"111011000",
  7165=>"000110110",
  7166=>"001000000",
  7167=>"000000000",
  7168=>"001000110",
  7169=>"001000110",
  7170=>"100100111",
  7171=>"001000001",
  7172=>"110100100",
  7173=>"011001000",
  7174=>"001001000",
  7175=>"001000001",
  7176=>"110000100",
  7177=>"000100110",
  7178=>"110000000",
  7179=>"110000100",
  7180=>"001001000",
  7181=>"001001000",
  7182=>"110100100",
  7183=>"110100100",
  7184=>"111011001",
  7185=>"111001001",
  7186=>"011100011",
  7187=>"010010000",
  7188=>"001111100",
  7189=>"100000000",
  7190=>"100111000",
  7191=>"110100010",
  7192=>"000100000",
  7193=>"100111101",
  7194=>"001011000",
  7195=>"000000011",
  7196=>"000000110",
  7197=>"011001011",
  7198=>"111101011",
  7199=>"000100000",
  7200=>"010000111",
  7201=>"011011000",
  7202=>"000100111",
  7203=>"000000011",
  7204=>"000000000",
  7205=>"001111110",
  7206=>"100101111",
  7207=>"010011000",
  7208=>"001001111",
  7209=>"000000100",
  7210=>"100100000",
  7211=>"000001000",
  7212=>"100101101",
  7213=>"110101011",
  7214=>"011100110",
  7215=>"000011000",
  7216=>"010011011",
  7217=>"111010010",
  7218=>"000010011",
  7219=>"011111111",
  7220=>"100100110",
  7221=>"100100101",
  7222=>"111011110",
  7223=>"010100010",
  7224=>"011011000",
  7225=>"111000111",
  7226=>"110100110",
  7227=>"010100110",
  7228=>"000001000",
  7229=>"111111110",
  7230=>"100001111",
  7231=>"111100000",
  7232=>"100110111",
  7233=>"001000000",
  7234=>"011011000",
  7235=>"110000010",
  7236=>"000001011",
  7237=>"111000100",
  7238=>"001000011",
  7239=>"111101111",
  7240=>"110110010",
  7241=>"111011011",
  7242=>"110100111",
  7243=>"110100100",
  7244=>"110100110",
  7245=>"001111111",
  7246=>"010011111",
  7247=>"100100111",
  7248=>"001011011",
  7249=>"111110111",
  7250=>"111110010",
  7251=>"000000000",
  7252=>"100111111",
  7253=>"111111111",
  7254=>"011110011",
  7255=>"100100001",
  7256=>"111000010",
  7257=>"111111111",
  7258=>"101111001",
  7259=>"010010100",
  7260=>"001011000",
  7261=>"001000000",
  7262=>"000011111",
  7263=>"100100110",
  7264=>"000100010",
  7265=>"010011011",
  7266=>"111001100",
  7267=>"100000000",
  7268=>"000110111",
  7269=>"001011011",
  7270=>"000000111",
  7271=>"110100100",
  7272=>"110000001",
  7273=>"011011001",
  7274=>"011000000",
  7275=>"100100110",
  7276=>"000101111",
  7277=>"111001011",
  7278=>"011000000",
  7279=>"010000110",
  7280=>"101111101",
  7281=>"111000000",
  7282=>"000100111",
  7283=>"100100111",
  7284=>"001000000",
  7285=>"110100010",
  7286=>"001001001",
  7287=>"011011011",
  7288=>"000000000",
  7289=>"011001000",
  7290=>"100010100",
  7291=>"010011100",
  7292=>"111111011",
  7293=>"111110000",
  7294=>"001011011",
  7295=>"000101111",
  7296=>"100000110",
  7297=>"001000000",
  7298=>"011000010",
  7299=>"000000010",
  7300=>"100000110",
  7301=>"110110101",
  7302=>"000100100",
  7303=>"000011111",
  7304=>"000000000",
  7305=>"011011111",
  7306=>"010010011",
  7307=>"011011000",
  7308=>"000000011",
  7309=>"000000000",
  7310=>"100101001",
  7311=>"110000001",
  7312=>"100111111",
  7313=>"100110110",
  7314=>"000100010",
  7315=>"001000111",
  7316=>"100001011",
  7317=>"000001000",
  7318=>"111110111",
  7319=>"001000000",
  7320=>"000110111",
  7321=>"111001001",
  7322=>"100100110",
  7323=>"000000110",
  7324=>"001011011",
  7325=>"100001001",
  7326=>"111000000",
  7327=>"110100110",
  7328=>"001000100",
  7329=>"111010000",
  7330=>"001011000",
  7331=>"110000100",
  7332=>"001101101",
  7333=>"100110111",
  7334=>"111111000",
  7335=>"011011001",
  7336=>"011111011",
  7337=>"011010100",
  7338=>"001001000",
  7339=>"100000100",
  7340=>"010011000",
  7341=>"101101111",
  7342=>"101100110",
  7343=>"001011010",
  7344=>"000010101",
  7345=>"000111111",
  7346=>"010011000",
  7347=>"000000000",
  7348=>"011000011",
  7349=>"100010100",
  7350=>"011010111",
  7351=>"001011010",
  7352=>"111011010",
  7353=>"100011001",
  7354=>"001001010",
  7355=>"111000111",
  7356=>"001111001",
  7357=>"001011011",
  7358=>"000000000",
  7359=>"001111001",
  7360=>"110000000",
  7361=>"000100000",
  7362=>"110111011",
  7363=>"010011010",
  7364=>"000110111",
  7365=>"100111111",
  7366=>"001000001",
  7367=>"100100100",
  7368=>"000010001",
  7369=>"100100100",
  7370=>"110111001",
  7371=>"101100111",
  7372=>"111110110",
  7373=>"010000110",
  7374=>"110110011",
  7375=>"100011111",
  7376=>"000100010",
  7377=>"110110110",
  7378=>"100000101",
  7379=>"101000100",
  7380=>"110100111",
  7381=>"011010011",
  7382=>"101100110",
  7383=>"111011000",
  7384=>"100100010",
  7385=>"000001011",
  7386=>"110010100",
  7387=>"101001001",
  7388=>"110100110",
  7389=>"001001100",
  7390=>"101100100",
  7391=>"111100000",
  7392=>"100111111",
  7393=>"000011000",
  7394=>"000001100",
  7395=>"101111011",
  7396=>"100100100",
  7397=>"000000000",
  7398=>"011101011",
  7399=>"011110010",
  7400=>"001001001",
  7401=>"100011010",
  7402=>"110100000",
  7403=>"001011011",
  7404=>"001011011",
  7405=>"111100101",
  7406=>"000100010",
  7407=>"001111110",
  7408=>"110100110",
  7409=>"010111100",
  7410=>"010100000",
  7411=>"111111101",
  7412=>"111111011",
  7413=>"001001000",
  7414=>"100000000",
  7415=>"011001000",
  7416=>"000001001",
  7417=>"011011000",
  7418=>"110100000",
  7419=>"000010110",
  7420=>"100100110",
  7421=>"001011000",
  7422=>"001010011",
  7423=>"100110110",
  7424=>"000000100",
  7425=>"110000000",
  7426=>"000001001",
  7427=>"111101101",
  7428=>"000110110",
  7429=>"001111111",
  7430=>"000000000",
  7431=>"000000111",
  7432=>"110111111",
  7433=>"000010000",
  7434=>"001000110",
  7435=>"000000000",
  7436=>"110100000",
  7437=>"000000010",
  7438=>"111010010",
  7439=>"111000000",
  7440=>"100111111",
  7441=>"101010111",
  7442=>"000111111",
  7443=>"101101000",
  7444=>"111000000",
  7445=>"111101101",
  7446=>"000111111",
  7447=>"101011111",
  7448=>"110001000",
  7449=>"111111111",
  7450=>"101101111",
  7451=>"001000000",
  7452=>"000000011",
  7453=>"001101000",
  7454=>"111111001",
  7455=>"111101100",
  7456=>"000010011",
  7457=>"111111100",
  7458=>"100000110",
  7459=>"000111111",
  7460=>"110110110",
  7461=>"000010000",
  7462=>"101000000",
  7463=>"100000001",
  7464=>"110100110",
  7465=>"010110100",
  7466=>"101000011",
  7467=>"110100010",
  7468=>"100100001",
  7469=>"111001000",
  7470=>"000111111",
  7471=>"000011000",
  7472=>"000010111",
  7473=>"011100100",
  7474=>"000000000",
  7475=>"000111111",
  7476=>"000111011",
  7477=>"000111001",
  7478=>"000111010",
  7479=>"100000000",
  7480=>"111111111",
  7481=>"111001001",
  7482=>"011000000",
  7483=>"111000000",
  7484=>"100010001",
  7485=>"000111011",
  7486=>"111000010",
  7487=>"000000000",
  7488=>"111000000",
  7489=>"011110100",
  7490=>"110111110",
  7491=>"000110011",
  7492=>"111000000",
  7493=>"111011000",
  7494=>"111000000",
  7495=>"101111000",
  7496=>"111111011",
  7497=>"110000000",
  7498=>"111000000",
  7499=>"001111100",
  7500=>"111000000",
  7501=>"000000110",
  7502=>"110001001",
  7503=>"110000000",
  7504=>"000101010",
  7505=>"101111010",
  7506=>"100000001",
  7507=>"100110000",
  7508=>"111001001",
  7509=>"000110100",
  7510=>"000001011",
  7511=>"000000101",
  7512=>"111001001",
  7513=>"011110110",
  7514=>"010010000",
  7515=>"111111110",
  7516=>"000111111",
  7517=>"010010001",
  7518=>"111100000",
  7519=>"000011000",
  7520=>"000000111",
  7521=>"000010000",
  7522=>"110000101",
  7523=>"011011000",
  7524=>"011001100",
  7525=>"011000111",
  7526=>"101110010",
  7527=>"000100111",
  7528=>"110000101",
  7529=>"111011001",
  7530=>"000100111",
  7531=>"111101111",
  7532=>"000111111",
  7533=>"111000010",
  7534=>"100000000",
  7535=>"000000000",
  7536=>"001011011",
  7537=>"100111111",
  7538=>"000110010",
  7539=>"111110010",
  7540=>"000001010",
  7541=>"110000000",
  7542=>"001001000",
  7543=>"111100000",
  7544=>"111111001",
  7545=>"000101001",
  7546=>"000000000",
  7547=>"000110000",
  7548=>"000000110",
  7549=>"101001100",
  7550=>"111101000",
  7551=>"010011000",
  7552=>"111110110",
  7553=>"001101010",
  7554=>"000000101",
  7555=>"111111110",
  7556=>"000001011",
  7557=>"111011110",
  7558=>"100011011",
  7559=>"101011110",
  7560=>"000111110",
  7561=>"000010010",
  7562=>"111010000",
  7563=>"101111000",
  7564=>"000000000",
  7565=>"111000011",
  7566=>"001111111",
  7567=>"111011111",
  7568=>"100000000",
  7569=>"111000000",
  7570=>"101000101",
  7571=>"101010001",
  7572=>"000001111",
  7573=>"000000111",
  7574=>"111111111",
  7575=>"010110100",
  7576=>"111000010",
  7577=>"010001111",
  7578=>"001011010",
  7579=>"111111001",
  7580=>"110111110",
  7581=>"000010110",
  7582=>"111111111",
  7583=>"000111110",
  7584=>"110110001",
  7585=>"011110000",
  7586=>"100111010",
  7587=>"110000001",
  7588=>"001000000",
  7589=>"111011000",
  7590=>"000111110",
  7591=>"111101011",
  7592=>"000000110",
  7593=>"000000111",
  7594=>"000111100",
  7595=>"000010110",
  7596=>"110111110",
  7597=>"000000000",
  7598=>"001001011",
  7599=>"111100000",
  7600=>"110000000",
  7601=>"110110010",
  7602=>"111000000",
  7603=>"110000000",
  7604=>"001110110",
  7605=>"100111110",
  7606=>"010111111",
  7607=>"101011110",
  7608=>"001010011",
  7609=>"000110010",
  7610=>"000000111",
  7611=>"111111001",
  7612=>"101111111",
  7613=>"011001111",
  7614=>"011100110",
  7615=>"010111111",
  7616=>"111100000",
  7617=>"001011011",
  7618=>"111000000",
  7619=>"000011000",
  7620=>"010011010",
  7621=>"001000110",
  7622=>"000000100",
  7623=>"010000111",
  7624=>"111000110",
  7625=>"111001000",
  7626=>"000000000",
  7627=>"111000100",
  7628=>"010000000",
  7629=>"001010011",
  7630=>"001111110",
  7631=>"000011001",
  7632=>"011000000",
  7633=>"100001011",
  7634=>"001011000",
  7635=>"101101101",
  7636=>"101011000",
  7637=>"001011110",
  7638=>"111111101",
  7639=>"000000001",
  7640=>"110101000",
  7641=>"110000101",
  7642=>"111111100",
  7643=>"111101001",
  7644=>"001011011",
  7645=>"000100111",
  7646=>"111011010",
  7647=>"101001100",
  7648=>"010000000",
  7649=>"000011101",
  7650=>"011111001",
  7651=>"111111011",
  7652=>"001000111",
  7653=>"011000101",
  7654=>"000000001",
  7655=>"000100110",
  7656=>"000000000",
  7657=>"101110011",
  7658=>"110000010",
  7659=>"001011111",
  7660=>"111101000",
  7661=>"101111111",
  7662=>"000110000",
  7663=>"000000010",
  7664=>"111000000",
  7665=>"100100110",
  7666=>"100000010",
  7667=>"110011011",
  7668=>"000000101",
  7669=>"110000000",
  7670=>"100000011",
  7671=>"010111111",
  7672=>"000000001",
  7673=>"111101000",
  7674=>"100111100",
  7675=>"111101100",
  7676=>"111011111",
  7677=>"001111111",
  7678=>"000011011",
  7679=>"010000010",
  7680=>"110011000",
  7681=>"001101111",
  7682=>"000000000",
  7683=>"111111111",
  7684=>"011101111",
  7685=>"111111001",
  7686=>"000000000",
  7687=>"111010111",
  7688=>"111110111",
  7689=>"000000000",
  7690=>"000000000",
  7691=>"111011111",
  7692=>"000000110",
  7693=>"001000000",
  7694=>"111100100",
  7695=>"111111100",
  7696=>"000001001",
  7697=>"111111110",
  7698=>"111111110",
  7699=>"011100000",
  7700=>"101101110",
  7701=>"000000000",
  7702=>"000010100",
  7703=>"001010010",
  7704=>"000101000",
  7705=>"011111000",
  7706=>"111111111",
  7707=>"110010010",
  7708=>"000000000",
  7709=>"000000000",
  7710=>"111000000",
  7711=>"111000111",
  7712=>"000000111",
  7713=>"000111111",
  7714=>"111011110",
  7715=>"111111111",
  7716=>"001001011",
  7717=>"000010001",
  7718=>"111111000",
  7719=>"110111110",
  7720=>"111011000",
  7721=>"111111111",
  7722=>"000001000",
  7723=>"111111000",
  7724=>"000000000",
  7725=>"000100010",
  7726=>"101011101",
  7727=>"001010000",
  7728=>"000000010",
  7729=>"011011011",
  7730=>"001111111",
  7731=>"111000000",
  7732=>"000000000",
  7733=>"000000000",
  7734=>"010000000",
  7735=>"111010111",
  7736=>"111101111",
  7737=>"000000000",
  7738=>"001101111",
  7739=>"000000111",
  7740=>"110010011",
  7741=>"000011010",
  7742=>"001110110",
  7743=>"111010011",
  7744=>"010000100",
  7745=>"000100111",
  7746=>"111111111",
  7747=>"111101110",
  7748=>"111111011",
  7749=>"000111111",
  7750=>"000000110",
  7751=>"110000000",
  7752=>"010110101",
  7753=>"000000000",
  7754=>"000000111",
  7755=>"000000000",
  7756=>"010110110",
  7757=>"110110111",
  7758=>"101111101",
  7759=>"111001000",
  7760=>"011111110",
  7761=>"011111000",
  7762=>"010111010",
  7763=>"011000000",
  7764=>"001110000",
  7765=>"000110110",
  7766=>"010011000",
  7767=>"100000000",
  7768=>"101110110",
  7769=>"100000010",
  7770=>"000000001",
  7771=>"000000000",
  7772=>"011111011",
  7773=>"001001111",
  7774=>"111111111",
  7775=>"011110011",
  7776=>"111110111",
  7777=>"111111111",
  7778=>"000010001",
  7779=>"001001000",
  7780=>"010001101",
  7781=>"000110111",
  7782=>"000001001",
  7783=>"111011010",
  7784=>"111001101",
  7785=>"000000000",
  7786=>"001011000",
  7787=>"010110111",
  7788=>"111111111",
  7789=>"000001001",
  7790=>"111110011",
  7791=>"000001111",
  7792=>"000000001",
  7793=>"000000110",
  7794=>"000000000",
  7795=>"000000000",
  7796=>"111111111",
  7797=>"000000000",
  7798=>"000001001",
  7799=>"111001001",
  7800=>"111000000",
  7801=>"000001111",
  7802=>"001000111",
  7803=>"101101111",
  7804=>"110000000",
  7805=>"110100000",
  7806=>"110000001",
  7807=>"100100000",
  7808=>"111000000",
  7809=>"000000001",
  7810=>"111111111",
  7811=>"111000100",
  7812=>"111110000",
  7813=>"000010000",
  7814=>"000000000",
  7815=>"000000111",
  7816=>"000000100",
  7817=>"010100001",
  7818=>"001011000",
  7819=>"111000000",
  7820=>"111111111",
  7821=>"011010010",
  7822=>"100111111",
  7823=>"011011001",
  7824=>"000111011",
  7825=>"000000000",
  7826=>"000110000",
  7827=>"111111010",
  7828=>"000001000",
  7829=>"111111111",
  7830=>"011111111",
  7831=>"111111111",
  7832=>"001111011",
  7833=>"011111111",
  7834=>"011010010",
  7835=>"100000101",
  7836=>"111111110",
  7837=>"000000100",
  7838=>"111111110",
  7839=>"000000000",
  7840=>"000101011",
  7841=>"000010000",
  7842=>"001011010",
  7843=>"001011110",
  7844=>"111000010",
  7845=>"011100001",
  7846=>"111110110",
  7847=>"000000111",
  7848=>"000100011",
  7849=>"110111111",
  7850=>"110111111",
  7851=>"000000000",
  7852=>"110010011",
  7853=>"111111010",
  7854=>"001011010",
  7855=>"111111101",
  7856=>"100111111",
  7857=>"111011011",
  7858=>"001110000",
  7859=>"100111111",
  7860=>"000011111",
  7861=>"000000000",
  7862=>"111111011",
  7863=>"111111100",
  7864=>"111110010",
  7865=>"100010000",
  7866=>"000000000",
  7867=>"001001111",
  7868=>"000000101",
  7869=>"111111011",
  7870=>"111111111",
  7871=>"000000000",
  7872=>"000011010",
  7873=>"111111010",
  7874=>"000110111",
  7875=>"100110111",
  7876=>"000010010",
  7877=>"110000000",
  7878=>"000001000",
  7879=>"000000001",
  7880=>"010111011",
  7881=>"110000000",
  7882=>"010111000",
  7883=>"000000001",
  7884=>"111111100",
  7885=>"110000000",
  7886=>"000000000",
  7887=>"110000101",
  7888=>"011010000",
  7889=>"101100111",
  7890=>"111001000",
  7891=>"111111101",
  7892=>"110111111",
  7893=>"000101111",
  7894=>"110111000",
  7895=>"001111110",
  7896=>"000000000",
  7897=>"110000100",
  7898=>"000001000",
  7899=>"000000000",
  7900=>"000011011",
  7901=>"111111111",
  7902=>"111111000",
  7903=>"111000000",
  7904=>"111100000",
  7905=>"000000000",
  7906=>"000111110",
  7907=>"111111011",
  7908=>"111010000",
  7909=>"111010110",
  7910=>"101111111",
  7911=>"000010000",
  7912=>"101001000",
  7913=>"110010111",
  7914=>"000000000",
  7915=>"110000000",
  7916=>"111111111",
  7917=>"111111111",
  7918=>"000000000",
  7919=>"101111111",
  7920=>"000000000",
  7921=>"011001000",
  7922=>"111111111",
  7923=>"001001000",
  7924=>"111110100",
  7925=>"000000100",
  7926=>"010100110",
  7927=>"000000000",
  7928=>"000011111",
  7929=>"011100111",
  7930=>"000000000",
  7931=>"001000000",
  7932=>"000000101",
  7933=>"111111001",
  7934=>"111101101",
  7935=>"000000000",
  7936=>"110010110",
  7937=>"110000000",
  7938=>"001001111",
  7939=>"111000101",
  7940=>"011001011",
  7941=>"010000001",
  7942=>"001000110",
  7943=>"101111111",
  7944=>"010000001",
  7945=>"001001001",
  7946=>"000100011",
  7947=>"000001000",
  7948=>"111000100",
  7949=>"000100000",
  7950=>"000001001",
  7951=>"111000110",
  7952=>"000111000",
  7953=>"000010110",
  7954=>"110000110",
  7955=>"011000000",
  7956=>"111101001",
  7957=>"111000100",
  7958=>"100110001",
  7959=>"101111110",
  7960=>"101000001",
  7961=>"011010101",
  7962=>"111000000",
  7963=>"001001011",
  7964=>"101000000",
  7965=>"110111000",
  7966=>"111101111",
  7967=>"111110000",
  7968=>"101111010",
  7969=>"001100100",
  7970=>"100111111",
  7971=>"110000000",
  7972=>"111001001",
  7973=>"100000011",
  7974=>"100000000",
  7975=>"001100110",
  7976=>"000111111",
  7977=>"110110110",
  7978=>"000000111",
  7979=>"000000010",
  7980=>"001001001",
  7981=>"100101101",
  7982=>"110101111",
  7983=>"111001110",
  7984=>"111000000",
  7985=>"111001001",
  7986=>"111111110",
  7987=>"001011111",
  7988=>"011001011",
  7989=>"110000111",
  7990=>"110001011",
  7991=>"111101000",
  7992=>"000000111",
  7993=>"000000000",
  7994=>"100001000",
  7995=>"111111111",
  7996=>"100111001",
  7997=>"110000000",
  7998=>"000000000",
  7999=>"010000000",
  8000=>"001010111",
  8001=>"101000001",
  8002=>"111011101",
  8003=>"100000001",
  8004=>"111000000",
  8005=>"111111101",
  8006=>"001000011",
  8007=>"101111101",
  8008=>"010011000",
  8009=>"000001000",
  8010=>"001000000",
  8011=>"001101111",
  8012=>"001000001",
  8013=>"011000101",
  8014=>"111100100",
  8015=>"111101100",
  8016=>"111000000",
  8017=>"100111010",
  8018=>"010010101",
  8019=>"001001000",
  8020=>"001000000",
  8021=>"110100000",
  8022=>"111110000",
  8023=>"001010011",
  8024=>"111111001",
  8025=>"101000000",
  8026=>"111001000",
  8027=>"000010100",
  8028=>"000000000",
  8029=>"011001000",
  8030=>"010010111",
  8031=>"010001000",
  8032=>"000000000",
  8033=>"001000000",
  8034=>"000000111",
  8035=>"100110001",
  8036=>"111000000",
  8037=>"000111000",
  8038=>"000000111",
  8039=>"010111000",
  8040=>"101010111",
  8041=>"000010000",
  8042=>"000110110",
  8043=>"011110000",
  8044=>"111111100",
  8045=>"001001101",
  8046=>"001101110",
  8047=>"000000000",
  8048=>"011011010",
  8049=>"000111111",
  8050=>"001100110",
  8051=>"000000100",
  8052=>"110100000",
  8053=>"011000101",
  8054=>"000000111",
  8055=>"000100101",
  8056=>"101001101",
  8057=>"010000010",
  8058=>"001000000",
  8059=>"010000000",
  8060=>"000001000",
  8061=>"101101011",
  8062=>"000110010",
  8063=>"101001000",
  8064=>"100000111",
  8065=>"111010010",
  8066=>"001001001",
  8067=>"110111000",
  8068=>"000001000",
  8069=>"000001110",
  8070=>"011000000",
  8071=>"001001101",
  8072=>"010101100",
  8073=>"110101101",
  8074=>"101101111",
  8075=>"110101111",
  8076=>"000010111",
  8077=>"000100011",
  8078=>"000000110",
  8079=>"000000101",
  8080=>"111101000",
  8081=>"101011000",
  8082=>"001001111",
  8083=>"111111001",
  8084=>"000000100",
  8085=>"000000111",
  8086=>"010011001",
  8087=>"001011000",
  8088=>"000100101",
  8089=>"000010001",
  8090=>"000000111",
  8091=>"100001111",
  8092=>"011011000",
  8093=>"101101111",
  8094=>"100000000",
  8095=>"000000010",
  8096=>"011011111",
  8097=>"101111111",
  8098=>"111111001",
  8099=>"101000000",
  8100=>"010101111",
  8101=>"001001001",
  8102=>"011010000",
  8103=>"110101000",
  8104=>"111000111",
  8105=>"110000000",
  8106=>"100100111",
  8107=>"001000111",
  8108=>"110100101",
  8109=>"000000001",
  8110=>"101111001",
  8111=>"000110111",
  8112=>"000100111",
  8113=>"111011100",
  8114=>"111101000",
  8115=>"000000000",
  8116=>"110010000",
  8117=>"011111111",
  8118=>"011111111",
  8119=>"000000100",
  8120=>"011101100",
  8121=>"010000000",
  8122=>"111000000",
  8123=>"011001000",
  8124=>"001111000",
  8125=>"100110111",
  8126=>"000000011",
  8127=>"101111110",
  8128=>"000000000",
  8129=>"000101111",
  8130=>"000000010",
  8131=>"010000100",
  8132=>"001000001",
  8133=>"100011110",
  8134=>"101111111",
  8135=>"000000011",
  8136=>"010101111",
  8137=>"111001101",
  8138=>"010111111",
  8139=>"000000101",
  8140=>"010000001",
  8141=>"000000001",
  8142=>"101101110",
  8143=>"110111110",
  8144=>"000000110",
  8145=>"110110100",
  8146=>"111001111",
  8147=>"011111000",
  8148=>"000000001",
  8149=>"111100000",
  8150=>"111000000",
  8151=>"001111000",
  8152=>"111110010",
  8153=>"010000000",
  8154=>"000101111",
  8155=>"001000111",
  8156=>"111011000",
  8157=>"000000111",
  8158=>"010111111",
  8159=>"111100111",
  8160=>"111011101",
  8161=>"101110000",
  8162=>"101110010",
  8163=>"011000001",
  8164=>"000011111",
  8165=>"000100101",
  8166=>"110111111",
  8167=>"011111000",
  8168=>"000110110",
  8169=>"101000000",
  8170=>"101001000",
  8171=>"000000111",
  8172=>"000000001",
  8173=>"011000000",
  8174=>"000000000",
  8175=>"111000000",
  8176=>"011000000",
  8177=>"011100111",
  8178=>"100010010",
  8179=>"111101000",
  8180=>"110110001",
  8181=>"110100101",
  8182=>"001101011",
  8183=>"000000111",
  8184=>"000111111",
  8185=>"111110000",
  8186=>"110000000",
  8187=>"010000001",
  8188=>"000000111",
  8189=>"000100111",
  8190=>"000100100",
  8191=>"101001100",
  8192=>"101001000",
  8193=>"110111001",
  8194=>"111011001",
  8195=>"101100110",
  8196=>"111011011",
  8197=>"111000000",
  8198=>"000110111",
  8199=>"010110010",
  8200=>"001000100",
  8201=>"110001001",
  8202=>"011000100",
  8203=>"000010100",
  8204=>"111001000",
  8205=>"000001100",
  8206=>"111001001",
  8207=>"100101101",
  8208=>"110100001",
  8209=>"111000111",
  8210=>"110000000",
  8211=>"110000000",
  8212=>"011110000",
  8213=>"111011000",
  8214=>"001101111",
  8215=>"111001000",
  8216=>"111011000",
  8217=>"011010011",
  8218=>"111001011",
  8219=>"100000001",
  8220=>"000001001",
  8221=>"000101101",
  8222=>"001011111",
  8223=>"000000111",
  8224=>"110111100",
  8225=>"001001001",
  8226=>"000000101",
  8227=>"111001000",
  8228=>"000110010",
  8229=>"001001001",
  8230=>"100011001",
  8231=>"000100110",
  8232=>"001111110",
  8233=>"000111011",
  8234=>"110111111",
  8235=>"111000000",
  8236=>"100001001",
  8237=>"100111111",
  8238=>"000001100",
  8239=>"000100100",
  8240=>"001000110",
  8241=>"101000111",
  8242=>"001010010",
  8243=>"001111111",
  8244=>"000110100",
  8245=>"101111100",
  8246=>"111001001",
  8247=>"101000001",
  8248=>"100110110",
  8249=>"111011011",
  8250=>"111111100",
  8251=>"011011011",
  8252=>"111000001",
  8253=>"111011001",
  8254=>"101001000",
  8255=>"010011001",
  8256=>"111101001",
  8257=>"101011011",
  8258=>"001000101",
  8259=>"110000011",
  8260=>"111011111",
  8261=>"011010000",
  8262=>"000100010",
  8263=>"000110111",
  8264=>"100100011",
  8265=>"110000000",
  8266=>"110010010",
  8267=>"111001101",
  8268=>"110001001",
  8269=>"010101111",
  8270=>"111001111",
  8271=>"110110110",
  8272=>"111000000",
  8273=>"100111001",
  8274=>"010100100",
  8275=>"000110100",
  8276=>"001001000",
  8277=>"001100100",
  8278=>"000010101",
  8279=>"011001001",
  8280=>"011000111",
  8281=>"000000111",
  8282=>"111001001",
  8283=>"001011110",
  8284=>"001001001",
  8285=>"100000001",
  8286=>"000111111",
  8287=>"111100011",
  8288=>"111001011",
  8289=>"000001000",
  8290=>"110001001",
  8291=>"111101111",
  8292=>"111011110",
  8293=>"000110110",
  8294=>"010000000",
  8295=>"000110100",
  8296=>"111001101",
  8297=>"110000110",
  8298=>"000110000",
  8299=>"001011111",
  8300=>"001011000",
  8301=>"101101100",
  8302=>"000000000",
  8303=>"111000110",
  8304=>"000100101",
  8305=>"001000100",
  8306=>"110000001",
  8307=>"011110100",
  8308=>"111100000",
  8309=>"010011011",
  8310=>"111000011",
  8311=>"000100011",
  8312=>"000100000",
  8313=>"000000011",
  8314=>"011011100",
  8315=>"000000101",
  8316=>"111010001",
  8317=>"110101000",
  8318=>"000101101",
  8319=>"110001001",
  8320=>"000000000",
  8321=>"110010000",
  8322=>"000111111",
  8323=>"000100100",
  8324=>"000111110",
  8325=>"000110100",
  8326=>"001001101",
  8327=>"111001001",
  8328=>"101011111",
  8329=>"110010100",
  8330=>"001101111",
  8331=>"001111001",
  8332=>"001000001",
  8333=>"110110000",
  8334=>"100000000",
  8335=>"110000001",
  8336=>"010111111",
  8337=>"111011010",
  8338=>"111001001",
  8339=>"111111011",
  8340=>"111000001",
  8341=>"001001001",
  8342=>"111001001",
  8343=>"000100100",
  8344=>"100110010",
  8345=>"000110111",
  8346=>"101001111",
  8347=>"000100000",
  8348=>"110100000",
  8349=>"111000010",
  8350=>"000111111",
  8351=>"010001000",
  8352=>"011000000",
  8353=>"001111111",
  8354=>"000110000",
  8355=>"100001110",
  8356=>"111110110",
  8357=>"000000100",
  8358=>"000101100",
  8359=>"011001110",
  8360=>"001111001",
  8361=>"111110000",
  8362=>"111001000",
  8363=>"110000000",
  8364=>"000001000",
  8365=>"100001001",
  8366=>"111111011",
  8367=>"110000110",
  8368=>"100110110",
  8369=>"100000001",
  8370=>"001011111",
  8371=>"010000100",
  8372=>"001110110",
  8373=>"101101101",
  8374=>"001111111",
  8375=>"100010000",
  8376=>"100000001",
  8377=>"100101001",
  8378=>"000110101",
  8379=>"000000011",
  8380=>"101000100",
  8381=>"110001001",
  8382=>"011000011",
  8383=>"100110111",
  8384=>"110100100",
  8385=>"111001000",
  8386=>"101000111",
  8387=>"000110110",
  8388=>"001100100",
  8389=>"000110001",
  8390=>"001100111",
  8391=>"001011011",
  8392=>"000000000",
  8393=>"010001011",
  8394=>"101111110",
  8395=>"010000100",
  8396=>"100010110",
  8397=>"111111001",
  8398=>"010001000",
  8399=>"111001110",
  8400=>"111000001",
  8401=>"001010010",
  8402=>"011011010",
  8403=>"001110111",
  8404=>"000000100",
  8405=>"111001000",
  8406=>"111011001",
  8407=>"100110100",
  8408=>"000100110",
  8409=>"110001000",
  8410=>"100100000",
  8411=>"100001000",
  8412=>"010010001",
  8413=>"100110110",
  8414=>"000111111",
  8415=>"001001111",
  8416=>"111110010",
  8417=>"101111011",
  8418=>"000100110",
  8419=>"011100100",
  8420=>"111001000",
  8421=>"001110011",
  8422=>"110111111",
  8423=>"100000000",
  8424=>"001110110",
  8425=>"111001101",
  8426=>"111011010",
  8427=>"000000001",
  8428=>"011110000",
  8429=>"001100000",
  8430=>"000000000",
  8431=>"101110010",
  8432=>"010001000",
  8433=>"000001011",
  8434=>"000011011",
  8435=>"000100100",
  8436=>"111011111",
  8437=>"111001001",
  8438=>"011001001",
  8439=>"000110110",
  8440=>"111001001",
  8441=>"100100100",
  8442=>"001011001",
  8443=>"100001011",
  8444=>"000110111",
  8445=>"001110110",
  8446=>"000010011",
  8447=>"010110010",
  8448=>"011011000",
  8449=>"101101100",
  8450=>"100000101",
  8451=>"000000100",
  8452=>"100111001",
  8453=>"110101101",
  8454=>"010111111",
  8455=>"010000001",
  8456=>"000101111",
  8457=>"000000101",
  8458=>"010110110",
  8459=>"010010000",
  8460=>"101000110",
  8461=>"111011101",
  8462=>"100100010",
  8463=>"111000000",
  8464=>"101101110",
  8465=>"000000111",
  8466=>"101100110",
  8467=>"000001000",
  8468=>"111110100",
  8469=>"001101111",
  8470=>"101000100",
  8471=>"001111000",
  8472=>"000001101",
  8473=>"011001000",
  8474=>"011011011",
  8475=>"000000101",
  8476=>"100101100",
  8477=>"111111011",
  8478=>"000101101",
  8479=>"000100000",
  8480=>"000000000",
  8481=>"111001110",
  8482=>"100111101",
  8483=>"000000100",
  8484=>"101000001",
  8485=>"011001011",
  8486=>"000010110",
  8487=>"111010000",
  8488=>"111111010",
  8489=>"011000011",
  8490=>"101101000",
  8491=>"001000000",
  8492=>"000100000",
  8493=>"000110111",
  8494=>"111111101",
  8495=>"101111111",
  8496=>"000001111",
  8497=>"100101111",
  8498=>"011110101",
  8499=>"101101111",
  8500=>"111010000",
  8501=>"100100000",
  8502=>"001001001",
  8503=>"000010011",
  8504=>"111100110",
  8505=>"000000000",
  8506=>"001111111",
  8507=>"000000100",
  8508=>"110001000",
  8509=>"111111000",
  8510=>"000000000",
  8511=>"011011101",
  8512=>"000110111",
  8513=>"001111111",
  8514=>"010000111",
  8515=>"110111011",
  8516=>"111101110",
  8517=>"100110111",
  8518=>"111100000",
  8519=>"000000110",
  8520=>"001100000",
  8521=>"010011000",
  8522=>"000000000",
  8523=>"110110011",
  8524=>"100100101",
  8525=>"100000010",
  8526=>"000100111",
  8527=>"000000111",
  8528=>"000001010",
  8529=>"111111111",
  8530=>"010010100",
  8531=>"101001000",
  8532=>"000010100",
  8533=>"110000100",
  8534=>"111111110",
  8535=>"000000001",
  8536=>"100111000",
  8537=>"000001000",
  8538=>"100000001",
  8539=>"100001100",
  8540=>"111101101",
  8541=>"001000000",
  8542=>"111000000",
  8543=>"011110111",
  8544=>"000000111",
  8545=>"111111000",
  8546=>"000000101",
  8547=>"110101000",
  8548=>"110000010",
  8549=>"101011110",
  8550=>"110111000",
  8551=>"001100010",
  8552=>"111000000",
  8553=>"110111101",
  8554=>"000011100",
  8555=>"110111001",
  8556=>"010000111",
  8557=>"110111101",
  8558=>"110000100",
  8559=>"100001010",
  8560=>"100110011",
  8561=>"000110111",
  8562=>"100100000",
  8563=>"001000000",
  8564=>"011010000",
  8565=>"000000000",
  8566=>"101010010",
  8567=>"010111000",
  8568=>"000000000",
  8569=>"100111011",
  8570=>"100010111",
  8571=>"000100001",
  8572=>"000011110",
  8573=>"000000000",
  8574=>"000000101",
  8575=>"110110000",
  8576=>"111111111",
  8577=>"101101111",
  8578=>"110000000",
  8579=>"100111010",
  8580=>"001101001",
  8581=>"111010001",
  8582=>"100101101",
  8583=>"000000000",
  8584=>"001010010",
  8585=>"110000000",
  8586=>"011011010",
  8587=>"000000111",
  8588=>"111111010",
  8589=>"000001011",
  8590=>"000101011",
  8591=>"000000000",
  8592=>"111111011",
  8593=>"100111010",
  8594=>"010010000",
  8595=>"111111111",
  8596=>"101110011",
  8597=>"001101101",
  8598=>"110011010",
  8599=>"001111111",
  8600=>"010001111",
  8601=>"000001000",
  8602=>"111110100",
  8603=>"101101101",
  8604=>"101100111",
  8605=>"001000000",
  8606=>"101101101",
  8607=>"000000000",
  8608=>"001000001",
  8609=>"001111111",
  8610=>"111010011",
  8611=>"000100111",
  8612=>"101111111",
  8613=>"110110011",
  8614=>"000100100",
  8615=>"000000000",
  8616=>"000000101",
  8617=>"100100111",
  8618=>"101101111",
  8619=>"000100010",
  8620=>"000111011",
  8621=>"000000100",
  8622=>"110111000",
  8623=>"011101010",
  8624=>"101101000",
  8625=>"101101001",
  8626=>"001111110",
  8627=>"000010010",
  8628=>"001011011",
  8629=>"100111000",
  8630=>"000111011",
  8631=>"110010111",
  8632=>"101100000",
  8633=>"111011010",
  8634=>"110011100",
  8635=>"000011110",
  8636=>"110100010",
  8637=>"101001000",
  8638=>"000000000",
  8639=>"000110101",
  8640=>"000101000",
  8641=>"111111011",
  8642=>"001000010",
  8643=>"101101101",
  8644=>"110010111",
  8645=>"101001111",
  8646=>"000101011",
  8647=>"001000000",
  8648=>"110010010",
  8649=>"111111111",
  8650=>"000111110",
  8651=>"000100110",
  8652=>"110111000",
  8653=>"101110001",
  8654=>"101111010",
  8655=>"101101101",
  8656=>"000000000",
  8657=>"111111110",
  8658=>"111110110",
  8659=>"010010111",
  8660=>"101001101",
  8661=>"100100110",
  8662=>"100000000",
  8663=>"110000110",
  8664=>"111000000",
  8665=>"010011111",
  8666=>"010010111",
  8667=>"101111101",
  8668=>"111001011",
  8669=>"000001111",
  8670=>"111111111",
  8671=>"010011110",
  8672=>"000010000",
  8673=>"100000100",
  8674=>"100111110",
  8675=>"001000011",
  8676=>"001101001",
  8677=>"110110010",
  8678=>"100000010",
  8679=>"011100010",
  8680=>"111110110",
  8681=>"000000000",
  8682=>"110011001",
  8683=>"000000111",
  8684=>"010010011",
  8685=>"110101100",
  8686=>"000000000",
  8687=>"011100100",
  8688=>"111110000",
  8689=>"100000101",
  8690=>"000000101",
  8691=>"101110010",
  8692=>"110001010",
  8693=>"001011000",
  8694=>"000000000",
  8695=>"000100000",
  8696=>"000000000",
  8697=>"000100100",
  8698=>"110010000",
  8699=>"101111100",
  8700=>"001101111",
  8701=>"111000000",
  8702=>"101100100",
  8703=>"001000000",
  8704=>"000001011",
  8705=>"100010011",
  8706=>"111001000",
  8707=>"111000000",
  8708=>"011010001",
  8709=>"111101000",
  8710=>"010101000",
  8711=>"000000010",
  8712=>"000000000",
  8713=>"111000000",
  8714=>"111101100",
  8715=>"001001111",
  8716=>"100000010",
  8717=>"000111111",
  8718=>"100100100",
  8719=>"100000101",
  8720=>"011000001",
  8721=>"111111000",
  8722=>"000000000",
  8723=>"100001000",
  8724=>"000111111",
  8725=>"000010000",
  8726=>"000010111",
  8727=>"000110110",
  8728=>"111001101",
  8729=>"100111110",
  8730=>"000110111",
  8731=>"000000001",
  8732=>"000001100",
  8733=>"001000000",
  8734=>"000000000",
  8735=>"001000010",
  8736=>"111100101",
  8737=>"101000001",
  8738=>"000010010",
  8739=>"101000000",
  8740=>"011110110",
  8741=>"010000010",
  8742=>"010010010",
  8743=>"000100100",
  8744=>"110110010",
  8745=>"010011111",
  8746=>"011001001",
  8747=>"000001000",
  8748=>"000111011",
  8749=>"111111110",
  8750=>"110110101",
  8751=>"001011001",
  8752=>"111000111",
  8753=>"000110111",
  8754=>"001001000",
  8755=>"111000011",
  8756=>"111101001",
  8757=>"110010010",
  8758=>"111110011",
  8759=>"000001001",
  8760=>"111000000",
  8761=>"001001101",
  8762=>"000111111",
  8763=>"000000110",
  8764=>"000011110",
  8765=>"010000011",
  8766=>"111001000",
  8767=>"100101000",
  8768=>"111000000",
  8769=>"111010001",
  8770=>"010111001",
  8771=>"000000001",
  8772=>"000000111",
  8773=>"101001001",
  8774=>"000001101",
  8775=>"111111110",
  8776=>"100000111",
  8777=>"110110111",
  8778=>"000000000",
  8779=>"001000001",
  8780=>"110001000",
  8781=>"011001111",
  8782=>"000000100",
  8783=>"000110111",
  8784=>"101111100",
  8785=>"111010000",
  8786=>"100110110",
  8787=>"001110011",
  8788=>"100000001",
  8789=>"111100011",
  8790=>"001011011",
  8791=>"001001000",
  8792=>"000101110",
  8793=>"000111111",
  8794=>"000111101",
  8795=>"000011010",
  8796=>"111001001",
  8797=>"000110000",
  8798=>"111010111",
  8799=>"010000101",
  8800=>"110111000",
  8801=>"000000111",
  8802=>"111001001",
  8803=>"000011011",
  8804=>"001001110",
  8805=>"010110110",
  8806=>"000010110",
  8807=>"111111001",
  8808=>"110111100",
  8809=>"010111000",
  8810=>"001000000",
  8811=>"000000111",
  8812=>"111111010",
  8813=>"111111001",
  8814=>"000000001",
  8815=>"000000111",
  8816=>"000111011",
  8817=>"010111110",
  8818=>"111111111",
  8819=>"111101000",
  8820=>"000001010",
  8821=>"000000000",
  8822=>"011000000",
  8823=>"011001000",
  8824=>"001111000",
  8825=>"000000110",
  8826=>"000111101",
  8827=>"000001010",
  8828=>"011000010",
  8829=>"000001110",
  8830=>"010001111",
  8831=>"001101000",
  8832=>"000010010",
  8833=>"111110000",
  8834=>"111001000",
  8835=>"001001110",
  8836=>"101000000",
  8837=>"001000110",
  8838=>"100110100",
  8839=>"000000010",
  8840=>"001010111",
  8841=>"000000111",
  8842=>"011111000",
  8843=>"000111111",
  8844=>"111001001",
  8845=>"111101111",
  8846=>"001111100",
  8847=>"000000000",
  8848=>"011111000",
  8849=>"010111111",
  8850=>"111101101",
  8851=>"000110110",
  8852=>"001100110",
  8853=>"111000000",
  8854=>"111100100",
  8855=>"000100100",
  8856=>"000000000",
  8857=>"000000000",
  8858=>"110100000",
  8859=>"101010010",
  8860=>"110001000",
  8861=>"111101101",
  8862=>"111001000",
  8863=>"000000010",
  8864=>"000011110",
  8865=>"111101001",
  8866=>"000000110",
  8867=>"101110110",
  8868=>"000000100",
  8869=>"000111110",
  8870=>"001001001",
  8871=>"000111101",
  8872=>"111111000",
  8873=>"010011000",
  8874=>"111100001",
  8875=>"000001001",
  8876=>"001110110",
  8877=>"010100101",
  8878=>"100110100",
  8879=>"011110110",
  8880=>"000010110",
  8881=>"000101011",
  8882=>"000001100",
  8883=>"000010011",
  8884=>"000110111",
  8885=>"101110100",
  8886=>"100100111",
  8887=>"001111011",
  8888=>"000000111",
  8889=>"000000110",
  8890=>"000001000",
  8891=>"100010010",
  8892=>"000000001",
  8893=>"111111001",
  8894=>"011001000",
  8895=>"111011001",
  8896=>"000010110",
  8897=>"010000000",
  8898=>"110110111",
  8899=>"000100110",
  8900=>"000000000",
  8901=>"101111011",
  8902=>"111110111",
  8903=>"000111001",
  8904=>"000100101",
  8905=>"001000110",
  8906=>"001111110",
  8907=>"111110000",
  8908=>"000001111",
  8909=>"100000010",
  8910=>"000101101",
  8911=>"111111000",
  8912=>"011111110",
  8913=>"001001111",
  8914=>"010000110",
  8915=>"001000011",
  8916=>"000000111",
  8917=>"101101101",
  8918=>"101001001",
  8919=>"110111001",
  8920=>"000110110",
  8921=>"010000000",
  8922=>"000110110",
  8923=>"111101000",
  8924=>"000100111",
  8925=>"000111001",
  8926=>"010000011",
  8927=>"000010000",
  8928=>"000110110",
  8929=>"101100011",
  8930=>"001111111",
  8931=>"011011011",
  8932=>"010111001",
  8933=>"110000011",
  8934=>"000000101",
  8935=>"000011101",
  8936=>"101111111",
  8937=>"111101001",
  8938=>"111001001",
  8939=>"111101001",
  8940=>"111010110",
  8941=>"001111000",
  8942=>"000000000",
  8943=>"000000110",
  8944=>"000001011",
  8945=>"101010000",
  8946=>"111000000",
  8947=>"000110110",
  8948=>"111001011",
  8949=>"111111001",
  8950=>"001001000",
  8951=>"010101000",
  8952=>"000000110",
  8953=>"100110111",
  8954=>"000000100",
  8955=>"000111111",
  8956=>"011010010",
  8957=>"000101101",
  8958=>"110100001",
  8959=>"010110110",
  8960=>"011011001",
  8961=>"010000111",
  8962=>"111101101",
  8963=>"000000010",
  8964=>"000001001",
  8965=>"111111110",
  8966=>"100110111",
  8967=>"000100111",
  8968=>"000000000",
  8969=>"001100010",
  8970=>"111100000",
  8971=>"101000000",
  8972=>"000010010",
  8973=>"111000100",
  8974=>"101001011",
  8975=>"000011100",
  8976=>"100100010",
  8977=>"100001011",
  8978=>"111101000",
  8979=>"111010000",
  8980=>"101101101",
  8981=>"111010000",
  8982=>"001101111",
  8983=>"000000111",
  8984=>"111111011",
  8985=>"000110110",
  8986=>"010111111",
  8987=>"000000001",
  8988=>"011011000",
  8989=>"111000000",
  8990=>"001101101",
  8991=>"000111000",
  8992=>"000010010",
  8993=>"010010011",
  8994=>"100000000",
  8995=>"000000000",
  8996=>"011101001",
  8997=>"110110111",
  8998=>"000000011",
  8999=>"000000101",
  9000=>"000000111",
  9001=>"000001011",
  9002=>"000101000",
  9003=>"000111111",
  9004=>"001000001",
  9005=>"101110000",
  9006=>"111111111",
  9007=>"001101010",
  9008=>"110111000",
  9009=>"010011011",
  9010=>"000111101",
  9011=>"111110111",
  9012=>"111111001",
  9013=>"010000000",
  9014=>"100001000",
  9015=>"100110010",
  9016=>"111010111",
  9017=>"111000000",
  9018=>"000000000",
  9019=>"000100010",
  9020=>"000110100",
  9021=>"111111000",
  9022=>"111101101",
  9023=>"110111001",
  9024=>"001101101",
  9025=>"100010111",
  9026=>"111100111",
  9027=>"111101000",
  9028=>"010010000",
  9029=>"100100000",
  9030=>"111101110",
  9031=>"000001010",
  9032=>"010000000",
  9033=>"010010000",
  9034=>"000000000",
  9035=>"010000000",
  9036=>"111101100",
  9037=>"001111101",
  9038=>"000111110",
  9039=>"110111000",
  9040=>"111000100",
  9041=>"111111110",
  9042=>"111011000",
  9043=>"010011100",
  9044=>"101101101",
  9045=>"001001110",
  9046=>"011011011",
  9047=>"111000010",
  9048=>"001110011",
  9049=>"000011011",
  9050=>"011001101",
  9051=>"000100100",
  9052=>"000110000",
  9053=>"010001001",
  9054=>"111101111",
  9055=>"011100001",
  9056=>"000101111",
  9057=>"100000010",
  9058=>"001000111",
  9059=>"100101101",
  9060=>"000000000",
  9061=>"100100100",
  9062=>"000000010",
  9063=>"011111100",
  9064=>"111011011",
  9065=>"111100111",
  9066=>"010101101",
  9067=>"001010000",
  9068=>"000011111",
  9069=>"101101111",
  9070=>"000110111",
  9071=>"101101100",
  9072=>"001001000",
  9073=>"000000010",
  9074=>"000000000",
  9075=>"000111110",
  9076=>"011010000",
  9077=>"101000000",
  9078=>"001101101",
  9079=>"000100101",
  9080=>"111000111",
  9081=>"000110111",
  9082=>"100000110",
  9083=>"100111000",
  9084=>"100100110",
  9085=>"011110100",
  9086=>"011111100",
  9087=>"101101001",
  9088=>"111000101",
  9089=>"111101000",
  9090=>"011000000",
  9091=>"101111011",
  9092=>"011010000",
  9093=>"001000010",
  9094=>"010011110",
  9095=>"000001011",
  9096=>"000110100",
  9097=>"110110011",
  9098=>"100100101",
  9099=>"011010000",
  9100=>"111101000",
  9101=>"111111111",
  9102=>"010011000",
  9103=>"100000100",
  9104=>"011101101",
  9105=>"000000000",
  9106=>"000000111",
  9107=>"111101111",
  9108=>"011001111",
  9109=>"000100101",
  9110=>"111011101",
  9111=>"001110111",
  9112=>"111001000",
  9113=>"010000001",
  9114=>"111000000",
  9115=>"110000001",
  9116=>"010100001",
  9117=>"101001000",
  9118=>"101111000",
  9119=>"000000010",
  9120=>"000110111",
  9121=>"101001001",
  9122=>"000011101",
  9123=>"000011111",
  9124=>"000111011",
  9125=>"000100101",
  9126=>"000000000",
  9127=>"000000000",
  9128=>"011111101",
  9129=>"000111111",
  9130=>"001011001",
  9131=>"111001101",
  9132=>"001111111",
  9133=>"111000111",
  9134=>"110101100",
  9135=>"000111111",
  9136=>"010111101",
  9137=>"000011111",
  9138=>"110000111",
  9139=>"001000100",
  9140=>"100011000",
  9141=>"101111101",
  9142=>"000011000",
  9143=>"000000001",
  9144=>"000011011",
  9145=>"010011111",
  9146=>"000000001",
  9147=>"010010010",
  9148=>"100010000",
  9149=>"010111110",
  9150=>"100111110",
  9151=>"000011000",
  9152=>"111000000",
  9153=>"000101111",
  9154=>"010010000",
  9155=>"110000000",
  9156=>"000011101",
  9157=>"010011101",
  9158=>"000000110",
  9159=>"101111111",
  9160=>"000010010",
  9161=>"001000000",
  9162=>"111111110",
  9163=>"111000000",
  9164=>"001100101",
  9165=>"001001110",
  9166=>"101101101",
  9167=>"000010010",
  9168=>"111100000",
  9169=>"101111111",
  9170=>"000010111",
  9171=>"011010000",
  9172=>"011101011",
  9173=>"000100111",
  9174=>"000000000",
  9175=>"000111111",
  9176=>"111000101",
  9177=>"111110010",
  9178=>"000000111",
  9179=>"111100110",
  9180=>"100101000",
  9181=>"010000011",
  9182=>"101101010",
  9183=>"001101111",
  9184=>"110000010",
  9185=>"111111000",
  9186=>"111000000",
  9187=>"010011001",
  9188=>"000001001",
  9189=>"100011010",
  9190=>"110110110",
  9191=>"001111011",
  9192=>"111000101",
  9193=>"000010000",
  9194=>"111001001",
  9195=>"000010010",
  9196=>"000000000",
  9197=>"110000000",
  9198=>"110010110",
  9199=>"001000000",
  9200=>"000010000",
  9201=>"000100001",
  9202=>"000111011",
  9203=>"000110001",
  9204=>"010110111",
  9205=>"011111111",
  9206=>"000010000",
  9207=>"000000101",
  9208=>"000111000",
  9209=>"110010001",
  9210=>"011101100",
  9211=>"100101010",
  9212=>"011101101",
  9213=>"100100000",
  9214=>"111100100",
  9215=>"110100111",
  9216=>"001000100",
  9217=>"100101100",
  9218=>"000000111",
  9219=>"000101111",
  9220=>"011110110",
  9221=>"000001111",
  9222=>"011111101",
  9223=>"101010111",
  9224=>"000101010",
  9225=>"000101010",
  9226=>"110100100",
  9227=>"000011011",
  9228=>"010001001",
  9229=>"000000101",
  9230=>"100001011",
  9231=>"011111100",
  9232=>"000000011",
  9233=>"000101101",
  9234=>"000000001",
  9235=>"100000100",
  9236=>"011101111",
  9237=>"110001010",
  9238=>"101101111",
  9239=>"010110111",
  9240=>"010000100",
  9241=>"111101001",
  9242=>"001101010",
  9243=>"101100011",
  9244=>"110100100",
  9245=>"000000000",
  9246=>"001000000",
  9247=>"000101100",
  9248=>"110000001",
  9249=>"010101111",
  9250=>"010010010",
  9251=>"111100101",
  9252=>"101100000",
  9253=>"111010111",
  9254=>"000111000",
  9255=>"011111111",
  9256=>"100111111",
  9257=>"111111000",
  9258=>"101101111",
  9259=>"111000000",
  9260=>"101100011",
  9261=>"101111000",
  9262=>"001110110",
  9263=>"000011101",
  9264=>"000010010",
  9265=>"101101000",
  9266=>"001000000",
  9267=>"001010010",
  9268=>"111101001",
  9269=>"001111111",
  9270=>"001001001",
  9271=>"010010111",
  9272=>"111111010",
  9273=>"000000100",
  9274=>"000000101",
  9275=>"101101111",
  9276=>"011000000",
  9277=>"111111111",
  9278=>"000000000",
  9279=>"001000100",
  9280=>"100111101",
  9281=>"110000001",
  9282=>"101100100",
  9283=>"100100100",
  9284=>"010000000",
  9285=>"000000000",
  9286=>"111110101",
  9287=>"000101111",
  9288=>"000000001",
  9289=>"101010010",
  9290=>"000000000",
  9291=>"101000110",
  9292=>"111001000",
  9293=>"001000000",
  9294=>"110011001",
  9295=>"110111111",
  9296=>"111000110",
  9297=>"000111111",
  9298=>"000000111",
  9299=>"100100100",
  9300=>"101111011",
  9301=>"100101000",
  9302=>"101100001",
  9303=>"100100100",
  9304=>"110010011",
  9305=>"001001001",
  9306=>"000010011",
  9307=>"010011010",
  9308=>"111000000",
  9309=>"000000101",
  9310=>"100001110",
  9311=>"001001001",
  9312=>"011011000",
  9313=>"010010011",
  9314=>"100100001",
  9315=>"010111110",
  9316=>"000001100",
  9317=>"101001000",
  9318=>"100111111",
  9319=>"101100111",
  9320=>"010001000",
  9321=>"111101101",
  9322=>"111111111",
  9323=>"000000011",
  9324=>"010001010",
  9325=>"000011110",
  9326=>"111011011",
  9327=>"001000011",
  9328=>"000000001",
  9329=>"111111111",
  9330=>"100100100",
  9331=>"111011000",
  9332=>"111101000",
  9333=>"010000000",
  9334=>"101010110",
  9335=>"000010000",
  9336=>"000000000",
  9337=>"101001101",
  9338=>"110010110",
  9339=>"010000111",
  9340=>"011110100",
  9341=>"001000001",
  9342=>"111000000",
  9343=>"000000110",
  9344=>"110000101",
  9345=>"000000011",
  9346=>"111010110",
  9347=>"111011110",
  9348=>"100000001",
  9349=>"111010010",
  9350=>"111110110",
  9351=>"110010000",
  9352=>"000001011",
  9353=>"100110010",
  9354=>"100010001",
  9355=>"011101110",
  9356=>"010111100",
  9357=>"110010000",
  9358=>"101101100",
  9359=>"001000010",
  9360=>"000100100",
  9361=>"111111111",
  9362=>"010010100",
  9363=>"110110110",
  9364=>"010011111",
  9365=>"101101101",
  9366=>"101101111",
  9367=>"001001001",
  9368=>"111111011",
  9369=>"011000001",
  9370=>"001011000",
  9371=>"000101001",
  9372=>"011111011",
  9373=>"011010010",
  9374=>"111101111",
  9375=>"111111011",
  9376=>"001100100",
  9377=>"001000000",
  9378=>"100001101",
  9379=>"111010111",
  9380=>"101011100",
  9381=>"011010000",
  9382=>"001110111",
  9383=>"110100100",
  9384=>"000111111",
  9385=>"111111111",
  9386=>"000000100",
  9387=>"101101101",
  9388=>"000100110",
  9389=>"000000001",
  9390=>"011011001",
  9391=>"010011010",
  9392=>"010000110",
  9393=>"011010100",
  9394=>"100101100",
  9395=>"111100100",
  9396=>"010011011",
  9397=>"100111010",
  9398=>"000010001",
  9399=>"100000001",
  9400=>"000000000",
  9401=>"001011000",
  9402=>"111010111",
  9403=>"011101100",
  9404=>"000000000",
  9405=>"111111000",
  9406=>"110100011",
  9407=>"100010000",
  9408=>"000101101",
  9409=>"010010010",
  9410=>"000101111",
  9411=>"100101110",
  9412=>"111101100",
  9413=>"110111011",
  9414=>"011011111",
  9415=>"010100101",
  9416=>"101100101",
  9417=>"000011010",
  9418=>"010101101",
  9419=>"001000001",
  9420=>"011101001",
  9421=>"110011001",
  9422=>"111100100",
  9423=>"001101111",
  9424=>"010111111",
  9425=>"110111100",
  9426=>"001010011",
  9427=>"011010010",
  9428=>"111101101",
  9429=>"110010111",
  9430=>"111101101",
  9431=>"001011001",
  9432=>"010010000",
  9433=>"000101111",
  9434=>"111001011",
  9435=>"011010010",
  9436=>"101101001",
  9437=>"101000000",
  9438=>"111000010",
  9439=>"000000010",
  9440=>"001100000",
  9441=>"000000010",
  9442=>"100110111",
  9443=>"011011110",
  9444=>"000000000",
  9445=>"010111110",
  9446=>"011000000",
  9447=>"100100000",
  9448=>"000000000",
  9449=>"111000000",
  9450=>"011011001",
  9451=>"001110100",
  9452=>"011001000",
  9453=>"011001001",
  9454=>"000000110",
  9455=>"000000011",
  9456=>"011000000",
  9457=>"101110100",
  9458=>"001010000",
  9459=>"100100000",
  9460=>"110101000",
  9461=>"111110110",
  9462=>"100000010",
  9463=>"101001011",
  9464=>"111000000",
  9465=>"101010000",
  9466=>"111100000",
  9467=>"001101101",
  9468=>"101101000",
  9469=>"001000101",
  9470=>"111111011",
  9471=>"110100110",
  9472=>"111100101",
  9473=>"000111000",
  9474=>"000001111",
  9475=>"101110110",
  9476=>"001001000",
  9477=>"111011000",
  9478=>"100001111",
  9479=>"110110000",
  9480=>"000101101",
  9481=>"000111000",
  9482=>"110111111",
  9483=>"001101111",
  9484=>"101111011",
  9485=>"000000010",
  9486=>"101111001",
  9487=>"000111110",
  9488=>"100001111",
  9489=>"001001111",
  9490=>"000001111",
  9491=>"100000010",
  9492=>"111001111",
  9493=>"010110100",
  9494=>"011000001",
  9495=>"111010000",
  9496=>"101000111",
  9497=>"011001111",
  9498=>"100100111",
  9499=>"000000000",
  9500=>"011110111",
  9501=>"110111111",
  9502=>"101001011",
  9503=>"000111111",
  9504=>"001010110",
  9505=>"000000001",
  9506=>"000110111",
  9507=>"110110000",
  9508=>"001000100",
  9509=>"010101111",
  9510=>"010111000",
  9511=>"011111000",
  9512=>"000101111",
  9513=>"111110000",
  9514=>"010000000",
  9515=>"000000111",
  9516=>"001001011",
  9517=>"000111111",
  9518=>"001111010",
  9519=>"100001101",
  9520=>"000000101",
  9521=>"111011111",
  9522=>"000000101",
  9523=>"001101111",
  9524=>"001000000",
  9525=>"111001011",
  9526=>"110010011",
  9527=>"010000000",
  9528=>"000000110",
  9529=>"101111101",
  9530=>"000101010",
  9531=>"100000111",
  9532=>"010001111",
  9533=>"111111000",
  9534=>"000000111",
  9535=>"111011100",
  9536=>"011111101",
  9537=>"101111010",
  9538=>"111111100",
  9539=>"011100000",
  9540=>"010011011",
  9541=>"010010000",
  9542=>"000101111",
  9543=>"110101001",
  9544=>"101111100",
  9545=>"101111111",
  9546=>"111000000",
  9547=>"000000111",
  9548=>"110010000",
  9549=>"100110000",
  9550=>"001110100",
  9551=>"101011111",
  9552=>"111000001",
  9553=>"011000000",
  9554=>"000011101",
  9555=>"001001000",
  9556=>"000001001",
  9557=>"101111111",
  9558=>"001000000",
  9559=>"001001111",
  9560=>"111111111",
  9561=>"000001011",
  9562=>"011111110",
  9563=>"000000101",
  9564=>"111000000",
  9565=>"000001011",
  9566=>"000001101",
  9567=>"001000100",
  9568=>"111110000",
  9569=>"010111010",
  9570=>"111011011",
  9571=>"001111001",
  9572=>"100100000",
  9573=>"100000000",
  9574=>"110110110",
  9575=>"001111110",
  9576=>"011101001",
  9577=>"110000000",
  9578=>"001000000",
  9579=>"101101000",
  9580=>"110111011",
  9581=>"000111001",
  9582=>"101111010",
  9583=>"010011111",
  9584=>"000011000",
  9585=>"000000110",
  9586=>"000100110",
  9587=>"111010000",
  9588=>"000001110",
  9589=>"000000000",
  9590=>"000000111",
  9591=>"001111010",
  9592=>"000000000",
  9593=>"010000000",
  9594=>"000000001",
  9595=>"101001011",
  9596=>"001011110",
  9597=>"100100100",
  9598=>"000011111",
  9599=>"111001011",
  9600=>"110010000",
  9601=>"100111111",
  9602=>"110100010",
  9603=>"010100101",
  9604=>"010111111",
  9605=>"101001000",
  9606=>"100100110",
  9607=>"100000000",
  9608=>"100101100",
  9609=>"000000011",
  9610=>"111100111",
  9611=>"111000000",
  9612=>"000000010",
  9613=>"011001000",
  9614=>"000000001",
  9615=>"000100001",
  9616=>"011111100",
  9617=>"111001000",
  9618=>"000010111",
  9619=>"110000000",
  9620=>"100101000",
  9621=>"001001000",
  9622=>"000010111",
  9623=>"011011000",
  9624=>"111111101",
  9625=>"000111111",
  9626=>"101110111",
  9627=>"111111000",
  9628=>"000000010",
  9629=>"111000000",
  9630=>"110000000",
  9631=>"110111000",
  9632=>"101111111",
  9633=>"000000100",
  9634=>"111110000",
  9635=>"101011111",
  9636=>"000110000",
  9637=>"010000011",
  9638=>"110010001",
  9639=>"110010000",
  9640=>"001100101",
  9641=>"000000000",
  9642=>"101111111",
  9643=>"111111010",
  9644=>"101010000",
  9645=>"011001111",
  9646=>"110011111",
  9647=>"001001011",
  9648=>"110000100",
  9649=>"001000001",
  9650=>"101111111",
  9651=>"000111111",
  9652=>"001100100",
  9653=>"000111111",
  9654=>"100111000",
  9655=>"000101110",
  9656=>"100100111",
  9657=>"111111011",
  9658=>"110101000",
  9659=>"101000000",
  9660=>"000101111",
  9661=>"111111111",
  9662=>"111110110",
  9663=>"000000010",
  9664=>"000000111",
  9665=>"000000111",
  9666=>"000111010",
  9667=>"000100100",
  9668=>"000000000",
  9669=>"100000000",
  9670=>"000110110",
  9671=>"110010000",
  9672=>"000000110",
  9673=>"000000000",
  9674=>"101000100",
  9675=>"001001111",
  9676=>"110100100",
  9677=>"001100110",
  9678=>"000010111",
  9679=>"111000010",
  9680=>"000010111",
  9681=>"110110010",
  9682=>"101010000",
  9683=>"010000001",
  9684=>"001011110",
  9685=>"100000000",
  9686=>"111111100",
  9687=>"000010100",
  9688=>"111100000",
  9689=>"100000111",
  9690=>"001001111",
  9691=>"101001000",
  9692=>"001100111",
  9693=>"001111111",
  9694=>"111110000",
  9695=>"000000101",
  9696=>"111001011",
  9697=>"000101101",
  9698=>"100111000",
  9699=>"011101010",
  9700=>"000000011",
  9701=>"000000000",
  9702=>"111110111",
  9703=>"111001100",
  9704=>"111111110",
  9705=>"001000110",
  9706=>"011011111",
  9707=>"000000001",
  9708=>"111000000",
  9709=>"111110010",
  9710=>"000000000",
  9711=>"001000010",
  9712=>"111010000",
  9713=>"001000000",
  9714=>"111000000",
  9715=>"000000000",
  9716=>"001001011",
  9717=>"100000011",
  9718=>"000000000",
  9719=>"100000000",
  9720=>"001000110",
  9721=>"101110101",
  9722=>"100100111",
  9723=>"010000000",
  9724=>"000000000",
  9725=>"101100111",
  9726=>"001001000",
  9727=>"111001000",
  9728=>"110010000",
  9729=>"110001110",
  9730=>"001001101",
  9731=>"110100100",
  9732=>"011010001",
  9733=>"110110000",
  9734=>"111001010",
  9735=>"100000111",
  9736=>"110110110",
  9737=>"000001111",
  9738=>"101001011",
  9739=>"110111001",
  9740=>"110100000",
  9741=>"100100110",
  9742=>"000100110",
  9743=>"000001000",
  9744=>"111000000",
  9745=>"001001111",
  9746=>"010000111",
  9747=>"011110110",
  9748=>"101111110",
  9749=>"110111011",
  9750=>"110110110",
  9751=>"000111111",
  9752=>"011001001",
  9753=>"111001001",
  9754=>"110110000",
  9755=>"011001001",
  9756=>"000001111",
  9757=>"000001111",
  9758=>"110110001",
  9759=>"000110110",
  9760=>"000000011",
  9761=>"110110111",
  9762=>"110001111",
  9763=>"100110110",
  9764=>"001001010",
  9765=>"011000000",
  9766=>"110110100",
  9767=>"110110110",
  9768=>"001001111",
  9769=>"100110100",
  9770=>"001001111",
  9771=>"100000011",
  9772=>"001011111",
  9773=>"001000001",
  9774=>"110110010",
  9775=>"000011111",
  9776=>"001000110",
  9777=>"111111011",
  9778=>"101001000",
  9779=>"001001011",
  9780=>"001001111",
  9781=>"111111101",
  9782=>"000110011",
  9783=>"000001001",
  9784=>"000110111",
  9785=>"001001001",
  9786=>"000101000",
  9787=>"000101111",
  9788=>"001010000",
  9789=>"110111000",
  9790=>"000000001",
  9791=>"110111000",
  9792=>"101111111",
  9793=>"110111011",
  9794=>"001000111",
  9795=>"100111000",
  9796=>"110110100",
  9797=>"000000101",
  9798=>"000000110",
  9799=>"010111001",
  9800=>"111010111",
  9801=>"000000000",
  9802=>"001001111",
  9803=>"100111111",
  9804=>"100110000",
  9805=>"111111100",
  9806=>"100100000",
  9807=>"000001111",
  9808=>"111111001",
  9809=>"100001000",
  9810=>"110110000",
  9811=>"110011101",
  9812=>"111001001",
  9813=>"111111111",
  9814=>"011000001",
  9815=>"001111111",
  9816=>"000110100",
  9817=>"001011111",
  9818=>"101001010",
  9819=>"110111000",
  9820=>"001000111",
  9821=>"000010010",
  9822=>"111001001",
  9823=>"111110000",
  9824=>"100110000",
  9825=>"110111111",
  9826=>"101000101",
  9827=>"011011111",
  9828=>"011001011",
  9829=>"110001000",
  9830=>"000001111",
  9831=>"000000110",
  9832=>"001100010",
  9833=>"110000000",
  9834=>"010000001",
  9835=>"110110001",
  9836=>"011001001",
  9837=>"001001001",
  9838=>"110110110",
  9839=>"101000000",
  9840=>"111111011",
  9841=>"000000111",
  9842=>"000000100",
  9843=>"110111000",
  9844=>"000000001",
  9845=>"001000000",
  9846=>"100000001",
  9847=>"110111100",
  9848=>"001001001",
  9849=>"110000000",
  9850=>"110100000",
  9851=>"100110110",
  9852=>"010000000",
  9853=>"111001000",
  9854=>"011011111",
  9855=>"110000000",
  9856=>"000001110",
  9857=>"110111000",
  9858=>"110110110",
  9859=>"110100000",
  9860=>"110110110",
  9861=>"001011111",
  9862=>"000010011",
  9863=>"000100000",
  9864=>"100101100",
  9865=>"000000100",
  9866=>"000000000",
  9867=>"110011000",
  9868=>"111001001",
  9869=>"010000100",
  9870=>"000000000",
  9871=>"000000111",
  9872=>"111101001",
  9873=>"011011111",
  9874=>"001001110",
  9875=>"110000000",
  9876=>"000000000",
  9877=>"100100111",
  9878=>"110110101",
  9879=>"110111000",
  9880=>"001000001",
  9881=>"001011110",
  9882=>"001001111",
  9883=>"100001101",
  9884=>"000010000",
  9885=>"000100100",
  9886=>"111111111",
  9887=>"000000000",
  9888=>"000011101",
  9889=>"000011011",
  9890=>"011001111",
  9891=>"000110001",
  9892=>"110110100",
  9893=>"111111101",
  9894=>"100110000",
  9895=>"001001111",
  9896=>"011000001",
  9897=>"101000000",
  9898=>"000000110",
  9899=>"010000110",
  9900=>"110000001",
  9901=>"110110000",
  9902=>"101111111",
  9903=>"100111100",
  9904=>"000000000",
  9905=>"110010011",
  9906=>"111001001",
  9907=>"111001000",
  9908=>"011110111",
  9909=>"000011111",
  9910=>"000011001",
  9911=>"000001000",
  9912=>"010110100",
  9913=>"010010001",
  9914=>"110110111",
  9915=>"111001001",
  9916=>"001011000",
  9917=>"111111010",
  9918=>"110110000",
  9919=>"000110110",
  9920=>"000000111",
  9921=>"001001001",
  9922=>"110110110",
  9923=>"000000000",
  9924=>"001001111",
  9925=>"111001110",
  9926=>"000101111",
  9927=>"000001111",
  9928=>"011111101",
  9929=>"000000000",
  9930=>"000011111",
  9931=>"110000110",
  9932=>"100000111",
  9933=>"000001001",
  9934=>"001001001",
  9935=>"110000011",
  9936=>"110110110",
  9937=>"110110110",
  9938=>"110000001",
  9939=>"110001000",
  9940=>"111001000",
  9941=>"101011001",
  9942=>"011110110",
  9943=>"001111111",
  9944=>"001001011",
  9945=>"110100001",
  9946=>"110100000",
  9947=>"001001011",
  9948=>"111111111",
  9949=>"110110110",
  9950=>"111110010",
  9951=>"011001011",
  9952=>"000001010",
  9953=>"011000000",
  9954=>"111000000",
  9955=>"011111001",
  9956=>"001001011",
  9957=>"110110000",
  9958=>"110110110",
  9959=>"100110010",
  9960=>"110001000",
  9961=>"010000000",
  9962=>"001001000",
  9963=>"000111111",
  9964=>"000000000",
  9965=>"110010000",
  9966=>"010010000",
  9967=>"000000000",
  9968=>"000000000",
  9969=>"001001111",
  9970=>"010000100",
  9971=>"000110100",
  9972=>"111111001",
  9973=>"001001001",
  9974=>"000011000",
  9975=>"111101101",
  9976=>"001001111",
  9977=>"000010110",
  9978=>"100001000",
  9979=>"010001101",
  9980=>"011001001",
  9981=>"000001000",
  9982=>"111100000",
  9983=>"001001101",
  9984=>"001000111",
  9985=>"111001000",
  9986=>"000000000",
  9987=>"111000001",
  9988=>"110100101",
  9989=>"111000101",
  9990=>"111111111",
  9991=>"000101000",
  9992=>"101101100",
  9993=>"111101111",
  9994=>"001100001",
  9995=>"001101110",
  9996=>"000011100",
  9997=>"111111000",
  9998=>"011011000",
  9999=>"110111111",
  10000=>"111000101",
  10001=>"010111000",
  10002=>"010100110",
  10003=>"000000111",
  10004=>"111001111",
  10005=>"111111001",
  10006=>"000111101",
  10007=>"010000000",
  10008=>"101000000",
  10009=>"011000011",
  10010=>"111101111",
  10011=>"001001101",
  10012=>"000000000",
  10013=>"000011011",
  10014=>"110000110",
  10015=>"000111111",
  10016=>"111100000",
  10017=>"101100011",
  10018=>"000001010",
  10019=>"000000000",
  10020=>"101000001",
  10021=>"100000111",
  10022=>"010001011",
  10023=>"110001001",
  10024=>"101111010",
  10025=>"000011011",
  10026=>"010101100",
  10027=>"100100000",
  10028=>"001011101",
  10029=>"110010111",
  10030=>"111101011",
  10031=>"011111010",
  10032=>"111101000",
  10033=>"100100101",
  10034=>"000010011",
  10035=>"110110110",
  10036=>"000000000",
  10037=>"010111110",
  10038=>"111111111",
  10039=>"011000001",
  10040=>"100001111",
  10041=>"101101111",
  10042=>"001111111",
  10043=>"000000101",
  10044=>"001100110",
  10045=>"110111000",
  10046=>"101101100",
  10047=>"101101000",
  10048=>"111111010",
  10049=>"100101111",
  10050=>"111010000",
  10051=>"011000100",
  10052=>"010111010",
  10053=>"101000101",
  10054=>"110000100",
  10055=>"100111011",
  10056=>"011111000",
  10057=>"110101000",
  10058=>"000000000",
  10059=>"000000111",
  10060=>"110000001",
  10061=>"100000101",
  10062=>"111001001",
  10063=>"100000101",
  10064=>"000110000",
  10065=>"111111010",
  10066=>"000111010",
  10067=>"000011011",
  10068=>"000010011",
  10069=>"100101101",
  10070=>"001101100",
  10071=>"101000111",
  10072=>"001111110",
  10073=>"000010101",
  10074=>"110011001",
  10075=>"101111011",
  10076=>"100000111",
  10077=>"100000100",
  10078=>"010111101",
  10079=>"111001001",
  10080=>"111101101",
  10081=>"001110010",
  10082=>"101101001",
  10083=>"011110100",
  10084=>"100000101",
  10085=>"101111010",
  10086=>"111010000",
  10087=>"000110111",
  10088=>"001111010",
  10089=>"110101010",
  10090=>"000000011",
  10091=>"111000001",
  10092=>"110001000",
  10093=>"000011110",
  10094=>"101101010",
  10095=>"111111011",
  10096=>"100000111",
  10097=>"000101001",
  10098=>"110111111",
  10099=>"101111010",
  10100=>"100111111",
  10101=>"111011101",
  10102=>"111011001",
  10103=>"111111001",
  10104=>"110110110",
  10105=>"000000111",
  10106=>"000000001",
  10107=>"101110000",
  10108=>"011100001",
  10109=>"000000110",
  10110=>"000010010",
  10111=>"001111111",
  10112=>"011001001",
  10113=>"111101000",
  10114=>"000000000",
  10115=>"000010000",
  10116=>"000100111",
  10117=>"111110000",
  10118=>"001001111",
  10119=>"011000000",
  10120=>"001001001",
  10121=>"111000011",
  10122=>"000010010",
  10123=>"010110100",
  10124=>"101000000",
  10125=>"001100001",
  10126=>"000111111",
  10127=>"110000010",
  10128=>"001000001",
  10129=>"111101100",
  10130=>"110000100",
  10131=>"011000000",
  10132=>"000001110",
  10133=>"101001000",
  10134=>"101001001",
  10135=>"001100100",
  10136=>"101000000",
  10137=>"001010010",
  10138=>"000111111",
  10139=>"010010000",
  10140=>"000001001",
  10141=>"111000100",
  10142=>"011111111",
  10143=>"100001001",
  10144=>"101000100",
  10145=>"111111101",
  10146=>"000110000",
  10147=>"000010010",
  10148=>"111111111",
  10149=>"000001001",
  10150=>"111111111",
  10151=>"101101011",
  10152=>"011111001",
  10153=>"110110111",
  10154=>"101101101",
  10155=>"001000000",
  10156=>"010010000",
  10157=>"111101001",
  10158=>"000000001",
  10159=>"101011000",
  10160=>"011000000",
  10161=>"110001001",
  10162=>"000000000",
  10163=>"000001000",
  10164=>"010111111",
  10165=>"011111011",
  10166=>"101101101",
  10167=>"000000011",
  10168=>"100000001",
  10169=>"010010000",
  10170=>"110010111",
  10171=>"000000101",
  10172=>"101111111",
  10173=>"011111101",
  10174=>"111000101",
  10175=>"000101110",
  10176=>"111000010",
  10177=>"001000111",
  10178=>"000110001",
  10179=>"100000111",
  10180=>"000010110",
  10181=>"001000101",
  10182=>"011111000",
  10183=>"111111101",
  10184=>"010000010",
  10185=>"001011001",
  10186=>"110111101",
  10187=>"111001001",
  10188=>"001100000",
  10189=>"111101101",
  10190=>"000000101",
  10191=>"111111101",
  10192=>"111110110",
  10193=>"000001001",
  10194=>"010010010",
  10195=>"110011010",
  10196=>"101101101",
  10197=>"100000000",
  10198=>"101101101",
  10199=>"000110011",
  10200=>"101101101",
  10201=>"111010010",
  10202=>"110011010",
  10203=>"111101000",
  10204=>"000111001",
  10205=>"111000000",
  10206=>"000101111",
  10207=>"101001000",
  10208=>"000010010",
  10209=>"111011101",
  10210=>"000010011",
  10211=>"110000000",
  10212=>"101000000",
  10213=>"111001010",
  10214=>"111001110",
  10215=>"000000000",
  10216=>"100111101",
  10217=>"100001000",
  10218=>"101001000",
  10219=>"101111101",
  10220=>"101001000",
  10221=>"000001101",
  10222=>"100101110",
  10223=>"101000000",
  10224=>"101100100",
  10225=>"100000111",
  10226=>"101101001",
  10227=>"011110110",
  10228=>"100010110",
  10229=>"101010011",
  10230=>"000000001",
  10231=>"011111010",
  10232=>"101101101",
  10233=>"010010000",
  10234=>"000000111",
  10235=>"111011110",
  10236=>"100101101",
  10237=>"000100000",
  10238=>"001100101",
  10239=>"001000010",
  10240=>"101001001",
  10241=>"000000000",
  10242=>"101100101",
  10243=>"000000110",
  10244=>"101111110",
  10245=>"011000000",
  10246=>"111110000",
  10247=>"110000111",
  10248=>"101011010",
  10249=>"000001000",
  10250=>"001100110",
  10251=>"110010000",
  10252=>"000100101",
  10253=>"100111110",
  10254=>"100001001",
  10255=>"000001111",
  10256=>"110111010",
  10257=>"100111000",
  10258=>"111010101",
  10259=>"000000011",
  10260=>"001001000",
  10261=>"010000100",
  10262=>"000111111",
  10263=>"111100111",
  10264=>"111100111",
  10265=>"011011001",
  10266=>"010000000",
  10267=>"011000000",
  10268=>"111110100",
  10269=>"111101010",
  10270=>"101111111",
  10271=>"100000000",
  10272=>"111111111",
  10273=>"111010010",
  10274=>"101101100",
  10275=>"010100110",
  10276=>"111100100",
  10277=>"001100000",
  10278=>"110010000",
  10279=>"000111110",
  10280=>"111000000",
  10281=>"110000001",
  10282=>"000111111",
  10283=>"010111111",
  10284=>"010001001",
  10285=>"100000111",
  10286=>"100000000",
  10287=>"101001111",
  10288=>"000000010",
  10289=>"111111111",
  10290=>"100001001",
  10291=>"000000001",
  10292=>"111110000",
  10293=>"000010101",
  10294=>"100011011",
  10295=>"110101101",
  10296=>"110000101",
  10297=>"000000000",
  10298=>"111010010",
  10299=>"111000000",
  10300=>"010111110",
  10301=>"111101101",
  10302=>"000000000",
  10303=>"001011111",
  10304=>"110010111",
  10305=>"111000000",
  10306=>"011100111",
  10307=>"000100110",
  10308=>"111111010",
  10309=>"111001101",
  10310=>"000111010",
  10311=>"000000000",
  10312=>"111110000",
  10313=>"000111010",
  10314=>"100001101",
  10315=>"010110110",
  10316=>"111011000",
  10317=>"000001000",
  10318=>"111111111",
  10319=>"000101111",
  10320=>"111111100",
  10321=>"100010001",
  10322=>"100000010",
  10323=>"111101101",
  10324=>"101101111",
  10325=>"010111111",
  10326=>"110110010",
  10327=>"000111111",
  10328=>"111111111",
  10329=>"011000010",
  10330=>"010110110",
  10331=>"011110000",
  10332=>"010000000",
  10333=>"001001011",
  10334=>"010000111",
  10335=>"000011011",
  10336=>"000000000",
  10337=>"010110000",
  10338=>"001101111",
  10339=>"001011000",
  10340=>"100101000",
  10341=>"101011011",
  10342=>"110000000",
  10343=>"000001111",
  10344=>"110010111",
  10345=>"010111101",
  10346=>"000000111",
  10347=>"111001000",
  10348=>"111100101",
  10349=>"000010111",
  10350=>"011010011",
  10351=>"010000000",
  10352=>"011100000",
  10353=>"111000000",
  10354=>"110110110",
  10355=>"000000111",
  10356=>"000000111",
  10357=>"001000000",
  10358=>"010000010",
  10359=>"000101000",
  10360=>"000000111",
  10361=>"000000111",
  10362=>"100000010",
  10363=>"001001000",
  10364=>"000110110",
  10365=>"101100110",
  10366=>"000001111",
  10367=>"101101000",
  10368=>"000000010",
  10369=>"111100100",
  10370=>"000000000",
  10371=>"001000111",
  10372=>"101000100",
  10373=>"100000000",
  10374=>"001001000",
  10375=>"010011000",
  10376=>"101001001",
  10377=>"110111000",
  10378=>"000001000",
  10379=>"001100111",
  10380=>"111100101",
  10381=>"000000100",
  10382=>"111111111",
  10383=>"000000001",
  10384=>"101101111",
  10385=>"111001000",
  10386=>"111011000",
  10387=>"110010110",
  10388=>"110111111",
  10389=>"000111111",
  10390=>"110111111",
  10391=>"000000000",
  10392=>"111111110",
  10393=>"000111111",
  10394=>"010100100",
  10395=>"100000110",
  10396=>"000011011",
  10397=>"101000000",
  10398=>"000000110",
  10399=>"001001000",
  10400=>"101011101",
  10401=>"010010011",
  10402=>"000101111",
  10403=>"111010111",
  10404=>"000000010",
  10405=>"110001000",
  10406=>"101001000",
  10407=>"010010100",
  10408=>"000000110",
  10409=>"010111111",
  10410=>"101000001",
  10411=>"110010000",
  10412=>"010011111",
  10413=>"100000000",
  10414=>"101111000",
  10415=>"000011000",
  10416=>"010010001",
  10417=>"011111110",
  10418=>"000000010",
  10419=>"001101100",
  10420=>"110100100",
  10421=>"000100111",
  10422=>"010100111",
  10423=>"000110111",
  10424=>"000001011",
  10425=>"111111111",
  10426=>"001010010",
  10427=>"000000111",
  10428=>"000000101",
  10429=>"111101111",
  10430=>"100100000",
  10431=>"110110101",
  10432=>"000000000",
  10433=>"111000000",
  10434=>"010000110",
  10435=>"111101100",
  10436=>"001000111",
  10437=>"111111010",
  10438=>"011000011",
  10439=>"111001000",
  10440=>"101111111",
  10441=>"111010000",
  10442=>"100101111",
  10443=>"111101011",
  10444=>"111011001",
  10445=>"010011011",
  10446=>"001111111",
  10447=>"001000010",
  10448=>"010000000",
  10449=>"101100000",
  10450=>"110010110",
  10451=>"101111101",
  10452=>"110000000",
  10453=>"111111001",
  10454=>"001000000",
  10455=>"111000011",
  10456=>"000000111",
  10457=>"100000000",
  10458=>"101011000",
  10459=>"111010111",
  10460=>"011111101",
  10461=>"000011111",
  10462=>"010000101",
  10463=>"000000000",
  10464=>"000000000",
  10465=>"101000010",
  10466=>"000000000",
  10467=>"011111100",
  10468=>"111100000",
  10469=>"111000101",
  10470=>"101101111",
  10471=>"101110010",
  10472=>"100000000",
  10473=>"010000100",
  10474=>"000100000",
  10475=>"010110111",
  10476=>"011001000",
  10477=>"100000000",
  10478=>"000000000",
  10479=>"000010000",
  10480=>"111011100",
  10481=>"111111100",
  10482=>"011000100",
  10483=>"111101100",
  10484=>"100110000",
  10485=>"100100100",
  10486=>"000000000",
  10487=>"111001011",
  10488=>"011110111",
  10489=>"000111111",
  10490=>"001000000",
  10491=>"111111000",
  10492=>"000000001",
  10493=>"000000110",
  10494=>"010010001",
  10495=>"000000000",
  10496=>"110011000",
  10497=>"000100111",
  10498=>"101000001",
  10499=>"000000110",
  10500=>"001001010",
  10501=>"100000000",
  10502=>"110111010",
  10503=>"010100000",
  10504=>"110110110",
  10505=>"001000100",
  10506=>"000000100",
  10507=>"000000000",
  10508=>"001000000",
  10509=>"111110110",
  10510=>"001011011",
  10511=>"110000000",
  10512=>"011001111",
  10513=>"000000001",
  10514=>"000000000",
  10515=>"000111111",
  10516=>"111001101",
  10517=>"000000000",
  10518=>"001111111",
  10519=>"100100111",
  10520=>"101000100",
  10521=>"000111001",
  10522=>"011000000",
  10523=>"111101000",
  10524=>"000001110",
  10525=>"000000101",
  10526=>"111001000",
  10527=>"010000000",
  10528=>"110101100",
  10529=>"011101000",
  10530=>"001100010",
  10531=>"000000000",
  10532=>"001011111",
  10533=>"111111111",
  10534=>"000000001",
  10535=>"000000111",
  10536=>"111111110",
  10537=>"111111100",
  10538=>"000000000",
  10539=>"110101111",
  10540=>"010111011",
  10541=>"000000111",
  10542=>"101111001",
  10543=>"000100000",
  10544=>"000000111",
  10545=>"001001001",
  10546=>"001100000",
  10547=>"111111111",
  10548=>"110000111",
  10549=>"111110111",
  10550=>"010100101",
  10551=>"000000000",
  10552=>"110000000",
  10553=>"000001101",
  10554=>"101000101",
  10555=>"000100100",
  10556=>"100010101",
  10557=>"111111111",
  10558=>"100000001",
  10559=>"110111010",
  10560=>"110001000",
  10561=>"001101000",
  10562=>"000001010",
  10563=>"110010100",
  10564=>"000110111",
  10565=>"110001111",
  10566=>"111000111",
  10567=>"011110000",
  10568=>"000000011",
  10569=>"010001000",
  10570=>"111001111",
  10571=>"110000000",
  10572=>"000100110",
  10573=>"011100011",
  10574=>"000111100",
  10575=>"011011011",
  10576=>"111111010",
  10577=>"010011010",
  10578=>"001110111",
  10579=>"011001001",
  10580=>"000000000",
  10581=>"111011111",
  10582=>"100100100",
  10583=>"000000000",
  10584=>"111100000",
  10585=>"000011010",
  10586=>"000000000",
  10587=>"110110000",
  10588=>"000010000",
  10589=>"011001001",
  10590=>"000010010",
  10591=>"000001001",
  10592=>"010111110",
  10593=>"111111101",
  10594=>"101000101",
  10595=>"000000000",
  10596=>"000001000",
  10597=>"111011011",
  10598=>"111110000",
  10599=>"000100000",
  10600=>"110000111",
  10601=>"000000000",
  10602=>"110000001",
  10603=>"100001000",
  10604=>"101111111",
  10605=>"000100001",
  10606=>"111011011",
  10607=>"110000000",
  10608=>"111111111",
  10609=>"010000111",
  10610=>"110100101",
  10611=>"100111111",
  10612=>"100110111",
  10613=>"000000100",
  10614=>"110110110",
  10615=>"111110010",
  10616=>"000000000",
  10617=>"111111010",
  10618=>"111111100",
  10619=>"001000001",
  10620=>"100100110",
  10621=>"111101001",
  10622=>"000001110",
  10623=>"011000000",
  10624=>"111111001",
  10625=>"110100000",
  10626=>"011011110",
  10627=>"001000011",
  10628=>"000000101",
  10629=>"111111111",
  10630=>"100111110",
  10631=>"011100000",
  10632=>"110111111",
  10633=>"101111111",
  10634=>"000000111",
  10635=>"010000000",
  10636=>"110110000",
  10637=>"110110000",
  10638=>"001000000",
  10639=>"000000100",
  10640=>"110100100",
  10641=>"000001101",
  10642=>"000000000",
  10643=>"111001000",
  10644=>"000001001",
  10645=>"000000000",
  10646=>"000001000",
  10647=>"110011011",
  10648=>"001110000",
  10649=>"000000111",
  10650=>"000000000",
  10651=>"101000000",
  10652=>"010111010",
  10653=>"111111111",
  10654=>"111000010",
  10655=>"000000000",
  10656=>"001101101",
  10657=>"111001111",
  10658=>"110111111",
  10659=>"000111111",
  10660=>"101001110",
  10661=>"110111000",
  10662=>"111111011",
  10663=>"110111111",
  10664=>"000111001",
  10665=>"110001110",
  10666=>"001000000",
  10667=>"000000001",
  10668=>"111100111",
  10669=>"110111011",
  10670=>"110101111",
  10671=>"010111010",
  10672=>"100010000",
  10673=>"100100000",
  10674=>"000000000",
  10675=>"011101010",
  10676=>"110110111",
  10677=>"111001000",
  10678=>"010111010",
  10679=>"111111001",
  10680=>"011110111",
  10681=>"110110001",
  10682=>"010010000",
  10683=>"110111010",
  10684=>"101111001",
  10685=>"111111111",
  10686=>"010011111",
  10687=>"110111011",
  10688=>"011000000",
  10689=>"111000001",
  10690=>"000000111",
  10691=>"011011001",
  10692=>"101110000",
  10693=>"001111111",
  10694=>"000000010",
  10695=>"000000000",
  10696=>"100101111",
  10697=>"010010000",
  10698=>"100110111",
  10699=>"001000000",
  10700=>"011000000",
  10701=>"001011110",
  10702=>"111000000",
  10703=>"111101111",
  10704=>"110101110",
  10705=>"111111111",
  10706=>"000110111",
  10707=>"110111111",
  10708=>"001000000",
  10709=>"011000100",
  10710=>"110110011",
  10711=>"110100000",
  10712=>"000000111",
  10713=>"000000010",
  10714=>"000000100",
  10715=>"001000000",
  10716=>"100111101",
  10717=>"000100000",
  10718=>"110111000",
  10719=>"110001000",
  10720=>"001000000",
  10721=>"111001101",
  10722=>"000000000",
  10723=>"110111111",
  10724=>"101011010",
  10725=>"000111010",
  10726=>"000110110",
  10727=>"010011001",
  10728=>"100111111",
  10729=>"010010111",
  10730=>"001000001",
  10731=>"110110110",
  10732=>"010010000",
  10733=>"000101010",
  10734=>"011000010",
  10735=>"001000010",
  10736=>"101100101",
  10737=>"100001111",
  10738=>"000001001",
  10739=>"011000010",
  10740=>"111100000",
  10741=>"010110111",
  10742=>"000000000",
  10743=>"100000000",
  10744=>"010000000",
  10745=>"000010010",
  10746=>"000000000",
  10747=>"001110000",
  10748=>"000000000",
  10749=>"011001000",
  10750=>"100100100",
  10751=>"001000000",
  10752=>"000100110",
  10753=>"000010001",
  10754=>"100000010",
  10755=>"000000000",
  10756=>"000010000",
  10757=>"100000110",
  10758=>"001001111",
  10759=>"000010010",
  10760=>"010011000",
  10761=>"001000111",
  10762=>"001001000",
  10763=>"000001000",
  10764=>"001000001",
  10765=>"111111101",
  10766=>"000011100",
  10767=>"000000000",
  10768=>"111000000",
  10769=>"110100010",
  10770=>"100000001",
  10771=>"110101111",
  10772=>"110011000",
  10773=>"111100110",
  10774=>"001000000",
  10775=>"101001000",
  10776=>"101000111",
  10777=>"011111011",
  10778=>"000000000",
  10779=>"111000101",
  10780=>"111000010",
  10781=>"100000001",
  10782=>"110111111",
  10783=>"001110000",
  10784=>"000010010",
  10785=>"100001101",
  10786=>"110101000",
  10787=>"111010000",
  10788=>"111000000",
  10789=>"000011111",
  10790=>"010110000",
  10791=>"011110000",
  10792=>"010110001",
  10793=>"010010001",
  10794=>"100110101",
  10795=>"111110111",
  10796=>"000000100",
  10797=>"111101111",
  10798=>"010010000",
  10799=>"000000000",
  10800=>"101111101",
  10801=>"000000111",
  10802=>"100010010",
  10803=>"000101111",
  10804=>"001000111",
  10805=>"001011000",
  10806=>"000001111",
  10807=>"111001101",
  10808=>"010000011",
  10809=>"001101111",
  10810=>"111101010",
  10811=>"011000110",
  10812=>"000011011",
  10813=>"110111111",
  10814=>"011000100",
  10815=>"110110010",
  10816=>"000010011",
  10817=>"000010111",
  10818=>"111010101",
  10819=>"010000110",
  10820=>"100101000",
  10821=>"001001101",
  10822=>"000001111",
  10823=>"111111101",
  10824=>"110000111",
  10825=>"111110000",
  10826=>"001001011",
  10827=>"011011000",
  10828=>"100000111",
  10829=>"100100100",
  10830=>"001000001",
  10831=>"010100101",
  10832=>"101101000",
  10833=>"111111111",
  10834=>"111111101",
  10835=>"010111010",
  10836=>"001100110",
  10837=>"000000000",
  10838=>"011000000",
  10839=>"000000011",
  10840=>"100000000",
  10841=>"111111000",
  10842=>"111011111",
  10843=>"111111000",
  10844=>"000000000",
  10845=>"000011110",
  10846=>"111111111",
  10847=>"110000011",
  10848=>"000010000",
  10849=>"100000100",
  10850=>"101001111",
  10851=>"001100111",
  10852=>"111111001",
  10853=>"000000100",
  10854=>"101111111",
  10855=>"010010000",
  10856=>"101001111",
  10857=>"101101011",
  10858=>"111010010",
  10859=>"001111111",
  10860=>"110110101",
  10861=>"111111111",
  10862=>"010000000",
  10863=>"000000100",
  10864=>"011011010",
  10865=>"000000001",
  10866=>"000000111",
  10867=>"001010000",
  10868=>"011000000",
  10869=>"001101110",
  10870=>"000000100",
  10871=>"110000111",
  10872=>"100001111",
  10873=>"010000110",
  10874=>"000001001",
  10875=>"101111101",
  10876=>"000000111",
  10877=>"011101010",
  10878=>"001010111",
  10879=>"101101100",
  10880=>"011001010",
  10881=>"111010011",
  10882=>"111101100",
  10883=>"111111100",
  10884=>"001001001",
  10885=>"111011011",
  10886=>"000111111",
  10887=>"100000100",
  10888=>"100101110",
  10889=>"011001101",
  10890=>"100000111",
  10891=>"111110010",
  10892=>"101101111",
  10893=>"000000010",
  10894=>"000000100",
  10895=>"001001000",
  10896=>"101101001",
  10897=>"101111111",
  10898=>"101000010",
  10899=>"000111010",
  10900=>"000000001",
  10901=>"010000111",
  10902=>"000100111",
  10903=>"001111100",
  10904=>"011010101",
  10905=>"101111110",
  10906=>"001000111",
  10907=>"000000101",
  10908=>"101111000",
  10909=>"111001011",
  10910=>"011000000",
  10911=>"110110000",
  10912=>"001001110",
  10913=>"001000001",
  10914=>"111011100",
  10915=>"000010000",
  10916=>"110111111",
  10917=>"110101000",
  10918=>"110110001",
  10919=>"111010111",
  10920=>"101000111",
  10921=>"000010000",
  10922=>"101100111",
  10923=>"000000111",
  10924=>"111111111",
  10925=>"000000000",
  10926=>"100001001",
  10927=>"010111101",
  10928=>"101000111",
  10929=>"001000100",
  10930=>"101101110",
  10931=>"000110001",
  10932=>"110111010",
  10933=>"111111111",
  10934=>"011100100",
  10935=>"000011101",
  10936=>"000100100",
  10937=>"011000010",
  10938=>"111010000",
  10939=>"111101000",
  10940=>"001011110",
  10941=>"010010101",
  10942=>"111111001",
  10943=>"101011010",
  10944=>"101001111",
  10945=>"101000111",
  10946=>"010010000",
  10947=>"000000011",
  10948=>"000000001",
  10949=>"110000110",
  10950=>"000011100",
  10951=>"101000000",
  10952=>"001111100",
  10953=>"001001001",
  10954=>"011011111",
  10955=>"000000111",
  10956=>"000000100",
  10957=>"000000001",
  10958=>"101101000",
  10959=>"101101010",
  10960=>"111101101",
  10961=>"110110001",
  10962=>"010000000",
  10963=>"000000000",
  10964=>"110000000",
  10965=>"100000000",
  10966=>"010000111",
  10967=>"001011011",
  10968=>"111010000",
  10969=>"011111111",
  10970=>"100101001",
  10971=>"111001111",
  10972=>"000000100",
  10973=>"101111010",
  10974=>"000100111",
  10975=>"001000101",
  10976=>"111101101",
  10977=>"101100111",
  10978=>"001010000",
  10979=>"000100000",
  10980=>"101000010",
  10981=>"000000000",
  10982=>"000000000",
  10983=>"000000000",
  10984=>"100100100",
  10985=>"000111111",
  10986=>"100000100",
  10987=>"000101101",
  10988=>"000000101",
  10989=>"010001001",
  10990=>"010000010",
  10991=>"101000001",
  10992=>"111001000",
  10993=>"011010001",
  10994=>"010111111",
  10995=>"000110100",
  10996=>"000011000",
  10997=>"101001100",
  10998=>"000100000",
  10999=>"000110110",
  11000=>"001101010",
  11001=>"010101010",
  11002=>"000000000",
  11003=>"011000000",
  11004=>"101001101",
  11005=>"010010010",
  11006=>"001111000",
  11007=>"001010111",
  11008=>"101100101",
  11009=>"011000010",
  11010=>"000010010",
  11011=>"011000000",
  11012=>"000001001",
  11013=>"001011010",
  11014=>"111111111",
  11015=>"010111000",
  11016=>"001001001",
  11017=>"101000010",
  11018=>"000000000",
  11019=>"000100110",
  11020=>"011010000",
  11021=>"000000011",
  11022=>"110101000",
  11023=>"101011100",
  11024=>"111111011",
  11025=>"111111010",
  11026=>"111110011",
  11027=>"000000000",
  11028=>"001000110",
  11029=>"111001001",
  11030=>"111100110",
  11031=>"010000000",
  11032=>"010000100",
  11033=>"011010010",
  11034=>"000000111",
  11035=>"001000110",
  11036=>"000000011",
  11037=>"001111100",
  11038=>"000010010",
  11039=>"101111101",
  11040=>"000000101",
  11041=>"000000000",
  11042=>"011101111",
  11043=>"000001000",
  11044=>"000000000",
  11045=>"000001111",
  11046=>"000010011",
  11047=>"001001101",
  11048=>"011111001",
  11049=>"000100011",
  11050=>"010000001",
  11051=>"001011011",
  11052=>"001100101",
  11053=>"100101110",
  11054=>"111001111",
  11055=>"111111111",
  11056=>"111111111",
  11057=>"000000001",
  11058=>"010111100",
  11059=>"000100110",
  11060=>"101001111",
  11061=>"111111110",
  11062=>"010000011",
  11063=>"001001101",
  11064=>"101000000",
  11065=>"000110000",
  11066=>"000011110",
  11067=>"011011111",
  11068=>"000111011",
  11069=>"011111011",
  11070=>"000000000",
  11071=>"100100110",
  11072=>"001000110",
  11073=>"000000011",
  11074=>"000100000",
  11075=>"101001011",
  11076=>"101001011",
  11077=>"111111011",
  11078=>"011000111",
  11079=>"111111011",
  11080=>"000001000",
  11081=>"111111111",
  11082=>"000000000",
  11083=>"001001101",
  11084=>"111011111",
  11085=>"000000001",
  11086=>"000000000",
  11087=>"101111111",
  11088=>"000000000",
  11089=>"111111000",
  11090=>"000101111",
  11091=>"000010011",
  11092=>"000000110",
  11093=>"001001111",
  11094=>"000000010",
  11095=>"000110101",
  11096=>"000111111",
  11097=>"000000011",
  11098=>"101011001",
  11099=>"000000011",
  11100=>"000000010",
  11101=>"001110100",
  11102=>"111111100",
  11103=>"111101000",
  11104=>"111000000",
  11105=>"000000010",
  11106=>"000000000",
  11107=>"111000100",
  11108=>"011111011",
  11109=>"000111000",
  11110=>"100011000",
  11111=>"111111111",
  11112=>"111010111",
  11113=>"111010111",
  11114=>"010111001",
  11115=>"111111011",
  11116=>"000111011",
  11117=>"110110000",
  11118=>"000000001",
  11119=>"000000011",
  11120=>"000000100",
  11121=>"000000000",
  11122=>"101000100",
  11123=>"010110100",
  11124=>"111001001",
  11125=>"001000010",
  11126=>"111111011",
  11127=>"111101101",
  11128=>"000110010",
  11129=>"000011101",
  11130=>"000100101",
  11131=>"101010110",
  11132=>"001001000",
  11133=>"000000100",
  11134=>"001111101",
  11135=>"000010001",
  11136=>"001000000",
  11137=>"001111011",
  11138=>"100000000",
  11139=>"111111011",
  11140=>"010010001",
  11141=>"101101101",
  11142=>"000000110",
  11143=>"000000101",
  11144=>"000000001",
  11145=>"000111111",
  11146=>"000011010",
  11147=>"111011010",
  11148=>"001001000",
  11149=>"001000011",
  11150=>"011000001",
  11151=>"101001001",
  11152=>"100100000",
  11153=>"111100000",
  11154=>"001000000",
  11155=>"000000000",
  11156=>"000000000",
  11157=>"110111100",
  11158=>"101000110",
  11159=>"000000001",
  11160=>"000000110",
  11161=>"000111111",
  11162=>"000011000",
  11163=>"000111001",
  11164=>"000101100",
  11165=>"111000101",
  11166=>"001000010",
  11167=>"000011011",
  11168=>"000000101",
  11169=>"111110000",
  11170=>"111111101",
  11171=>"001000000",
  11172=>"010000000",
  11173=>"000000111",
  11174=>"000000000",
  11175=>"111001111",
  11176=>"000000111",
  11177=>"000001000",
  11178=>"111000010",
  11179=>"000000000",
  11180=>"111111111",
  11181=>"111111111",
  11182=>"000101011",
  11183=>"011111000",
  11184=>"001111101",
  11185=>"001001100",
  11186=>"001110000",
  11187=>"000011011",
  11188=>"111111011",
  11189=>"111000101",
  11190=>"000000001",
  11191=>"000011111",
  11192=>"000100100",
  11193=>"001000001",
  11194=>"010111101",
  11195=>"100000111",
  11196=>"111010111",
  11197=>"001000000",
  11198=>"100111011",
  11199=>"000111111",
  11200=>"011001010",
  11201=>"000000111",
  11202=>"111101101",
  11203=>"000010010",
  11204=>"000111000",
  11205=>"000000100",
  11206=>"000000000",
  11207=>"000000101",
  11208=>"001101101",
  11209=>"001101001",
  11210=>"111001001",
  11211=>"000101000",
  11212=>"000100000",
  11213=>"100000001",
  11214=>"110101000",
  11215=>"001111111",
  11216=>"111111110",
  11217=>"000000111",
  11218=>"001000000",
  11219=>"111111010",
  11220=>"000000000",
  11221=>"111001001",
  11222=>"001000000",
  11223=>"100111111",
  11224=>"000111111",
  11225=>"000100111",
  11226=>"000001001",
  11227=>"000000000",
  11228=>"111010111",
  11229=>"111111111",
  11230=>"111011111",
  11231=>"111111010",
  11232=>"000000110",
  11233=>"110111010",
  11234=>"111111000",
  11235=>"100101111",
  11236=>"010000000",
  11237=>"011001000",
  11238=>"001000101",
  11239=>"000000001",
  11240=>"110000000",
  11241=>"000000001",
  11242=>"100100111",
  11243=>"110000000",
  11244=>"111111111",
  11245=>"100111011",
  11246=>"000001000",
  11247=>"111011011",
  11248=>"001111111",
  11249=>"000000011",
  11250=>"001000010",
  11251=>"100101101",
  11252=>"011001011",
  11253=>"000000000",
  11254=>"010000010",
  11255=>"111001001",
  11256=>"010000001",
  11257=>"111101101",
  11258=>"000000000",
  11259=>"001001001",
  11260=>"000010010",
  11261=>"000010000",
  11262=>"001000000",
  11263=>"111001011",
  11264=>"111011101",
  11265=>"111111111",
  11266=>"000010010",
  11267=>"100000000",
  11268=>"110111111",
  11269=>"111000111",
  11270=>"110010111",
  11271=>"000111011",
  11272=>"100100000",
  11273=>"000000000",
  11274=>"100100100",
  11275=>"001101111",
  11276=>"111010000",
  11277=>"110100101",
  11278=>"100101100",
  11279=>"111111101",
  11280=>"000000000",
  11281=>"000000100",
  11282=>"011001000",
  11283=>"011101111",
  11284=>"000000100",
  11285=>"000111111",
  11286=>"011011001",
  11287=>"101001100",
  11288=>"000000000",
  11289=>"000000010",
  11290=>"100100101",
  11291=>"111100000",
  11292=>"100001111",
  11293=>"001111111",
  11294=>"001000000",
  11295=>"000010111",
  11296=>"000111011",
  11297=>"100100000",
  11298=>"000010110",
  11299=>"100000010",
  11300=>"000100111",
  11301=>"011011101",
  11302=>"001011111",
  11303=>"111010000",
  11304=>"111111111",
  11305=>"111111110",
  11306=>"100000100",
  11307=>"011111010",
  11308=>"111110011",
  11309=>"100000110",
  11310=>"111001000",
  11311=>"111000000",
  11312=>"000000111",
  11313=>"010101111",
  11314=>"101111100",
  11315=>"000111110",
  11316=>"011011001",
  11317=>"111111000",
  11318=>"011011001",
  11319=>"000111011",
  11320=>"111001000",
  11321=>"000000000",
  11322=>"101100100",
  11323=>"000000111",
  11324=>"100000000",
  11325=>"010111011",
  11326=>"001001111",
  11327=>"010111110",
  11328=>"111010000",
  11329=>"000100000",
  11330=>"111000000",
  11331=>"111110000",
  11332=>"000100011",
  11333=>"101000100",
  11334=>"100111011",
  11335=>"100010111",
  11336=>"000000011",
  11337=>"101001011",
  11338=>"101000000",
  11339=>"000000000",
  11340=>"111111011",
  11341=>"000100110",
  11342=>"000010110",
  11343=>"000110111",
  11344=>"000011111",
  11345=>"110101000",
  11346=>"011111111",
  11347=>"111111111",
  11348=>"111110010",
  11349=>"011011011",
  11350=>"000110101",
  11351=>"101111111",
  11352=>"100111110",
  11353=>"000111000",
  11354=>"100111111",
  11355=>"101111110",
  11356=>"100000000",
  11357=>"000000001",
  11358=>"111111111",
  11359=>"111111100",
  11360=>"111111111",
  11361=>"000000001",
  11362=>"111110011",
  11363=>"000001101",
  11364=>"000100000",
  11365=>"010011100",
  11366=>"111010010",
  11367=>"000111111",
  11368=>"001000100",
  11369=>"010100100",
  11370=>"011000000",
  11371=>"010011111",
  11372=>"000100000",
  11373=>"000100111",
  11374=>"000000010",
  11375=>"111000111",
  11376=>"000001011",
  11377=>"000000000",
  11378=>"110110110",
  11379=>"001011000",
  11380=>"000111011",
  11381=>"011000111",
  11382=>"111010000",
  11383=>"111111111",
  11384=>"000000000",
  11385=>"000000111",
  11386=>"111100000",
  11387=>"101111000",
  11388=>"000000000",
  11389=>"101100111",
  11390=>"001001001",
  11391=>"000000000",
  11392=>"101100000",
  11393=>"010000000",
  11394=>"111100000",
  11395=>"011001000",
  11396=>"000100011",
  11397=>"101111010",
  11398=>"110110110",
  11399=>"000000110",
  11400=>"010110110",
  11401=>"000001001",
  11402=>"000100110",
  11403=>"111000100",
  11404=>"101101101",
  11405=>"100111111",
  11406=>"111000000",
  11407=>"111101001",
  11408=>"101011111",
  11409=>"111111000",
  11410=>"000000001",
  11411=>"000000000",
  11412=>"001001111",
  11413=>"101000000",
  11414=>"111100000",
  11415=>"000001001",
  11416=>"111101101",
  11417=>"101100000",
  11418=>"000101110",
  11419=>"111101111",
  11420=>"001011101",
  11421=>"000000000",
  11422=>"000000110",
  11423=>"001101111",
  11424=>"100010011",
  11425=>"011111111",
  11426=>"100000110",
  11427=>"000110000",
  11428=>"111000000",
  11429=>"001111111",
  11430=>"001000101",
  11431=>"111111010",
  11432=>"000000101",
  11433=>"011001101",
  11434=>"010000100",
  11435=>"010011101",
  11436=>"100010000",
  11437=>"111111110",
  11438=>"110110110",
  11439=>"100000010",
  11440=>"111010000",
  11441=>"000001011",
  11442=>"110000101",
  11443=>"000000100",
  11444=>"101101010",
  11445=>"111010110",
  11446=>"001000000",
  11447=>"000000110",
  11448=>"001000000",
  11449=>"000000111",
  11450=>"111011111",
  11451=>"101000111",
  11452=>"000100110",
  11453=>"111000010",
  11454=>"000000000",
  11455=>"000111000",
  11456=>"000010010",
  11457=>"101000100",
  11458=>"111100010",
  11459=>"000100000",
  11460=>"101101100",
  11461=>"000001111",
  11462=>"111101010",
  11463=>"001000101",
  11464=>"011010111",
  11465=>"111100000",
  11466=>"010101110",
  11467=>"101100000",
  11468=>"100111111",
  11469=>"000000000",
  11470=>"101101101",
  11471=>"000000101",
  11472=>"010100000",
  11473=>"110110111",
  11474=>"011000100",
  11475=>"110111101",
  11476=>"010111001",
  11477=>"000101111",
  11478=>"010101000",
  11479=>"000011101",
  11480=>"011111010",
  11481=>"000110110",
  11482=>"010111100",
  11483=>"000000111",
  11484=>"110110010",
  11485=>"100101000",
  11486=>"010010100",
  11487=>"111111111",
  11488=>"100000000",
  11489=>"010000000",
  11490=>"111001110",
  11491=>"000111101",
  11492=>"000101101",
  11493=>"000000000",
  11494=>"010001000",
  11495=>"001011111",
  11496=>"111101001",
  11497=>"000001001",
  11498=>"001001001",
  11499=>"111000100",
  11500=>"110000000",
  11501=>"000100100",
  11502=>"000000000",
  11503=>"110100000",
  11504=>"000100011",
  11505=>"000100111",
  11506=>"011111011",
  11507=>"000111111",
  11508=>"111110011",
  11509=>"000000111",
  11510=>"000110111",
  11511=>"001010000",
  11512=>"100000000",
  11513=>"111111101",
  11514=>"000100100",
  11515=>"000000010",
  11516=>"100111000",
  11517=>"000100101",
  11518=>"010010111",
  11519=>"111110000",
  11520=>"111100110",
  11521=>"010110011",
  11522=>"101001101",
  11523=>"100101111",
  11524=>"100110110",
  11525=>"100100101",
  11526=>"111111011",
  11527=>"111011010",
  11528=>"110100000",
  11529=>"100000000",
  11530=>"101011101",
  11531=>"100110100",
  11532=>"110100100",
  11533=>"110111001",
  11534=>"100110000",
  11535=>"010100111",
  11536=>"100000100",
  11537=>"111100111",
  11538=>"000100111",
  11539=>"000000001",
  11540=>"111001111",
  11541=>"110110011",
  11542=>"111001000",
  11543=>"001110000",
  11544=>"100110110",
  11545=>"000101011",
  11546=>"110100110",
  11547=>"100100000",
  11548=>"011110110",
  11549=>"011011001",
  11550=>"110100011",
  11551=>"101001000",
  11552=>"110001101",
  11553=>"100100110",
  11554=>"000100110",
  11555=>"110000010",
  11556=>"000110111",
  11557=>"110100110",
  11558=>"000010111",
  11559=>"100000100",
  11560=>"010011100",
  11561=>"000111100",
  11562=>"111110110",
  11563=>"001001000",
  11564=>"001110110",
  11565=>"001110111",
  11566=>"001110110",
  11567=>"110111111",
  11568=>"011001001",
  11569=>"110001000",
  11570=>"000100100",
  11571=>"111100011",
  11572=>"100011011",
  11573=>"110010000",
  11574=>"000001011",
  11575=>"110110100",
  11576=>"011010110",
  11577=>"100100100",
  11578=>"111110010",
  11579=>"101001000",
  11580=>"000100100",
  11581=>"110011011",
  11582=>"100100000",
  11583=>"000010011",
  11584=>"101011100",
  11585=>"010100110",
  11586=>"011110000",
  11587=>"100100100",
  11588=>"011000000",
  11589=>"110110000",
  11590=>"000001010",
  11591=>"001011101",
  11592=>"101111110",
  11593=>"110100100",
  11594=>"110000011",
  11595=>"100111111",
  11596=>"000100000",
  11597=>"111111111",
  11598=>"101011001",
  11599=>"011100000",
  11600=>"100010010",
  11601=>"101011111",
  11602=>"111110001",
  11603=>"001000000",
  11604=>"111110111",
  11605=>"110000110",
  11606=>"111001001",
  11607=>"101001001",
  11608=>"001111111",
  11609=>"000000001",
  11610=>"100001001",
  11611=>"101001001",
  11612=>"101100100",
  11613=>"100000000",
  11614=>"000011011",
  11615=>"100100111",
  11616=>"100100100",
  11617=>"000000000",
  11618=>"100100100",
  11619=>"111110110",
  11620=>"011000000",
  11621=>"101001100",
  11622=>"100100100",
  11623=>"001011011",
  11624=>"110100010",
  11625=>"100100000",
  11626=>"000100110",
  11627=>"011111010",
  11628=>"111100100",
  11629=>"001011000",
  11630=>"010100100",
  11631=>"101110110",
  11632=>"111111011",
  11633=>"100110110",
  11634=>"111111101",
  11635=>"001001000",
  11636=>"011110111",
  11637=>"100100000",
  11638=>"100100001",
  11639=>"000010111",
  11640=>"011010111",
  11641=>"001100111",
  11642=>"000100010",
  11643=>"011011000",
  11644=>"011000000",
  11645=>"001010010",
  11646=>"011011011",
  11647=>"100001000",
  11648=>"101100111",
  11649=>"101000100",
  11650=>"001111011",
  11651=>"111100100",
  11652=>"111011011",
  11653=>"011011111",
  11654=>"000100100",
  11655=>"100100100",
  11656=>"100101111",
  11657=>"111111100",
  11658=>"001011000",
  11659=>"010000000",
  11660=>"100011011",
  11661=>"100100000",
  11662=>"000100100",
  11663=>"100100100",
  11664=>"010010000",
  11665=>"100101100",
  11666=>"100100110",
  11667=>"111110110",
  11668=>"011000000",
  11669=>"101100100",
  11670=>"110100100",
  11671=>"100110010",
  11672=>"011001000",
  11673=>"001011011",
  11674=>"100101011",
  11675=>"011011001",
  11676=>"111110110",
  11677=>"100001100",
  11678=>"011110011",
  11679=>"110110110",
  11680=>"101011101",
  11681=>"000110000",
  11682=>"011000001",
  11683=>"100100111",
  11684=>"011110110",
  11685=>"111111110",
  11686=>"010010010",
  11687=>"011100100",
  11688=>"001011111",
  11689=>"111111111",
  11690=>"100100100",
  11691=>"100100100",
  11692=>"000000111",
  11693=>"100000000",
  11694=>"000101010",
  11695=>"001001011",
  11696=>"100100110",
  11697=>"111100100",
  11698=>"101110000",
  11699=>"110110011",
  11700=>"001001001",
  11701=>"110111111",
  11702=>"110110110",
  11703=>"001000000",
  11704=>"110100110",
  11705=>"111100100",
  11706=>"100110100",
  11707=>"011111111",
  11708=>"111111111",
  11709=>"011001000",
  11710=>"110110110",
  11711=>"011001001",
  11712=>"101110101",
  11713=>"110010000",
  11714=>"100110001",
  11715=>"100000101",
  11716=>"100100110",
  11717=>"000101100",
  11718=>"110010000",
  11719=>"111111110",
  11720=>"011011110",
  11721=>"011001000",
  11722=>"010000100",
  11723=>"011011001",
  11724=>"000011001",
  11725=>"001010100",
  11726=>"011011001",
  11727=>"100101111",
  11728=>"000011000",
  11729=>"000000010",
  11730=>"111110010",
  11731=>"110100100",
  11732=>"110000100",
  11733=>"111110110",
  11734=>"111100100",
  11735=>"000100100",
  11736=>"001001001",
  11737=>"000000010",
  11738=>"110110110",
  11739=>"011011011",
  11740=>"001110000",
  11741=>"111011111",
  11742=>"100100011",
  11743=>"110110100",
  11744=>"011111011",
  11745=>"101111110",
  11746=>"011011011",
  11747=>"110111110",
  11748=>"000001010",
  11749=>"111101100",
  11750=>"001110100",
  11751=>"001010111",
  11752=>"000110100",
  11753=>"001000111",
  11754=>"100001001",
  11755=>"111100000",
  11756=>"111100100",
  11757=>"100000000",
  11758=>"000000000",
  11759=>"100000111",
  11760=>"010111111",
  11761=>"000100100",
  11762=>"000110000",
  11763=>"011011010",
  11764=>"011100100",
  11765=>"000001011",
  11766=>"000100010",
  11767=>"001011011",
  11768=>"110100111",
  11769=>"011011111",
  11770=>"010010110",
  11771=>"000000000",
  11772=>"011101111",
  11773=>"001011110",
  11774=>"000000010",
  11775=>"000000000",
  11776=>"000000100",
  11777=>"000000000",
  11778=>"101101101",
  11779=>"111000111",
  11780=>"111011110",
  11781=>"101111000",
  11782=>"100100010",
  11783=>"111110111",
  11784=>"111101101",
  11785=>"010000000",
  11786=>"011011000",
  11787=>"101101100",
  11788=>"000100000",
  11789=>"111000000",
  11790=>"001111110",
  11791=>"010111100",
  11792=>"111011001",
  11793=>"100101101",
  11794=>"000000011",
  11795=>"000000000",
  11796=>"000000000",
  11797=>"011111000",
  11798=>"110101111",
  11799=>"001011111",
  11800=>"000000111",
  11801=>"011111111",
  11802=>"100000101",
  11803=>"111001101",
  11804=>"010111000",
  11805=>"010000000",
  11806=>"111000001",
  11807=>"011111000",
  11808=>"010101111",
  11809=>"111000111",
  11810=>"011011111",
  11811=>"010010000",
  11812=>"111111010",
  11813=>"000100000",
  11814=>"111111111",
  11815=>"100110000",
  11816=>"000001101",
  11817=>"101100111",
  11818=>"001111000",
  11819=>"011000001",
  11820=>"110010011",
  11821=>"010011101",
  11822=>"111111011",
  11823=>"000010100",
  11824=>"100000000",
  11825=>"110011001",
  11826=>"001000111",
  11827=>"111110111",
  11828=>"110000000",
  11829=>"111111111",
  11830=>"110110100",
  11831=>"010001111",
  11832=>"000100000",
  11833=>"101000000",
  11834=>"000000000",
  11835=>"111111111",
  11836=>"111111110",
  11837=>"001011011",
  11838=>"101000000",
  11839=>"101111011",
  11840=>"111001011",
  11841=>"111110010",
  11842=>"000000000",
  11843=>"110111110",
  11844=>"011001000",
  11845=>"000010010",
  11846=>"000111100",
  11847=>"101100110",
  11848=>"101110010",
  11849=>"000000001",
  11850=>"100100111",
  11851=>"110000111",
  11852=>"111000111",
  11853=>"001001000",
  11854=>"111110111",
  11855=>"010101111",
  11856=>"110111111",
  11857=>"000100111",
  11858=>"111111111",
  11859=>"110010010",
  11860=>"101111100",
  11861=>"110100111",
  11862=>"111110111",
  11863=>"111101101",
  11864=>"000000001",
  11865=>"111111111",
  11866=>"011111110",
  11867=>"111111010",
  11868=>"011100111",
  11869=>"001011000",
  11870=>"000100101",
  11871=>"111111011",
  11872=>"111111000",
  11873=>"111111111",
  11874=>"101000111",
  11875=>"110111000",
  11876=>"111111100",
  11877=>"010010010",
  11878=>"001000010",
  11879=>"000000000",
  11880=>"000011000",
  11881=>"000000000",
  11882=>"000000000",
  11883=>"110111000",
  11884=>"011111111",
  11885=>"000111000",
  11886=>"011111111",
  11887=>"010111010",
  11888=>"110111111",
  11889=>"000000000",
  11890=>"111111001",
  11891=>"000110000",
  11892=>"111100000",
  11893=>"000101000",
  11894=>"000000011",
  11895=>"101000000",
  11896=>"111101000",
  11897=>"010011111",
  11898=>"000100001",
  11899=>"001001001",
  11900=>"001000111",
  11901=>"100100000",
  11902=>"000001001",
  11903=>"110111000",
  11904=>"111010010",
  11905=>"100000000",
  11906=>"111000111",
  11907=>"111000101",
  11908=>"011111111",
  11909=>"000000010",
  11910=>"011011000",
  11911=>"010110110",
  11912=>"111111111",
  11913=>"111111100",
  11914=>"000111011",
  11915=>"110010111",
  11916=>"111101001",
  11917=>"100111111",
  11918=>"000110111",
  11919=>"110110000",
  11920=>"000011110",
  11921=>"111111010",
  11922=>"100111111",
  11923=>"001001011",
  11924=>"111011111",
  11925=>"111111111",
  11926=>"101111000",
  11927=>"111000001",
  11928=>"000000000",
  11929=>"000100111",
  11930=>"111011111",
  11931=>"100111000",
  11932=>"010101111",
  11933=>"110100111",
  11934=>"000000000",
  11935=>"111001111",
  11936=>"000010001",
  11937=>"111000111",
  11938=>"100001000",
  11939=>"000000111",
  11940=>"000000010",
  11941=>"111111110",
  11942=>"000001011",
  11943=>"000000000",
  11944=>"111101111",
  11945=>"111100111",
  11946=>"000000000",
  11947=>"101101101",
  11948=>"001010110",
  11949=>"111111111",
  11950=>"000111011",
  11951=>"011111110",
  11952=>"100101111",
  11953=>"000101010",
  11954=>"111101111",
  11955=>"001001111",
  11956=>"000010000",
  11957=>"000011000",
  11958=>"010000100",
  11959=>"011000110",
  11960=>"100110110",
  11961=>"011010111",
  11962=>"000000111",
  11963=>"111000111",
  11964=>"101100111",
  11965=>"111000000",
  11966=>"010111100",
  11967=>"000000101",
  11968=>"011111000",
  11969=>"010000111",
  11970=>"100101000",
  11971=>"111111010",
  11972=>"101111111",
  11973=>"000101101",
  11974=>"100101111",
  11975=>"111111111",
  11976=>"110110000",
  11977=>"111111111",
  11978=>"011010101",
  11979=>"010111110",
  11980=>"010111011",
  11981=>"000000111",
  11982=>"100101100",
  11983=>"111111111",
  11984=>"111111000",
  11985=>"001111100",
  11986=>"111111111",
  11987=>"101011111",
  11988=>"000000000",
  11989=>"000110000",
  11990=>"101001000",
  11991=>"100101010",
  11992=>"111111011",
  11993=>"110001000",
  11994=>"000000010",
  11995=>"101000101",
  11996=>"111101011",
  11997=>"000111111",
  11998=>"111110111",
  11999=>"011100010",
  12000=>"010011111",
  12001=>"001000111",
  12002=>"110111111",
  12003=>"011111011",
  12004=>"011111001",
  12005=>"111011101",
  12006=>"110111000",
  12007=>"111111101",
  12008=>"101100000",
  12009=>"000000100",
  12010=>"001011100",
  12011=>"111001111",
  12012=>"101001001",
  12013=>"110101111",
  12014=>"000000111",
  12015=>"000100011",
  12016=>"111100000",
  12017=>"010011111",
  12018=>"111111111",
  12019=>"110111000",
  12020=>"110100011",
  12021=>"010110111",
  12022=>"111000000",
  12023=>"111001111",
  12024=>"111111111",
  12025=>"111011000",
  12026=>"011010111",
  12027=>"101110000",
  12028=>"111111101",
  12029=>"010110111",
  12030=>"110110000",
  12031=>"001111110",
  12032=>"011011001",
  12033=>"000100111",
  12034=>"101000000",
  12035=>"000101110",
  12036=>"100111001",
  12037=>"111110010",
  12038=>"100111111",
  12039=>"010000000",
  12040=>"000110100",
  12041=>"110010110",
  12042=>"011111011",
  12043=>"000000011",
  12044=>"101100000",
  12045=>"011101111",
  12046=>"111111111",
  12047=>"000001001",
  12048=>"110110111",
  12049=>"110111110",
  12050=>"111111000",
  12051=>"011011111",
  12052=>"101000000",
  12053=>"011111010",
  12054=>"011001000",
  12055=>"000000111",
  12056=>"111111100",
  12057=>"111111101",
  12058=>"000111000",
  12059=>"000000010",
  12060=>"101000111",
  12061=>"000000100",
  12062=>"111111000",
  12063=>"110010010",
  12064=>"010010000",
  12065=>"010011011",
  12066=>"011000111",
  12067=>"000000000",
  12068=>"100101111",
  12069=>"111101001",
  12070=>"000011011",
  12071=>"000011010",
  12072=>"101000100",
  12073=>"001000100",
  12074=>"001111111",
  12075=>"111100100",
  12076=>"000100001",
  12077=>"000001010",
  12078=>"011111001",
  12079=>"110111111",
  12080=>"000110000",
  12081=>"111001000",
  12082=>"001000011",
  12083=>"111110111",
  12084=>"111111101",
  12085=>"111111010",
  12086=>"111100110",
  12087=>"000011111",
  12088=>"111111000",
  12089=>"111111111",
  12090=>"000000100",
  12091=>"100011000",
  12092=>"111111001",
  12093=>"001101111",
  12094=>"010000100",
  12095=>"111111111",
  12096=>"111101101",
  12097=>"000110110",
  12098=>"111100000",
  12099=>"011011110",
  12100=>"000110110",
  12101=>"111001001",
  12102=>"010110000",
  12103=>"000110101",
  12104=>"000000000",
  12105=>"110111111",
  12106=>"111101110",
  12107=>"001110111",
  12108=>"111111111",
  12109=>"000111111",
  12110=>"011101110",
  12111=>"000000000",
  12112=>"111110111",
  12113=>"011011111",
  12114=>"010111100",
  12115=>"011001000",
  12116=>"000000000",
  12117=>"111111100",
  12118=>"001001001",
  12119=>"111111111",
  12120=>"000100101",
  12121=>"001111111",
  12122=>"111111101",
  12123=>"111111111",
  12124=>"010111110",
  12125=>"000001001",
  12126=>"000000000",
  12127=>"111110110",
  12128=>"000010010",
  12129=>"001111000",
  12130=>"110000000",
  12131=>"110100000",
  12132=>"111111111",
  12133=>"111001000",
  12134=>"000100101",
  12135=>"110111111",
  12136=>"111111010",
  12137=>"000111111",
  12138=>"000010110",
  12139=>"000000101",
  12140=>"010100010",
  12141=>"010110111",
  12142=>"010011000",
  12143=>"010010111",
  12144=>"010110110",
  12145=>"000001000",
  12146=>"111011011",
  12147=>"000110111",
  12148=>"110000111",
  12149=>"000000001",
  12150=>"101111111",
  12151=>"111111000",
  12152=>"000000000",
  12153=>"101010110",
  12154=>"010111111",
  12155=>"001001001",
  12156=>"000110111",
  12157=>"110100000",
  12158=>"000101000",
  12159=>"111111111",
  12160=>"110111000",
  12161=>"111101111",
  12162=>"010111111",
  12163=>"000100111",
  12164=>"010111111",
  12165=>"101110101",
  12166=>"111101101",
  12167=>"011111111",
  12168=>"111111001",
  12169=>"100000010",
  12170=>"000000011",
  12171=>"000000000",
  12172=>"000000000",
  12173=>"110111111",
  12174=>"111111010",
  12175=>"101001111",
  12176=>"100001011",
  12177=>"110010001",
  12178=>"111111101",
  12179=>"000000001",
  12180=>"111011001",
  12181=>"111111110",
  12182=>"011110011",
  12183=>"101101011",
  12184=>"000110111",
  12185=>"000000001",
  12186=>"010111111",
  12187=>"000000000",
  12188=>"111011001",
  12189=>"110110010",
  12190=>"000000111",
  12191=>"000000000",
  12192=>"001001001",
  12193=>"111111000",
  12194=>"001101100",
  12195=>"010000101",
  12196=>"110110000",
  12197=>"100110100",
  12198=>"001111111",
  12199=>"010001010",
  12200=>"010111111",
  12201=>"111111111",
  12202=>"000000000",
  12203=>"111101110",
  12204=>"001001000",
  12205=>"111111111",
  12206=>"111100000",
  12207=>"001000010",
  12208=>"000001010",
  12209=>"000110110",
  12210=>"010001000",
  12211=>"000100110",
  12212=>"000110111",
  12213=>"010111000",
  12214=>"111111111",
  12215=>"101111011",
  12216=>"011110001",
  12217=>"010111100",
  12218=>"111110110",
  12219=>"010110110",
  12220=>"001000100",
  12221=>"111111111",
  12222=>"010010001",
  12223=>"111111000",
  12224=>"010111000",
  12225=>"010111110",
  12226=>"110111111",
  12227=>"001101111",
  12228=>"000000000",
  12229=>"100100100",
  12230=>"111111101",
  12231=>"010111111",
  12232=>"000000101",
  12233=>"111111000",
  12234=>"111111111",
  12235=>"000111010",
  12236=>"000011011",
  12237=>"000010111",
  12238=>"001010110",
  12239=>"000010111",
  12240=>"010010110",
  12241=>"001101100",
  12242=>"111001000",
  12243=>"000110001",
  12244=>"111001111",
  12245=>"011100100",
  12246=>"110000111",
  12247=>"110111111",
  12248=>"000000000",
  12249=>"110110000",
  12250=>"111100100",
  12251=>"110000010",
  12252=>"111101000",
  12253=>"000011111",
  12254=>"000111111",
  12255=>"111110110",
  12256=>"010000000",
  12257=>"110000000",
  12258=>"101100001",
  12259=>"000100100",
  12260=>"000010111",
  12261=>"010100010",
  12262=>"000000111",
  12263=>"010001100",
  12264=>"110100101",
  12265=>"000110100",
  12266=>"101110111",
  12267=>"000111110",
  12268=>"111000000",
  12269=>"101010110",
  12270=>"011001001",
  12271=>"010000101",
  12272=>"000000000",
  12273=>"011011001",
  12274=>"000010010",
  12275=>"010011011",
  12276=>"111111100",
  12277=>"101001000",
  12278=>"111111110",
  12279=>"000110011",
  12280=>"111000000",
  12281=>"111000010",
  12282=>"011111111",
  12283=>"111111111",
  12284=>"010111111",
  12285=>"000110101",
  12286=>"001101111",
  12287=>"000000111",
  12288=>"011011000",
  12289=>"001011011",
  12290=>"100100100",
  12291=>"100100001",
  12292=>"110110110",
  12293=>"000100100",
  12294=>"101100100",
  12295=>"000000000",
  12296=>"000000000",
  12297=>"100000110",
  12298=>"001010010",
  12299=>"100100100",
  12300=>"000000100",
  12301=>"100011111",
  12302=>"111100110",
  12303=>"011100111",
  12304=>"111101111",
  12305=>"111100110",
  12306=>"100100110",
  12307=>"001011011",
  12308=>"111111101",
  12309=>"111100000",
  12310=>"000101001",
  12311=>"100010110",
  12312=>"100100100",
  12313=>"101011011",
  12314=>"111011111",
  12315=>"000001111",
  12316=>"011011001",
  12317=>"011011000",
  12318=>"111100100",
  12319=>"000011011",
  12320=>"011011001",
  12321=>"100000100",
  12322=>"000111110",
  12323=>"011011000",
  12324=>"100010100",
  12325=>"001011011",
  12326=>"000011011",
  12327=>"000000000",
  12328=>"110011011",
  12329=>"000011111",
  12330=>"100000000",
  12331=>"011000000",
  12332=>"010011011",
  12333=>"111110111",
  12334=>"110111100",
  12335=>"110000000",
  12336=>"010011000",
  12337=>"111101000",
  12338=>"010000000",
  12339=>"011011001",
  12340=>"000011011",
  12341=>"001000111",
  12342=>"001011011",
  12343=>"000000000",
  12344=>"111100011",
  12345=>"111100000",
  12346=>"010000000",
  12347=>"010010011",
  12348=>"010010010",
  12349=>"111011110",
  12350=>"001100000",
  12351=>"100111101",
  12352=>"111111010",
  12353=>"001001000",
  12354=>"011100100",
  12355=>"111000000",
  12356=>"011101101",
  12357=>"000100100",
  12358=>"011111111",
  12359=>"000011011",
  12360=>"001111101",
  12361=>"111100111",
  12362=>"111100100",
  12363=>"011110111",
  12364=>"000000000",
  12365=>"100000000",
  12366=>"011110111",
  12367=>"010011011",
  12368=>"101000100",
  12369=>"111111111",
  12370=>"001000000",
  12371=>"011101000",
  12372=>"000000001",
  12373=>"011011010",
  12374=>"000001000",
  12375=>"111000100",
  12376=>"011110111",
  12377=>"011011001",
  12378=>"000101001",
  12379=>"100101111",
  12380=>"010100000",
  12381=>"111101100",
  12382=>"111011010",
  12383=>"110100100",
  12384=>"011001000",
  12385=>"010000000",
  12386=>"111100100",
  12387=>"000110010",
  12388=>"100000100",
  12389=>"111111111",
  12390=>"000111111",
  12391=>"100011011",
  12392=>"100010101",
  12393=>"011000100",
  12394=>"100111011",
  12395=>"000011000",
  12396=>"000101010",
  12397=>"111101001",
  12398=>"111100101",
  12399=>"000101111",
  12400=>"110011111",
  12401=>"111000000",
  12402=>"110100000",
  12403=>"000100000",
  12404=>"000101011",
  12405=>"100100001",
  12406=>"100000000",
  12407=>"000100000",
  12408=>"011011000",
  12409=>"100110011",
  12410=>"100000011",
  12411=>"000000000",
  12412=>"010110011",
  12413=>"010110000",
  12414=>"010000101",
  12415=>"100100100",
  12416=>"011011000",
  12417=>"101100110",
  12418=>"100000000",
  12419=>"000111110",
  12420=>"100000100",
  12421=>"011011111",
  12422=>"110011000",
  12423=>"000001001",
  12424=>"001101101",
  12425=>"111100000",
  12426=>"111100100",
  12427=>"100000000",
  12428=>"100100001",
  12429=>"000000100",
  12430=>"111100000",
  12431=>"001000000",
  12432=>"100101101",
  12433=>"000000011",
  12434=>"000011001",
  12435=>"000101101",
  12436=>"000011011",
  12437=>"111100101",
  12438=>"111011000",
  12439=>"110100000",
  12440=>"000000000",
  12441=>"011011111",
  12442=>"010011011",
  12443=>"100000000",
  12444=>"011010100",
  12445=>"100000000",
  12446=>"111100000",
  12447=>"111100100",
  12448=>"011011000",
  12449=>"111000011",
  12450=>"110011000",
  12451=>"000010111",
  12452=>"101100000",
  12453=>"100110000",
  12454=>"000111011",
  12455=>"100111010",
  12456=>"111000000",
  12457=>"100100101",
  12458=>"111100101",
  12459=>"111100100",
  12460=>"000010010",
  12461=>"000000100",
  12462=>"011110010",
  12463=>"100101111",
  12464=>"101000000",
  12465=>"111110110",
  12466=>"011100100",
  12467=>"001110110",
  12468=>"000011111",
  12469=>"000010001",
  12470=>"000101100",
  12471=>"000000001",
  12472=>"000001001",
  12473=>"010001001",
  12474=>"000011111",
  12475=>"011111111",
  12476=>"001011110",
  12477=>"111111100",
  12478=>"000000000",
  12479=>"000000000",
  12480=>"110000100",
  12481=>"100100100",
  12482=>"111111000",
  12483=>"111000111",
  12484=>"000000100",
  12485=>"011011100",
  12486=>"011011110",
  12487=>"111111111",
  12488=>"000100100",
  12489=>"000000011",
  12490=>"110101100",
  12491=>"000000000",
  12492=>"000011011",
  12493=>"100001000",
  12494=>"000111001",
  12495=>"100000010",
  12496=>"000000011",
  12497=>"001111101",
  12498=>"100001011",
  12499=>"111100111",
  12500=>"100000101",
  12501=>"000100000",
  12502=>"100100000",
  12503=>"100100011",
  12504=>"010011000",
  12505=>"000100011",
  12506=>"000111110",
  12507=>"100100100",
  12508=>"001011110",
  12509=>"100100111",
  12510=>"101110111",
  12511=>"000000011",
  12512=>"111000000",
  12513=>"111100100",
  12514=>"011000100",
  12515=>"011000011",
  12516=>"111100001",
  12517=>"100100100",
  12518=>"101000011",
  12519=>"000011011",
  12520=>"111100101",
  12521=>"010011011",
  12522=>"110101101",
  12523=>"011100110",
  12524=>"111100100",
  12525=>"001000001",
  12526=>"111100001",
  12527=>"110100110",
  12528=>"011011011",
  12529=>"111111000",
  12530=>"000100000",
  12531=>"010111000",
  12532=>"000100000",
  12533=>"101100100",
  12534=>"100000011",
  12535=>"000001011",
  12536=>"010110010",
  12537=>"100101111",
  12538=>"000011000",
  12539=>"101111101",
  12540=>"111011000",
  12541=>"110100100",
  12542=>"001011011",
  12543=>"111100100",
  12544=>"011001000",
  12545=>"100110110",
  12546=>"000000000",
  12547=>"000111101",
  12548=>"100000101",
  12549=>"000000101",
  12550=>"000000100",
  12551=>"110000111",
  12552=>"101100001",
  12553=>"000000000",
  12554=>"100000101",
  12555=>"100110000",
  12556=>"110110000",
  12557=>"010011111",
  12558=>"010011101",
  12559=>"101111111",
  12560=>"111111000",
  12561=>"100000001",
  12562=>"001101001",
  12563=>"101111111",
  12564=>"111001000",
  12565=>"101111010",
  12566=>"111101010",
  12567=>"111110111",
  12568=>"000001101",
  12569=>"111111001",
  12570=>"000000101",
  12571=>"000000111",
  12572=>"101101111",
  12573=>"000111111",
  12574=>"111000000",
  12575=>"000110111",
  12576=>"000000001",
  12577=>"011111000",
  12578=>"000110010",
  12579=>"100110000",
  12580=>"000001000",
  12581=>"111001001",
  12582=>"001111111",
  12583=>"000000000",
  12584=>"111111010",
  12585=>"011110001",
  12586=>"111101101",
  12587=>"101001111",
  12588=>"111111100",
  12589=>"000101111",
  12590=>"000000100",
  12591=>"010000100",
  12592=>"000001101",
  12593=>"101001001",
  12594=>"000000000",
  12595=>"101001001",
  12596=>"000110101",
  12597=>"110000000",
  12598=>"011111110",
  12599=>"000000001",
  12600=>"111001000",
  12601=>"000000111",
  12602=>"101100101",
  12603=>"000001110",
  12604=>"100100100",
  12605=>"110111101",
  12606=>"000100111",
  12607=>"011001010",
  12608=>"101101001",
  12609=>"111001001",
  12610=>"000010000",
  12611=>"100110101",
  12612=>"011000001",
  12613=>"000001000",
  12614=>"111111101",
  12615=>"111111111",
  12616=>"110110011",
  12617=>"111110001",
  12618=>"000000111",
  12619=>"010101000",
  12620=>"000000111",
  12621=>"001101110",
  12622=>"011001000",
  12623=>"101010111",
  12624=>"010010110",
  12625=>"111000000",
  12626=>"111111110",
  12627=>"001001011",
  12628=>"010010000",
  12629=>"100010011",
  12630=>"000000100",
  12631=>"110001001",
  12632=>"000000000",
  12633=>"100100000",
  12634=>"000110111",
  12635=>"101100001",
  12636=>"101000101",
  12637=>"000001011",
  12638=>"111011000",
  12639=>"010000000",
  12640=>"010110111",
  12641=>"010000100",
  12642=>"010010000",
  12643=>"100001111",
  12644=>"100101001",
  12645=>"011001101",
  12646=>"111001000",
  12647=>"001111111",
  12648=>"000000000",
  12649=>"101000000",
  12650=>"111110111",
  12651=>"111101000",
  12652=>"001000000",
  12653=>"010011111",
  12654=>"000000101",
  12655=>"110000001",
  12656=>"110110101",
  12657=>"111001000",
  12658=>"111111010",
  12659=>"001001111",
  12660=>"100000000",
  12661=>"000001001",
  12662=>"000100111",
  12663=>"111110000",
  12664=>"011001000",
  12665=>"010000111",
  12666=>"000001111",
  12667=>"111000010",
  12668=>"100110110",
  12669=>"100000100",
  12670=>"010111010",
  12671=>"000000010",
  12672=>"001000000",
  12673=>"111000000",
  12674=>"111111000",
  12675=>"001111000",
  12676=>"111110000",
  12677=>"001000111",
  12678=>"110001000",
  12679=>"000000100",
  12680=>"011011011",
  12681=>"010010000",
  12682=>"000001111",
  12683=>"100001000",
  12684=>"010110000",
  12685=>"101010000",
  12686=>"111111101",
  12687=>"000000001",
  12688=>"110110111",
  12689=>"011111011",
  12690=>"101101101",
  12691=>"101100000",
  12692=>"001111101",
  12693=>"000000000",
  12694=>"111101000",
  12695=>"000011110",
  12696=>"111111001",
  12697=>"000110110",
  12698=>"011111001",
  12699=>"000010000",
  12700=>"001111010",
  12701=>"010000001",
  12702=>"000100111",
  12703=>"000000101",
  12704=>"000100110",
  12705=>"100000000",
  12706=>"010101111",
  12707=>"111000000",
  12708=>"010000011",
  12709=>"001001010",
  12710=>"011110100",
  12711=>"000101111",
  12712=>"000111111",
  12713=>"000110110",
  12714=>"000110011",
  12715=>"010000000",
  12716=>"111010000",
  12717=>"000000111",
  12718=>"100100101",
  12719=>"110110111",
  12720=>"000000010",
  12721=>"010011001",
  12722=>"111000000",
  12723=>"000100110",
  12724=>"111111011",
  12725=>"111000000",
  12726=>"111111011",
  12727=>"111111000",
  12728=>"001001001",
  12729=>"000010010",
  12730=>"111111111",
  12731=>"111100111",
  12732=>"000000100",
  12733=>"110110111",
  12734=>"011000000",
  12735=>"110110000",
  12736=>"001011000",
  12737=>"001000111",
  12738=>"101111111",
  12739=>"101001010",
  12740=>"011011001",
  12741=>"000001101",
  12742=>"000000011",
  12743=>"111100110",
  12744=>"111101000",
  12745=>"010110110",
  12746=>"101111000",
  12747=>"111000000",
  12748=>"000000111",
  12749=>"001011111",
  12750=>"000000111",
  12751=>"000000111",
  12752=>"000000000",
  12753=>"011000011",
  12754=>"101000011",
  12755=>"000000101",
  12756=>"110110000",
  12757=>"110100111",
  12758=>"001000111",
  12759=>"110000111",
  12760=>"111111010",
  12761=>"000101001",
  12762=>"111010001",
  12763=>"000010000",
  12764=>"101100111",
  12765=>"101111000",
  12766=>"111110000",
  12767=>"111111000",
  12768=>"000000100",
  12769=>"000000101",
  12770=>"111110010",
  12771=>"000111011",
  12772=>"101001111",
  12773=>"000010000",
  12774=>"000000101",
  12775=>"001000000",
  12776=>"000000000",
  12777=>"000010111",
  12778=>"001000101",
  12779=>"111111110",
  12780=>"000010111",
  12781=>"000001001",
  12782=>"000000000",
  12783=>"111000000",
  12784=>"100100011",
  12785=>"000011111",
  12786=>"011000101",
  12787=>"111000100",
  12788=>"100110101",
  12789=>"000000010",
  12790=>"000001000",
  12791=>"001000101",
  12792=>"111111000",
  12793=>"110000010",
  12794=>"101000110",
  12795=>"001011001",
  12796=>"111101000",
  12797=>"111010001",
  12798=>"100100111",
  12799=>"111111001",
  12800=>"111011000",
  12801=>"110011111",
  12802=>"100000000",
  12803=>"000000111",
  12804=>"001011011",
  12805=>"000001001",
  12806=>"000010000",
  12807=>"011011111",
  12808=>"001011110",
  12809=>"011010000",
  12810=>"011011000",
  12811=>"000100111",
  12812=>"000000111",
  12813=>"000000101",
  12814=>"100011001",
  12815=>"000001111",
  12816=>"011010000",
  12817=>"011111000",
  12818=>"101111100",
  12819=>"000111101",
  12820=>"111011000",
  12821=>"111110000",
  12822=>"010011001",
  12823=>"111111010",
  12824=>"010010110",
  12825=>"111111111",
  12826=>"111011000",
  12827=>"011010000",
  12828=>"100100101",
  12829=>"111010000",
  12830=>"000011011",
  12831=>"000000010",
  12832=>"000000101",
  12833=>"011000111",
  12834=>"111011010",
  12835=>"111011011",
  12836=>"001001000",
  12837=>"000110001",
  12838=>"110010000",
  12839=>"111000000",
  12840=>"111011000",
  12841=>"011000001",
  12842=>"011000000",
  12843=>"000000010",
  12844=>"110100000",
  12845=>"111011011",
  12846=>"111011000",
  12847=>"010000000",
  12848=>"000111111",
  12849=>"001001001",
  12850=>"111111011",
  12851=>"000010111",
  12852=>"111011000",
  12853=>"111111111",
  12854=>"010011100",
  12855=>"000110000",
  12856=>"011111110",
  12857=>"001101111",
  12858=>"000100101",
  12859=>"100000000",
  12860=>"000100101",
  12861=>"111111010",
  12862=>"000000000",
  12863=>"111111000",
  12864=>"001000111",
  12865=>"010011000",
  12866=>"000010000",
  12867=>"111111010",
  12868=>"101100101",
  12869=>"010000100",
  12870=>"000000101",
  12871=>"000000100",
  12872=>"001111111",
  12873=>"010111000",
  12874=>"010000101",
  12875=>"000000101",
  12876=>"111111000",
  12877=>"100100110",
  12878=>"100100100",
  12879=>"001000101",
  12880=>"101011011",
  12881=>"000111010",
  12882=>"000010011",
  12883=>"011111000",
  12884=>"000011010",
  12885=>"110110011",
  12886=>"000100110",
  12887=>"011111000",
  12888=>"111001010",
  12889=>"111001001",
  12890=>"100100000",
  12891=>"000000000",
  12892=>"010011000",
  12893=>"001001001",
  12894=>"010000011",
  12895=>"111001000",
  12896=>"100010000",
  12897=>"111111000",
  12898=>"100000100",
  12899=>"100100110",
  12900=>"000100001",
  12901=>"111010100",
  12902=>"111010000",
  12903=>"011111000",
  12904=>"000011111",
  12905=>"000010011",
  12906=>"000000000",
  12907=>"000000111",
  12908=>"100111110",
  12909=>"111111010",
  12910=>"101100100",
  12911=>"111101111",
  12912=>"000001101",
  12913=>"000000010",
  12914=>"011010000",
  12915=>"010000000",
  12916=>"010000000",
  12917=>"000000111",
  12918=>"111111101",
  12919=>"000000000",
  12920=>"111001010",
  12921=>"000100111",
  12922=>"010000000",
  12923=>"100101100",
  12924=>"110000000",
  12925=>"111100000",
  12926=>"111110000",
  12927=>"111111001",
  12928=>"011010000",
  12929=>"000111111",
  12930=>"010010000",
  12931=>"111001011",
  12932=>"001010010",
  12933=>"000000100",
  12934=>"000010100",
  12935=>"000001001",
  12936=>"101111111",
  12937=>"100101010",
  12938=>"011001100",
  12939=>"000010000",
  12940=>"111011000",
  12941=>"101100101",
  12942=>"010011000",
  12943=>"000000001",
  12944=>"011011000",
  12945=>"000111001",
  12946=>"010010000",
  12947=>"000000011",
  12948=>"100000011",
  12949=>"011011000",
  12950=>"000000001",
  12951=>"011001100",
  12952=>"000000000",
  12953=>"000000111",
  12954=>"000000000",
  12955=>"000000110",
  12956=>"111110000",
  12957=>"101000100",
  12958=>"011000000",
  12959=>"010010000",
  12960=>"111111001",
  12961=>"010111010",
  12962=>"010011000",
  12963=>"000111111",
  12964=>"001101111",
  12965=>"111101100",
  12966=>"111110000",
  12967=>"001111010",
  12968=>"010010010",
  12969=>"001111111",
  12970=>"000100100",
  12971=>"111010000",
  12972=>"011010111",
  12973=>"111010000",
  12974=>"100111000",
  12975=>"000100111",
  12976=>"001010100",
  12977=>"001111111",
  12978=>"000000110",
  12979=>"110100010",
  12980=>"111110011",
  12981=>"010111000",
  12982=>"111011001",
  12983=>"100000101",
  12984=>"100100100",
  12985=>"100000010",
  12986=>"000000100",
  12987=>"001111001",
  12988=>"000000000",
  12989=>"100111111",
  12990=>"110011001",
  12991=>"011010000",
  12992=>"111000001",
  12993=>"101101011",
  12994=>"010110011",
  12995=>"101100100",
  12996=>"100101000",
  12997=>"100000001",
  12998=>"000001011",
  12999=>"111000100",
  13000=>"111111111",
  13001=>"010011010",
  13002=>"000000000",
  13003=>"100000101",
  13004=>"000011000",
  13005=>"011110100",
  13006=>"000000000",
  13007=>"010010000",
  13008=>"000000000",
  13009=>"111100100",
  13010=>"000100111",
  13011=>"111111011",
  13012=>"100101111",
  13013=>"100111110",
  13014=>"000000000",
  13015=>"100111111",
  13016=>"000011010",
  13017=>"010011111",
  13018=>"010000100",
  13019=>"000000000",
  13020=>"000111101",
  13021=>"000111111",
  13022=>"111101111",
  13023=>"000000111",
  13024=>"111111010",
  13025=>"000100110",
  13026=>"111100010",
  13027=>"111110000",
  13028=>"000000000",
  13029=>"000000110",
  13030=>"010000111",
  13031=>"100100111",
  13032=>"000111111",
  13033=>"011011111",
  13034=>"110011001",
  13035=>"111101011",
  13036=>"011111010",
  13037=>"100000011",
  13038=>"000110000",
  13039=>"110000000",
  13040=>"000000010",
  13041=>"001000101",
  13042=>"001001010",
  13043=>"011011000",
  13044=>"111110001",
  13045=>"110001010",
  13046=>"000000000",
  13047=>"000011111",
  13048=>"000000010",
  13049=>"001111111",
  13050=>"111101111",
  13051=>"011111111",
  13052=>"000000101",
  13053=>"000100000",
  13054=>"100111111",
  13055=>"000000000",
  13056=>"100000000",
  13057=>"000100000",
  13058=>"110000000",
  13059=>"000000111",
  13060=>"000001011",
  13061=>"110000001",
  13062=>"111101010",
  13063=>"111000001",
  13064=>"000101101",
  13065=>"010110000",
  13066=>"111111010",
  13067=>"000110000",
  13068=>"000111101",
  13069=>"000010000",
  13070=>"111011010",
  13071=>"000111111",
  13072=>"000010110",
  13073=>"000111111",
  13074=>"000000000",
  13075=>"110111111",
  13076=>"101000010",
  13077=>"001111111",
  13078=>"011100000",
  13079=>"000111111",
  13080=>"001001000",
  13081=>"000100111",
  13082=>"000000111",
  13083=>"001000000",
  13084=>"000111111",
  13085=>"000100000",
  13086=>"111110000",
  13087=>"101000000",
  13088=>"001100001",
  13089=>"000000000",
  13090=>"111010010",
  13091=>"000000111",
  13092=>"111000001",
  13093=>"000000001",
  13094=>"000000111",
  13095=>"111111111",
  13096=>"000111010",
  13097=>"000000000",
  13098=>"111011111",
  13099=>"000111000",
  13100=>"111011111",
  13101=>"000111111",
  13102=>"101001001",
  13103=>"000001110",
  13104=>"000101111",
  13105=>"010000001",
  13106=>"000000101",
  13107=>"110011111",
  13108=>"001000000",
  13109=>"000110101",
  13110=>"100111011",
  13111=>"111000100",
  13112=>"110000000",
  13113=>"111000100",
  13114=>"001101011",
  13115=>"001000000",
  13116=>"000010011",
  13117=>"011001010",
  13118=>"110100000",
  13119=>"111110000",
  13120=>"000000111",
  13121=>"111010000",
  13122=>"111111101",
  13123=>"011100110",
  13124=>"111111001",
  13125=>"001111101",
  13126=>"100000000",
  13127=>"011000000",
  13128=>"100111100",
  13129=>"110111000",
  13130=>"111111010",
  13131=>"111010000",
  13132=>"010000000",
  13133=>"010010110",
  13134=>"111101100",
  13135=>"110110111",
  13136=>"111000000",
  13137=>"101000000",
  13138=>"011111111",
  13139=>"011000000",
  13140=>"000000010",
  13141=>"011000000",
  13142=>"111011000",
  13143=>"111111110",
  13144=>"111111011",
  13145=>"010011001",
  13146=>"111110000",
  13147=>"111010001",
  13148=>"000000000",
  13149=>"111100000",
  13150=>"001111111",
  13151=>"100001111",
  13152=>"101111101",
  13153=>"111110000",
  13154=>"000000000",
  13155=>"011101000",
  13156=>"010000000",
  13157=>"110000000",
  13158=>"000001111",
  13159=>"111101111",
  13160=>"111101000",
  13161=>"101110111",
  13162=>"011000000",
  13163=>"001001001",
  13164=>"000000000",
  13165=>"111111111",
  13166=>"010111011",
  13167=>"111111100",
  13168=>"101000001",
  13169=>"000000111",
  13170=>"001111111",
  13171=>"000000111",
  13172=>"100111010",
  13173=>"000000100",
  13174=>"111111000",
  13175=>"000001000",
  13176=>"000101100",
  13177=>"110010111",
  13178=>"111110011",
  13179=>"000000100",
  13180=>"111111100",
  13181=>"100000001",
  13182=>"001111010",
  13183=>"111000000",
  13184=>"010011000",
  13185=>"010010000",
  13186=>"000000111",
  13187=>"000111000",
  13188=>"000000111",
  13189=>"111000000",
  13190=>"000000100",
  13191=>"110000100",
  13192=>"110111010",
  13193=>"111100111",
  13194=>"111011111",
  13195=>"000000100",
  13196=>"111101000",
  13197=>"101101111",
  13198=>"111000000",
  13199=>"000010000",
  13200=>"101101011",
  13201=>"010011000",
  13202=>"111010010",
  13203=>"001100000",
  13204=>"000000010",
  13205=>"001011000",
  13206=>"111110101",
  13207=>"000000001",
  13208=>"001101111",
  13209=>"101000110",
  13210=>"000000111",
  13211=>"010000000",
  13212=>"111010001",
  13213=>"000000000",
  13214=>"000000110",
  13215=>"111000000",
  13216=>"011001101",
  13217=>"010111000",
  13218=>"000101111",
  13219=>"111000000",
  13220=>"001111100",
  13221=>"111110110",
  13222=>"111001001",
  13223=>"110010111",
  13224=>"010111111",
  13225=>"010000000",
  13226=>"000000000",
  13227=>"111001000",
  13228=>"000110010",
  13229=>"111000000",
  13230=>"010100000",
  13231=>"111110101",
  13232=>"000110111",
  13233=>"111110001",
  13234=>"010000101",
  13235=>"011011100",
  13236=>"100110111",
  13237=>"001111101",
  13238=>"000111111",
  13239=>"000101101",
  13240=>"100000110",
  13241=>"110000100",
  13242=>"000000110",
  13243=>"001111110",
  13244=>"000001111",
  13245=>"111111111",
  13246=>"001011010",
  13247=>"101000111",
  13248=>"110000011",
  13249=>"111000000",
  13250=>"000111111",
  13251=>"011001000",
  13252=>"001000100",
  13253=>"101000000",
  13254=>"100111111",
  13255=>"101001000",
  13256=>"110000000",
  13257=>"000111010",
  13258=>"000110010",
  13259=>"000000111",
  13260=>"000111000",
  13261=>"001001110",
  13262=>"111001000",
  13263=>"000000110",
  13264=>"000011111",
  13265=>"110000001",
  13266=>"111000110",
  13267=>"000110111",
  13268=>"101000000",
  13269=>"111000000",
  13270=>"000000000",
  13271=>"000000000",
  13272=>"000111111",
  13273=>"000111110",
  13274=>"010100000",
  13275=>"111111000",
  13276=>"000010001",
  13277=>"100111111",
  13278=>"100110010",
  13279=>"000000101",
  13280=>"010111000",
  13281=>"111000000",
  13282=>"001000100",
  13283=>"111000000",
  13284=>"011000000",
  13285=>"110000000",
  13286=>"010000000",
  13287=>"110000100",
  13288=>"000010110",
  13289=>"001111100",
  13290=>"111110010",
  13291=>"000111111",
  13292=>"000111111",
  13293=>"000100111",
  13294=>"111000000",
  13295=>"000000100",
  13296=>"000010010",
  13297=>"111110010",
  13298=>"001011000",
  13299=>"111111000",
  13300=>"011010000",
  13301=>"111101000",
  13302=>"010000011",
  13303=>"011100110",
  13304=>"000000001",
  13305=>"001111111",
  13306=>"000000111",
  13307=>"111000000",
  13308=>"010010001",
  13309=>"000000000",
  13310=>"111101111",
  13311=>"000101101",
  13312=>"100100111",
  13313=>"111100110",
  13314=>"010111111",
  13315=>"111000000",
  13316=>"110011111",
  13317=>"100001000",
  13318=>"100111111",
  13319=>"000000010",
  13320=>"000011011",
  13321=>"000111000",
  13322=>"111101111",
  13323=>"010011010",
  13324=>"000010000",
  13325=>"000000000",
  13326=>"110110100",
  13327=>"111000100",
  13328=>"000001011",
  13329=>"000100101",
  13330=>"001111111",
  13331=>"111100111",
  13332=>"100011000",
  13333=>"010000101",
  13334=>"111011101",
  13335=>"111000000",
  13336=>"000011011",
  13337=>"000010010",
  13338=>"000001000",
  13339=>"110111111",
  13340=>"011011111",
  13341=>"000100000",
  13342=>"000000111",
  13343=>"000101000",
  13344=>"110001000",
  13345=>"000000000",
  13346=>"111100111",
  13347=>"111001010",
  13348=>"111010100",
  13349=>"000001011",
  13350=>"110110010",
  13351=>"001000000",
  13352=>"000000000",
  13353=>"100000111",
  13354=>"111111111",
  13355=>"111011111",
  13356=>"111011000",
  13357=>"000000000",
  13358=>"100000111",
  13359=>"000000101",
  13360=>"000000100",
  13361=>"110110110",
  13362=>"111011111",
  13363=>"111100100",
  13364=>"111100111",
  13365=>"000110110",
  13366=>"110111011",
  13367=>"110100100",
  13368=>"100100110",
  13369=>"000100000",
  13370=>"011111011",
  13371=>"100101100",
  13372=>"000000001",
  13373=>"000100111",
  13374=>"000111010",
  13375=>"011000100",
  13376=>"000111111",
  13377=>"000000110",
  13378=>"000111010",
  13379=>"001110111",
  13380=>"010111011",
  13381=>"000000010",
  13382=>"110010010",
  13383=>"010011110",
  13384=>"010110010",
  13385=>"110010001",
  13386=>"100100111",
  13387=>"101101101",
  13388=>"010010000",
  13389=>"011011011",
  13390=>"011011001",
  13391=>"000100000",
  13392=>"101000000",
  13393=>"011111111",
  13394=>"110000010",
  13395=>"100010011",
  13396=>"000000000",
  13397=>"000011011",
  13398=>"011110010",
  13399=>"110000000",
  13400=>"000110000",
  13401=>"010011000",
  13402=>"010000000",
  13403=>"011010110",
  13404=>"000000000",
  13405=>"111010000",
  13406=>"000000000",
  13407=>"111111111",
  13408=>"000010000",
  13409=>"010010000",
  13410=>"011111010",
  13411=>"011000000",
  13412=>"001010011",
  13413=>"000001000",
  13414=>"010110000",
  13415=>"010011011",
  13416=>"000100000",
  13417=>"000000000",
  13418=>"111011000",
  13419=>"000011000",
  13420=>"000101011",
  13421=>"101111111",
  13422=>"111000100",
  13423=>"111111000",
  13424=>"011000000",
  13425=>"100100100",
  13426=>"011111110",
  13427=>"110011010",
  13428=>"010100000",
  13429=>"000000010",
  13430=>"000000101",
  13431=>"000010000",
  13432=>"111000110",
  13433=>"011011000",
  13434=>"111111111",
  13435=>"111010111",
  13436=>"010000100",
  13437=>"011011011",
  13438=>"011101111",
  13439=>"010110111",
  13440=>"010111010",
  13441=>"011101100",
  13442=>"000101111",
  13443=>"000111100",
  13444=>"100111111",
  13445=>"011111010",
  13446=>"000100010",
  13447=>"011110110",
  13448=>"011010010",
  13449=>"000111011",
  13450=>"001000000",
  13451=>"000000110",
  13452=>"000000000",
  13453=>"010010000",
  13454=>"101000001",
  13455=>"011010110",
  13456=>"011010010",
  13457=>"110000000",
  13458=>"101000000",
  13459=>"010111011",
  13460=>"010110000",
  13461=>"000111011",
  13462=>"111111100",
  13463=>"010110011",
  13464=>"011101110",
  13465=>"000000000",
  13466=>"110100110",
  13467=>"111111111",
  13468=>"011011010",
  13469=>"010011011",
  13470=>"011101111",
  13471=>"000011010",
  13472=>"011011011",
  13473=>"000000000",
  13474=>"111010000",
  13475=>"111111000",
  13476=>"101100000",
  13477=>"011010010",
  13478=>"011000111",
  13479=>"000000100",
  13480=>"100100101",
  13481=>"111110110",
  13482=>"000000000",
  13483=>"101101111",
  13484=>"001001000",
  13485=>"010111011",
  13486=>"001000000",
  13487=>"101111010",
  13488=>"000001111",
  13489=>"010011111",
  13490=>"000011010",
  13491=>"111111000",
  13492=>"001000000",
  13493=>"111100110",
  13494=>"000001011",
  13495=>"111000010",
  13496=>"001110000",
  13497=>"001001001",
  13498=>"000000010",
  13499=>"111111110",
  13500=>"000000000",
  13501=>"111111111",
  13502=>"110010010",
  13503=>"000110000",
  13504=>"010111010",
  13505=>"001000000",
  13506=>"000000100",
  13507=>"111000011",
  13508=>"111111111",
  13509=>"011000111",
  13510=>"011110000",
  13511=>"001011111",
  13512=>"111000000",
  13513=>"000011111",
  13514=>"101111100",
  13515=>"000010000",
  13516=>"010011010",
  13517=>"010100100",
  13518=>"111010111",
  13519=>"000000001",
  13520=>"100011001",
  13521=>"011010000",
  13522=>"111111000",
  13523=>"000010011",
  13524=>"000000101",
  13525=>"000000010",
  13526=>"000010000",
  13527=>"010000100",
  13528=>"011000000",
  13529=>"111100000",
  13530=>"011011011",
  13531=>"000111111",
  13532=>"001111110",
  13533=>"000101100",
  13534=>"111111010",
  13535=>"111101110",
  13536=>"100111110",
  13537=>"000000111",
  13538=>"000000010",
  13539=>"011011111",
  13540=>"101100000",
  13541=>"010111011",
  13542=>"111110100",
  13543=>"100000000",
  13544=>"011000000",
  13545=>"111100101",
  13546=>"101101100",
  13547=>"101000100",
  13548=>"100100111",
  13549=>"100111111",
  13550=>"001111111",
  13551=>"101000000",
  13552=>"010100000",
  13553=>"010111111",
  13554=>"111111100",
  13555=>"110000000",
  13556=>"101011011",
  13557=>"000000000",
  13558=>"000010000",
  13559=>"011011111",
  13560=>"111111000",
  13561=>"101100100",
  13562=>"111110111",
  13563=>"001000000",
  13564=>"011111111",
  13565=>"100000000",
  13566=>"011011111",
  13567=>"100000000",
  13568=>"000001110",
  13569=>"001000111",
  13570=>"000001111",
  13571=>"011000101",
  13572=>"100100111",
  13573=>"001000001",
  13574=>"010000010",
  13575=>"111100111",
  13576=>"100111110",
  13577=>"000010000",
  13578=>"110001000",
  13579=>"001001101",
  13580=>"000000011",
  13581=>"000001000",
  13582=>"000100000",
  13583=>"101101111",
  13584=>"010100001",
  13585=>"111000111",
  13586=>"101000010",
  13587=>"110000000",
  13588=>"111111110",
  13589=>"001101111",
  13590=>"111011000",
  13591=>"111111101",
  13592=>"010001101",
  13593=>"000000111",
  13594=>"111110100",
  13595=>"001000000",
  13596=>"101101010",
  13597=>"101000000",
  13598=>"000010111",
  13599=>"110101101",
  13600=>"000000001",
  13601=>"001001001",
  13602=>"000000001",
  13603=>"100100110",
  13604=>"100000111",
  13605=>"001000100",
  13606=>"001111110",
  13607=>"110010000",
  13608=>"100111000",
  13609=>"001110100",
  13610=>"001101100",
  13611=>"001101111",
  13612=>"010000000",
  13613=>"111000111",
  13614=>"101000000",
  13615=>"011111011",
  13616=>"110000000",
  13617=>"000110111",
  13618=>"111111001",
  13619=>"111110100",
  13620=>"111010000",
  13621=>"111000000",
  13622=>"011000001",
  13623=>"101111111",
  13624=>"000001101",
  13625=>"100000000",
  13626=>"111011000",
  13627=>"111010100",
  13628=>"010011001",
  13629=>"011000000",
  13630=>"111001000",
  13631=>"111001110",
  13632=>"001010100",
  13633=>"001111111",
  13634=>"000010011",
  13635=>"100000001",
  13636=>"000111111",
  13637=>"100101001",
  13638=>"001000111",
  13639=>"111001000",
  13640=>"011101101",
  13641=>"111001001",
  13642=>"001011111",
  13643=>"111111100",
  13644=>"001001010",
  13645=>"001001011",
  13646=>"011111110",
  13647=>"111000110",
  13648=>"011011111",
  13649=>"110000011",
  13650=>"110000001",
  13651=>"010000000",
  13652=>"001001000",
  13653=>"011000011",
  13654=>"100110110",
  13655=>"101101011",
  13656=>"001111111",
  13657=>"011101100",
  13658=>"011011111",
  13659=>"011001000",
  13660=>"110110111",
  13661=>"010110110",
  13662=>"110111000",
  13663=>"111100011",
  13664=>"000111000",
  13665=>"111111001",
  13666=>"000101111",
  13667=>"001100100",
  13668=>"101101111",
  13669=>"111010000",
  13670=>"111000000",
  13671=>"011111110",
  13672=>"000110110",
  13673=>"001010000",
  13674=>"110110110",
  13675=>"001101111",
  13676=>"001001111",
  13677=>"000000011",
  13678=>"001011111",
  13679=>"011001000",
  13680=>"101111001",
  13681=>"110111100",
  13682=>"110110000",
  13683=>"010000001",
  13684=>"001111111",
  13685=>"101111100",
  13686=>"100011010",
  13687=>"001001111",
  13688=>"110110001",
  13689=>"110110000",
  13690=>"000101111",
  13691=>"010111111",
  13692=>"110000011",
  13693=>"101010110",
  13694=>"111001001",
  13695=>"000000000",
  13696=>"001000000",
  13697=>"000000111",
  13698=>"100100100",
  13699=>"000100001",
  13700=>"000100111",
  13701=>"110100001",
  13702=>"000110010",
  13703=>"000001010",
  13704=>"001011111",
  13705=>"110110000",
  13706=>"111111000",
  13707=>"000101011",
  13708=>"001111111",
  13709=>"001101111",
  13710=>"001100000",
  13711=>"001100100",
  13712=>"100000011",
  13713=>"111110011",
  13714=>"001000000",
  13715=>"001000000",
  13716=>"101001000",
  13717=>"101110000",
  13718=>"110000000",
  13719=>"100100111",
  13720=>"000000001",
  13721=>"000111111",
  13722=>"100111111",
  13723=>"111000010",
  13724=>"110010000",
  13725=>"101100000",
  13726=>"000000000",
  13727=>"011000100",
  13728=>"111011110",
  13729=>"111000101",
  13730=>"111000011",
  13731=>"110010000",
  13732=>"110111011",
  13733=>"100100100",
  13734=>"011111001",
  13735=>"000101011",
  13736=>"111110010",
  13737=>"111111111",
  13738=>"001111111",
  13739=>"111001101",
  13740=>"110011011",
  13741=>"101111111",
  13742=>"110100111",
  13743=>"000000000",
  13744=>"001000001",
  13745=>"000010111",
  13746=>"111000000",
  13747=>"001101110",
  13748=>"111010110",
  13749=>"010010000",
  13750=>"010101100",
  13751=>"000001001",
  13752=>"110110100",
  13753=>"010000100",
  13754=>"110110000",
  13755=>"110000000",
  13756=>"011010000",
  13757=>"101001111",
  13758=>"000010010",
  13759=>"011110000",
  13760=>"001000010",
  13761=>"111010100",
  13762=>"001000000",
  13763=>"000110100",
  13764=>"010110000",
  13765=>"100101110",
  13766=>"001111101",
  13767=>"111101000",
  13768=>"110101000",
  13769=>"011011011",
  13770=>"001001001",
  13771=>"001111111",
  13772=>"000000100",
  13773=>"111001101",
  13774=>"000001001",
  13775=>"011111101",
  13776=>"110001001",
  13777=>"010111110",
  13778=>"110100110",
  13779=>"110100000",
  13780=>"000000000",
  13781=>"001001111",
  13782=>"101000000",
  13783=>"110000000",
  13784=>"101111111",
  13785=>"110100000",
  13786=>"010010000",
  13787=>"101110111",
  13788=>"010010000",
  13789=>"001101111",
  13790=>"000110000",
  13791=>"110001001",
  13792=>"000010010",
  13793=>"111101101",
  13794=>"110110010",
  13795=>"111100100",
  13796=>"111010000",
  13797=>"001000100",
  13798=>"100000000",
  13799=>"000111111",
  13800=>"001001001",
  13801=>"000011001",
  13802=>"011000000",
  13803=>"111101001",
  13804=>"001111011",
  13805=>"000001101",
  13806=>"001000010",
  13807=>"111111110",
  13808=>"000001100",
  13809=>"011011001",
  13810=>"110111000",
  13811=>"100000000",
  13812=>"000000011",
  13813=>"010110110",
  13814=>"000000000",
  13815=>"000010000",
  13816=>"000000110",
  13817=>"000000000",
  13818=>"000001110",
  13819=>"111001000",
  13820=>"111110010",
  13821=>"000110010",
  13822=>"011101001",
  13823=>"000000011",
  13824=>"011111100",
  13825=>"111000010",
  13826=>"000000001",
  13827=>"000000000",
  13828=>"000111000",
  13829=>"011001111",
  13830=>"000001111",
  13831=>"011000010",
  13832=>"001000010",
  13833=>"000000001",
  13834=>"100110011",
  13835=>"100001100",
  13836=>"000000101",
  13837=>"010111101",
  13838=>"100011110",
  13839=>"111110100",
  13840=>"001000001",
  13841=>"010010000",
  13842=>"000000010",
  13843=>"010110111",
  13844=>"000001000",
  13845=>"000000101",
  13846=>"010111001",
  13847=>"111111110",
  13848=>"000000000",
  13849=>"111011111",
  13850=>"110011111",
  13851=>"111011001",
  13852=>"111000001",
  13853=>"111000000",
  13854=>"000101101",
  13855=>"000001011",
  13856=>"001111111",
  13857=>"000011111",
  13858=>"111000001",
  13859=>"000000000",
  13860=>"110100100",
  13861=>"111111011",
  13862=>"011010111",
  13863=>"101100000",
  13864=>"110010111",
  13865=>"100000011",
  13866=>"000111110",
  13867=>"111011000",
  13868=>"011000000",
  13869=>"000000000",
  13870=>"010001110",
  13871=>"111001111",
  13872=>"111001000",
  13873=>"110101001",
  13874=>"100000000",
  13875=>"111000111",
  13876=>"101000111",
  13877=>"111111011",
  13878=>"110011011",
  13879=>"111001000",
  13880=>"001001111",
  13881=>"000101010",
  13882=>"001001000",
  13883=>"010000101",
  13884=>"111011010",
  13885=>"011010000",
  13886=>"000001011",
  13887=>"100001000",
  13888=>"111111111",
  13889=>"111111001",
  13890=>"101001011",
  13891=>"000000011",
  13892=>"110110000",
  13893=>"101110110",
  13894=>"011111010",
  13895=>"101100111",
  13896=>"000000110",
  13897=>"111000111",
  13898=>"101001001",
  13899=>"001100111",
  13900=>"000000111",
  13901=>"011111001",
  13902=>"001001101",
  13903=>"111000011",
  13904=>"101111001",
  13905=>"000111011",
  13906=>"000111111",
  13907=>"001001000",
  13908=>"101100000",
  13909=>"111110011",
  13910=>"001001100",
  13911=>"100000000",
  13912=>"111011111",
  13913=>"000000011",
  13914=>"110101000",
  13915=>"000010110",
  13916=>"111111010",
  13917=>"100100100",
  13918=>"110110000",
  13919=>"001010100",
  13920=>"111111111",
  13921=>"000000000",
  13922=>"001111111",
  13923=>"111110010",
  13924=>"000001011",
  13925=>"000000111",
  13926=>"001111111",
  13927=>"000000111",
  13928=>"001101000",
  13929=>"111000111",
  13930=>"000110110",
  13931=>"001111111",
  13932=>"111001001",
  13933=>"111111100",
  13934=>"101101000",
  13935=>"101001001",
  13936=>"000010000",
  13937=>"000111111",
  13938=>"000110110",
  13939=>"000000100",
  13940=>"000000110",
  13941=>"000000000",
  13942=>"001001000",
  13943=>"000000101",
  13944=>"000100110",
  13945=>"111000000",
  13946=>"000000111",
  13947=>"000101000",
  13948=>"111001000",
  13949=>"101000011",
  13950=>"000000111",
  13951=>"001001001",
  13952=>"111101101",
  13953=>"001011001",
  13954=>"000110111",
  13955=>"000000011",
  13956=>"000000000",
  13957=>"000111010",
  13958=>"111100100",
  13959=>"110000011",
  13960=>"000000111",
  13961=>"000000001",
  13962=>"010010011",
  13963=>"000110101",
  13964=>"010110000",
  13965=>"111111101",
  13966=>"000111111",
  13967=>"000000001",
  13968=>"111100111",
  13969=>"101000000",
  13970=>"000000101",
  13971=>"001000101",
  13972=>"000000100",
  13973=>"000001010",
  13974=>"111010110",
  13975=>"000110110",
  13976=>"000001101",
  13977=>"111001000",
  13978=>"011011000",
  13979=>"000000010",
  13980=>"000000111",
  13981=>"000111000",
  13982=>"000111010",
  13983=>"000001000",
  13984=>"000011011",
  13985=>"010111111",
  13986=>"001111010",
  13987=>"000011111",
  13988=>"000110010",
  13989=>"001001110",
  13990=>"000010111",
  13991=>"101101101",
  13992=>"110010001",
  13993=>"101101011",
  13994=>"110111111",
  13995=>"000000001",
  13996=>"011000101",
  13997=>"001000011",
  13998=>"111111010",
  13999=>"000111101",
  14000=>"111101000",
  14001=>"111110100",
  14002=>"010000000",
  14003=>"011100000",
  14004=>"100111110",
  14005=>"100110000",
  14006=>"010000111",
  14007=>"111111000",
  14008=>"111110110",
  14009=>"001001000",
  14010=>"111001110",
  14011=>"111001101",
  14012=>"001000001",
  14013=>"000110000",
  14014=>"101110101",
  14015=>"111000110",
  14016=>"110000000",
  14017=>"000010010",
  14018=>"000100100",
  14019=>"111011110",
  14020=>"000111000",
  14021=>"110001011",
  14022=>"101001001",
  14023=>"000111100",
  14024=>"000000100",
  14025=>"110001000",
  14026=>"000111100",
  14027=>"000000111",
  14028=>"101111010",
  14029=>"110101000",
  14030=>"111101000",
  14031=>"110111101",
  14032=>"011111111",
  14033=>"000111011",
  14034=>"000000100",
  14035=>"101111010",
  14036=>"000000100",
  14037=>"111110000",
  14038=>"000000101",
  14039=>"110101000",
  14040=>"010110000",
  14041=>"000001111",
  14042=>"001000101",
  14043=>"001000111",
  14044=>"110010110",
  14045=>"000001000",
  14046=>"000011100",
  14047=>"011001011",
  14048=>"000000001",
  14049=>"000000011",
  14050=>"000100110",
  14051=>"111000101",
  14052=>"000000111",
  14053=>"111111000",
  14054=>"001101010",
  14055=>"111111000",
  14056=>"101000111",
  14057=>"111000000",
  14058=>"011010110",
  14059=>"111001101",
  14060=>"000010111",
  14061=>"000010000",
  14062=>"100000000",
  14063=>"000111000",
  14064=>"000110101",
  14065=>"010001100",
  14066=>"000000000",
  14067=>"010111111",
  14068=>"100111001",
  14069=>"000001111",
  14070=>"010000110",
  14071=>"110011011",
  14072=>"011111000",
  14073=>"001000000",
  14074=>"111111111",
  14075=>"000000101",
  14076=>"111111001",
  14077=>"001010011",
  14078=>"101001000",
  14079=>"000110110",
  14080=>"011111011",
  14081=>"000000001",
  14082=>"101101101",
  14083=>"000000000",
  14084=>"011101100",
  14085=>"011111000",
  14086=>"111001001",
  14087=>"111111111",
  14088=>"111111000",
  14089=>"001000111",
  14090=>"000100110",
  14091=>"000000000",
  14092=>"110111000",
  14093=>"000000000",
  14094=>"111111011",
  14095=>"000000111",
  14096=>"010010000",
  14097=>"100111111",
  14098=>"100100111",
  14099=>"111101111",
  14100=>"000000111",
  14101=>"000000101",
  14102=>"100000000",
  14103=>"101100001",
  14104=>"111111011",
  14105=>"000111110",
  14106=>"110000000",
  14107=>"000000000",
  14108=>"101000000",
  14109=>"000111110",
  14110=>"111000000",
  14111=>"010100000",
  14112=>"001100100",
  14113=>"101000000",
  14114=>"000000000",
  14115=>"111110000",
  14116=>"000001000",
  14117=>"110111111",
  14118=>"010010000",
  14119=>"111000000",
  14120=>"100100000",
  14121=>"101111110",
  14122=>"100100100",
  14123=>"111000111",
  14124=>"101101001",
  14125=>"111010011",
  14126=>"111001000",
  14127=>"011001011",
  14128=>"100111000",
  14129=>"100100000",
  14130=>"001111011",
  14131=>"000000001",
  14132=>"000000000",
  14133=>"000000010",
  14134=>"000000000",
  14135=>"101000000",
  14136=>"111010010",
  14137=>"000100110",
  14138=>"100100000",
  14139=>"101101101",
  14140=>"100010110",
  14141=>"111010111",
  14142=>"000000111",
  14143=>"011001001",
  14144=>"100111111",
  14145=>"010111100",
  14146=>"110111010",
  14147=>"000111100",
  14148=>"010000000",
  14149=>"110010000",
  14150=>"101101111",
  14151=>"000000001",
  14152=>"011001000",
  14153=>"000111010",
  14154=>"110010001",
  14155=>"000100111",
  14156=>"101101111",
  14157=>"010111010",
  14158=>"001001001",
  14159=>"111111111",
  14160=>"000000101",
  14161=>"010111111",
  14162=>"000011100",
  14163=>"000111011",
  14164=>"000111111",
  14165=>"000000010",
  14166=>"011111000",
  14167=>"000000101",
  14168=>"111000000",
  14169=>"100100100",
  14170=>"100100000",
  14171=>"010100100",
  14172=>"010000000",
  14173=>"001001000",
  14174=>"111111000",
  14175=>"010001011",
  14176=>"111000000",
  14177=>"100001000",
  14178=>"110000111",
  14179=>"001001011",
  14180=>"000000110",
  14181=>"101111000",
  14182=>"101001100",
  14183=>"101000100",
  14184=>"000000000",
  14185=>"001100000",
  14186=>"111010111",
  14187=>"110110100",
  14188=>"110111010",
  14189=>"001111111",
  14190=>"011001111",
  14191=>"000111111",
  14192=>"011011110",
  14193=>"000000000",
  14194=>"000000100",
  14195=>"111101111",
  14196=>"101010101",
  14197=>"011000000",
  14198=>"010111100",
  14199=>"010111111",
  14200=>"110001001",
  14201=>"111111000",
  14202=>"000100111",
  14203=>"111111011",
  14204=>"101000101",
  14205=>"100100100",
  14206=>"000000011",
  14207=>"110110001",
  14208=>"000100111",
  14209=>"101111111",
  14210=>"000111100",
  14211=>"010000110",
  14212=>"000110111",
  14213=>"110111011",
  14214=>"000100000",
  14215=>"011001000",
  14216=>"100100001",
  14217=>"000000110",
  14218=>"110010000",
  14219=>"111010011",
  14220=>"001001101",
  14221=>"101101111",
  14222=>"111110010",
  14223=>"100110111",
  14224=>"100110000",
  14225=>"100000000",
  14226=>"101111111",
  14227=>"101000110",
  14228=>"101010111",
  14229=>"000000000",
  14230=>"111011010",
  14231=>"011111111",
  14232=>"111111011",
  14233=>"100010000",
  14234=>"110111111",
  14235=>"101111010",
  14236=>"110111000",
  14237=>"010010000",
  14238=>"111111010",
  14239=>"001001000",
  14240=>"110110000",
  14241=>"000111101",
  14242=>"111111010",
  14243=>"111000000",
  14244=>"001110111",
  14245=>"110001001",
  14246=>"110010001",
  14247=>"000010010",
  14248=>"000110111",
  14249=>"111111110",
  14250=>"101101000",
  14251=>"000000100",
  14252=>"111111000",
  14253=>"001111111",
  14254=>"000001001",
  14255=>"011011010",
  14256=>"001000000",
  14257=>"111011001",
  14258=>"111111000",
  14259=>"100000000",
  14260=>"101011000",
  14261=>"100000111",
  14262=>"100100000",
  14263=>"111010110",
  14264=>"001100000",
  14265=>"101100111",
  14266=>"101110110",
  14267=>"010010000",
  14268=>"101111111",
  14269=>"110110000",
  14270=>"111011000",
  14271=>"000000000",
  14272=>"000000101",
  14273=>"111101111",
  14274=>"101111001",
  14275=>"110111000",
  14276=>"000010010",
  14277=>"001101110",
  14278=>"010010000",
  14279=>"100100101",
  14280=>"111010010",
  14281=>"111011011",
  14282=>"101000000",
  14283=>"001001011",
  14284=>"111101101",
  14285=>"001101101",
  14286=>"101101101",
  14287=>"010000000",
  14288=>"010001111",
  14289=>"110110110",
  14290=>"100111111",
  14291=>"110000110",
  14292=>"000000111",
  14293=>"110110000",
  14294=>"111111000",
  14295=>"111000000",
  14296=>"000000111",
  14297=>"001000000",
  14298=>"111111000",
  14299=>"001111111",
  14300=>"001001100",
  14301=>"111111000",
  14302=>"000101101",
  14303=>"100001001",
  14304=>"110010000",
  14305=>"010111101",
  14306=>"000000101",
  14307=>"111011000",
  14308=>"111100001",
  14309=>"000000000",
  14310=>"000000010",
  14311=>"000000000",
  14312=>"111101111",
  14313=>"000000000",
  14314=>"000001011",
  14315=>"100000001",
  14316=>"010111000",
  14317=>"000000000",
  14318=>"010010000",
  14319=>"000101111",
  14320=>"101000000",
  14321=>"100001001",
  14322=>"101101110",
  14323=>"111101000",
  14324=>"010011001",
  14325=>"000000101",
  14326=>"000000100",
  14327=>"100101001",
  14328=>"000000000",
  14329=>"001011110",
  14330=>"000111111",
  14331=>"100101101",
  14332=>"110110000",
  14333=>"000000001",
  14334=>"011111001",
  14335=>"110110111",
  14336=>"101111110",
  14337=>"111111010",
  14338=>"111111100",
  14339=>"111101000",
  14340=>"111110100",
  14341=>"111111000",
  14342=>"100000000",
  14343=>"000000000",
  14344=>"001001001",
  14345=>"111111100",
  14346=>"000001011",
  14347=>"111000001",
  14348=>"000000001",
  14349=>"111010010",
  14350=>"100100000",
  14351=>"010010001",
  14352=>"001010001",
  14353=>"100000100",
  14354=>"001000000",
  14355=>"000111111",
  14356=>"000100110",
  14357=>"000000000",
  14358=>"111111011",
  14359=>"010111111",
  14360=>"101101111",
  14361=>"000000000",
  14362=>"111100111",
  14363=>"000000000",
  14364=>"000101000",
  14365=>"101101010",
  14366=>"000001000",
  14367=>"100000110",
  14368=>"111111011",
  14369=>"111111111",
  14370=>"110000000",
  14371=>"101100000",
  14372=>"010110110",
  14373=>"001000001",
  14374=>"000000111",
  14375=>"000100101",
  14376=>"111111111",
  14377=>"001001010",
  14378=>"000010011",
  14379=>"101111111",
  14380=>"000000011",
  14381=>"000000110",
  14382=>"011111110",
  14383=>"111111111",
  14384=>"111111010",
  14385=>"001000011",
  14386=>"010110000",
  14387=>"000001001",
  14388=>"111001000",
  14389=>"000000001",
  14390=>"001011011",
  14391=>"000001000",
  14392=>"000000000",
  14393=>"000001000",
  14394=>"111111110",
  14395=>"011101100",
  14396=>"011011011",
  14397=>"010111111",
  14398=>"000111111",
  14399=>"101111101",
  14400=>"000111000",
  14401=>"101111101",
  14402=>"111101111",
  14403=>"111000110",
  14404=>"000000111",
  14405=>"001101101",
  14406=>"000001000",
  14407=>"011101110",
  14408=>"100000011",
  14409=>"111000000",
  14410=>"111111111",
  14411=>"000110000",
  14412=>"000000000",
  14413=>"110100110",
  14414=>"010011011",
  14415=>"001000000",
  14416=>"111101100",
  14417=>"111111100",
  14418=>"101111110",
  14419=>"110011111",
  14420=>"111001111",
  14421=>"001000011",
  14422=>"100111111",
  14423=>"000000111",
  14424=>"111111001",
  14425=>"000100010",
  14426=>"111110011",
  14427=>"000110111",
  14428=>"111101011",
  14429=>"110110110",
  14430=>"000111000",
  14431=>"110000001",
  14432=>"001001111",
  14433=>"010000010",
  14434=>"111101101",
  14435=>"111111011",
  14436=>"011111011",
  14437=>"000000000",
  14438=>"010010000",
  14439=>"000101111",
  14440=>"101110111",
  14441=>"000000011",
  14442=>"111111010",
  14443=>"011111111",
  14444=>"000011011",
  14445=>"000111000",
  14446=>"100100000",
  14447=>"000001000",
  14448=>"110110110",
  14449=>"000010000",
  14450=>"001111011",
  14451=>"000001111",
  14452=>"111111111",
  14453=>"111110110",
  14454=>"111101000",
  14455=>"001001110",
  14456=>"111101000",
  14457=>"111101100",
  14458=>"000010010",
  14459=>"111110010",
  14460=>"011001001",
  14461=>"011111111",
  14462=>"000101111",
  14463=>"000001111",
  14464=>"111111111",
  14465=>"011111110",
  14466=>"001010010",
  14467=>"001101111",
  14468=>"111000000",
  14469=>"100111100",
  14470=>"100100110",
  14471=>"000011100",
  14472=>"000010111",
  14473=>"001001001",
  14474=>"000101111",
  14475=>"000100110",
  14476=>"011111001",
  14477=>"001000100",
  14478=>"111111011",
  14479=>"111110000",
  14480=>"100100110",
  14481=>"111000000",
  14482=>"110111001",
  14483=>"110000000",
  14484=>"000000000",
  14485=>"111111111",
  14486=>"000010000",
  14487=>"101111100",
  14488=>"000000000",
  14489=>"000011101",
  14490=>"111111110",
  14491=>"111111111",
  14492=>"000000000",
  14493=>"101011101",
  14494=>"100111111",
  14495=>"000000110",
  14496=>"100111110",
  14497=>"111011101",
  14498=>"001101011",
  14499=>"000000000",
  14500=>"111111110",
  14501=>"000110111",
  14502=>"000000110",
  14503=>"100111111",
  14504=>"010101000",
  14505=>"000001001",
  14506=>"111111000",
  14507=>"001000001",
  14508=>"111101111",
  14509=>"000000000",
  14510=>"001011011",
  14511=>"100101000",
  14512=>"111111000",
  14513=>"110110010",
  14514=>"111111111",
  14515=>"111000000",
  14516=>"000001111",
  14517=>"000010011",
  14518=>"000001110",
  14519=>"010111000",
  14520=>"110100010",
  14521=>"000001001",
  14522=>"111111111",
  14523=>"111110000",
  14524=>"000000010",
  14525=>"111111111",
  14526=>"100100101",
  14527=>"010011000",
  14528=>"000111010",
  14529=>"001001111",
  14530=>"000000001",
  14531=>"001001001",
  14532=>"000000001",
  14533=>"111000110",
  14534=>"000001110",
  14535=>"111110000",
  14536=>"000000111",
  14537=>"000001011",
  14538=>"000111011",
  14539=>"000101111",
  14540=>"101000100",
  14541=>"111000000",
  14542=>"011101101",
  14543=>"111010101",
  14544=>"111011011",
  14545=>"111110010",
  14546=>"000000000",
  14547=>"000101111",
  14548=>"010000000",
  14549=>"011111011",
  14550=>"110110000",
  14551=>"000001110",
  14552=>"000000111",
  14553=>"000000000",
  14554=>"010111111",
  14555=>"111111101",
  14556=>"000111100",
  14557=>"111101111",
  14558=>"011010000",
  14559=>"000000010",
  14560=>"000000000",
  14561=>"111000000",
  14562=>"111000001",
  14563=>"001011011",
  14564=>"001101111",
  14565=>"111000000",
  14566=>"111111110",
  14567=>"100101010",
  14568=>"111100110",
  14569=>"011000000",
  14570=>"000000100",
  14571=>"110011011",
  14572=>"000000000",
  14573=>"001111111",
  14574=>"111111000",
  14575=>"111111010",
  14576=>"000000011",
  14577=>"010110110",
  14578=>"111111111",
  14579=>"000001111",
  14580=>"001111011",
  14581=>"111111000",
  14582=>"010010010",
  14583=>"111000100",
  14584=>"000110110",
  14585=>"100001101",
  14586=>"011110000",
  14587=>"000100000",
  14588=>"000000010",
  14589=>"101000000",
  14590=>"101011010",
  14591=>"000000000",
  14592=>"000000011",
  14593=>"111111001",
  14594=>"000111010",
  14595=>"000000000",
  14596=>"000000000",
  14597=>"000010010",
  14598=>"101111000",
  14599=>"000000000",
  14600=>"000001001",
  14601=>"000011001",
  14602=>"000000001",
  14603=>"000000110",
  14604=>"110000000",
  14605=>"100111111",
  14606=>"100100000",
  14607=>"000011111",
  14608=>"000000111",
  14609=>"111100000",
  14610=>"001000010",
  14611=>"101111101",
  14612=>"000000000",
  14613=>"110111100",
  14614=>"000111111",
  14615=>"111000111",
  14616=>"010000000",
  14617=>"000000000",
  14618=>"111100000",
  14619=>"111111111",
  14620=>"101000100",
  14621=>"001000000",
  14622=>"000000110",
  14623=>"101101001",
  14624=>"000010110",
  14625=>"111110011",
  14626=>"010101100",
  14627=>"010111011",
  14628=>"111011011",
  14629=>"100001000",
  14630=>"110100000",
  14631=>"000000000",
  14632=>"111111101",
  14633=>"000101111",
  14634=>"000000001",
  14635=>"000000110",
  14636=>"000010111",
  14637=>"000000000",
  14638=>"000000000",
  14639=>"000000000",
  14640=>"101111010",
  14641=>"111011110",
  14642=>"010001101",
  14643=>"111001100",
  14644=>"000000000",
  14645=>"000000010",
  14646=>"000000000",
  14647=>"001000001",
  14648=>"111000000",
  14649=>"111101000",
  14650=>"000000011",
  14651=>"110110000",
  14652=>"111111110",
  14653=>"111111111",
  14654=>"111100010",
  14655=>"101111111",
  14656=>"100010010",
  14657=>"000001010",
  14658=>"110111000",
  14659=>"111011111",
  14660=>"000000010",
  14661=>"101001111",
  14662=>"100110011",
  14663=>"001001110",
  14664=>"110111000",
  14665=>"110000000",
  14666=>"111101111",
  14667=>"010001000",
  14668=>"111100000",
  14669=>"101110100",
  14670=>"011110011",
  14671=>"000000000",
  14672=>"101101101",
  14673=>"111101111",
  14674=>"111111100",
  14675=>"100000000",
  14676=>"111111110",
  14677=>"100011001",
  14678=>"001000001",
  14679=>"000000000",
  14680=>"001111111",
  14681=>"011001000",
  14682=>"010111110",
  14683=>"100111111",
  14684=>"000001011",
  14685=>"000110100",
  14686=>"011110000",
  14687=>"110100000",
  14688=>"000000000",
  14689=>"000101101",
  14690=>"111010010",
  14691=>"001001001",
  14692=>"100000010",
  14693=>"101111111",
  14694=>"000000000",
  14695=>"000000001",
  14696=>"111010010",
  14697=>"000000110",
  14698=>"010110110",
  14699=>"001111111",
  14700=>"000000111",
  14701=>"000001101",
  14702=>"001000000",
  14703=>"000000000",
  14704=>"110111101",
  14705=>"010111111",
  14706=>"000000000",
  14707=>"000000101",
  14708=>"000111101",
  14709=>"000010000",
  14710=>"100000111",
  14711=>"011101101",
  14712=>"111111111",
  14713=>"111110101",
  14714=>"010000111",
  14715=>"111111000",
  14716=>"000001100",
  14717=>"000011010",
  14718=>"010111100",
  14719=>"011111010",
  14720=>"000101101",
  14721=>"101000000",
  14722=>"000001011",
  14723=>"001001001",
  14724=>"111000000",
  14725=>"000111000",
  14726=>"111110100",
  14727=>"011100000",
  14728=>"001011000",
  14729=>"111111000",
  14730=>"001000111",
  14731=>"000000110",
  14732=>"001000000",
  14733=>"111010000",
  14734=>"100000010",
  14735=>"000000000",
  14736=>"010100000",
  14737=>"111111111",
  14738=>"000000101",
  14739=>"000000000",
  14740=>"111111100",
  14741=>"001000010",
  14742=>"011011000",
  14743=>"110100110",
  14744=>"000010111",
  14745=>"000000101",
  14746=>"100111111",
  14747=>"000011000",
  14748=>"010010000",
  14749=>"110111011",
  14750=>"010111111",
  14751=>"000000000",
  14752=>"000111000",
  14753=>"111000011",
  14754=>"000000000",
  14755=>"001000000",
  14756=>"100000000",
  14757=>"000101111",
  14758=>"011001011",
  14759=>"000000111",
  14760=>"111111001",
  14761=>"000000101",
  14762=>"111110110",
  14763=>"010010000",
  14764=>"001101111",
  14765=>"100100111",
  14766=>"010110000",
  14767=>"000011011",
  14768=>"100111110",
  14769=>"111101000",
  14770=>"111101000",
  14771=>"000000001",
  14772=>"000001100",
  14773=>"000000011",
  14774=>"000000000",
  14775=>"000111111",
  14776=>"111111001",
  14777=>"100101100",
  14778=>"111111111",
  14779=>"100111111",
  14780=>"000000001",
  14781=>"111111000",
  14782=>"100100000",
  14783=>"000011111",
  14784=>"101101010",
  14785=>"001000000",
  14786=>"111101001",
  14787=>"000001001",
  14788=>"000000000",
  14789=>"001010000",
  14790=>"000000001",
  14791=>"111101001",
  14792=>"001000001",
  14793=>"111001000",
  14794=>"000000101",
  14795=>"010111110",
  14796=>"010011111",
  14797=>"010000001",
  14798=>"000000101",
  14799=>"111111110",
  14800=>"000111000",
  14801=>"000100110",
  14802=>"011101000",
  14803=>"000000101",
  14804=>"111110000",
  14805=>"100100000",
  14806=>"001000000",
  14807=>"000111111",
  14808=>"000000000",
  14809=>"000000000",
  14810=>"011010001",
  14811=>"000110111",
  14812=>"000110111",
  14813=>"000111111",
  14814=>"000000000",
  14815=>"111111101",
  14816=>"110111110",
  14817=>"111011010",
  14818=>"111111101",
  14819=>"000001101",
  14820=>"000000100",
  14821=>"100110111",
  14822=>"111111010",
  14823=>"000100111",
  14824=>"111111111",
  14825=>"000001101",
  14826=>"000000110",
  14827=>"000000000",
  14828=>"001000000",
  14829=>"001000101",
  14830=>"000111000",
  14831=>"010111101",
  14832=>"000000101",
  14833=>"000000000",
  14834=>"000101111",
  14835=>"010110101",
  14836=>"000001000",
  14837=>"000110101",
  14838=>"111111000",
  14839=>"000010000",
  14840=>"000000101",
  14841=>"000000000",
  14842=>"000000100",
  14843=>"000000011",
  14844=>"111011000",
  14845=>"111111111",
  14846=>"000110011",
  14847=>"100100010",
  14848=>"001000001",
  14849=>"000000000",
  14850=>"010111010",
  14851=>"101000000",
  14852=>"000000100",
  14853=>"000000001",
  14854=>"101111101",
  14855=>"110000000",
  14856=>"000000000",
  14857=>"110001000",
  14858=>"000100100",
  14859=>"110111111",
  14860=>"001011011",
  14861=>"111001001",
  14862=>"000111011",
  14863=>"000000000",
  14864=>"111000100",
  14865=>"001110000",
  14866=>"000000000",
  14867=>"110000111",
  14868=>"000000000",
  14869=>"010111111",
  14870=>"001111100",
  14871=>"010010110",
  14872=>"000000000",
  14873=>"011000100",
  14874=>"000000101",
  14875=>"111111001",
  14876=>"101010110",
  14877=>"001111000",
  14878=>"101000000",
  14879=>"111111001",
  14880=>"111111111",
  14881=>"111000111",
  14882=>"110111000",
  14883=>"111111111",
  14884=>"111001001",
  14885=>"001011101",
  14886=>"000111000",
  14887=>"110001101",
  14888=>"111001111",
  14889=>"010000000",
  14890=>"111111111",
  14891=>"000111000",
  14892=>"111110110",
  14893=>"101000001",
  14894=>"101111111",
  14895=>"111000100",
  14896=>"000000010",
  14897=>"000000000",
  14898=>"000000000",
  14899=>"110110000",
  14900=>"000001001",
  14901=>"000000000",
  14902=>"110111111",
  14903=>"111001000",
  14904=>"001000000",
  14905=>"100000101",
  14906=>"000000000",
  14907=>"000000010",
  14908=>"110011100",
  14909=>"111111111",
  14910=>"000000101",
  14911=>"000000000",
  14912=>"111000110",
  14913=>"111111111",
  14914=>"110100000",
  14915=>"001101001",
  14916=>"000000100",
  14917=>"000000000",
  14918=>"111101110",
  14919=>"000111111",
  14920=>"111111111",
  14921=>"000000101",
  14922=>"101000101",
  14923=>"111111110",
  14924=>"000100110",
  14925=>"011000000",
  14926=>"011001000",
  14927=>"100011111",
  14928=>"100101111",
  14929=>"111111010",
  14930=>"001000000",
  14931=>"001010100",
  14932=>"000000000",
  14933=>"000111100",
  14934=>"111001001",
  14935=>"010000010",
  14936=>"010010010",
  14937=>"110110111",
  14938=>"010111101",
  14939=>"001000100",
  14940=>"101101101",
  14941=>"000000001",
  14942=>"010111111",
  14943=>"100100111",
  14944=>"111101111",
  14945=>"101111111",
  14946=>"000000010",
  14947=>"000111110",
  14948=>"000001100",
  14949=>"101000011",
  14950=>"100110111",
  14951=>"111000000",
  14952=>"000000000",
  14953=>"000000000",
  14954=>"101000001",
  14955=>"100110111",
  14956=>"111101000",
  14957=>"101000000",
  14958=>"111000000",
  14959=>"111000000",
  14960=>"101001000",
  14961=>"000000000",
  14962=>"111111111",
  14963=>"111100101",
  14964=>"010100000",
  14965=>"101000000",
  14966=>"010000000",
  14967=>"110101000",
  14968=>"010111011",
  14969=>"111111111",
  14970=>"000011111",
  14971=>"011001000",
  14972=>"000100100",
  14973=>"100000000",
  14974=>"111111111",
  14975=>"000111111",
  14976=>"101101000",
  14977=>"000111011",
  14978=>"000000000",
  14979=>"111000111",
  14980=>"101000000",
  14981=>"100000000",
  14982=>"011111011",
  14983=>"100110111",
  14984=>"000000001",
  14985=>"111111111",
  14986=>"111101100",
  14987=>"111101010",
  14988=>"010010000",
  14989=>"101111100",
  14990=>"110111111",
  14991=>"001001000",
  14992=>"000000000",
  14993=>"111111101",
  14994=>"111101101",
  14995=>"111010000",
  14996=>"001011111",
  14997=>"111000000",
  14998=>"011111111",
  14999=>"000000011",
  15000=>"001000000",
  15001=>"000000000",
  15002=>"111111111",
  15003=>"110010001",
  15004=>"000000000",
  15005=>"000000000",
  15006=>"000000101",
  15007=>"000000111",
  15008=>"110111110",
  15009=>"111011111",
  15010=>"111111111",
  15011=>"110000000",
  15012=>"110101000",
  15013=>"010001001",
  15014=>"100100100",
  15015=>"000000010",
  15016=>"111111000",
  15017=>"110101100",
  15018=>"111010000",
  15019=>"000000111",
  15020=>"101100111",
  15021=>"111000000",
  15022=>"000000100",
  15023=>"100111111",
  15024=>"000100000",
  15025=>"111111111",
  15026=>"000001011",
  15027=>"000010100",
  15028=>"100100000",
  15029=>"110111010",
  15030=>"000000000",
  15031=>"000000010",
  15032=>"011010001",
  15033=>"001000101",
  15034=>"111111001",
  15035=>"111001000",
  15036=>"000100000",
  15037=>"000011010",
  15038=>"000000000",
  15039=>"011000000",
  15040=>"111101000",
  15041=>"000110000",
  15042=>"111101000",
  15043=>"001001001",
  15044=>"100000000",
  15045=>"100110001",
  15046=>"111100000",
  15047=>"000000110",
  15048=>"001000010",
  15049=>"111111111",
  15050=>"000000000",
  15051=>"111101111",
  15052=>"011000100",
  15053=>"000001010",
  15054=>"101000011",
  15055=>"000000000",
  15056=>"111111111",
  15057=>"111011011",
  15058=>"100011000",
  15059=>"001000000",
  15060=>"001001111",
  15061=>"100101100",
  15062=>"000000000",
  15063=>"000000000",
  15064=>"111000011",
  15065=>"010010111",
  15066=>"011001001",
  15067=>"000010000",
  15068=>"001111011",
  15069=>"000000000",
  15070=>"010110110",
  15071=>"111001100",
  15072=>"011100001",
  15073=>"000011101",
  15074=>"001000101",
  15075=>"000011000",
  15076=>"101001101",
  15077=>"011111100",
  15078=>"000001111",
  15079=>"001101001",
  15080=>"000000000",
  15081=>"100000100",
  15082=>"000000001",
  15083=>"010011000",
  15084=>"000001000",
  15085=>"100000100",
  15086=>"000010000",
  15087=>"111100000",
  15088=>"111000000",
  15089=>"011111110",
  15090=>"111111000",
  15091=>"011001011",
  15092=>"110110100",
  15093=>"000111111",
  15094=>"000000000",
  15095=>"000010000",
  15096=>"011010011",
  15097=>"001000001",
  15098=>"101100100",
  15099=>"101010010",
  15100=>"011111011",
  15101=>"110111111",
  15102=>"100000000",
  15103=>"001000000",
  15104=>"011101100",
  15105=>"111000000",
  15106=>"000000000",
  15107=>"111010110",
  15108=>"110110000",
  15109=>"101110110",
  15110=>"010111000",
  15111=>"000000001",
  15112=>"111011110",
  15113=>"000001110",
  15114=>"000011011",
  15115=>"000010000",
  15116=>"000000111",
  15117=>"110000000",
  15118=>"110100010",
  15119=>"111101100",
  15120=>"110010011",
  15121=>"111011000",
  15122=>"010000000",
  15123=>"000000000",
  15124=>"111000000",
  15125=>"111111111",
  15126=>"001111111",
  15127=>"111111000",
  15128=>"000000011",
  15129=>"111111111",
  15130=>"000000000",
  15131=>"000111000",
  15132=>"110100000",
  15133=>"000100001",
  15134=>"000110100",
  15135=>"000000111",
  15136=>"101001000",
  15137=>"111001001",
  15138=>"111101101",
  15139=>"100111110",
  15140=>"110111100",
  15141=>"100001011",
  15142=>"000000010",
  15143=>"010100010",
  15144=>"000000001",
  15145=>"011001111",
  15146=>"100110110",
  15147=>"110100110",
  15148=>"000000011",
  15149=>"000000111",
  15150=>"111101110",
  15151=>"111011111",
  15152=>"010010000",
  15153=>"000110100",
  15154=>"110001000",
  15155=>"111000000",
  15156=>"111111101",
  15157=>"000000000",
  15158=>"000000101",
  15159=>"011111011",
  15160=>"001000000",
  15161=>"111000000",
  15162=>"111000000",
  15163=>"011111100",
  15164=>"111101000",
  15165=>"000111111",
  15166=>"000000000",
  15167=>"010001111",
  15168=>"111110111",
  15169=>"000101111",
  15170=>"101111111",
  15171=>"000111111",
  15172=>"000110110",
  15173=>"001010000",
  15174=>"000111011",
  15175=>"111111111",
  15176=>"110001111",
  15177=>"000101111",
  15178=>"101000000",
  15179=>"111111011",
  15180=>"000011110",
  15181=>"011111111",
  15182=>"000111011",
  15183=>"010000001",
  15184=>"000001000",
  15185=>"101010111",
  15186=>"110101100",
  15187=>"101000000",
  15188=>"000100111",
  15189=>"011001001",
  15190=>"010011101",
  15191=>"100111000",
  15192=>"000000111",
  15193=>"000110100",
  15194=>"111000100",
  15195=>"011100010",
  15196=>"000111111",
  15197=>"111101100",
  15198=>"111001000",
  15199=>"000011111",
  15200=>"000110111",
  15201=>"000111111",
  15202=>"000000111",
  15203=>"111000010",
  15204=>"111001100",
  15205=>"010011001",
  15206=>"000110110",
  15207=>"101011111",
  15208=>"110111111",
  15209=>"000010111",
  15210=>"000010111",
  15211=>"111001111",
  15212=>"111111011",
  15213=>"111111000",
  15214=>"011000001",
  15215=>"111111011",
  15216=>"001011011",
  15217=>"000010000",
  15218=>"000000110",
  15219=>"001001000",
  15220=>"000000110",
  15221=>"100111111",
  15222=>"111111011",
  15223=>"000001100",
  15224=>"000001010",
  15225=>"110111101",
  15226=>"010111101",
  15227=>"110111101",
  15228=>"001001000",
  15229=>"111000011",
  15230=>"001101110",
  15231=>"000000111",
  15232=>"110111110",
  15233=>"111011000",
  15234=>"000111111",
  15235=>"111111111",
  15236=>"010000111",
  15237=>"000000100",
  15238=>"001000110",
  15239=>"000110100",
  15240=>"010110110",
  15241=>"100111111",
  15242=>"010110100",
  15243=>"101111000",
  15244=>"111000001",
  15245=>"101111111",
  15246=>"111000000",
  15247=>"000101000",
  15248=>"110100100",
  15249=>"001101111",
  15250=>"111001101",
  15251=>"000000100",
  15252=>"111110000",
  15253=>"111000000",
  15254=>"111111111",
  15255=>"010010011",
  15256=>"000111010",
  15257=>"100101011",
  15258=>"000001111",
  15259=>"010011101",
  15260=>"100001111",
  15261=>"000110111",
  15262=>"001010100",
  15263=>"000111111",
  15264=>"011110000",
  15265=>"111111000",
  15266=>"000000101",
  15267=>"100001100",
  15268=>"111101010",
  15269=>"000010010",
  15270=>"111101100",
  15271=>"000001000",
  15272=>"111110000",
  15273=>"100101111",
  15274=>"111000000",
  15275=>"011010000",
  15276=>"111101111",
  15277=>"000000111",
  15278=>"100000001",
  15279=>"110011011",
  15280=>"000110010",
  15281=>"001000100",
  15282=>"101111011",
  15283=>"000011011",
  15284=>"010100110",
  15285=>"111101000",
  15286=>"010000011",
  15287=>"111000000",
  15288=>"111001100",
  15289=>"000000001",
  15290=>"111000000",
  15291=>"111001110",
  15292=>"101100111",
  15293=>"000000111",
  15294=>"100110111",
  15295=>"000000100",
  15296=>"101000111",
  15297=>"111100000",
  15298=>"111011000",
  15299=>"110100110",
  15300=>"000101010",
  15301=>"111111001",
  15302=>"110111111",
  15303=>"111101111",
  15304=>"101110101",
  15305=>"000001111",
  15306=>"000100110",
  15307=>"000101111",
  15308=>"000000111",
  15309=>"101100100",
  15310=>"000000000",
  15311=>"110110111",
  15312=>"000000100",
  15313=>"001111100",
  15314=>"111111001",
  15315=>"011001000",
  15316=>"000101111",
  15317=>"001011000",
  15318=>"111000111",
  15319=>"111000000",
  15320=>"000000100",
  15321=>"000111000",
  15322=>"111111011",
  15323=>"000111010",
  15324=>"011111111",
  15325=>"111111111",
  15326=>"010001100",
  15327=>"000111010",
  15328=>"000110111",
  15329=>"111001101",
  15330=>"111000000",
  15331=>"011011011",
  15332=>"000000000",
  15333=>"011011111",
  15334=>"111000001",
  15335=>"000011000",
  15336=>"010111110",
  15337=>"000100101",
  15338=>"000000110",
  15339=>"000101010",
  15340=>"000000000",
  15341=>"000000111",
  15342=>"000000010",
  15343=>"101000000",
  15344=>"111111111",
  15345=>"111110100",
  15346=>"101000110",
  15347=>"000011000",
  15348=>"001101011",
  15349=>"000000000",
  15350=>"100100110",
  15351=>"111111000",
  15352=>"111000000",
  15353=>"001001000",
  15354=>"111100100",
  15355=>"111011100",
  15356=>"101111010",
  15357=>"000000000",
  15358=>"000011000",
  15359=>"111000111",
  15360=>"111011001",
  15361=>"011011000",
  15362=>"000000000",
  15363=>"011011011",
  15364=>"100100000",
  15365=>"100111111",
  15366=>"001111000",
  15367=>"000011111",
  15368=>"100110110",
  15369=>"000001011",
  15370=>"001001000",
  15371=>"101110110",
  15372=>"111101111",
  15373=>"000000000",
  15374=>"111111110",
  15375=>"110110101",
  15376=>"100000001",
  15377=>"110111011",
  15378=>"000000000",
  15379=>"011001001",
  15380=>"111111001",
  15381=>"000000000",
  15382=>"111101001",
  15383=>"111111111",
  15384=>"000001101",
  15385=>"100000001",
  15386=>"110111001",
  15387=>"000010001",
  15388=>"000100000",
  15389=>"111010011",
  15390=>"111100000",
  15391=>"000100100",
  15392=>"101111001",
  15393=>"111010011",
  15394=>"110101010",
  15395=>"101101001",
  15396=>"101101001",
  15397=>"000000000",
  15398=>"000011011",
  15399=>"101111111",
  15400=>"101110100",
  15401=>"010001001",
  15402=>"000000000",
  15403=>"110111101",
  15404=>"100011000",
  15405=>"110001011",
  15406=>"111010011",
  15407=>"101110000",
  15408=>"011001111",
  15409=>"111111100",
  15410=>"110000101",
  15411=>"110010000",
  15412=>"111110011",
  15413=>"111001010",
  15414=>"111011111",
  15415=>"101011111",
  15416=>"100001111",
  15417=>"000001111",
  15418=>"001101111",
  15419=>"111000010",
  15420=>"000101100",
  15421=>"110110110",
  15422=>"000000000",
  15423=>"101111000",
  15424=>"000010111",
  15425=>"000000010",
  15426=>"111101000",
  15427=>"001001001",
  15428=>"001110110",
  15429=>"111000101",
  15430=>"001010000",
  15431=>"110100110",
  15432=>"011001101",
  15433=>"100000011",
  15434=>"001001111",
  15435=>"110110010",
  15436=>"100010000",
  15437=>"111001001",
  15438=>"111111100",
  15439=>"011110111",
  15440=>"010110110",
  15441=>"100110111",
  15442=>"111010001",
  15443=>"011001100",
  15444=>"000010010",
  15445=>"101100000",
  15446=>"011101101",
  15447=>"000000001",
  15448=>"000100010",
  15449=>"001001000",
  15450=>"001111111",
  15451=>"011011010",
  15452=>"000011111",
  15453=>"000000101",
  15454=>"111011111",
  15455=>"111110011",
  15456=>"000111110",
  15457=>"000011000",
  15458=>"001111011",
  15459=>"001000000",
  15460=>"000101101",
  15461=>"011001000",
  15462=>"111111111",
  15463=>"000101110",
  15464=>"111000011",
  15465=>"111001011",
  15466=>"110111111",
  15467=>"111110111",
  15468=>"000100101",
  15469=>"100000100",
  15470=>"001011011",
  15471=>"111111110",
  15472=>"001101101",
  15473=>"111111111",
  15474=>"011001000",
  15475=>"111100000",
  15476=>"100000000",
  15477=>"111000001",
  15478=>"110000010",
  15479=>"111000000",
  15480=>"000000000",
  15481=>"000001010",
  15482=>"110010000",
  15483=>"000000000",
  15484=>"110101101",
  15485=>"100000001",
  15486=>"101111111",
  15487=>"000000000",
  15488=>"110000000",
  15489=>"010011000",
  15490=>"110000001",
  15491=>"111110110",
  15492=>"101111111",
  15493=>"101010110",
  15494=>"011100101",
  15495=>"000110000",
  15496=>"001001001",
  15497=>"000000000",
  15498=>"000000001",
  15499=>"111000111",
  15500=>"000110100",
  15501=>"101110010",
  15502=>"101111111",
  15503=>"100100110",
  15504=>"000100100",
  15505=>"101000110",
  15506=>"000010001",
  15507=>"001100111",
  15508=>"011011010",
  15509=>"100001011",
  15510=>"010010010",
  15511=>"011101110",
  15512=>"110100010",
  15513=>"000010100",
  15514=>"000110000",
  15515=>"000001111",
  15516=>"111011000",
  15517=>"000100010",
  15518=>"110110011",
  15519=>"000000000",
  15520=>"000011111",
  15521=>"010001000",
  15522=>"110000001",
  15523=>"110000110",
  15524=>"111001110",
  15525=>"000110111",
  15526=>"110000001",
  15527=>"000100000",
  15528=>"100000000",
  15529=>"010011111",
  15530=>"001100100",
  15531=>"010001111",
  15532=>"111100000",
  15533=>"111110111",
  15534=>"000000000",
  15535=>"001001111",
  15536=>"100000001",
  15537=>"011011110",
  15538=>"010010100",
  15539=>"101100110",
  15540=>"101111111",
  15541=>"011001110",
  15542=>"111000001",
  15543=>"100100100",
  15544=>"110000000",
  15545=>"000000000",
  15546=>"000100000",
  15547=>"111111100",
  15548=>"101000001",
  15549=>"111110100",
  15550=>"110000011",
  15551=>"000001000",
  15552=>"111110000",
  15553=>"000000100",
  15554=>"111101101",
  15555=>"011001100",
  15556=>"001001001",
  15557=>"100110000",
  15558=>"000000111",
  15559=>"011101101",
  15560=>"100100000",
  15561=>"000010010",
  15562=>"111001111",
  15563=>"000000010",
  15564=>"010011000",
  15565=>"000100111",
  15566=>"011111111",
  15567=>"001001111",
  15568=>"010010110",
  15569=>"101111111",
  15570=>"000100110",
  15571=>"010111101",
  15572=>"100110100",
  15573=>"000100101",
  15574=>"100000001",
  15575=>"110100011",
  15576=>"011011000",
  15577=>"000000111",
  15578=>"011101001",
  15579=>"000000000",
  15580=>"111111111",
  15581=>"000000000",
  15582=>"110010111",
  15583=>"000000110",
  15584=>"000000111",
  15585=>"111111101",
  15586=>"111111000",
  15587=>"001011110",
  15588=>"000010000",
  15589=>"100101011",
  15590=>"110111111",
  15591=>"111111111",
  15592=>"011011011",
  15593=>"010001101",
  15594=>"111111111",
  15595=>"110100001",
  15596=>"011001111",
  15597=>"111111001",
  15598=>"100001000",
  15599=>"100001001",
  15600=>"000001000",
  15601=>"110011100",
  15602=>"001001000",
  15603=>"001101001",
  15604=>"000000000",
  15605=>"001111101",
  15606=>"000000001",
  15607=>"001110110",
  15608=>"001011001",
  15609=>"111111111",
  15610=>"111111111",
  15611=>"111110111",
  15612=>"010010000",
  15613=>"010010000",
  15614=>"010110100",
  15615=>"010111000",
  15616=>"000110011",
  15617=>"000000010",
  15618=>"111000000",
  15619=>"011000101",
  15620=>"100110110",
  15621=>"111000000",
  15622=>"000010010",
  15623=>"101110111",
  15624=>"000011111",
  15625=>"000110011",
  15626=>"110001001",
  15627=>"111001111",
  15628=>"101101101",
  15629=>"000110111",
  15630=>"101000000",
  15631=>"100000101",
  15632=>"111000010",
  15633=>"101000010",
  15634=>"000111101",
  15635=>"100111011",
  15636=>"101000000",
  15637=>"111100100",
  15638=>"011011011",
  15639=>"000111011",
  15640=>"111000001",
  15641=>"111101101",
  15642=>"010100100",
  15643=>"010100111",
  15644=>"000000100",
  15645=>"111100111",
  15646=>"111011111",
  15647=>"101110100",
  15648=>"100000000",
  15649=>"000010111",
  15650=>"010111000",
  15651=>"100110010",
  15652=>"000110100",
  15653=>"011011001",
  15654=>"000000110",
  15655=>"000000100",
  15656=>"111001111",
  15657=>"110011010",
  15658=>"110100111",
  15659=>"011111001",
  15660=>"000110010",
  15661=>"101000100",
  15662=>"010001100",
  15663=>"111010101",
  15664=>"101011000",
  15665=>"110010011",
  15666=>"110011111",
  15667=>"100001100",
  15668=>"011000100",
  15669=>"101010111",
  15670=>"000011011",
  15671=>"000011111",
  15672=>"111011100",
  15673=>"000101111",
  15674=>"100000100",
  15675=>"100011101",
  15676=>"001111001",
  15677=>"111111011",
  15678=>"010000100",
  15679=>"000001111",
  15680=>"111111100",
  15681=>"010111010",
  15682=>"000000000",
  15683=>"111101100",
  15684=>"100010011",
  15685=>"000000100",
  15686=>"000001111",
  15687=>"111101000",
  15688=>"000100001",
  15689=>"101101101",
  15690=>"010000000",
  15691=>"111101101",
  15692=>"110100110",
  15693=>"011111100",
  15694=>"010000100",
  15695=>"100101011",
  15696=>"100101100",
  15697=>"111111111",
  15698=>"111011010",
  15699=>"110011001",
  15700=>"111100000",
  15701=>"000000101",
  15702=>"000111110",
  15703=>"000000000",
  15704=>"111101111",
  15705=>"000011011",
  15706=>"110110010",
  15707=>"000001000",
  15708=>"100111111",
  15709=>"010000000",
  15710=>"010111010",
  15711=>"111100000",
  15712=>"000001111",
  15713=>"001101101",
  15714=>"011000100",
  15715=>"100001001",
  15716=>"000000000",
  15717=>"000111011",
  15718=>"101000101",
  15719=>"110100000",
  15720=>"000011011",
  15721=>"011111100",
  15722=>"000001010",
  15723=>"111101010",
  15724=>"100111011",
  15725=>"111100000",
  15726=>"000000100",
  15727=>"000000000",
  15728=>"001010100",
  15729=>"100000010",
  15730=>"000011010",
  15731=>"111101101",
  15732=>"011111100",
  15733=>"110000100",
  15734=>"000001110",
  15735=>"111111111",
  15736=>"000100000",
  15737=>"000110111",
  15738=>"111101000",
  15739=>"101101111",
  15740=>"001110100",
  15741=>"000110100",
  15742=>"110011000",
  15743=>"111000000",
  15744=>"000011011",
  15745=>"111111000",
  15746=>"100100011",
  15747=>"111000111",
  15748=>"101111000",
  15749=>"001010000",
  15750=>"100110010",
  15751=>"000000000",
  15752=>"101011000",
  15753=>"111000000",
  15754=>"011000001",
  15755=>"100100100",
  15756=>"000000101",
  15757=>"111000111",
  15758=>"000000111",
  15759=>"011000001",
  15760=>"111011101",
  15761=>"000011111",
  15762=>"100000011",
  15763=>"000000000",
  15764=>"000000000",
  15765=>"001101111",
  15766=>"101110000",
  15767=>"000110011",
  15768=>"100110111",
  15769=>"011000010",
  15770=>"111000100",
  15771=>"111101100",
  15772=>"000000011",
  15773=>"011000101",
  15774=>"111011100",
  15775=>"111101101",
  15776=>"000011111",
  15777=>"111010010",
  15778=>"101111010",
  15779=>"011000111",
  15780=>"011111010",
  15781=>"000100111",
  15782=>"011001101",
  15783=>"000001010",
  15784=>"000101111",
  15785=>"010101101",
  15786=>"101110100",
  15787=>"010100100",
  15788=>"001100001",
  15789=>"000000000",
  15790=>"000011111",
  15791=>"111001100",
  15792=>"101101001",
  15793=>"111110100",
  15794=>"111000011",
  15795=>"000101000",
  15796=>"110101111",
  15797=>"100011001",
  15798=>"000101100",
  15799=>"111111000",
  15800=>"000101100",
  15801=>"011101000",
  15802=>"000010000",
  15803=>"000111000",
  15804=>"110000000",
  15805=>"111000000",
  15806=>"000110111",
  15807=>"111000010",
  15808=>"111100000",
  15809=>"000100100",
  15810=>"111111100",
  15811=>"110011001",
  15812=>"000000101",
  15813=>"111100000",
  15814=>"001010010",
  15815=>"000000000",
  15816=>"000010111",
  15817=>"011000000",
  15818=>"101011111",
  15819=>"000110011",
  15820=>"000011011",
  15821=>"110011001",
  15822=>"010000010",
  15823=>"000000100",
  15824=>"111011110",
  15825=>"000111111",
  15826=>"111000100",
  15827=>"000111111",
  15828=>"110000111",
  15829=>"011101000",
  15830=>"110100000",
  15831=>"111110110",
  15832=>"000011000",
  15833=>"110000111",
  15834=>"000010111",
  15835=>"111000100",
  15836=>"110000101",
  15837=>"111101101",
  15838=>"111110101",
  15839=>"101011000",
  15840=>"111000000",
  15841=>"111100000",
  15842=>"111110100",
  15843=>"111010000",
  15844=>"111101000",
  15845=>"011011011",
  15846=>"000001101",
  15847=>"000110110",
  15848=>"011001111",
  15849=>"101101000",
  15850=>"001100100",
  15851=>"111101100",
  15852=>"111100110",
  15853=>"110111000",
  15854=>"000000001",
  15855=>"100000001",
  15856=>"000010111",
  15857=>"011001000",
  15858=>"000100000",
  15859=>"000010111",
  15860=>"000011010",
  15861=>"111001000",
  15862=>"110100010",
  15863=>"111000000",
  15864=>"000010011",
  15865=>"000000000",
  15866=>"111100111",
  15867=>"000000000",
  15868=>"100111010",
  15869=>"111000111",
  15870=>"000011001",
  15871=>"110000001",
  15872=>"010111001",
  15873=>"100000010",
  15874=>"000110010",
  15875=>"100000010",
  15876=>"011111110",
  15877=>"100000110",
  15878=>"001101111",
  15879=>"100101011",
  15880=>"000111111",
  15881=>"000000000",
  15882=>"011001110",
  15883=>"111111111",
  15884=>"111010000",
  15885=>"100010111",
  15886=>"111100001",
  15887=>"100000000",
  15888=>"000111111",
  15889=>"000000011",
  15890=>"000000000",
  15891=>"000000111",
  15892=>"101011111",
  15893=>"110111101",
  15894=>"000100011",
  15895=>"000010111",
  15896=>"000000000",
  15897=>"111110000",
  15898=>"111111111",
  15899=>"000111111",
  15900=>"111000111",
  15901=>"101010010",
  15902=>"111111110",
  15903=>"011101000",
  15904=>"000000000",
  15905=>"111111011",
  15906=>"111010111",
  15907=>"010000010",
  15908=>"011101111",
  15909=>"000001101",
  15910=>"000000000",
  15911=>"100111110",
  15912=>"111101111",
  15913=>"000111000",
  15914=>"000111111",
  15915=>"001101000",
  15916=>"111110001",
  15917=>"111010000",
  15918=>"101000001",
  15919=>"001000001",
  15920=>"000000000",
  15921=>"001000000",
  15922=>"010111101",
  15923=>"111010010",
  15924=>"000000100",
  15925=>"011000000",
  15926=>"110000011",
  15927=>"000000010",
  15928=>"001001001",
  15929=>"001111101",
  15930=>"100000000",
  15931=>"010000000",
  15932=>"011011001",
  15933=>"111101101",
  15934=>"000000110",
  15935=>"000101101",
  15936=>"111000110",
  15937=>"111111101",
  15938=>"000101101",
  15939=>"001001110",
  15940=>"000111010",
  15941=>"000000100",
  15942=>"000001101",
  15943=>"111000111",
  15944=>"111100110",
  15945=>"111011100",
  15946=>"101101111",
  15947=>"101010111",
  15948=>"000000111",
  15949=>"001011111",
  15950=>"110111000",
  15951=>"101010111",
  15952=>"101000000",
  15953=>"000111111",
  15954=>"010000110",
  15955=>"001000011",
  15956=>"110111111",
  15957=>"000100111",
  15958=>"111001001",
  15959=>"011010000",
  15960=>"010001010",
  15961=>"011110001",
  15962=>"110100100",
  15963=>"001001010",
  15964=>"110011000",
  15965=>"000000001",
  15966=>"010011111",
  15967=>"100010111",
  15968=>"000011010",
  15969=>"101111110",
  15970=>"000000000",
  15971=>"111101011",
  15972=>"110101100",
  15973=>"111011000",
  15974=>"110000000",
  15975=>"000000000",
  15976=>"111111000",
  15977=>"000111111",
  15978=>"000000111",
  15979=>"111001111",
  15980=>"111001111",
  15981=>"010010001",
  15982=>"111000010",
  15983=>"000000010",
  15984=>"110110100",
  15985=>"001101101",
  15986=>"001000100",
  15987=>"111100000",
  15988=>"000000111",
  15989=>"001000001",
  15990=>"111111000",
  15991=>"010000101",
  15992=>"001111111",
  15993=>"010000000",
  15994=>"110111111",
  15995=>"000001110",
  15996=>"001001100",
  15997=>"100100100",
  15998=>"000111011",
  15999=>"111000000",
  16000=>"000000111",
  16001=>"000000000",
  16002=>"000010111",
  16003=>"000000111",
  16004=>"010000000",
  16005=>"100111110",
  16006=>"001101101",
  16007=>"010011001",
  16008=>"011011001",
  16009=>"000000001",
  16010=>"111000100",
  16011=>"001010111",
  16012=>"000111111",
  16013=>"000000010",
  16014=>"000111111",
  16015=>"101000110",
  16016=>"110100100",
  16017=>"111101111",
  16018=>"000010111",
  16019=>"100000010",
  16020=>"111000101",
  16021=>"000010111",
  16022=>"001111011",
  16023=>"000001001",
  16024=>"111111111",
  16025=>"000000110",
  16026=>"000000100",
  16027=>"000000100",
  16028=>"000001001",
  16029=>"010010111",
  16030=>"000100001",
  16031=>"101000000",
  16032=>"101111111",
  16033=>"100100000",
  16034=>"001111111",
  16035=>"000011111",
  16036=>"010000100",
  16037=>"100000000",
  16038=>"111000110",
  16039=>"010111111",
  16040=>"100010111",
  16041=>"000000000",
  16042=>"100110110",
  16043=>"000000000",
  16044=>"110000100",
  16045=>"111111000",
  16046=>"111101000",
  16047=>"111000000",
  16048=>"111011010",
  16049=>"011111011",
  16050=>"000010101",
  16051=>"000001110",
  16052=>"111101101",
  16053=>"100100101",
  16054=>"000000000",
  16055=>"010110101",
  16056=>"100110100",
  16057=>"111001000",
  16058=>"011000111",
  16059=>"101000000",
  16060=>"101111101",
  16061=>"000111101",
  16062=>"110011100",
  16063=>"000000001",
  16064=>"111000000",
  16065=>"001001000",
  16066=>"111000010",
  16067=>"011000001",
  16068=>"010010000",
  16069=>"110000101",
  16070=>"100000001",
  16071=>"011000111",
  16072=>"000111111",
  16073=>"000000101",
  16074=>"000001101",
  16075=>"000010000",
  16076=>"000000001",
  16077=>"100101001",
  16078=>"000000010",
  16079=>"010010000",
  16080=>"000111011",
  16081=>"111101110",
  16082=>"000000010",
  16083=>"011011001",
  16084=>"111000010",
  16085=>"001111100",
  16086=>"000111000",
  16087=>"000100000",
  16088=>"100000000",
  16089=>"110010000",
  16090=>"100101101",
  16091=>"000000110",
  16092=>"001011111",
  16093=>"000011000",
  16094=>"111011000",
  16095=>"000000000",
  16096=>"000011001",
  16097=>"111010100",
  16098=>"000011010",
  16099=>"111111000",
  16100=>"111000000",
  16101=>"101101100",
  16102=>"100110000",
  16103=>"111011011",
  16104=>"111010101",
  16105=>"000100111",
  16106=>"100100010",
  16107=>"001010000",
  16108=>"000001000",
  16109=>"000111111",
  16110=>"001000000",
  16111=>"101000101",
  16112=>"000000010",
  16113=>"011000101",
  16114=>"111000000",
  16115=>"011011001",
  16116=>"110110110",
  16117=>"100001101",
  16118=>"000000000",
  16119=>"111111111",
  16120=>"000111011",
  16121=>"000000000",
  16122=>"000101101",
  16123=>"111001001",
  16124=>"000111111",
  16125=>"000000110",
  16126=>"100101111",
  16127=>"101001100",
  16128=>"011010100",
  16129=>"110010110",
  16130=>"101000001",
  16131=>"111000000",
  16132=>"100000000",
  16133=>"110111001",
  16134=>"100010111",
  16135=>"010111111",
  16136=>"000000000",
  16137=>"001000110",
  16138=>"001110110",
  16139=>"111111000",
  16140=>"010100000",
  16141=>"111110110",
  16142=>"111111100",
  16143=>"111110111",
  16144=>"001000000",
  16145=>"000000100",
  16146=>"111101111",
  16147=>"011010100",
  16148=>"101111000",
  16149=>"111111000",
  16150=>"001000000",
  16151=>"000000101",
  16152=>"000000101",
  16153=>"111111001",
  16154=>"111101000",
  16155=>"011000000",
  16156=>"110000000",
  16157=>"101110111",
  16158=>"010000111",
  16159=>"000110000",
  16160=>"111101000",
  16161=>"001011000",
  16162=>"000000111",
  16163=>"010010010",
  16164=>"100101000",
  16165=>"110000010",
  16166=>"111001110",
  16167=>"000000111",
  16168=>"011110010",
  16169=>"001011011",
  16170=>"111001001",
  16171=>"111100010",
  16172=>"111111011",
  16173=>"111110000",
  16174=>"110011101",
  16175=>"000000011",
  16176=>"110001000",
  16177=>"001001101",
  16178=>"000000000",
  16179=>"010000010",
  16180=>"000111111",
  16181=>"010110110",
  16182=>"100100111",
  16183=>"111100000",
  16184=>"001000001",
  16185=>"111101001",
  16186=>"100101000",
  16187=>"000000000",
  16188=>"101000000",
  16189=>"010101111",
  16190=>"100000000",
  16191=>"111100100",
  16192=>"001000000",
  16193=>"111000000",
  16194=>"111111000",
  16195=>"001111010",
  16196=>"110100000",
  16197=>"000000101",
  16198=>"110010111",
  16199=>"000111111",
  16200=>"001011111",
  16201=>"000111111",
  16202=>"101101000",
  16203=>"111101111",
  16204=>"111000111",
  16205=>"011101001",
  16206=>"100100101",
  16207=>"000000101",
  16208=>"000111110",
  16209=>"110111111",
  16210=>"111111010",
  16211=>"011100010",
  16212=>"110110000",
  16213=>"001000000",
  16214=>"101000110",
  16215=>"000000000",
  16216=>"111111110",
  16217=>"000101111",
  16218=>"101100111",
  16219=>"000111111",
  16220=>"110000100",
  16221=>"001101000",
  16222=>"111100000",
  16223=>"101101111",
  16224=>"111010000",
  16225=>"000100010",
  16226=>"100000000",
  16227=>"001101110",
  16228=>"111011000",
  16229=>"111111110",
  16230=>"111000001",
  16231=>"101011111",
  16232=>"000000000",
  16233=>"001000000",
  16234=>"010000000",
  16235=>"111111111",
  16236=>"001111111",
  16237=>"110110000",
  16238=>"010110100",
  16239=>"011001111",
  16240=>"001000001",
  16241=>"000000001",
  16242=>"001001011",
  16243=>"000010000",
  16244=>"111011011",
  16245=>"000000101",
  16246=>"101000000",
  16247=>"010010010",
  16248=>"111000101",
  16249=>"110000000",
  16250=>"111101000",
  16251=>"000000110",
  16252=>"100010110",
  16253=>"000001001",
  16254=>"000101111",
  16255=>"100101011",
  16256=>"000000000",
  16257=>"100111101",
  16258=>"110010000",
  16259=>"101110111",
  16260=>"000110111",
  16261=>"101111111",
  16262=>"011011111",
  16263=>"101100000",
  16264=>"100100000",
  16265=>"000011111",
  16266=>"111010010",
  16267=>"101111000",
  16268=>"110000000",
  16269=>"000100110",
  16270=>"111111101",
  16271=>"100000000",
  16272=>"100101101",
  16273=>"111001010",
  16274=>"010000000",
  16275=>"011000000",
  16276=>"100000000",
  16277=>"110000000",
  16278=>"010111000",
  16279=>"110100100",
  16280=>"010000110",
  16281=>"100111010",
  16282=>"001001100",
  16283=>"000000000",
  16284=>"111110100",
  16285=>"000000100",
  16286=>"010001101",
  16287=>"101101000",
  16288=>"001100100",
  16289=>"000000010",
  16290=>"000101101",
  16291=>"000000000",
  16292=>"110111011",
  16293=>"110111001",
  16294=>"001110001",
  16295=>"111011111",
  16296=>"011010000",
  16297=>"111000000",
  16298=>"111000000",
  16299=>"000001111",
  16300=>"000100000",
  16301=>"100100000",
  16302=>"100111110",
  16303=>"000110101",
  16304=>"101101101",
  16305=>"101011001",
  16306=>"000000100",
  16307=>"000010011",
  16308=>"000001100",
  16309=>"000100100",
  16310=>"111011011",
  16311=>"010000101",
  16312=>"101000000",
  16313=>"110000000",
  16314=>"010111001",
  16315=>"011100010",
  16316=>"010000010",
  16317=>"111111111",
  16318=>"011010000",
  16319=>"000000011",
  16320=>"000111100",
  16321=>"011001001",
  16322=>"110111010",
  16323=>"011001000",
  16324=>"111000100",
  16325=>"110110101",
  16326=>"110010111",
  16327=>"000000000",
  16328=>"111011101",
  16329=>"111010000",
  16330=>"111111111",
  16331=>"111101100",
  16332=>"010100110",
  16333=>"001011011",
  16334=>"000000111",
  16335=>"000111010",
  16336=>"110110111",
  16337=>"110001001",
  16338=>"111000001",
  16339=>"110111011",
  16340=>"111101001",
  16341=>"101100010",
  16342=>"111111000",
  16343=>"100000010",
  16344=>"010000000",
  16345=>"111111010",
  16346=>"100000111",
  16347=>"000000111",
  16348=>"000001000",
  16349=>"111111000",
  16350=>"011111101",
  16351=>"000000000",
  16352=>"101000101",
  16353=>"001001111",
  16354=>"010000011",
  16355=>"111001101",
  16356=>"111000000",
  16357=>"001111010",
  16358=>"111011010",
  16359=>"111101100",
  16360=>"111011010",
  16361=>"000000110",
  16362=>"000011011",
  16363=>"111001000",
  16364=>"000000010",
  16365=>"000010110",
  16366=>"111000010",
  16367=>"000111111",
  16368=>"010111010",
  16369=>"001001001",
  16370=>"111000010",
  16371=>"000110111",
  16372=>"110110001",
  16373=>"000101111",
  16374=>"000111110",
  16375=>"000100111",
  16376=>"010000100",
  16377=>"000010111",
  16378=>"111111111",
  16379=>"111101000",
  16380=>"000101111",
  16381=>"111010000",
  16382=>"001011000",
  16383=>"000111111",
  16384=>"001001111",
  16385=>"000001000",
  16386=>"011000100",
  16387=>"000111000",
  16388=>"111011111",
  16389=>"001001000",
  16390=>"000000011",
  16391=>"111110111",
  16392=>"101000111",
  16393=>"000000001",
  16394=>"110011011",
  16395=>"000111101",
  16396=>"111001000",
  16397=>"111101100",
  16398=>"110000100",
  16399=>"000010010",
  16400=>"111100011",
  16401=>"111000011",
  16402=>"110111100",
  16403=>"001000001",
  16404=>"000001101",
  16405=>"011001000",
  16406=>"000000100",
  16407=>"001111110",
  16408=>"100000110",
  16409=>"000000000",
  16410=>"000111111",
  16411=>"000000100",
  16412=>"000111010",
  16413=>"000111100",
  16414=>"101111101",
  16415=>"000000000",
  16416=>"000000000",
  16417=>"100111111",
  16418=>"010110001",
  16419=>"000000000",
  16420=>"110111100",
  16421=>"000011010",
  16422=>"000111110",
  16423=>"110000111",
  16424=>"000001000",
  16425=>"001111111",
  16426=>"000000010",
  16427=>"000000100",
  16428=>"100000111",
  16429=>"111111111",
  16430=>"000000111",
  16431=>"110111110",
  16432=>"101111110",
  16433=>"111111100",
  16434=>"011100010",
  16435=>"000101101",
  16436=>"111111000",
  16437=>"001101111",
  16438=>"000000101",
  16439=>"111111110",
  16440=>"000001100",
  16441=>"000000111",
  16442=>"001000000",
  16443=>"000001000",
  16444=>"001100011",
  16445=>"111111011",
  16446=>"101001001",
  16447=>"111111100",
  16448=>"001010011",
  16449=>"111111100",
  16450=>"110111001",
  16451=>"101101111",
  16452=>"000000111",
  16453=>"101101101",
  16454=>"000000011",
  16455=>"110011011",
  16456=>"100111111",
  16457=>"100111111",
  16458=>"000000000",
  16459=>"000000000",
  16460=>"111111111",
  16461=>"111000010",
  16462=>"111111001",
  16463=>"111000000",
  16464=>"111000000",
  16465=>"111111000",
  16466=>"101111000",
  16467=>"000100101",
  16468=>"000000111",
  16469=>"010110110",
  16470=>"110010000",
  16471=>"000000110",
  16472=>"000001100",
  16473=>"111111110",
  16474=>"110000101",
  16475=>"111111011",
  16476=>"110010111",
  16477=>"000000001",
  16478=>"100110000",
  16479=>"001000110",
  16480=>"000111011",
  16481=>"000000001",
  16482=>"011011001",
  16483=>"111011000",
  16484=>"000000001",
  16485=>"010111101",
  16486=>"000111111",
  16487=>"000101000",
  16488=>"000111111",
  16489=>"111111111",
  16490=>"000010111",
  16491=>"101000101",
  16492=>"111110111",
  16493=>"111110010",
  16494=>"101000001",
  16495=>"000111111",
  16496=>"111111111",
  16497=>"110000110",
  16498=>"000001100",
  16499=>"111111011",
  16500=>"111111000",
  16501=>"001011001",
  16502=>"110010001",
  16503=>"000001000",
  16504=>"000000111",
  16505=>"000000111",
  16506=>"111111011",
  16507=>"101111100",
  16508=>"011001001",
  16509=>"000001011",
  16510=>"000001000",
  16511=>"001001001",
  16512=>"000000100",
  16513=>"000000011",
  16514=>"100111111",
  16515=>"111000000",
  16516=>"111111000",
  16517=>"100100110",
  16518=>"000100110",
  16519=>"111000000",
  16520=>"110110000",
  16521=>"000101111",
  16522=>"000111000",
  16523=>"111011000",
  16524=>"000000110",
  16525=>"001001001",
  16526=>"000000000",
  16527=>"000000000",
  16528=>"111111000",
  16529=>"100100000",
  16530=>"000001010",
  16531=>"000000010",
  16532=>"111000000",
  16533=>"000000111",
  16534=>"111110000",
  16535=>"100101100",
  16536=>"111001000",
  16537=>"001000000",
  16538=>"000010010",
  16539=>"010010000",
  16540=>"010001101",
  16541=>"000000000",
  16542=>"000001101",
  16543=>"000000111",
  16544=>"111011100",
  16545=>"111110000",
  16546=>"000000111",
  16547=>"111000000",
  16548=>"100100000",
  16549=>"111000000",
  16550=>"000000011",
  16551=>"000000111",
  16552=>"001000011",
  16553=>"110010000",
  16554=>"111111011",
  16555=>"001000000",
  16556=>"111001110",
  16557=>"111111100",
  16558=>"010011011",
  16559=>"111000001",
  16560=>"100000000",
  16561=>"111000110",
  16562=>"000000001",
  16563=>"111001001",
  16564=>"111100100",
  16565=>"000111110",
  16566=>"011011010",
  16567=>"100000010",
  16568=>"000001110",
  16569=>"110000010",
  16570=>"000000000",
  16571=>"000101111",
  16572=>"101000000",
  16573=>"010010100",
  16574=>"111111011",
  16575=>"111110101",
  16576=>"000100111",
  16577=>"100000110",
  16578=>"101000010",
  16579=>"101101000",
  16580=>"000111111",
  16581=>"011111111",
  16582=>"100000000",
  16583=>"000000111",
  16584=>"111101110",
  16585=>"001000000",
  16586=>"101110000",
  16587=>"110101100",
  16588=>"011110110",
  16589=>"100000100",
  16590=>"110000000",
  16591=>"000011000",
  16592=>"010110110",
  16593=>"111111001",
  16594=>"000000101",
  16595=>"110010011",
  16596=>"111000001",
  16597=>"111000011",
  16598=>"000011111",
  16599=>"000110111",
  16600=>"000110111",
  16601=>"000000001",
  16602=>"111100011",
  16603=>"111000000",
  16604=>"000000100",
  16605=>"111010000",
  16606=>"000000000",
  16607=>"101001000",
  16608=>"111000100",
  16609=>"111100001",
  16610=>"101110010",
  16611=>"011110110",
  16612=>"111100000",
  16613=>"111110101",
  16614=>"000001110",
  16615=>"000000100",
  16616=>"101001000",
  16617=>"000000100",
  16618=>"101100110",
  16619=>"000000001",
  16620=>"000000100",
  16621=>"111111001",
  16622=>"111000000",
  16623=>"000000000",
  16624=>"000001111",
  16625=>"100111111",
  16626=>"101111101",
  16627=>"111011011",
  16628=>"000000001",
  16629=>"111000000",
  16630=>"111000000",
  16631=>"111111001",
  16632=>"000000111",
  16633=>"111111111",
  16634=>"000000000",
  16635=>"000000000",
  16636=>"111111000",
  16637=>"000111111",
  16638=>"111000001",
  16639=>"111111110",
  16640=>"110100000",
  16641=>"000101101",
  16642=>"111101100",
  16643=>"010110000",
  16644=>"111000110",
  16645=>"110000000",
  16646=>"010110010",
  16647=>"011001110",
  16648=>"010000100",
  16649=>"111101100",
  16650=>"010000000",
  16651=>"000010011",
  16652=>"111100000",
  16653=>"000000011",
  16654=>"110100100",
  16655=>"110111100",
  16656=>"000011011",
  16657=>"010000000",
  16658=>"011111000",
  16659=>"010000000",
  16660=>"110111101",
  16661=>"111001100",
  16662=>"001101111",
  16663=>"010111101",
  16664=>"010010000",
  16665=>"000100111",
  16666=>"000000000",
  16667=>"000001111",
  16668=>"001000000",
  16669=>"010011010",
  16670=>"001100010",
  16671=>"111010001",
  16672=>"101000010",
  16673=>"000010011",
  16674=>"111000100",
  16675=>"000101000",
  16676=>"000100111",
  16677=>"011011111",
  16678=>"111100100",
  16679=>"000100110",
  16680=>"010011011",
  16681=>"011101100",
  16682=>"000010100",
  16683=>"000000000",
  16684=>"100001011",
  16685=>"110011110",
  16686=>"000011101",
  16687=>"101011100",
  16688=>"111100000",
  16689=>"011001011",
  16690=>"000000000",
  16691=>"111100000",
  16692=>"010001101",
  16693=>"111111111",
  16694=>"001111111",
  16695=>"111010100",
  16696=>"010111000",
  16697=>"011001100",
  16698=>"011000100",
  16699=>"001101100",
  16700=>"010001011",
  16701=>"010111100",
  16702=>"000000000",
  16703=>"001011111",
  16704=>"001101011",
  16705=>"000101111",
  16706=>"111110111",
  16707=>"100000000",
  16708=>"111000000",
  16709=>"111100000",
  16710=>"010000111",
  16711=>"010010000",
  16712=>"000001110",
  16713=>"000011011",
  16714=>"000100000",
  16715=>"111111011",
  16716=>"111101101",
  16717=>"110001101",
  16718=>"100100111",
  16719=>"001111100",
  16720=>"100100111",
  16721=>"010010111",
  16722=>"101111111",
  16723=>"000011000",
  16724=>"111101101",
  16725=>"111011011",
  16726=>"000000000",
  16727=>"000100000",
  16728=>"000010110",
  16729=>"001001101",
  16730=>"110001001",
  16731=>"100100110",
  16732=>"010000111",
  16733=>"010000001",
  16734=>"111100000",
  16735=>"100100100",
  16736=>"000000010",
  16737=>"000010011",
  16738=>"001000100",
  16739=>"001001101",
  16740=>"011000000",
  16741=>"010100011",
  16742=>"000010011",
  16743=>"111100100",
  16744=>"001011011",
  16745=>"111110111",
  16746=>"001001010",
  16747=>"111111111",
  16748=>"110110000",
  16749=>"111111101",
  16750=>"000000000",
  16751=>"010001001",
  16752=>"000110110",
  16753=>"000100010",
  16754=>"011111110",
  16755=>"000001000",
  16756=>"010101110",
  16757=>"111100100",
  16758=>"011111010",
  16759=>"000011010",
  16760=>"110000100",
  16761=>"111000100",
  16762=>"011111010",
  16763=>"011100100",
  16764=>"011111100",
  16765=>"011110000",
  16766=>"000100000",
  16767=>"001001000",
  16768=>"111111000",
  16769=>"000010000",
  16770=>"010001000",
  16771=>"111011111",
  16772=>"101101110",
  16773=>"111000000",
  16774=>"100110100",
  16775=>"000100111",
  16776=>"000001001",
  16777=>"001000000",
  16778=>"000001011",
  16779=>"100100000",
  16780=>"110010000",
  16781=>"111101100",
  16782=>"001000000",
  16783=>"000100000",
  16784=>"111100111",
  16785=>"011111111",
  16786=>"011101100",
  16787=>"000111111",
  16788=>"000111111",
  16789=>"111000000",
  16790=>"101011110",
  16791=>"010010100",
  16792=>"000001011",
  16793=>"111000001",
  16794=>"000000111",
  16795=>"000000000",
  16796=>"110100100",
  16797=>"000011011",
  16798=>"111111000",
  16799=>"100100000",
  16800=>"001000100",
  16801=>"010000000",
  16802=>"101010100",
  16803=>"011000000",
  16804=>"111101101",
  16805=>"010000001",
  16806=>"011011001",
  16807=>"000011111",
  16808=>"010001101",
  16809=>"000000000",
  16810=>"111000100",
  16811=>"000111010",
  16812=>"111111011",
  16813=>"010000000",
  16814=>"110011111",
  16815=>"011011011",
  16816=>"000100001",
  16817=>"000011000",
  16818=>"011111111",
  16819=>"000101000",
  16820=>"000000110",
  16821=>"111110111",
  16822=>"011111011",
  16823=>"111100000",
  16824=>"001100011",
  16825=>"001111111",
  16826=>"000010011",
  16827=>"000110010",
  16828=>"111110000",
  16829=>"010111111",
  16830=>"010000000",
  16831=>"011111001",
  16832=>"000001000",
  16833=>"010110100",
  16834=>"000000100",
  16835=>"011001000",
  16836=>"000010010",
  16837=>"110111011",
  16838=>"111010100",
  16839=>"001101101",
  16840=>"000100010",
  16841=>"010010010",
  16842=>"101000101",
  16843=>"000100111",
  16844=>"000011011",
  16845=>"100001011",
  16846=>"111110110",
  16847=>"110100000",
  16848=>"000010010",
  16849=>"110100101",
  16850=>"000000010",
  16851=>"011111111",
  16852=>"000000011",
  16853=>"011100100",
  16854=>"011101000",
  16855=>"100111000",
  16856=>"000100100",
  16857=>"001011111",
  16858=>"010110100",
  16859=>"110000000",
  16860=>"110111101",
  16861=>"110010001",
  16862=>"011010101",
  16863=>"000010010",
  16864=>"111101001",
  16865=>"111111101",
  16866=>"111101101",
  16867=>"000001001",
  16868=>"100100000",
  16869=>"011001100",
  16870=>"100110100",
  16871=>"010000000",
  16872=>"000000111",
  16873=>"110111010",
  16874=>"000000000",
  16875=>"111100000",
  16876=>"010010011",
  16877=>"111100000",
  16878=>"000000000",
  16879=>"111110000",
  16880=>"001100100",
  16881=>"001111100",
  16882=>"010111100",
  16883=>"000000100",
  16884=>"010110101",
  16885=>"101100100",
  16886=>"100000000",
  16887=>"110000100",
  16888=>"000111111",
  16889=>"101001100",
  16890=>"111101111",
  16891=>"100000101",
  16892=>"101011001",
  16893=>"000000010",
  16894=>"011011101",
  16895=>"000100000",
  16896=>"000011011",
  16897=>"011011111",
  16898=>"101100000",
  16899=>"000100010",
  16900=>"000000100",
  16901=>"111111100",
  16902=>"100000110",
  16903=>"001000011",
  16904=>"000000011",
  16905=>"000111111",
  16906=>"101100000",
  16907=>"010011001",
  16908=>"000000110",
  16909=>"000000000",
  16910=>"101101001",
  16911=>"000000011",
  16912=>"011111111",
  16913=>"010010011",
  16914=>"110100000",
  16915=>"011100000",
  16916=>"101111110",
  16917=>"000011010",
  16918=>"100100100",
  16919=>"111111110",
  16920=>"000000011",
  16921=>"010111101",
  16922=>"010111100",
  16923=>"010010110",
  16924=>"111100100",
  16925=>"000100100",
  16926=>"111010000",
  16927=>"000111111",
  16928=>"000110000",
  16929=>"011111011",
  16930=>"100010011",
  16931=>"000101111",
  16932=>"010011001",
  16933=>"001101100",
  16934=>"000000000",
  16935=>"100001000",
  16936=>"001111101",
  16937=>"001111011",
  16938=>"100000000",
  16939=>"000000000",
  16940=>"000001001",
  16941=>"011000011",
  16942=>"110000100",
  16943=>"001110100",
  16944=>"100101111",
  16945=>"001011111",
  16946=>"111011011",
  16947=>"100100100",
  16948=>"111000000",
  16949=>"101000001",
  16950=>"110100001",
  16951=>"000000010",
  16952=>"111000110",
  16953=>"111101000",
  16954=>"111100100",
  16955=>"111101101",
  16956=>"011010001",
  16957=>"111111110",
  16958=>"000000110",
  16959=>"001111111",
  16960=>"000111010",
  16961=>"011111100",
  16962=>"000000110",
  16963=>"111011001",
  16964=>"111100010",
  16965=>"001010011",
  16966=>"101000000",
  16967=>"111111000",
  16968=>"010110111",
  16969=>"001011011",
  16970=>"101000000",
  16971=>"011100001",
  16972=>"111111000",
  16973=>"001110100",
  16974=>"000110111",
  16975=>"111101111",
  16976=>"101111000",
  16977=>"110111101",
  16978=>"000100010",
  16979=>"011001000",
  16980=>"111000000",
  16981=>"110110111",
  16982=>"011011001",
  16983=>"010001111",
  16984=>"111101001",
  16985=>"001110001",
  16986=>"000111111",
  16987=>"010111111",
  16988=>"000000000",
  16989=>"110001001",
  16990=>"111111100",
  16991=>"111100000",
  16992=>"000011111",
  16993=>"111111101",
  16994=>"111100111",
  16995=>"100000000",
  16996=>"111111111",
  16997=>"111110110",
  16998=>"111110111",
  16999=>"000000111",
  17000=>"101000010",
  17001=>"011010000",
  17002=>"010000111",
  17003=>"111111000",
  17004=>"111111111",
  17005=>"000000010",
  17006=>"000111010",
  17007=>"011010111",
  17008=>"101111001",
  17009=>"000100110",
  17010=>"111001000",
  17011=>"000011001",
  17012=>"000001001",
  17013=>"110000000",
  17014=>"000000000",
  17015=>"000001000",
  17016=>"000000000",
  17017=>"111011100",
  17018=>"110111111",
  17019=>"000000100",
  17020=>"000110111",
  17021=>"011110000",
  17022=>"000000000",
  17023=>"111000101",
  17024=>"000010100",
  17025=>"111100000",
  17026=>"001111111",
  17027=>"000000011",
  17028=>"011011011",
  17029=>"111111100",
  17030=>"100011001",
  17031=>"000000001",
  17032=>"101100100",
  17033=>"001000000",
  17034=>"000000001",
  17035=>"011011000",
  17036=>"000100111",
  17037=>"000000000",
  17038=>"100000000",
  17039=>"100000101",
  17040=>"111111001",
  17041=>"100111101",
  17042=>"101000001",
  17043=>"110000000",
  17044=>"001010011",
  17045=>"111000010",
  17046=>"111111111",
  17047=>"000011011",
  17048=>"011011111",
  17049=>"000000111",
  17050=>"111000100",
  17051=>"000100110",
  17052=>"111100100",
  17053=>"010111011",
  17054=>"100000100",
  17055=>"111000000",
  17056=>"001000001",
  17057=>"110000010",
  17058=>"100010110",
  17059=>"000000111",
  17060=>"011011001",
  17061=>"100011111",
  17062=>"001110111",
  17063=>"010111111",
  17064=>"111011111",
  17065=>"000010011",
  17066=>"101110110",
  17067=>"111100100",
  17068=>"010000000",
  17069=>"001001001",
  17070=>"001100100",
  17071=>"000000011",
  17072=>"100011111",
  17073=>"000011001",
  17074=>"111111111",
  17075=>"000010010",
  17076=>"010111011",
  17077=>"000000011",
  17078=>"000111011",
  17079=>"001000000",
  17080=>"110101011",
  17081=>"100000110",
  17082=>"111111001",
  17083=>"101111010",
  17084=>"010110010",
  17085=>"111111111",
  17086=>"000110011",
  17087=>"101001111",
  17088=>"111100100",
  17089=>"111101110",
  17090=>"111101111",
  17091=>"000110010",
  17092=>"101101000",
  17093=>"011000101",
  17094=>"110100000",
  17095=>"000100000",
  17096=>"000010010",
  17097=>"000100001",
  17098=>"000011111",
  17099=>"000011011",
  17100=>"100101111",
  17101=>"100001011",
  17102=>"100100110",
  17103=>"010111000",
  17104=>"000100000",
  17105=>"000110000",
  17106=>"000011011",
  17107=>"001011001",
  17108=>"011100100",
  17109=>"010110110",
  17110=>"100000010",
  17111=>"000011011",
  17112=>"001011000",
  17113=>"111000101",
  17114=>"100100100",
  17115=>"100000000",
  17116=>"001111011",
  17117=>"010011111",
  17118=>"101111111",
  17119=>"111010000",
  17120=>"101000100",
  17121=>"101100100",
  17122=>"000000000",
  17123=>"000000110",
  17124=>"101000000",
  17125=>"000000000",
  17126=>"000001000",
  17127=>"000001001",
  17128=>"000000010",
  17129=>"000001010",
  17130=>"111001000",
  17131=>"000000001",
  17132=>"000000111",
  17133=>"000000001",
  17134=>"000100000",
  17135=>"000101010",
  17136=>"111111000",
  17137=>"010100101",
  17138=>"010010011",
  17139=>"000111011",
  17140=>"100110100",
  17141=>"000000101",
  17142=>"010000010",
  17143=>"000111011",
  17144=>"111010010",
  17145=>"100111111",
  17146=>"000000000",
  17147=>"011101101",
  17148=>"101000010",
  17149=>"100111011",
  17150=>"000000001",
  17151=>"101000000",
  17152=>"011001000",
  17153=>"010000111",
  17154=>"010011010",
  17155=>"101000000",
  17156=>"111110111",
  17157=>"000001000",
  17158=>"110100010",
  17159=>"000000111",
  17160=>"111111111",
  17161=>"001000000",
  17162=>"110110110",
  17163=>"001101001",
  17164=>"101101101",
  17165=>"000001000",
  17166=>"001011011",
  17167=>"111110010",
  17168=>"111111001",
  17169=>"110000000",
  17170=>"110000000",
  17171=>"000000111",
  17172=>"110000100",
  17173=>"111100100",
  17174=>"011011101",
  17175=>"110111111",
  17176=>"100100110",
  17177=>"001001101",
  17178=>"101101101",
  17179=>"111010010",
  17180=>"000000000",
  17181=>"000000010",
  17182=>"000000000",
  17183=>"101001101",
  17184=>"100101111",
  17185=>"111111011",
  17186=>"010110110",
  17187=>"110000110",
  17188=>"110110100",
  17189=>"011011111",
  17190=>"010000000",
  17191=>"111111111",
  17192=>"111111011",
  17193=>"011011001",
  17194=>"000000111",
  17195=>"101000100",
  17196=>"010111011",
  17197=>"000000000",
  17198=>"000000000",
  17199=>"000100000",
  17200=>"000000100",
  17201=>"111111011",
  17202=>"000000100",
  17203=>"000000000",
  17204=>"011110110",
  17205=>"101011110",
  17206=>"111111111",
  17207=>"000100011",
  17208=>"000000000",
  17209=>"000000111",
  17210=>"000010100",
  17211=>"111000000",
  17212=>"000000001",
  17213=>"011101001",
  17214=>"100100100",
  17215=>"111111111",
  17216=>"000000000",
  17217=>"101111111",
  17218=>"000100000",
  17219=>"010001001",
  17220=>"000000110",
  17221=>"001101101",
  17222=>"100101100",
  17223=>"001001001",
  17224=>"000000000",
  17225=>"101101101",
  17226=>"101101100",
  17227=>"101011101",
  17228=>"000000000",
  17229=>"111111111",
  17230=>"111111011",
  17231=>"111101110",
  17232=>"001101000",
  17233=>"111001000",
  17234=>"000000100",
  17235=>"011000010",
  17236=>"010111111",
  17237=>"100100100",
  17238=>"111111001",
  17239=>"000100100",
  17240=>"101111111",
  17241=>"001011111",
  17242=>"111111110",
  17243=>"001000101",
  17244=>"101000111",
  17245=>"011011011",
  17246=>"010111011",
  17247=>"000100100",
  17248=>"111111111",
  17249=>"101000101",
  17250=>"100000000",
  17251=>"111111011",
  17252=>"101111110",
  17253=>"111111111",
  17254=>"111111100",
  17255=>"011000111",
  17256=>"000000000",
  17257=>"000000011",
  17258=>"000000001",
  17259=>"010011001",
  17260=>"010101001",
  17261=>"111011011",
  17262=>"111000000",
  17263=>"000000000",
  17264=>"100100100",
  17265=>"000000010",
  17266=>"111011111",
  17267=>"011111010",
  17268=>"000000000",
  17269=>"000101101",
  17270=>"000000000",
  17271=>"011111000",
  17272=>"000010011",
  17273=>"000000000",
  17274=>"000011010",
  17275=>"111111111",
  17276=>"001000110",
  17277=>"110110110",
  17278=>"111000000",
  17279=>"010111010",
  17280=>"000000000",
  17281=>"000000100",
  17282=>"000000000",
  17283=>"000000000",
  17284=>"000000000",
  17285=>"000000100",
  17286=>"110110110",
  17287=>"011011011",
  17288=>"011011001",
  17289=>"010011010",
  17290=>"011011010",
  17291=>"110100100",
  17292=>"101111011",
  17293=>"111101110",
  17294=>"101001110",
  17295=>"101101100",
  17296=>"111110110",
  17297=>"111111110",
  17298=>"001010000",
  17299=>"000000000",
  17300=>"101110110",
  17301=>"110100101",
  17302=>"110111011",
  17303=>"001101111",
  17304=>"000100111",
  17305=>"000000111",
  17306=>"000010011",
  17307=>"000000000",
  17308=>"000000000",
  17309=>"000000010",
  17310=>"000000000",
  17311=>"110011000",
  17312=>"011111011",
  17313=>"000000000",
  17314=>"111011000",
  17315=>"000000000",
  17316=>"000000000",
  17317=>"110101110",
  17318=>"101011111",
  17319=>"111111111",
  17320=>"000000001",
  17321=>"000001010",
  17322=>"000001111",
  17323=>"000000000",
  17324=>"111111111",
  17325=>"000000000",
  17326=>"110101010",
  17327=>"101101100",
  17328=>"000000100",
  17329=>"000001111",
  17330=>"111010111",
  17331=>"100000100",
  17332=>"111111111",
  17333=>"011010000",
  17334=>"000100100",
  17335=>"011000000",
  17336=>"000000100",
  17337=>"001111010",
  17338=>"000000000",
  17339=>"000000000",
  17340=>"111101010",
  17341=>"000110111",
  17342=>"110100110",
  17343=>"000000000",
  17344=>"111100110",
  17345=>"000000101",
  17346=>"000100001",
  17347=>"001001011",
  17348=>"000000000",
  17349=>"100000001",
  17350=>"000000101",
  17351=>"000000111",
  17352=>"111111111",
  17353=>"010010000",
  17354=>"101101110",
  17355=>"111111110",
  17356=>"001000000",
  17357=>"110100111",
  17358=>"111111001",
  17359=>"000000000",
  17360=>"010010000",
  17361=>"111111111",
  17362=>"010010010",
  17363=>"111110100",
  17364=>"001000101",
  17365=>"111111111",
  17366=>"010111010",
  17367=>"000000000",
  17368=>"111111111",
  17369=>"111011011",
  17370=>"110111111",
  17371=>"010011000",
  17372=>"000000000",
  17373=>"000001000",
  17374=>"011100101",
  17375=>"000000000",
  17376=>"010010000",
  17377=>"000000000",
  17378=>"100011011",
  17379=>"111100001",
  17380=>"001000101",
  17381=>"001100111",
  17382=>"000010000",
  17383=>"010001111",
  17384=>"001000000",
  17385=>"111111111",
  17386=>"011111101",
  17387=>"111111100",
  17388=>"100111000",
  17389=>"000000000",
  17390=>"100000000",
  17391=>"100101111",
  17392=>"010010010",
  17393=>"101000001",
  17394=>"000110000",
  17395=>"111111111",
  17396=>"110000001",
  17397=>"111111111",
  17398=>"001001000",
  17399=>"000000000",
  17400=>"111111111",
  17401=>"000000000",
  17402=>"111000101",
  17403=>"111111010",
  17404=>"111001011",
  17405=>"111010111",
  17406=>"111101110",
  17407=>"011110000",
  17408=>"011111001",
  17409=>"001000000",
  17410=>"111101100",
  17411=>"010000000",
  17412=>"000111011",
  17413=>"000000000",
  17414=>"111000101",
  17415=>"101101110",
  17416=>"010010011",
  17417=>"000000000",
  17418=>"111001111",
  17419=>"000011111",
  17420=>"000101010",
  17421=>"010001000",
  17422=>"000111111",
  17423=>"111111000",
  17424=>"010100000",
  17425=>"000100101",
  17426=>"000000100",
  17427=>"000010010",
  17428=>"101000000",
  17429=>"101100000",
  17430=>"111111000",
  17431=>"111110111",
  17432=>"000000000",
  17433=>"101001111",
  17434=>"111110011",
  17435=>"110000000",
  17436=>"011000000",
  17437=>"001101001",
  17438=>"011010000",
  17439=>"000000111",
  17440=>"110101001",
  17441=>"100101010",
  17442=>"000000110",
  17443=>"000111111",
  17444=>"111101101",
  17445=>"011111110",
  17446=>"100000010",
  17447=>"101000000",
  17448=>"111000111",
  17449=>"101010000",
  17450=>"001010000",
  17451=>"101100000",
  17452=>"001011001",
  17453=>"110000011",
  17454=>"001011000",
  17455=>"010111101",
  17456=>"001111100",
  17457=>"000111011",
  17458=>"011000111",
  17459=>"000000000",
  17460=>"000110000",
  17461=>"100111111",
  17462=>"011110000",
  17463=>"010111111",
  17464=>"111101111",
  17465=>"111101001",
  17466=>"100101110",
  17467=>"001010010",
  17468=>"000011111",
  17469=>"100011111",
  17470=>"011101000",
  17471=>"110011011",
  17472=>"100111111",
  17473=>"001111111",
  17474=>"000000101",
  17475=>"110000110",
  17476=>"010010000",
  17477=>"101101010",
  17478=>"100100000",
  17479=>"010001111",
  17480=>"110110110",
  17481=>"000111111",
  17482=>"101100100",
  17483=>"111100100",
  17484=>"000110000",
  17485=>"111101100",
  17486=>"000010110",
  17487=>"011111101",
  17488=>"111100000",
  17489=>"010010000",
  17490=>"000010011",
  17491=>"000011011",
  17492=>"000000111",
  17493=>"010010000",
  17494=>"010011011",
  17495=>"100001101",
  17496=>"000001111",
  17497=>"100100011",
  17498=>"111110100",
  17499=>"000011111",
  17500=>"010001000",
  17501=>"111001001",
  17502=>"111111000",
  17503=>"001010110",
  17504=>"000000011",
  17505=>"000000011",
  17506=>"010000000",
  17507=>"011000000",
  17508=>"000111010",
  17509=>"000000100",
  17510=>"000000000",
  17511=>"100111011",
  17512=>"100001010",
  17513=>"000001111",
  17514=>"111000111",
  17515=>"000101111",
  17516=>"010010010",
  17517=>"111101101",
  17518=>"000000000",
  17519=>"110101001",
  17520=>"011011111",
  17521=>"111001111",
  17522=>"110001000",
  17523=>"000001011",
  17524=>"011111000",
  17525=>"000100001",
  17526=>"000111010",
  17527=>"000000011",
  17528=>"010000000",
  17529=>"110101110",
  17530=>"111001100",
  17531=>"000100011",
  17532=>"011100100",
  17533=>"000110000",
  17534=>"111000000",
  17535=>"000000111",
  17536=>"010010011",
  17537=>"100110101",
  17538=>"000000011",
  17539=>"000111111",
  17540=>"101100000",
  17541=>"000111111",
  17542=>"100110011",
  17543=>"110000011",
  17544=>"011111111",
  17545=>"111111001",
  17546=>"100111000",
  17547=>"000010110",
  17548=>"111000100",
  17549=>"000101101",
  17550=>"110111100",
  17551=>"001101100",
  17552=>"000111111",
  17553=>"111100101",
  17554=>"110100101",
  17555=>"010010111",
  17556=>"100000111",
  17557=>"111000000",
  17558=>"111000101",
  17559=>"100101110",
  17560=>"000000001",
  17561=>"010110111",
  17562=>"111000100",
  17563=>"000100110",
  17564=>"011011110",
  17565=>"000000011",
  17566=>"011111001",
  17567=>"000111111",
  17568=>"111011000",
  17569=>"111000000",
  17570=>"000111111",
  17571=>"111010000",
  17572=>"100111111",
  17573=>"000110110",
  17574=>"000110110",
  17575=>"011111100",
  17576=>"100000000",
  17577=>"000000001",
  17578=>"111000000",
  17579=>"111000000",
  17580=>"100101111",
  17581=>"011000111",
  17582=>"111101001",
  17583=>"111001000",
  17584=>"100101101",
  17585=>"011100111",
  17586=>"000000000",
  17587=>"011001100",
  17588=>"111111111",
  17589=>"100000010",
  17590=>"000100101",
  17591=>"010010011",
  17592=>"000100011",
  17593=>"010000111",
  17594=>"000010010",
  17595=>"011111101",
  17596=>"000011111",
  17597=>"111111111",
  17598=>"000011110",
  17599=>"001000100",
  17600=>"111001000",
  17601=>"001011011",
  17602=>"111111000",
  17603=>"011111110",
  17604=>"000111110",
  17605=>"000100100",
  17606=>"000011111",
  17607=>"111101100",
  17608=>"001000101",
  17609=>"101000000",
  17610=>"000001000",
  17611=>"000010111",
  17612=>"011010000",
  17613=>"111111000",
  17614=>"011101011",
  17615=>"111000000",
  17616=>"110111111",
  17617=>"000111010",
  17618=>"111101110",
  17619=>"101111100",
  17620=>"000000010",
  17621=>"101001010",
  17622=>"010000000",
  17623=>"111001101",
  17624=>"000011011",
  17625=>"100000111",
  17626=>"111111000",
  17627=>"000000000",
  17628=>"111111000",
  17629=>"111000110",
  17630=>"101111111",
  17631=>"010001000",
  17632=>"111000000",
  17633=>"111101100",
  17634=>"100000110",
  17635=>"100110100",
  17636=>"001000100",
  17637=>"000111111",
  17638=>"000111111",
  17639=>"111111001",
  17640=>"000111111",
  17641=>"011110110",
  17642=>"110110111",
  17643=>"001000000",
  17644=>"100000111",
  17645=>"000001000",
  17646=>"000001011",
  17647=>"010010111",
  17648=>"000011111",
  17649=>"010001011",
  17650=>"000000010",
  17651=>"000010110",
  17652=>"010110000",
  17653=>"100100000",
  17654=>"000000010",
  17655=>"000000111",
  17656=>"111010000",
  17657=>"001010000",
  17658=>"011111000",
  17659=>"000101101",
  17660=>"111111000",
  17661=>"000011111",
  17662=>"000111001",
  17663=>"001111000",
  17664=>"010101111",
  17665=>"000010010",
  17666=>"111110000",
  17667=>"000011011",
  17668=>"010000111",
  17669=>"001111111",
  17670=>"100000101",
  17671=>"100000000",
  17672=>"000011111",
  17673=>"110000000",
  17674=>"111100010",
  17675=>"000100100",
  17676=>"000000111",
  17677=>"000111111",
  17678=>"000100011",
  17679=>"111100100",
  17680=>"111000000",
  17681=>"010000000",
  17682=>"111010011",
  17683=>"000000000",
  17684=>"101111001",
  17685=>"110000010",
  17686=>"101111111",
  17687=>"111111010",
  17688=>"000000000",
  17689=>"111001001",
  17690=>"000000000",
  17691=>"000000111",
  17692=>"011000000",
  17693=>"101111110",
  17694=>"010000101",
  17695=>"101001111",
  17696=>"111111001",
  17697=>"101111111",
  17698=>"101101110",
  17699=>"110111111",
  17700=>"110111101",
  17701=>"111001011",
  17702=>"000000000",
  17703=>"011001000",
  17704=>"111000000",
  17705=>"110110000",
  17706=>"000110111",
  17707=>"001000110",
  17708=>"000111111",
  17709=>"000010000",
  17710=>"101111111",
  17711=>"010001100",
  17712=>"000000000",
  17713=>"001110100",
  17714=>"111000111",
  17715=>"000100001",
  17716=>"011000111",
  17717=>"000001110",
  17718=>"110110111",
  17719=>"011111111",
  17720=>"000000110",
  17721=>"110110101",
  17722=>"111010101",
  17723=>"111000111",
  17724=>"000100111",
  17725=>"111001001",
  17726=>"000000100",
  17727=>"001000001",
  17728=>"001000000",
  17729=>"101111011",
  17730=>"001110111",
  17731=>"100110110",
  17732=>"111110100",
  17733=>"001001100",
  17734=>"100100100",
  17735=>"000010110",
  17736=>"111111111",
  17737=>"111000000",
  17738=>"111111001",
  17739=>"000000000",
  17740=>"111000000",
  17741=>"010000111",
  17742=>"001001000",
  17743=>"000000110",
  17744=>"101101100",
  17745=>"111000000",
  17746=>"000000011",
  17747=>"110000001",
  17748=>"000000111",
  17749=>"111010100",
  17750=>"111100101",
  17751=>"111000000",
  17752=>"000001000",
  17753=>"000000011",
  17754=>"000000010",
  17755=>"111000000",
  17756=>"101010000",
  17757=>"110110001",
  17758=>"111000000",
  17759=>"011011011",
  17760=>"000000111",
  17761=>"000101111",
  17762=>"000000001",
  17763=>"001000100",
  17764=>"000000100",
  17765=>"111011111",
  17766=>"111110000",
  17767=>"110110010",
  17768=>"000000000",
  17769=>"111000101",
  17770=>"000000111",
  17771=>"111101110",
  17772=>"000011111",
  17773=>"111000010",
  17774=>"000000010",
  17775=>"000000001",
  17776=>"100011011",
  17777=>"011110111",
  17778=>"011011100",
  17779=>"001101110",
  17780=>"110000000",
  17781=>"100000000",
  17782=>"000000000",
  17783=>"000010111",
  17784=>"001110111",
  17785=>"111101011",
  17786=>"000000000",
  17787=>"011111011",
  17788=>"011011101",
  17789=>"100000100",
  17790=>"101010001",
  17791=>"111111000",
  17792=>"101000001",
  17793=>"111000111",
  17794=>"111010010",
  17795=>"000000110",
  17796=>"000000000",
  17797=>"001111110",
  17798=>"111101111",
  17799=>"111111110",
  17800=>"101100100",
  17801=>"001101000",
  17802=>"000100010",
  17803=>"111111001",
  17804=>"000000000",
  17805=>"111110001",
  17806=>"000000111",
  17807=>"000001001",
  17808=>"000000011",
  17809=>"000000111",
  17810=>"111000000",
  17811=>"000111101",
  17812=>"000110100",
  17813=>"000010111",
  17814=>"111111111",
  17815=>"000000011",
  17816=>"101100111",
  17817=>"111001110",
  17818=>"111011000",
  17819=>"100110000",
  17820=>"000001101",
  17821=>"111011000",
  17822=>"000000111",
  17823=>"000000111",
  17824=>"111010011",
  17825=>"011111010",
  17826=>"111111011",
  17827=>"111100111",
  17828=>"011010111",
  17829=>"100110110",
  17830=>"001001000",
  17831=>"000010110",
  17832=>"111010000",
  17833=>"000000111",
  17834=>"010111111",
  17835=>"100000101",
  17836=>"000001000",
  17837=>"000000111",
  17838=>"111110110",
  17839=>"000100111",
  17840=>"000000111",
  17841=>"110111111",
  17842=>"111000100",
  17843=>"010001110",
  17844=>"000011011",
  17845=>"001011010",
  17846=>"001000100",
  17847=>"000000111",
  17848=>"000010011",
  17849=>"001111111",
  17850=>"000000110",
  17851=>"111111000",
  17852=>"000100010",
  17853=>"110000101",
  17854=>"000000100",
  17855=>"000010101",
  17856=>"111111010",
  17857=>"111111000",
  17858=>"111001010",
  17859=>"101100111",
  17860=>"000000000",
  17861=>"111111011",
  17862=>"000001111",
  17863=>"111111110",
  17864=>"001010110",
  17865=>"000111100",
  17866=>"111111110",
  17867=>"111000101",
  17868=>"111000000",
  17869=>"000100110",
  17870=>"111111000",
  17871=>"110111001",
  17872=>"000000111",
  17873=>"011110111",
  17874=>"110110100",
  17875=>"000000111",
  17876=>"000000111",
  17877=>"111110100",
  17878=>"111111111",
  17879=>"101001100",
  17880=>"000000000",
  17881=>"010001000",
  17882=>"001100110",
  17883=>"110101000",
  17884=>"111101100",
  17885=>"000001111",
  17886=>"000001111",
  17887=>"000000011",
  17888=>"111000000",
  17889=>"000000110",
  17890=>"001000010",
  17891=>"010011001",
  17892=>"010000000",
  17893=>"000000000",
  17894=>"000111111",
  17895=>"111001111",
  17896=>"000110111",
  17897=>"101101111",
  17898=>"111011110",
  17899=>"000010000",
  17900=>"101000000",
  17901=>"100001111",
  17902=>"111000000",
  17903=>"000000110",
  17904=>"010000001",
  17905=>"111111111",
  17906=>"000111110",
  17907=>"010011100",
  17908=>"100100101",
  17909=>"000001000",
  17910=>"101000000",
  17911=>"000001010",
  17912=>"111110000",
  17913=>"001000010",
  17914=>"110101111",
  17915=>"000011011",
  17916=>"011000010",
  17917=>"000110111",
  17918=>"001001111",
  17919=>"100101000",
  17920=>"011001000",
  17921=>"000000101",
  17922=>"000000000",
  17923=>"111101111",
  17924=>"100000000",
  17925=>"001100100",
  17926=>"111111000",
  17927=>"111111111",
  17928=>"111001000",
  17929=>"110111011",
  17930=>"100100110",
  17931=>"001101111",
  17932=>"000000001",
  17933=>"111001000",
  17934=>"101011011",
  17935=>"101111101",
  17936=>"011101011",
  17937=>"000111000",
  17938=>"000010010",
  17939=>"101111111",
  17940=>"111010000",
  17941=>"000000111",
  17942=>"011001111",
  17943=>"010111111",
  17944=>"101000000",
  17945=>"011000111",
  17946=>"111101111",
  17947=>"111011110",
  17948=>"110010111",
  17949=>"000100000",
  17950=>"111000010",
  17951=>"000111011",
  17952=>"101000100",
  17953=>"101001001",
  17954=>"101000010",
  17955=>"111111011",
  17956=>"111110100",
  17957=>"010111000",
  17958=>"101000111",
  17959=>"000110111",
  17960=>"101001111",
  17961=>"111111111",
  17962=>"000000111",
  17963=>"111000010",
  17964=>"111111010",
  17965=>"011000111",
  17966=>"011000000",
  17967=>"111111000",
  17968=>"111000101",
  17969=>"111101100",
  17970=>"111101010",
  17971=>"111000001",
  17972=>"101111100",
  17973=>"011101100",
  17974=>"110111111",
  17975=>"110000111",
  17976=>"000000001",
  17977=>"111010110",
  17978=>"000000111",
  17979=>"111000110",
  17980=>"111110011",
  17981=>"010111010",
  17982=>"000000000",
  17983=>"011001001",
  17984=>"001000000",
  17985=>"111111000",
  17986=>"000001111",
  17987=>"100110100",
  17988=>"100000000",
  17989=>"010000001",
  17990=>"010010000",
  17991=>"110100000",
  17992=>"000010000",
  17993=>"111111000",
  17994=>"000000111",
  17995=>"010110000",
  17996=>"000000000",
  17997=>"111101000",
  17998=>"101101000",
  17999=>"111100111",
  18000=>"111101101",
  18001=>"010111000",
  18002=>"111010000",
  18003=>"011011000",
  18004=>"000000010",
  18005=>"001100110",
  18006=>"111111110",
  18007=>"010110000",
  18008=>"001000100",
  18009=>"101001001",
  18010=>"111110100",
  18011=>"000001000",
  18012=>"010111111",
  18013=>"001000001",
  18014=>"101000011",
  18015=>"101111000",
  18016=>"101001111",
  18017=>"000010111",
  18018=>"000111000",
  18019=>"010001001",
  18020=>"111001000",
  18021=>"111011010",
  18022=>"001000010",
  18023=>"010111001",
  18024=>"000100101",
  18025=>"000000000",
  18026=>"101001000",
  18027=>"000010111",
  18028=>"000000110",
  18029=>"110000000",
  18030=>"000000111",
  18031=>"000000111",
  18032=>"001001100",
  18033=>"111000011",
  18034=>"011011110",
  18035=>"001000100",
  18036=>"101110000",
  18037=>"000000110",
  18038=>"000111111",
  18039=>"000000001",
  18040=>"010000011",
  18041=>"110010111",
  18042=>"101000000",
  18043=>"001000000",
  18044=>"110110110",
  18045=>"100100010",
  18046=>"010001101",
  18047=>"010110100",
  18048=>"000000101",
  18049=>"010000110",
  18050=>"111010000",
  18051=>"111111111",
  18052=>"111101111",
  18053=>"010110111",
  18054=>"011110000",
  18055=>"011010000",
  18056=>"000100000",
  18057=>"011111111",
  18058=>"111111111",
  18059=>"000000010",
  18060=>"000000001",
  18061=>"000000100",
  18062=>"001000000",
  18063=>"000001101",
  18064=>"100100100",
  18065=>"000111000",
  18066=>"000111111",
  18067=>"011000000",
  18068=>"000000111",
  18069=>"111111001",
  18070=>"101001010",
  18071=>"110100100",
  18072=>"010101000",
  18073=>"100010111",
  18074=>"001000111",
  18075=>"000000010",
  18076=>"001011111",
  18077=>"000000000",
  18078=>"111001000",
  18079=>"011111010",
  18080=>"000001000",
  18081=>"101010011",
  18082=>"000000001",
  18083=>"111110111",
  18084=>"000111111",
  18085=>"000100110",
  18086=>"001101001",
  18087=>"001001000",
  18088=>"111111011",
  18089=>"000000000",
  18090=>"100000000",
  18091=>"000111011",
  18092=>"011001000",
  18093=>"000000110",
  18094=>"110110010",
  18095=>"111001010",
  18096=>"000000111",
  18097=>"111000011",
  18098=>"000000000",
  18099=>"000100110",
  18100=>"111110111",
  18101=>"101110111",
  18102=>"111100011",
  18103=>"111111111",
  18104=>"111011011",
  18105=>"010011111",
  18106=>"000000010",
  18107=>"111010000",
  18108=>"000000101",
  18109=>"000000000",
  18110=>"100111001",
  18111=>"000000101",
  18112=>"011010010",
  18113=>"111110111",
  18114=>"000110111",
  18115=>"010101001",
  18116=>"000000101",
  18117=>"001101000",
  18118=>"000000111",
  18119=>"110111000",
  18120=>"101110111",
  18121=>"111000000",
  18122=>"100000000",
  18123=>"111111000",
  18124=>"000000001",
  18125=>"110111011",
  18126=>"010010000",
  18127=>"110111101",
  18128=>"011000000",
  18129=>"011011000",
  18130=>"111110011",
  18131=>"110101111",
  18132=>"110000000",
  18133=>"100000000",
  18134=>"111111111",
  18135=>"111111001",
  18136=>"010110101",
  18137=>"000000111",
  18138=>"001110000",
  18139=>"001001000",
  18140=>"100000111",
  18141=>"000000100",
  18142=>"011100111",
  18143=>"111001011",
  18144=>"010000000",
  18145=>"101000000",
  18146=>"110111000",
  18147=>"101101110",
  18148=>"000110000",
  18149=>"110101101",
  18150=>"000000000",
  18151=>"011111101",
  18152=>"000000001",
  18153=>"111010000",
  18154=>"001001011",
  18155=>"111101110",
  18156=>"000000011",
  18157=>"101101001",
  18158=>"000000000",
  18159=>"000100001",
  18160=>"111111101",
  18161=>"010111010",
  18162=>"101101111",
  18163=>"111101111",
  18164=>"111001011",
  18165=>"111111101",
  18166=>"000000000",
  18167=>"101000111",
  18168=>"111010010",
  18169=>"000000010",
  18170=>"111110010",
  18171=>"111111111",
  18172=>"011001111",
  18173=>"011010111",
  18174=>"001001001",
  18175=>"000010111",
  18176=>"011011001",
  18177=>"000101111",
  18178=>"001100100",
  18179=>"000000101",
  18180=>"110111111",
  18181=>"010010000",
  18182=>"101000001",
  18183=>"000000111",
  18184=>"011111010",
  18185=>"111111011",
  18186=>"100100000",
  18187=>"010010101",
  18188=>"100000111",
  18189=>"010011111",
  18190=>"010100001",
  18191=>"001000100",
  18192=>"000000000",
  18193=>"100100100",
  18194=>"000111001",
  18195=>"010000000",
  18196=>"100000011",
  18197=>"000010000",
  18198=>"000101100",
  18199=>"111010101",
  18200=>"111100111",
  18201=>"111111110",
  18202=>"011011001",
  18203=>"100111010",
  18204=>"000101111",
  18205=>"000100100",
  18206=>"111111000",
  18207=>"100000000",
  18208=>"011000111",
  18209=>"000011011",
  18210=>"100100000",
  18211=>"000010000",
  18212=>"111011011",
  18213=>"011111111",
  18214=>"010000010",
  18215=>"100101101",
  18216=>"011011011",
  18217=>"100111001",
  18218=>"001011000",
  18219=>"000111111",
  18220=>"000100100",
  18221=>"010100100",
  18222=>"010111111",
  18223=>"000110110",
  18224=>"000100100",
  18225=>"001111011",
  18226=>"000011011",
  18227=>"101101100",
  18228=>"101110010",
  18229=>"100000010",
  18230=>"011010111",
  18231=>"011011111",
  18232=>"011111001",
  18233=>"100100000",
  18234=>"111000011",
  18235=>"100010100",
  18236=>"110011111",
  18237=>"110111111",
  18238=>"000000100",
  18239=>"100111101",
  18240=>"100100000",
  18241=>"010100111",
  18242=>"001011111",
  18243=>"000001000",
  18244=>"001001111",
  18245=>"100101111",
  18246=>"000000111",
  18247=>"111011000",
  18248=>"000110111",
  18249=>"000000100",
  18250=>"101100000",
  18251=>"111001010",
  18252=>"011111111",
  18253=>"011111110",
  18254=>"111111111",
  18255=>"101100100",
  18256=>"101100100",
  18257=>"011111111",
  18258=>"010100101",
  18259=>"011101100",
  18260=>"100100110",
  18261=>"101001011",
  18262=>"001001001",
  18263=>"000000000",
  18264=>"111110101",
  18265=>"001100110",
  18266=>"101111011",
  18267=>"110110110",
  18268=>"000000000",
  18269=>"000000001",
  18270=>"001011011",
  18271=>"010000000",
  18272=>"000010000",
  18273=>"000000000",
  18274=>"001000000",
  18275=>"111111001",
  18276=>"110010110",
  18277=>"000100100",
  18278=>"000000000",
  18279=>"011011011",
  18280=>"111011111",
  18281=>"011011000",
  18282=>"000011001",
  18283=>"010010000",
  18284=>"010110111",
  18285=>"100000000",
  18286=>"111110111",
  18287=>"101100111",
  18288=>"111111011",
  18289=>"000000000",
  18290=>"110010001",
  18291=>"100100000",
  18292=>"111011010",
  18293=>"100000000",
  18294=>"111111011",
  18295=>"000100011",
  18296=>"111100101",
  18297=>"100000000",
  18298=>"101000010",
  18299=>"101111101",
  18300=>"110110111",
  18301=>"010010100",
  18302=>"100101101",
  18303=>"010010010",
  18304=>"000000000",
  18305=>"111100000",
  18306=>"011011010",
  18307=>"000000111",
  18308=>"011101000",
  18309=>"000000001",
  18310=>"010111111",
  18311=>"000100110",
  18312=>"100000001",
  18313=>"000000110",
  18314=>"111100100",
  18315=>"111010000",
  18316=>"111111011",
  18317=>"111001101",
  18318=>"100011111",
  18319=>"101000000",
  18320=>"111011011",
  18321=>"010111111",
  18322=>"000000000",
  18323=>"111101100",
  18324=>"101111011",
  18325=>"011011000",
  18326=>"111011010",
  18327=>"001001111",
  18328=>"111011111",
  18329=>"101101011",
  18330=>"010010000",
  18331=>"000010000",
  18332=>"011011011",
  18333=>"000011010",
  18334=>"011001010",
  18335=>"100100100",
  18336=>"101111111",
  18337=>"100100001",
  18338=>"000000000",
  18339=>"101000001",
  18340=>"111111111",
  18341=>"001011001",
  18342=>"111111000",
  18343=>"010111111",
  18344=>"100111111",
  18345=>"000111101",
  18346=>"010010010",
  18347=>"000100000",
  18348=>"111111111",
  18349=>"111000100",
  18350=>"110010001",
  18351=>"000000011",
  18352=>"001111110",
  18353=>"001001011",
  18354=>"111000011",
  18355=>"000100010",
  18356=>"100100000",
  18357=>"000000110",
  18358=>"110100100",
  18359=>"010000010",
  18360=>"011111111",
  18361=>"101011011",
  18362=>"011000111",
  18363=>"011000000",
  18364=>"111110111",
  18365=>"111111011",
  18366=>"111011001",
  18367=>"011011110",
  18368=>"100000100",
  18369=>"000000000",
  18370=>"111000010",
  18371=>"100111110",
  18372=>"101000000",
  18373=>"111011110",
  18374=>"101111111",
  18375=>"010111011",
  18376=>"010010000",
  18377=>"100101000",
  18378=>"000000101",
  18379=>"011110111",
  18380=>"011011011",
  18381=>"001011111",
  18382=>"010000010",
  18383=>"111111011",
  18384=>"010000000",
  18385=>"110110110",
  18386=>"000110111",
  18387=>"100100000",
  18388=>"000000111",
  18389=>"000010111",
  18390=>"000000000",
  18391=>"000000001",
  18392=>"100000100",
  18393=>"010000000",
  18394=>"101101101",
  18395=>"101100100",
  18396=>"100110110",
  18397=>"111111111",
  18398=>"100101101",
  18399=>"010000000",
  18400=>"111100110",
  18401=>"101000100",
  18402=>"101001111",
  18403=>"000000101",
  18404=>"000000000",
  18405=>"011111111",
  18406=>"010011010",
  18407=>"000100110",
  18408=>"011111011",
  18409=>"010000111",
  18410=>"100000000",
  18411=>"000000000",
  18412=>"000000000",
  18413=>"000000011",
  18414=>"111111000",
  18415=>"000111111",
  18416=>"010011000",
  18417=>"111011000",
  18418=>"010000100",
  18419=>"001000001",
  18420=>"110000110",
  18421=>"000100000",
  18422=>"000000100",
  18423=>"010111111",
  18424=>"000000010",
  18425=>"100101000",
  18426=>"100100100",
  18427=>"111110101",
  18428=>"010011010",
  18429=>"111011111",
  18430=>"110111010",
  18431=>"000100100",
  18432=>"011011110",
  18433=>"110111110",
  18434=>"000000010",
  18435=>"000110110",
  18436=>"000000100",
  18437=>"000111111",
  18438=>"111001101",
  18439=>"000000111",
  18440=>"000000000",
  18441=>"000000000",
  18442=>"111111011",
  18443=>"111111111",
  18444=>"000110100",
  18445=>"101000101",
  18446=>"101011001",
  18447=>"111010001",
  18448=>"110000000",
  18449=>"111110111",
  18450=>"111010000",
  18451=>"110111111",
  18452=>"111011010",
  18453=>"111110110",
  18454=>"110110110",
  18455=>"111000000",
  18456=>"000000000",
  18457=>"111101111",
  18458=>"111111111",
  18459=>"111110110",
  18460=>"111111111",
  18461=>"101100111",
  18462=>"010000001",
  18463=>"000000001",
  18464=>"111110111",
  18465=>"111111111",
  18466=>"001000000",
  18467=>"000101000",
  18468=>"110111011",
  18469=>"111110101",
  18470=>"010000010",
  18471=>"000011000",
  18472=>"010010110",
  18473=>"000110110",
  18474=>"111111100",
  18475=>"111111010",
  18476=>"111011111",
  18477=>"000110110",
  18478=>"111111111",
  18479=>"000001000",
  18480=>"000000000",
  18481=>"110110110",
  18482=>"011100000",
  18483=>"111111001",
  18484=>"111001101",
  18485=>"111111101",
  18486=>"111111110",
  18487=>"000000000",
  18488=>"110111110",
  18489=>"110111010",
  18490=>"000000000",
  18491=>"010011111",
  18492=>"101010010",
  18493=>"111011011",
  18494=>"000101101",
  18495=>"000000000",
  18496=>"010110110",
  18497=>"111110110",
  18498=>"010000000",
  18499=>"000010110",
  18500=>"100000001",
  18501=>"001001000",
  18502=>"111001111",
  18503=>"011001111",
  18504=>"111111010",
  18505=>"111110101",
  18506=>"000110010",
  18507=>"001000000",
  18508=>"000111101",
  18509=>"111011100",
  18510=>"000111100",
  18511=>"000111110",
  18512=>"111110111",
  18513=>"000010010",
  18514=>"000000000",
  18515=>"001000100",
  18516=>"010000010",
  18517=>"110010110",
  18518=>"111000000",
  18519=>"101111111",
  18520=>"100110110",
  18521=>"110100001",
  18522=>"111111111",
  18523=>"111000011",
  18524=>"000000000",
  18525=>"001001001",
  18526=>"010010000",
  18527=>"110110111",
  18528=>"000000101",
  18529=>"101111111",
  18530=>"000110110",
  18531=>"110000000",
  18532=>"101111101",
  18533=>"000000000",
  18534=>"111111101",
  18535=>"000000000",
  18536=>"000000000",
  18537=>"111100100",
  18538=>"010011101",
  18539=>"111110110",
  18540=>"000000000",
  18541=>"111111010",
  18542=>"100000000",
  18543=>"111111101",
  18544=>"101101101",
  18545=>"111110100",
  18546=>"110111111",
  18547=>"001101000",
  18548=>"100000011",
  18549=>"110000001",
  18550=>"111111111",
  18551=>"000000110",
  18552=>"000111011",
  18553=>"111111101",
  18554=>"000000011",
  18555=>"000000011",
  18556=>"100110100",
  18557=>"000000001",
  18558=>"000000001",
  18559=>"101000111",
  18560=>"111111000",
  18561=>"111111000",
  18562=>"000000000",
  18563=>"010111111",
  18564=>"000000000",
  18565=>"010001111",
  18566=>"110011011",
  18567=>"101110110",
  18568=>"011001111",
  18569=>"111100001",
  18570=>"000000000",
  18571=>"001000000",
  18572=>"000000100",
  18573=>"011101101",
  18574=>"000000011",
  18575=>"001001000",
  18576=>"011011001",
  18577=>"110110101",
  18578=>"111011111",
  18579=>"111101000",
  18580=>"111101101",
  18581=>"111111111",
  18582=>"110110000",
  18583=>"000001111",
  18584=>"011111101",
  18585=>"010101111",
  18586=>"111011111",
  18587=>"000000010",
  18588=>"101001001",
  18589=>"000000001",
  18590=>"100110111",
  18591=>"111110110",
  18592=>"011110000",
  18593=>"110111111",
  18594=>"110100010",
  18595=>"110111011",
  18596=>"111000001",
  18597=>"110011110",
  18598=>"011010000",
  18599=>"111111111",
  18600=>"111111110",
  18601=>"000000010",
  18602=>"000000110",
  18603=>"111111000",
  18604=>"000101011",
  18605=>"111011111",
  18606=>"111111111",
  18607=>"000111111",
  18608=>"000000100",
  18609=>"111111110",
  18610=>"000101001",
  18611=>"001001000",
  18612=>"111100001",
  18613=>"000000000",
  18614=>"110000111",
  18615=>"111111111",
  18616=>"011000111",
  18617=>"100100111",
  18618=>"010010111",
  18619=>"100110111",
  18620=>"101101010",
  18621=>"111001001",
  18622=>"000000000",
  18623=>"110000111",
  18624=>"100010000",
  18625=>"011000001",
  18626=>"111111110",
  18627=>"000010110",
  18628=>"000000000",
  18629=>"110100010",
  18630=>"100000000",
  18631=>"011111101",
  18632=>"010011011",
  18633=>"110110010",
  18634=>"001111111",
  18635=>"000010110",
  18636=>"110110111",
  18637=>"001011001",
  18638=>"110110100",
  18639=>"000000000",
  18640=>"111111111",
  18641=>"110001001",
  18642=>"101111100",
  18643=>"111010000",
  18644=>"000000000",
  18645=>"110110000",
  18646=>"011110101",
  18647=>"010000000",
  18648=>"000000000",
  18649=>"111101001",
  18650=>"111011111",
  18651=>"101011000",
  18652=>"110110011",
  18653=>"000001001",
  18654=>"110100100",
  18655=>"011000000",
  18656=>"000000000",
  18657=>"000010010",
  18658=>"000000000",
  18659=>"110111000",
  18660=>"000000000",
  18661=>"000110111",
  18662=>"000000101",
  18663=>"101111110",
  18664=>"000101111",
  18665=>"000000000",
  18666=>"111101111",
  18667=>"001111101",
  18668=>"000100000",
  18669=>"000000000",
  18670=>"001110000",
  18671=>"001001111",
  18672=>"111000110",
  18673=>"111110001",
  18674=>"010000000",
  18675=>"011111100",
  18676=>"100100111",
  18677=>"101111000",
  18678=>"000000000",
  18679=>"001000001",
  18680=>"111110000",
  18681=>"000001000",
  18682=>"111111110",
  18683=>"001011111",
  18684=>"010110000",
  18685=>"100100111",
  18686=>"110110111",
  18687=>"110111010",
  18688=>"111100010",
  18689=>"101000000",
  18690=>"000000111",
  18691=>"111111000",
  18692=>"001011000",
  18693=>"001000001",
  18694=>"000111100",
  18695=>"111111111",
  18696=>"111101000",
  18697=>"110110111",
  18698=>"000000101",
  18699=>"111110100",
  18700=>"010110000",
  18701=>"001101000",
  18702=>"011000000",
  18703=>"111001101",
  18704=>"111001111",
  18705=>"010000000",
  18706=>"001110101",
  18707=>"111111000",
  18708=>"010111101",
  18709=>"111000000",
  18710=>"111011001",
  18711=>"001010000",
  18712=>"101111000",
  18713=>"110111000",
  18714=>"111011000",
  18715=>"000010000",
  18716=>"111001000",
  18717=>"110110110",
  18718=>"000110111",
  18719=>"010000000",
  18720=>"111001011",
  18721=>"010000001",
  18722=>"001000000",
  18723=>"111101000",
  18724=>"101000000",
  18725=>"111011000",
  18726=>"111110000",
  18727=>"111101001",
  18728=>"000000101",
  18729=>"111111001",
  18730=>"011011000",
  18731=>"001000101",
  18732=>"111000000",
  18733=>"001111000",
  18734=>"000000011",
  18735=>"011011001",
  18736=>"000110000",
  18737=>"111000000",
  18738=>"111111000",
  18739=>"101111001",
  18740=>"111000111",
  18741=>"000000000",
  18742=>"111010001",
  18743=>"110111000",
  18744=>"000000111",
  18745=>"000011000",
  18746=>"001111000",
  18747=>"100011000",
  18748=>"111011010",
  18749=>"111000111",
  18750=>"011000000",
  18751=>"111000000",
  18752=>"000101000",
  18753=>"000001110",
  18754=>"111111000",
  18755=>"100100111",
  18756=>"000000100",
  18757=>"000010111",
  18758=>"110111010",
  18759=>"000010111",
  18760=>"011111000",
  18761=>"001000000",
  18762=>"111001011",
  18763=>"110000001",
  18764=>"000110111",
  18765=>"101000000",
  18766=>"101000000",
  18767=>"111101000",
  18768=>"101000101",
  18769=>"000111111",
  18770=>"111011000",
  18771=>"110000000",
  18772=>"011110000",
  18773=>"100111011",
  18774=>"111000010",
  18775=>"010111000",
  18776=>"111110000",
  18777=>"111010000",
  18778=>"111001000",
  18779=>"100111001",
  18780=>"111101001",
  18781=>"011000000",
  18782=>"011101111",
  18783=>"011001001",
  18784=>"111000000",
  18785=>"111101001",
  18786=>"000111111",
  18787=>"111000000",
  18788=>"111000000",
  18789=>"101000101",
  18790=>"010011000",
  18791=>"111000000",
  18792=>"111111000",
  18793=>"101000111",
  18794=>"111111111",
  18795=>"111111110",
  18796=>"111101010",
  18797=>"010110000",
  18798=>"000101111",
  18799=>"111111100",
  18800=>"111000000",
  18801=>"101111101",
  18802=>"111010000",
  18803=>"010010000",
  18804=>"111101000",
  18805=>"010011110",
  18806=>"111111000",
  18807=>"010000001",
  18808=>"011111111",
  18809=>"000100100",
  18810=>"101101011",
  18811=>"001000001",
  18812=>"011011000",
  18813=>"000000000",
  18814=>"011000111",
  18815=>"111000010",
  18816=>"010011001",
  18817=>"000000100",
  18818=>"010001000",
  18819=>"000111111",
  18820=>"010111100",
  18821=>"111010010",
  18822=>"100100000",
  18823=>"001100000",
  18824=>"110000000",
  18825=>"101000111",
  18826=>"111011000",
  18827=>"000111111",
  18828=>"000000110",
  18829=>"100000111",
  18830=>"001111111",
  18831=>"000000011",
  18832=>"100000000",
  18833=>"111101000",
  18834=>"110111110",
  18835=>"001101001",
  18836=>"111101000",
  18837=>"000111101",
  18838=>"011010100",
  18839=>"111000000",
  18840=>"101111000",
  18841=>"000110110",
  18842=>"100111100",
  18843=>"111111000",
  18844=>"000111111",
  18845=>"101100000",
  18846=>"111110011",
  18847=>"000010000",
  18848=>"000111000",
  18849=>"100111110",
  18850=>"000000000",
  18851=>"001101000",
  18852=>"111111000",
  18853=>"001001000",
  18854=>"110001111",
  18855=>"111000000",
  18856=>"111111101",
  18857=>"110001000",
  18858=>"000001001",
  18859=>"111000101",
  18860=>"000111111",
  18861=>"001010000",
  18862=>"110001000",
  18863=>"001000001",
  18864=>"011000111",
  18865=>"111001000",
  18866=>"000110111",
  18867=>"100000000",
  18868=>"111000000",
  18869=>"101101000",
  18870=>"011011100",
  18871=>"111111000",
  18872=>"111111010",
  18873=>"101001001",
  18874=>"000101111",
  18875=>"000001110",
  18876=>"111110101",
  18877=>"000110111",
  18878=>"001000000",
  18879=>"000000000",
  18880=>"001101000",
  18881=>"111011001",
  18882=>"010010000",
  18883=>"111100000",
  18884=>"000000000",
  18885=>"000000111",
  18886=>"111111001",
  18887=>"111111111",
  18888=>"000111111",
  18889=>"010110101",
  18890=>"000001000",
  18891=>"000110010",
  18892=>"011010000",
  18893=>"110111000",
  18894=>"110000110",
  18895=>"000111000",
  18896=>"110111000",
  18897=>"110000000",
  18898=>"000111100",
  18899=>"000111000",
  18900=>"111010111",
  18901=>"101000000",
  18902=>"101111000",
  18903=>"111111000",
  18904=>"000000000",
  18905=>"110111001",
  18906=>"000000000",
  18907=>"000101111",
  18908=>"101111100",
  18909=>"011111011",
  18910=>"101110110",
  18911=>"110111111",
  18912=>"000001000",
  18913=>"000000111",
  18914=>"100000000",
  18915=>"111001000",
  18916=>"111000000",
  18917=>"110100000",
  18918=>"111111000",
  18919=>"011010000",
  18920=>"111111000",
  18921=>"111111000",
  18922=>"010000000",
  18923=>"001000011",
  18924=>"110000000",
  18925=>"111111110",
  18926=>"000000111",
  18927=>"001011000",
  18928=>"000000000",
  18929=>"000000011",
  18930=>"111111010",
  18931=>"111000000",
  18932=>"111001001",
  18933=>"101000111",
  18934=>"111111111",
  18935=>"010000100",
  18936=>"000111101",
  18937=>"010001000",
  18938=>"000111111",
  18939=>"110000000",
  18940=>"101000100",
  18941=>"111000000",
  18942=>"011001001",
  18943=>"110110000",
  18944=>"101101100",
  18945=>"011011000",
  18946=>"100000111",
  18947=>"101000000",
  18948=>"111000000",
  18949=>"111111010",
  18950=>"111110111",
  18951=>"011010000",
  18952=>"000011000",
  18953=>"000000110",
  18954=>"001000001",
  18955=>"011111000",
  18956=>"001101011",
  18957=>"000000000",
  18958=>"111101000",
  18959=>"001000010",
  18960=>"111000000",
  18961=>"000011011",
  18962=>"100101111",
  18963=>"010000000",
  18964=>"100111111",
  18965=>"000000000",
  18966=>"111010100",
  18967=>"010111010",
  18968=>"000100111",
  18969=>"110101011",
  18970=>"100100000",
  18971=>"101100111",
  18972=>"000000000",
  18973=>"101110100",
  18974=>"111100000",
  18975=>"010111000",
  18976=>"111000000",
  18977=>"000000001",
  18978=>"101111111",
  18979=>"110111111",
  18980=>"010110000",
  18981=>"111110000",
  18982=>"010000000",
  18983=>"000110110",
  18984=>"100101111",
  18985=>"010010000",
  18986=>"101101000",
  18987=>"000000111",
  18988=>"010011001",
  18989=>"100101111",
  18990=>"010010110",
  18991=>"001111110",
  18992=>"111010000",
  18993=>"011001000",
  18994=>"000010111",
  18995=>"000100111",
  18996=>"101100111",
  18997=>"111111111",
  18998=>"011001001",
  18999=>"100000000",
  19000=>"000000111",
  19001=>"000100011",
  19002=>"100111010",
  19003=>"000011010",
  19004=>"111011001",
  19005=>"111000111",
  19006=>"000000101",
  19007=>"001001000",
  19008=>"000111111",
  19009=>"111010100",
  19010=>"111010111",
  19011=>"101001100",
  19012=>"000010110",
  19013=>"000000100",
  19014=>"101111111",
  19015=>"000010111",
  19016=>"101111111",
  19017=>"000101111",
  19018=>"101011111",
  19019=>"000000000",
  19020=>"110000000",
  19021=>"000001110",
  19022=>"010110100",
  19023=>"101000000",
  19024=>"011001100",
  19025=>"000111011",
  19026=>"110010010",
  19027=>"001100000",
  19028=>"000010001",
  19029=>"111110010",
  19030=>"111001000",
  19031=>"111010111",
  19032=>"101111010",
  19033=>"000011001",
  19034=>"001011000",
  19035=>"011110000",
  19036=>"000000010",
  19037=>"001111000",
  19038=>"111000111",
  19039=>"100100001",
  19040=>"111010000",
  19041=>"111110000",
  19042=>"000000111",
  19043=>"100100001",
  19044=>"100001101",
  19045=>"100011011",
  19046=>"111001000",
  19047=>"101101100",
  19048=>"101000000",
  19049=>"101110111",
  19050=>"101101111",
  19051=>"010010000",
  19052=>"011000000",
  19053=>"000111011",
  19054=>"111000000",
  19055=>"100111111",
  19056=>"001001000",
  19057=>"000010010",
  19058=>"010110100",
  19059=>"011010000",
  19060=>"000101101",
  19061=>"000111110",
  19062=>"010000001",
  19063=>"011000100",
  19064=>"000000101",
  19065=>"101000011",
  19066=>"101101111",
  19067=>"000111010",
  19068=>"111100100",
  19069=>"110100000",
  19070=>"000000111",
  19071=>"010000001",
  19072=>"001101000",
  19073=>"010010001",
  19074=>"010001000",
  19075=>"000011110",
  19076=>"111111110",
  19077=>"111111111",
  19078=>"010111000",
  19079=>"110000001",
  19080=>"110100000",
  19081=>"111111000",
  19082=>"111000000",
  19083=>"011110110",
  19084=>"111100101",
  19085=>"101001101",
  19086=>"111111100",
  19087=>"010100111",
  19088=>"010000110",
  19089=>"100000111",
  19090=>"000000000",
  19091=>"101000000",
  19092=>"111011011",
  19093=>"101000111",
  19094=>"111111111",
  19095=>"011101000",
  19096=>"101100000",
  19097=>"000010000",
  19098=>"000011010",
  19099=>"101000111",
  19100=>"000011000",
  19101=>"101100000",
  19102=>"010000000",
  19103=>"110100111",
  19104=>"100111011",
  19105=>"110010010",
  19106=>"011000000",
  19107=>"111111111",
  19108=>"101111111",
  19109=>"000101000",
  19110=>"110011000",
  19111=>"101101000",
  19112=>"000000011",
  19113=>"111010000",
  19114=>"101101011",
  19115=>"111000001",
  19116=>"001101111",
  19117=>"000000111",
  19118=>"011111001",
  19119=>"000010001",
  19120=>"001000111",
  19121=>"001011100",
  19122=>"010001000",
  19123=>"111100100",
  19124=>"010111000",
  19125=>"111111000",
  19126=>"000111111",
  19127=>"000100000",
  19128=>"111110100",
  19129=>"000011110",
  19130=>"010010000",
  19131=>"110010100",
  19132=>"111110110",
  19133=>"100000000",
  19134=>"010110000",
  19135=>"000110111",
  19136=>"000000111",
  19137=>"100000000",
  19138=>"101111000",
  19139=>"110101100",
  19140=>"000111010",
  19141=>"100100111",
  19142=>"001000000",
  19143=>"111111010",
  19144=>"000100101",
  19145=>"000000000",
  19146=>"000111101",
  19147=>"000100111",
  19148=>"011000100",
  19149=>"011000001",
  19150=>"000000000",
  19151=>"000000111",
  19152=>"110010000",
  19153=>"110110000",
  19154=>"000000101",
  19155=>"110000100",
  19156=>"111001111",
  19157=>"110000000",
  19158=>"111001111",
  19159=>"001001001",
  19160=>"000000000",
  19161=>"000010110",
  19162=>"100110111",
  19163=>"001101111",
  19164=>"001000001",
  19165=>"010011000",
  19166=>"011110101",
  19167=>"100001111",
  19168=>"000000000",
  19169=>"111001111",
  19170=>"000010100",
  19171=>"111011000",
  19172=>"111000111",
  19173=>"000000101",
  19174=>"011111000",
  19175=>"101111000",
  19176=>"101001000",
  19177=>"001000101",
  19178=>"100000100",
  19179=>"010000101",
  19180=>"010000010",
  19181=>"010000011",
  19182=>"000000000",
  19183=>"001000000",
  19184=>"111101000",
  19185=>"000001111",
  19186=>"010011000",
  19187=>"001100000",
  19188=>"100010000",
  19189=>"100000101",
  19190=>"000000001",
  19191=>"001100000",
  19192=>"101011010",
  19193=>"101111000",
  19194=>"011111110",
  19195=>"111100101",
  19196=>"001111000",
  19197=>"111100101",
  19198=>"001000000",
  19199=>"001100101",
  19200=>"010000000",
  19201=>"100000110",
  19202=>"010100001",
  19203=>"100000011",
  19204=>"000111111",
  19205=>"000100100",
  19206=>"100110101",
  19207=>"000010110",
  19208=>"100001000",
  19209=>"010110100",
  19210=>"111111011",
  19211=>"110100100",
  19212=>"110100000",
  19213=>"010111101",
  19214=>"011011111",
  19215=>"011101001",
  19216=>"110110110",
  19217=>"010010100",
  19218=>"010000000",
  19219=>"000010110",
  19220=>"100000100",
  19221=>"110110111",
  19222=>"111000001",
  19223=>"000110110",
  19224=>"100000000",
  19225=>"110100001",
  19226=>"100000110",
  19227=>"110000001",
  19228=>"110110110",
  19229=>"011000100",
  19230=>"100101000",
  19231=>"011010000",
  19232=>"110000100",
  19233=>"001101101",
  19234=>"101100100",
  19235=>"111111100",
  19236=>"011011010",
  19237=>"100000000",
  19238=>"010110100",
  19239=>"001000000",
  19240=>"011111110",
  19241=>"010000000",
  19242=>"001100100",
  19243=>"010000010",
  19244=>"111011111",
  19245=>"100100000",
  19246=>"111011001",
  19247=>"000000100",
  19248=>"111110000",
  19249=>"000000011",
  19250=>"000100000",
  19251=>"101001110",
  19252=>"110000001",
  19253=>"110001010",
  19254=>"111110010",
  19255=>"111001000",
  19256=>"001001001",
  19257=>"100001010",
  19258=>"000001001",
  19259=>"111111011",
  19260=>"000000000",
  19261=>"111011010",
  19262=>"000100000",
  19263=>"111111000",
  19264=>"100100001",
  19265=>"000000000",
  19266=>"001011110",
  19267=>"000010000",
  19268=>"001001001",
  19269=>"000001101",
  19270=>"111110010",
  19271=>"111111111",
  19272=>"011101001",
  19273=>"110100000",
  19274=>"110100100",
  19275=>"010111111",
  19276=>"000001001",
  19277=>"101011111",
  19278=>"111011000",
  19279=>"110001111",
  19280=>"000100000",
  19281=>"011011111",
  19282=>"100110111",
  19283=>"011101000",
  19284=>"100111010",
  19285=>"000000011",
  19286=>"101000001",
  19287=>"110110101",
  19288=>"100110111",
  19289=>"011011011",
  19290=>"101101001",
  19291=>"111111111",
  19292=>"110100000",
  19293=>"001001001",
  19294=>"010110110",
  19295=>"010000000",
  19296=>"001001100",
  19297=>"100110100",
  19298=>"010110111",
  19299=>"001011010",
  19300=>"000000001",
  19301=>"011111100",
  19302=>"011111000",
  19303=>"011010010",
  19304=>"000010101",
  19305=>"101001111",
  19306=>"011111110",
  19307=>"011110110",
  19308=>"111000011",
  19309=>"111111100",
  19310=>"010100100",
  19311=>"001001011",
  19312=>"011011111",
  19313=>"010001101",
  19314=>"111101001",
  19315=>"111000000",
  19316=>"111101110",
  19317=>"000101100",
  19318=>"000001100",
  19319=>"001001011",
  19320=>"110100100",
  19321=>"010001011",
  19322=>"001111110",
  19323=>"110100111",
  19324=>"111101101",
  19325=>"000000000",
  19326=>"011010110",
  19327=>"000100110",
  19328=>"100100101",
  19329=>"001001111",
  19330=>"100000000",
  19331=>"001100000",
  19332=>"000110100",
  19333=>"111100010",
  19334=>"000101111",
  19335=>"111000001",
  19336=>"001011011",
  19337=>"000100000",
  19338=>"111110010",
  19339=>"111000000",
  19340=>"000000110",
  19341=>"000111110",
  19342=>"111101000",
  19343=>"110001001",
  19344=>"111001011",
  19345=>"000010110",
  19346=>"000011010",
  19347=>"001000000",
  19348=>"111010110",
  19349=>"010100100",
  19350=>"000010011",
  19351=>"000001001",
  19352=>"110100110",
  19353=>"011111101",
  19354=>"010000010",
  19355=>"011010000",
  19356=>"000100111",
  19357=>"000000111",
  19358=>"010000010",
  19359=>"001001101",
  19360=>"101111001",
  19361=>"000101100",
  19362=>"010001001",
  19363=>"011110001",
  19364=>"001111111",
  19365=>"010010001",
  19366=>"101001001",
  19367=>"111001110",
  19368=>"100100111",
  19369=>"100001001",
  19370=>"101001001",
  19371=>"000000100",
  19372=>"100000001",
  19373=>"100010010",
  19374=>"010111111",
  19375=>"111110000",
  19376=>"000000100",
  19377=>"011101100",
  19378=>"000001001",
  19379=>"001001001",
  19380=>"010111111",
  19381=>"101010000",
  19382=>"000000101",
  19383=>"011000000",
  19384=>"000100111",
  19385=>"010010100",
  19386=>"010010100",
  19387=>"110011110",
  19388=>"101000000",
  19389=>"001011101",
  19390=>"100000101",
  19391=>"010110000",
  19392=>"100110101",
  19393=>"000110010",
  19394=>"110001011",
  19395=>"011011011",
  19396=>"001000001",
  19397=>"000000001",
  19398=>"000011011",
  19399=>"010000100",
  19400=>"000001001",
  19401=>"001000001",
  19402=>"011111011",
  19403=>"110000101",
  19404=>"010010011",
  19405=>"001001111",
  19406=>"110100000",
  19407=>"110111010",
  19408=>"001011011",
  19409=>"101001010",
  19410=>"111000000",
  19411=>"011111000",
  19412=>"000001001",
  19413=>"100100000",
  19414=>"110100001",
  19415=>"000010000",
  19416=>"100101000",
  19417=>"111000110",
  19418=>"000101011",
  19419=>"110100100",
  19420=>"000000011",
  19421=>"001011111",
  19422=>"001001111",
  19423=>"101000001",
  19424=>"110110100",
  19425=>"111001000",
  19426=>"101111100",
  19427=>"110110001",
  19428=>"000000000",
  19429=>"000011011",
  19430=>"101000111",
  19431=>"110000001",
  19432=>"011101011",
  19433=>"110101100",
  19434=>"110110000",
  19435=>"001011001",
  19436=>"110110000",
  19437=>"101001011",
  19438=>"010000000",
  19439=>"100001011",
  19440=>"000100110",
  19441=>"111011001",
  19442=>"110100101",
  19443=>"010000000",
  19444=>"000000011",
  19445=>"001011010",
  19446=>"001100000",
  19447=>"011011110",
  19448=>"100100101",
  19449=>"100000000",
  19450=>"110110110",
  19451=>"001011011",
  19452=>"111011011",
  19453=>"011010000",
  19454=>"111111110",
  19455=>"011111111",
  19456=>"000000000",
  19457=>"000100111",
  19458=>"010000000",
  19459=>"000101101",
  19460=>"001001001",
  19461=>"000000000",
  19462=>"000000000",
  19463=>"000111110",
  19464=>"010000101",
  19465=>"001000001",
  19466=>"111000000",
  19467=>"111100001",
  19468=>"000111000",
  19469=>"000000000",
  19470=>"001011000",
  19471=>"010000110",
  19472=>"001000000",
  19473=>"111111000",
  19474=>"000000000",
  19475=>"101101100",
  19476=>"111101000",
  19477=>"101001111",
  19478=>"101101001",
  19479=>"110110110",
  19480=>"000000001",
  19481=>"111000001",
  19482=>"101111111",
  19483=>"110010000",
  19484=>"011100001",
  19485=>"010000100",
  19486=>"000000000",
  19487=>"111000101",
  19488=>"111000111",
  19489=>"000000000",
  19490=>"110110001",
  19491=>"111111000",
  19492=>"110101001",
  19493=>"000100100",
  19494=>"111011000",
  19495=>"000100000",
  19496=>"000111111",
  19497=>"111110000",
  19498=>"101011111",
  19499=>"000110111",
  19500=>"000011111",
  19501=>"111111111",
  19502=>"000000000",
  19503=>"001001110",
  19504=>"000000011",
  19505=>"101111001",
  19506=>"111111111",
  19507=>"111000101",
  19508=>"000000000",
  19509=>"001101111",
  19510=>"110001000",
  19511=>"110000000",
  19512=>"000010101",
  19513=>"111100000",
  19514=>"000000111",
  19515=>"111101110",
  19516=>"110110100",
  19517=>"000000010",
  19518=>"110000000",
  19519=>"001001000",
  19520=>"010010001",
  19521=>"110000000",
  19522=>"111111110",
  19523=>"000110000",
  19524=>"111111111",
  19525=>"110111111",
  19526=>"010111001",
  19527=>"110100111",
  19528=>"001011111",
  19529=>"111111000",
  19530=>"001111011",
  19531=>"000111010",
  19532=>"000010000",
  19533=>"101101101",
  19534=>"011111100",
  19535=>"111100001",
  19536=>"110000000",
  19537=>"011001111",
  19538=>"100101000",
  19539=>"000100110",
  19540=>"000110000",
  19541=>"110101001",
  19542=>"001011100",
  19543=>"101000000",
  19544=>"010000111",
  19545=>"001000110",
  19546=>"110010011",
  19547=>"011110000",
  19548=>"111001000",
  19549=>"001000111",
  19550=>"001111011",
  19551=>"000011000",
  19552=>"101111010",
  19553=>"000000111",
  19554=>"111001000",
  19555=>"100000011",
  19556=>"000100000",
  19557=>"111010010",
  19558=>"110111000",
  19559=>"111001000",
  19560=>"001111110",
  19561=>"111001000",
  19562=>"111111111",
  19563=>"111100111",
  19564=>"101001000",
  19565=>"010010110",
  19566=>"100000000",
  19567=>"111010011",
  19568=>"000000000",
  19569=>"010010111",
  19570=>"011100000",
  19571=>"111110000",
  19572=>"111111010",
  19573=>"000000000",
  19574=>"000111111",
  19575=>"001110000",
  19576=>"010010111",
  19577=>"100000000",
  19578=>"000001000",
  19579=>"000101111",
  19580=>"100110110",
  19581=>"100000000",
  19582=>"110000000",
  19583=>"000000000",
  19584=>"110010000",
  19585=>"000000000",
  19586=>"000000111",
  19587=>"101000111",
  19588=>"111111011",
  19589=>"100000000",
  19590=>"000000101",
  19591=>"001100000",
  19592=>"000100010",
  19593=>"000000000",
  19594=>"111101001",
  19595=>"111101100",
  19596=>"000000101",
  19597=>"111001001",
  19598=>"000000010",
  19599=>"010001000",
  19600=>"100111011",
  19601=>"111111000",
  19602=>"100100110",
  19603=>"000001000",
  19604=>"000111001",
  19605=>"000000001",
  19606=>"001001001",
  19607=>"000001011",
  19608=>"111000000",
  19609=>"000111111",
  19610=>"001000111",
  19611=>"111001001",
  19612=>"000001000",
  19613=>"000001001",
  19614=>"010101111",
  19615=>"000010011",
  19616=>"111100101",
  19617=>"111010111",
  19618=>"101001000",
  19619=>"111111111",
  19620=>"010000000",
  19621=>"011001001",
  19622=>"100100101",
  19623=>"001111011",
  19624=>"111110111",
  19625=>"000111111",
  19626=>"000100100",
  19627=>"000110000",
  19628=>"110111111",
  19629=>"111110010",
  19630=>"000001100",
  19631=>"111111000",
  19632=>"010101010",
  19633=>"111000000",
  19634=>"000000100",
  19635=>"110100100",
  19636=>"110110111",
  19637=>"111101101",
  19638=>"110100100",
  19639=>"101111111",
  19640=>"011011001",
  19641=>"000100101",
  19642=>"111000100",
  19643=>"000000000",
  19644=>"111111111",
  19645=>"111110010",
  19646=>"000000000",
  19647=>"111000110",
  19648=>"111000101",
  19649=>"111010000",
  19650=>"000110110",
  19651=>"000100110",
  19652=>"010111111",
  19653=>"011001001",
  19654=>"010010111",
  19655=>"110111111",
  19656=>"011011000",
  19657=>"000010000",
  19658=>"100000000",
  19659=>"111010000",
  19660=>"110110000",
  19661=>"001011111",
  19662=>"000000000",
  19663=>"000000011",
  19664=>"000010110",
  19665=>"000111110",
  19666=>"111000000",
  19667=>"010000010",
  19668=>"000000000",
  19669=>"100000111",
  19670=>"101101001",
  19671=>"000111111",
  19672=>"101101111",
  19673=>"011011011",
  19674=>"100011001",
  19675=>"000000000",
  19676=>"111001100",
  19677=>"000111110",
  19678=>"111101000",
  19679=>"010000000",
  19680=>"111110000",
  19681=>"001101001",
  19682=>"111101111",
  19683=>"000110010",
  19684=>"111010000",
  19685=>"000101101",
  19686=>"011011001",
  19687=>"010000100",
  19688=>"010111111",
  19689=>"111001011",
  19690=>"011000000",
  19691=>"100101101",
  19692=>"000111010",
  19693=>"010100001",
  19694=>"000000000",
  19695=>"111000100",
  19696=>"010000010",
  19697=>"110101000",
  19698=>"101000101",
  19699=>"000001111",
  19700=>"100010001",
  19701=>"101000000",
  19702=>"000000000",
  19703=>"101111111",
  19704=>"000001111",
  19705=>"000111111",
  19706=>"111000100",
  19707=>"111101100",
  19708=>"111010000",
  19709=>"010011001",
  19710=>"101101100",
  19711=>"000111010",
  19712=>"000011011",
  19713=>"000001101",
  19714=>"111101000",
  19715=>"000000001",
  19716=>"011000111",
  19717=>"101100000",
  19718=>"111101000",
  19719=>"000000111",
  19720=>"111111000",
  19721=>"111101000",
  19722=>"001111111",
  19723=>"001011011",
  19724=>"000000010",
  19725=>"010111110",
  19726=>"000101111",
  19727=>"000001000",
  19728=>"111101010",
  19729=>"111101111",
  19730=>"010010100",
  19731=>"000000110",
  19732=>"000010001",
  19733=>"000010010",
  19734=>"110101101",
  19735=>"000111111",
  19736=>"001000000",
  19737=>"000110110",
  19738=>"101000000",
  19739=>"000000000",
  19740=>"000010111",
  19741=>"000000000",
  19742=>"111010000",
  19743=>"000000001",
  19744=>"011010001",
  19745=>"000010011",
  19746=>"000000010",
  19747=>"000100110",
  19748=>"001011110",
  19749=>"001110101",
  19750=>"000010010",
  19751=>"011100001",
  19752=>"010110111",
  19753=>"000010110",
  19754=>"111101001",
  19755=>"000000101",
  19756=>"000100111",
  19757=>"000111111",
  19758=>"001000111",
  19759=>"000000001",
  19760=>"110111001",
  19761=>"000100111",
  19762=>"001000001",
  19763=>"001111110",
  19764=>"000100111",
  19765=>"111010110",
  19766=>"110001111",
  19767=>"001001001",
  19768=>"111111001",
  19769=>"000000001",
  19770=>"111001110",
  19771=>"000101101",
  19772=>"001111111",
  19773=>"111000010",
  19774=>"000000001",
  19775=>"000011001",
  19776=>"001100000",
  19777=>"000010000",
  19778=>"011101001",
  19779=>"111001000",
  19780=>"101001000",
  19781=>"000000001",
  19782=>"101000001",
  19783=>"000000010",
  19784=>"000111111",
  19785=>"000110111",
  19786=>"100000000",
  19787=>"010011111",
  19788=>"010010000",
  19789=>"000110111",
  19790=>"001001111",
  19791=>"001100000",
  19792=>"000010110",
  19793=>"011010000",
  19794=>"100110111",
  19795=>"000001000",
  19796=>"100111010",
  19797=>"101110111",
  19798=>"011011011",
  19799=>"111000000",
  19800=>"001110111",
  19801=>"000100101",
  19802=>"011001000",
  19803=>"010100111",
  19804=>"111001101",
  19805=>"000001011",
  19806=>"111111110",
  19807=>"111001000",
  19808=>"111111000",
  19809=>"111111111",
  19810=>"110000000",
  19811=>"011000000",
  19812=>"001111110",
  19813=>"111111010",
  19814=>"110110010",
  19815=>"111000000",
  19816=>"111100000",
  19817=>"000000101",
  19818=>"000100111",
  19819=>"100011011",
  19820=>"000000111",
  19821=>"011001000",
  19822=>"110110100",
  19823=>"000000000",
  19824=>"100111111",
  19825=>"000000101",
  19826=>"100100101",
  19827=>"111000000",
  19828=>"000000100",
  19829=>"010001001",
  19830=>"000000111",
  19831=>"111111110",
  19832=>"111000000",
  19833=>"001000000",
  19834=>"111111101",
  19835=>"011101101",
  19836=>"001000111",
  19837=>"000100100",
  19838=>"111101000",
  19839=>"111111000",
  19840=>"000111011",
  19841=>"000000100",
  19842=>"000000001",
  19843=>"000000000",
  19844=>"001010000",
  19845=>"000000000",
  19846=>"000100111",
  19847=>"000000011",
  19848=>"001111111",
  19849=>"000100111",
  19850=>"111111000",
  19851=>"000011001",
  19852=>"110100000",
  19853=>"011111101",
  19854=>"111011001",
  19855=>"111001100",
  19856=>"001111111",
  19857=>"011110011",
  19858=>"000001000",
  19859=>"111110101",
  19860=>"000000000",
  19861=>"111101001",
  19862=>"000111111",
  19863=>"000000011",
  19864=>"001101111",
  19865=>"111001010",
  19866=>"111010111",
  19867=>"111101000",
  19868=>"111011111",
  19869=>"010000000",
  19870=>"000111110",
  19871=>"000000011",
  19872=>"000111111",
  19873=>"111111100",
  19874=>"000000001",
  19875=>"111100010",
  19876=>"111111111",
  19877=>"001111111",
  19878=>"110010110",
  19879=>"000001001",
  19880=>"000110011",
  19881=>"000111111",
  19882=>"111000000",
  19883=>"110101101",
  19884=>"010011111",
  19885=>"110111000",
  19886=>"011000100",
  19887=>"111010110",
  19888=>"110000000",
  19889=>"101110111",
  19890=>"111111000",
  19891=>"100000000",
  19892=>"000000011",
  19893=>"101110011",
  19894=>"000000111",
  19895=>"000111111",
  19896=>"000010111",
  19897=>"000000110",
  19898=>"001001011",
  19899=>"111111011",
  19900=>"000010110",
  19901=>"111111110",
  19902=>"111011000",
  19903=>"000110111",
  19904=>"100010110",
  19905=>"000011101",
  19906=>"001111111",
  19907=>"000000100",
  19908=>"011110111",
  19909=>"001010011",
  19910=>"111100101",
  19911=>"111000011",
  19912=>"100000111",
  19913=>"101001100",
  19914=>"000110111",
  19915=>"110110010",
  19916=>"011001101",
  19917=>"000000100",
  19918=>"111111110",
  19919=>"111000000",
  19920=>"111000000",
  19921=>"000100111",
  19922=>"101000110",
  19923=>"000101001",
  19924=>"111000111",
  19925=>"000110110",
  19926=>"000011111",
  19927=>"101001001",
  19928=>"000000110",
  19929=>"011000000",
  19930=>"000000100",
  19931=>"111100000",
  19932=>"001001101",
  19933=>"111010111",
  19934=>"000111111",
  19935=>"101011000",
  19936=>"111101000",
  19937=>"111101100",
  19938=>"111000000",
  19939=>"100001111",
  19940=>"111101000",
  19941=>"101101111",
  19942=>"000001111",
  19943=>"100010110",
  19944=>"111101001",
  19945=>"111000000",
  19946=>"100110111",
  19947=>"111000000",
  19948=>"111010000",
  19949=>"000000000",
  19950=>"010100000",
  19951=>"001000111",
  19952=>"000000000",
  19953=>"000010001",
  19954=>"111111111",
  19955=>"001001110",
  19956=>"000000110",
  19957=>"111111000",
  19958=>"001000010",
  19959=>"111000000",
  19960=>"000000111",
  19961=>"000001101",
  19962=>"000111111",
  19963=>"001010110",
  19964=>"000111111",
  19965=>"101001000",
  19966=>"000100111",
  19967=>"111000111",
  19968=>"011011000",
  19969=>"111100000",
  19970=>"100000000",
  19971=>"000000110",
  19972=>"100111110",
  19973=>"111101101",
  19974=>"100111111",
  19975=>"000110010",
  19976=>"000110110",
  19977=>"000000100",
  19978=>"110000101",
  19979=>"010010111",
  19980=>"000000101",
  19981=>"011101101",
  19982=>"100100010",
  19983=>"001100100",
  19984=>"111111000",
  19985=>"000111001",
  19986=>"100110000",
  19987=>"010111000",
  19988=>"001011011",
  19989=>"101010111",
  19990=>"011111111",
  19991=>"010101011",
  19992=>"000010000",
  19993=>"000110110",
  19994=>"011000100",
  19995=>"000000000",
  19996=>"111111111",
  19997=>"000000110",
  19998=>"101010010",
  19999=>"000000100",
  20000=>"111000011",
  20001=>"111101101",
  20002=>"100000000",
  20003=>"111111000",
  20004=>"000101001",
  20005=>"110110100",
  20006=>"000000001",
  20007=>"000000000",
  20008=>"111110110",
  20009=>"000010010",
  20010=>"000000111",
  20011=>"011001111",
  20012=>"110101001",
  20013=>"001111101",
  20014=>"111100100",
  20015=>"011101111",
  20016=>"110100000",
  20017=>"000001000",
  20018=>"111101101",
  20019=>"000010010",
  20020=>"101100000",
  20021=>"000110101",
  20022=>"100100000",
  20023=>"000110111",
  20024=>"111010010",
  20025=>"000001001",
  20026=>"000101111",
  20027=>"000000001",
  20028=>"000100100",
  20029=>"111111000",
  20030=>"000000000",
  20031=>"100000111",
  20032=>"111000111",
  20033=>"101010010",
  20034=>"111000000",
  20035=>"001001100",
  20036=>"111101010",
  20037=>"000010100",
  20038=>"000000101",
  20039=>"111010111",
  20040=>"010000100",
  20041=>"101001110",
  20042=>"000000111",
  20043=>"000010000",
  20044=>"000000010",
  20045=>"011101100",
  20046=>"000100000",
  20047=>"111111111",
  20048=>"010000000",
  20049=>"110100000",
  20050=>"001000110",
  20051=>"011001000",
  20052=>"100000000",
  20053=>"001100000",
  20054=>"011000000",
  20055=>"011010010",
  20056=>"001101001",
  20057=>"001111101",
  20058=>"101000111",
  20059=>"000011011",
  20060=>"000010010",
  20061=>"000100000",
  20062=>"111000010",
  20063=>"100000000",
  20064=>"000010010",
  20065=>"110111001",
  20066=>"000000000",
  20067=>"000100111",
  20068=>"000000101",
  20069=>"000000001",
  20070=>"010100000",
  20071=>"000010111",
  20072=>"000001111",
  20073=>"101000110",
  20074=>"101111111",
  20075=>"110000000",
  20076=>"000101110",
  20077=>"000101111",
  20078=>"000000111",
  20079=>"110010101",
  20080=>"011111100",
  20081=>"001001011",
  20082=>"001001001",
  20083=>"000111010",
  20084=>"111100000",
  20085=>"111000001",
  20086=>"101000001",
  20087=>"011110110",
  20088=>"001000011",
  20089=>"000011000",
  20090=>"101111000",
  20091=>"101101101",
  20092=>"001001101",
  20093=>"100000000",
  20094=>"010000011",
  20095=>"100101101",
  20096=>"010000010",
  20097=>"111101000",
  20098=>"111111010",
  20099=>"000000011",
  20100=>"001010111",
  20101=>"000100101",
  20102=>"101011000",
  20103=>"000100000",
  20104=>"100111101",
  20105=>"001101100",
  20106=>"000011111",
  20107=>"000110010",
  20108=>"001000100",
  20109=>"010110111",
  20110=>"111100000",
  20111=>"000000000",
  20112=>"100111101",
  20113=>"111001001",
  20114=>"100000101",
  20115=>"111010010",
  20116=>"001101000",
  20117=>"111010010",
  20118=>"111101111",
  20119=>"100000000",
  20120=>"010010111",
  20121=>"001111111",
  20122=>"100100000",
  20123=>"100000000",
  20124=>"010101111",
  20125=>"111100000",
  20126=>"010010100",
  20127=>"000010000",
  20128=>"000011001",
  20129=>"111111010",
  20130=>"101000100",
  20131=>"101111101",
  20132=>"111000000",
  20133=>"010110110",
  20134=>"110110000",
  20135=>"110110000",
  20136=>"100001000",
  20137=>"000000101",
  20138=>"100000000",
  20139=>"110111101",
  20140=>"100000000",
  20141=>"001101111",
  20142=>"110110100",
  20143=>"000000110",
  20144=>"010000010",
  20145=>"000101100",
  20146=>"010101101",
  20147=>"001001000",
  20148=>"000101111",
  20149=>"110111010",
  20150=>"011011011",
  20151=>"000000000",
  20152=>"000001001",
  20153=>"000001101",
  20154=>"011111101",
  20155=>"111001000",
  20156=>"010100010",
  20157=>"101001011",
  20158=>"011101001",
  20159=>"000010110",
  20160=>"001001000",
  20161=>"000000000",
  20162=>"001010000",
  20163=>"000110110",
  20164=>"000001101",
  20165=>"111111100",
  20166=>"000000011",
  20167=>"111001001",
  20168=>"000000111",
  20169=>"000010000",
  20170=>"100110110",
  20171=>"000111010",
  20172=>"000111101",
  20173=>"100100000",
  20174=>"000101000",
  20175=>"010110110",
  20176=>"011111110",
  20177=>"100101011",
  20178=>"000111111",
  20179=>"000010110",
  20180=>"010010000",
  20181=>"000100100",
  20182=>"111100000",
  20183=>"111111011",
  20184=>"000111111",
  20185=>"010111000",
  20186=>"010110110",
  20187=>"000000111",
  20188=>"110101000",
  20189=>"000111111",
  20190=>"111111101",
  20191=>"111111111",
  20192=>"000000010",
  20193=>"111100011",
  20194=>"000000101",
  20195=>"001011000",
  20196=>"001000000",
  20197=>"000111110",
  20198=>"010001111",
  20199=>"011011101",
  20200=>"111001000",
  20201=>"111101111",
  20202=>"111001001",
  20203=>"111000111",
  20204=>"110000000",
  20205=>"010000100",
  20206=>"001000000",
  20207=>"100000000",
  20208=>"110110010",
  20209=>"111111000",
  20210=>"100010010",
  20211=>"100111000",
  20212=>"110110011",
  20213=>"000000111",
  20214=>"100000111",
  20215=>"101000010",
  20216=>"111000000",
  20217=>"000100011",
  20218=>"000001001",
  20219=>"111111101",
  20220=>"111100000",
  20221=>"000000000",
  20222=>"001111001",
  20223=>"001010111",
  20224=>"111000000",
  20225=>"110000101",
  20226=>"100100100",
  20227=>"000111001",
  20228=>"011010110",
  20229=>"000110110",
  20230=>"110111111",
  20231=>"100110100",
  20232=>"010000010",
  20233=>"100100110",
  20234=>"000101001",
  20235=>"011001011",
  20236=>"110110000",
  20237=>"011000011",
  20238=>"001011001",
  20239=>"110111111",
  20240=>"110100110",
  20241=>"110110110",
  20242=>"100100110",
  20243=>"110110001",
  20244=>"110100111",
  20245=>"111111111",
  20246=>"101111110",
  20247=>"110110111",
  20248=>"000010010",
  20249=>"111111111",
  20250=>"000001111",
  20251=>"110110110",
  20252=>"000011110",
  20253=>"001110000",
  20254=>"110110100",
  20255=>"001011001",
  20256=>"001100101",
  20257=>"101100001",
  20258=>"000011011",
  20259=>"111111101",
  20260=>"011101111",
  20261=>"000001011",
  20262=>"001011011",
  20263=>"110100100",
  20264=>"011011101",
  20265=>"001110111",
  20266=>"110100100",
  20267=>"001001001",
  20268=>"000101111",
  20269=>"110100000",
  20270=>"010100100",
  20271=>"000000000",
  20272=>"000110110",
  20273=>"001000000",
  20274=>"100111101",
  20275=>"010110111",
  20276=>"111001100",
  20277=>"000000110",
  20278=>"100100100",
  20279=>"110110010",
  20280=>"100000111",
  20281=>"000110000",
  20282=>"001001111",
  20283=>"011000110",
  20284=>"011101111",
  20285=>"011001011",
  20286=>"000000100",
  20287=>"000000111",
  20288=>"100111111",
  20289=>"000000011",
  20290=>"110110010",
  20291=>"110010100",
  20292=>"011001001",
  20293=>"000000010",
  20294=>"000100110",
  20295=>"000110111",
  20296=>"001000011",
  20297=>"011101101",
  20298=>"110100110",
  20299=>"111101001",
  20300=>"110101111",
  20301=>"001101000",
  20302=>"111111111",
  20303=>"001100011",
  20304=>"001001001",
  20305=>"001100111",
  20306=>"101100111",
  20307=>"100110010",
  20308=>"001001001",
  20309=>"110100110",
  20310=>"011001100",
  20311=>"110110110",
  20312=>"111111111",
  20313=>"000000000",
  20314=>"001001001",
  20315=>"111010000",
  20316=>"110110110",
  20317=>"001001000",
  20318=>"110110110",
  20319=>"000100110",
  20320=>"011011011",
  20321=>"110011111",
  20322=>"000100110",
  20323=>"011011001",
  20324=>"010111110",
  20325=>"111111111",
  20326=>"000001001",
  20327=>"001000001",
  20328=>"111101111",
  20329=>"000100111",
  20330=>"001100110",
  20331=>"011011101",
  20332=>"111001101",
  20333=>"001001101",
  20334=>"110110010",
  20335=>"100110100",
  20336=>"000000000",
  20337=>"110110110",
  20338=>"110110000",
  20339=>"001001001",
  20340=>"100111111",
  20341=>"000000010",
  20342=>"110110110",
  20343=>"000011111",
  20344=>"110110100",
  20345=>"110111110",
  20346=>"111011011",
  20347=>"011101111",
  20348=>"001100110",
  20349=>"000000000",
  20350=>"010100000",
  20351=>"111011011",
  20352=>"000100110",
  20353=>"110110110",
  20354=>"011000111",
  20355=>"001011000",
  20356=>"111111001",
  20357=>"000110110",
  20358=>"000110001",
  20359=>"001001001",
  20360=>"001001101",
  20361=>"001001001",
  20362=>"111110111",
  20363=>"110100100",
  20364=>"110010001",
  20365=>"110111110",
  20366=>"110110110",
  20367=>"010000000",
  20368=>"000000000",
  20369=>"111011010",
  20370=>"101000000",
  20371=>"011000010",
  20372=>"001000000",
  20373=>"110110110",
  20374=>"011111101",
  20375=>"000111101",
  20376=>"011011011",
  20377=>"100100101",
  20378=>"001111111",
  20379=>"100110000",
  20380=>"111110110",
  20381=>"111111111",
  20382=>"110111111",
  20383=>"001100111",
  20384=>"001001101",
  20385=>"110111110",
  20386=>"111110011",
  20387=>"100110001",
  20388=>"011110110",
  20389=>"010001010",
  20390=>"111100000",
  20391=>"010001001",
  20392=>"110110110",
  20393=>"111111111",
  20394=>"001010010",
  20395=>"110000100",
  20396=>"000101000",
  20397=>"001001000",
  20398=>"100100010",
  20399=>"011011011",
  20400=>"110100100",
  20401=>"001000000",
  20402=>"111011000",
  20403=>"000000100",
  20404=>"000001000",
  20405=>"010000001",
  20406=>"000011001",
  20407=>"001010000",
  20408=>"100100100",
  20409=>"011000000",
  20410=>"111101111",
  20411=>"110110000",
  20412=>"011011001",
  20413=>"111011011",
  20414=>"111101001",
  20415=>"000000011",
  20416=>"011001001",
  20417=>"111011010",
  20418=>"110000111",
  20419=>"111011000",
  20420=>"000000011",
  20421=>"000100001",
  20422=>"110100110",
  20423=>"110110100",
  20424=>"001000000",
  20425=>"101111111",
  20426=>"000100001",
  20427=>"000000000",
  20428=>"011111001",
  20429=>"000100000",
  20430=>"001001001",
  20431=>"000110000",
  20432=>"001001111",
  20433=>"001001000",
  20434=>"111111011",
  20435=>"001000001",
  20436=>"101000110",
  20437=>"001011111",
  20438=>"101100110",
  20439=>"110100100",
  20440=>"000000000",
  20441=>"110000101",
  20442=>"010101001",
  20443=>"001011001",
  20444=>"100110100",
  20445=>"001001001",
  20446=>"011001010",
  20447=>"110000000",
  20448=>"111110100",
  20449=>"000011111",
  20450=>"001101011",
  20451=>"001000000",
  20452=>"100000000",
  20453=>"100000011",
  20454=>"011011011",
  20455=>"110110110",
  20456=>"110010111",
  20457=>"110010010",
  20458=>"011001000",
  20459=>"110101100",
  20460=>"100110010",
  20461=>"001001011",
  20462=>"110000010",
  20463=>"110000110",
  20464=>"000000000",
  20465=>"111110010",
  20466=>"111110110",
  20467=>"110111000",
  20468=>"100100110",
  20469=>"001011001",
  20470=>"000000000",
  20471=>"000001110",
  20472=>"110110110",
  20473=>"100000000",
  20474=>"011011111",
  20475=>"110100000",
  20476=>"111001000",
  20477=>"000100010",
  20478=>"010011101",
  20479=>"011111011",
  20480=>"011011001",
  20481=>"000001110",
  20482=>"000100000",
  20483=>"001001111",
  20484=>"010101100",
  20485=>"110110010",
  20486=>"100110111",
  20487=>"110001010",
  20488=>"000000001",
  20489=>"110001100",
  20490=>"010110010",
  20491=>"100100111",
  20492=>"001110111",
  20493=>"000010010",
  20494=>"010001011",
  20495=>"101001101",
  20496=>"011111001",
  20497=>"100111111",
  20498=>"001011110",
  20499=>"000001011",
  20500=>"111111000",
  20501=>"100110110",
  20502=>"011000001",
  20503=>"110100101",
  20504=>"010000001",
  20505=>"100111111",
  20506=>"111111010",
  20507=>"110000000",
  20508=>"100000100",
  20509=>"000000011",
  20510=>"111000000",
  20511=>"001001011",
  20512=>"000110010",
  20513=>"000001011",
  20514=>"110101001",
  20515=>"110011011",
  20516=>"011001011",
  20517=>"001001010",
  20518=>"011011001",
  20519=>"000010011",
  20520=>"010111111",
  20521=>"100000101",
  20522=>"110011000",
  20523=>"111100100",
  20524=>"111111111",
  20525=>"100000111",
  20526=>"111101000",
  20527=>"011001101",
  20528=>"011000010",
  20529=>"001001001",
  20530=>"000111110",
  20531=>"111111100",
  20532=>"100110111",
  20533=>"001000000",
  20534=>"000001011",
  20535=>"111110000",
  20536=>"011101110",
  20537=>"000100000",
  20538=>"100000001",
  20539=>"110000000",
  20540=>"000000011",
  20541=>"010001001",
  20542=>"000010001",
  20543=>"111111110",
  20544=>"111110111",
  20545=>"001111101",
  20546=>"000110011",
  20547=>"000000011",
  20548=>"110000000",
  20549=>"000100101",
  20550=>"000100001",
  20551=>"001011111",
  20552=>"011001001",
  20553=>"011010001",
  20554=>"001001001",
  20555=>"101111111",
  20556=>"100110100",
  20557=>"111011001",
  20558=>"011001001",
  20559=>"000100011",
  20560=>"001010010",
  20561=>"111000100",
  20562=>"111110001",
  20563=>"011000000",
  20564=>"111111101",
  20565=>"011000000",
  20566=>"001001001",
  20567=>"110100100",
  20568=>"110000110",
  20569=>"000001001",
  20570=>"001001001",
  20571=>"101101100",
  20572=>"110101110",
  20573=>"100000101",
  20574=>"110011110",
  20575=>"000111100",
  20576=>"110110110",
  20577=>"000010110",
  20578=>"100110110",
  20579=>"001001011",
  20580=>"000000000",
  20581=>"010001001",
  20582=>"100011011",
  20583=>"000011011",
  20584=>"010001111",
  20585=>"110000000",
  20586=>"111001011",
  20587=>"010111111",
  20588=>"111001111",
  20589=>"100100100",
  20590=>"000110010",
  20591=>"111100000",
  20592=>"001001001",
  20593=>"010111001",
  20594=>"011011000",
  20595=>"001001111",
  20596=>"001000110",
  20597=>"000100100",
  20598=>"000100100",
  20599=>"110111000",
  20600=>"110110000",
  20601=>"110101100",
  20602=>"010011011",
  20603=>"110000000",
  20604=>"110010000",
  20605=>"000000011",
  20606=>"110010110",
  20607=>"000110011",
  20608=>"101110010",
  20609=>"011000010",
  20610=>"110111000",
  20611=>"000000000",
  20612=>"001001000",
  20613=>"110110101",
  20614=>"111001110",
  20615=>"110100100",
  20616=>"011001001",
  20617=>"000001001",
  20618=>"001011111",
  20619=>"100110111",
  20620=>"100101000",
  20621=>"100110100",
  20622=>"000111101",
  20623=>"000000001",
  20624=>"101001001",
  20625=>"001000000",
  20626=>"111111011",
  20627=>"001000000",
  20628=>"100111001",
  20629=>"000010110",
  20630=>"001110010",
  20631=>"101101111",
  20632=>"000001100",
  20633=>"011110111",
  20634=>"111101111",
  20635=>"100111011",
  20636=>"100110111",
  20637=>"100110110",
  20638=>"010001111",
  20639=>"101100101",
  20640=>"001110100",
  20641=>"110100100",
  20642=>"001001111",
  20643=>"011110111",
  20644=>"111001111",
  20645=>"100110010",
  20646=>"000000111",
  20647=>"111011001",
  20648=>"110100000",
  20649=>"100010111",
  20650=>"011111111",
  20651=>"000000000",
  20652=>"010100110",
  20653=>"111101100",
  20654=>"000000010",
  20655=>"100010011",
  20656=>"000100010",
  20657=>"110100101",
  20658=>"001000000",
  20659=>"010000010",
  20660=>"100100000",
  20661=>"000000111",
  20662=>"011110111",
  20663=>"001001101",
  20664=>"111000000",
  20665=>"000100000",
  20666=>"011001100",
  20667=>"111000011",
  20668=>"000101111",
  20669=>"110111111",
  20670=>"111101000",
  20671=>"010111011",
  20672=>"100100110",
  20673=>"111010110",
  20674=>"000110011",
  20675=>"011001000",
  20676=>"100100000",
  20677=>"000110101",
  20678=>"110100000",
  20679=>"110010100",
  20680=>"100110001",
  20681=>"010000000",
  20682=>"011111000",
  20683=>"010011011",
  20684=>"111000001",
  20685=>"100101101",
  20686=>"111100100",
  20687=>"100000111",
  20688=>"110001111",
  20689=>"011111111",
  20690=>"100100110",
  20691=>"000001001",
  20692=>"000110111",
  20693=>"000000000",
  20694=>"001111111",
  20695=>"111011111",
  20696=>"011001011",
  20697=>"000011011",
  20698=>"000101110",
  20699=>"100110110",
  20700=>"011011011",
  20701=>"100001011",
  20702=>"000101111",
  20703=>"100000000",
  20704=>"000011011",
  20705=>"010110110",
  20706=>"110111110",
  20707=>"100100001",
  20708=>"010010010",
  20709=>"001001001",
  20710=>"100001001",
  20711=>"111001001",
  20712=>"110111011",
  20713=>"100110111",
  20714=>"110110110",
  20715=>"110111101",
  20716=>"010110010",
  20717=>"000000011",
  20718=>"000100000",
  20719=>"111110001",
  20720=>"011001111",
  20721=>"101000100",
  20722=>"111101100",
  20723=>"011001011",
  20724=>"000000010",
  20725=>"110110111",
  20726=>"100110100",
  20727=>"010110101",
  20728=>"110100100",
  20729=>"010011010",
  20730=>"100100100",
  20731=>"010000000",
  20732=>"111111011",
  20733=>"011111111",
  20734=>"000001101",
  20735=>"110111001",
  20736=>"011011011",
  20737=>"000110110",
  20738=>"101000000",
  20739=>"010111111",
  20740=>"011000000",
  20741=>"110010000",
  20742=>"100010101",
  20743=>"000101111",
  20744=>"010110100",
  20745=>"100111101",
  20746=>"000001001",
  20747=>"000000010",
  20748=>"111011000",
  20749=>"011000111",
  20750=>"110110110",
  20751=>"000110101",
  20752=>"110110000",
  20753=>"001101111",
  20754=>"101000010",
  20755=>"000010110",
  20756=>"111000010",
  20757=>"111000000",
  20758=>"000101101",
  20759=>"010111011",
  20760=>"000000000",
  20761=>"010000010",
  20762=>"000000010",
  20763=>"000111101",
  20764=>"000100010",
  20765=>"010010000",
  20766=>"000000000",
  20767=>"101000101",
  20768=>"011101111",
  20769=>"110110111",
  20770=>"001000101",
  20771=>"000000000",
  20772=>"001100101",
  20773=>"000000000",
  20774=>"110111111",
  20775=>"111111011",
  20776=>"011010011",
  20777=>"110111111",
  20778=>"110011110",
  20779=>"000100110",
  20780=>"011111011",
  20781=>"000111011",
  20782=>"010111101",
  20783=>"011000000",
  20784=>"110111001",
  20785=>"101110100",
  20786=>"101110000",
  20787=>"110101010",
  20788=>"000001001",
  20789=>"010110110",
  20790=>"000100100",
  20791=>"000010111",
  20792=>"011111000",
  20793=>"111010000",
  20794=>"101101100",
  20795=>"110111111",
  20796=>"100001001",
  20797=>"001101000",
  20798=>"001000000",
  20799=>"000101001",
  20800=>"001101110",
  20801=>"111111011",
  20802=>"100010110",
  20803=>"001001101",
  20804=>"111000000",
  20805=>"011000000",
  20806=>"000100100",
  20807=>"111111010",
  20808=>"010100000",
  20809=>"011111111",
  20810=>"000110100",
  20811=>"000101111",
  20812=>"101000111",
  20813=>"100001001",
  20814=>"101001000",
  20815=>"100110000",
  20816=>"001101111",
  20817=>"011000000",
  20818=>"111111010",
  20819=>"011011000",
  20820=>"111111110",
  20821=>"000101100",
  20822=>"100101100",
  20823=>"000000000",
  20824=>"011101010",
  20825=>"101100101",
  20826=>"001000011",
  20827=>"000000111",
  20828=>"010011001",
  20829=>"000000000",
  20830=>"111111111",
  20831=>"100100100",
  20832=>"111110111",
  20833=>"111111011",
  20834=>"101000011",
  20835=>"000100110",
  20836=>"100000000",
  20837=>"000001000",
  20838=>"010011010",
  20839=>"000000000",
  20840=>"011101101",
  20841=>"111111101",
  20842=>"001101000",
  20843=>"111111100",
  20844=>"111001000",
  20845=>"111000110",
  20846=>"000000010",
  20847=>"110111111",
  20848=>"001001100",
  20849=>"000111101",
  20850=>"000001011",
  20851=>"101000111",
  20852=>"111111111",
  20853=>"111000100",
  20854=>"000110111",
  20855=>"111111111",
  20856=>"110010110",
  20857=>"000001000",
  20858=>"101110010",
  20859=>"111000000",
  20860=>"000011001",
  20861=>"110110000",
  20862=>"110101111",
  20863=>"111000001",
  20864=>"010010000",
  20865=>"010000010",
  20866=>"110010100",
  20867=>"011110001",
  20868=>"011111000",
  20869=>"000010111",
  20870=>"010001000",
  20871=>"001000000",
  20872=>"100101001",
  20873=>"001010010",
  20874=>"001000111",
  20875=>"111011111",
  20876=>"110000000",
  20877=>"010010110",
  20878=>"000110111",
  20879=>"000110000",
  20880=>"101111001",
  20881=>"110000100",
  20882=>"011000001",
  20883=>"010100101",
  20884=>"000100011",
  20885=>"101111111",
  20886=>"000010110",
  20887=>"000000110",
  20888=>"111010000",
  20889=>"111001011",
  20890=>"111101000",
  20891=>"000010000",
  20892=>"011110000",
  20893=>"000111010",
  20894=>"011111000",
  20895=>"000111000",
  20896=>"000100000",
  20897=>"000100111",
  20898=>"101001000",
  20899=>"000000110",
  20900=>"110111010",
  20901=>"100000010",
  20902=>"000000100",
  20903=>"101100000",
  20904=>"010011111",
  20905=>"000000010",
  20906=>"111101000",
  20907=>"000101110",
  20908=>"010111010",
  20909=>"000001101",
  20910=>"000110110",
  20911=>"100000011",
  20912=>"111010010",
  20913=>"101001100",
  20914=>"111000000",
  20915=>"001001001",
  20916=>"001001101",
  20917=>"010010111",
  20918=>"111111010",
  20919=>"000000010",
  20920=>"001100010",
  20921=>"011011110",
  20922=>"000000110",
  20923=>"000111000",
  20924=>"111010111",
  20925=>"111011111",
  20926=>"000011000",
  20927=>"101001100",
  20928=>"000111010",
  20929=>"000111101",
  20930=>"010110111",
  20931=>"000001001",
  20932=>"111010000",
  20933=>"011101110",
  20934=>"010111110",
  20935=>"111110110",
  20936=>"111010111",
  20937=>"000000111",
  20938=>"111111011",
  20939=>"100101101",
  20940=>"000001010",
  20941=>"000100110",
  20942=>"000101111",
  20943=>"110101101",
  20944=>"010010011",
  20945=>"010011011",
  20946=>"100001111",
  20947=>"010010101",
  20948=>"111011111",
  20949=>"000101011",
  20950=>"100001010",
  20951=>"000110000",
  20952=>"000011100",
  20953=>"011000000",
  20954=>"000001000",
  20955=>"111000000",
  20956=>"100101001",
  20957=>"000000111",
  20958=>"010010001",
  20959=>"010010010",
  20960=>"101000000",
  20961=>"111100010",
  20962=>"110001000",
  20963=>"001001010",
  20964=>"000000010",
  20965=>"101100000",
  20966=>"010000011",
  20967=>"000011110",
  20968=>"111101111",
  20969=>"100101101",
  20970=>"000100100",
  20971=>"111011101",
  20972=>"010010000",
  20973=>"000100100",
  20974=>"111010010",
  20975=>"000001001",
  20976=>"000101111",
  20977=>"000111011",
  20978=>"010011011",
  20979=>"001001100",
  20980=>"000110110",
  20981=>"111000111",
  20982=>"000000010",
  20983=>"010000000",
  20984=>"010111011",
  20985=>"111101111",
  20986=>"011111110",
  20987=>"111111110",
  20988=>"000110101",
  20989=>"000000101",
  20990=>"101101000",
  20991=>"000000110",
  20992=>"011001110",
  20993=>"000000000",
  20994=>"111000100",
  20995=>"000100010",
  20996=>"000000000",
  20997=>"001000100",
  20998=>"000111110",
  20999=>"000000111",
  21000=>"101011000",
  21001=>"000011111",
  21002=>"000110001",
  21003=>"000010011",
  21004=>"001101101",
  21005=>"000010111",
  21006=>"000000011",
  21007=>"110000000",
  21008=>"111000100",
  21009=>"111000000",
  21010=>"111000000",
  21011=>"000000010",
  21012=>"110100000",
  21013=>"111100000",
  21014=>"101101111",
  21015=>"100000111",
  21016=>"000000000",
  21017=>"011111101",
  21018=>"001011111",
  21019=>"011000100",
  21020=>"010000001",
  21021=>"110011000",
  21022=>"010010000",
  21023=>"000000011",
  21024=>"001110111",
  21025=>"110000000",
  21026=>"010111000",
  21027=>"000111000",
  21028=>"100110110",
  21029=>"001000000",
  21030=>"000110111",
  21031=>"000100010",
  21032=>"011101101",
  21033=>"100000001",
  21034=>"000000011",
  21035=>"000100000",
  21036=>"111111111",
  21037=>"010111100",
  21038=>"111111111",
  21039=>"111101101",
  21040=>"000010000",
  21041=>"010001011",
  21042=>"000001001",
  21043=>"000100000",
  21044=>"000011010",
  21045=>"100000110",
  21046=>"011011110",
  21047=>"101000000",
  21048=>"000000000",
  21049=>"110110111",
  21050=>"000000101",
  21051=>"000000010",
  21052=>"000110111",
  21053=>"111111010",
  21054=>"000010000",
  21055=>"011001001",
  21056=>"100110111",
  21057=>"101010000",
  21058=>"000111000",
  21059=>"000101110",
  21060=>"111111001",
  21061=>"000000000",
  21062=>"101111111",
  21063=>"111111000",
  21064=>"000010110",
  21065=>"111100000",
  21066=>"000000000",
  21067=>"110010111",
  21068=>"111101000",
  21069=>"100001001",
  21070=>"000100110",
  21071=>"111111001",
  21072=>"101001000",
  21073=>"111000000",
  21074=>"110110111",
  21075=>"001001000",
  21076=>"010110000",
  21077=>"111011001",
  21078=>"010000011",
  21079=>"001000100",
  21080=>"000110110",
  21081=>"000001001",
  21082=>"111000000",
  21083=>"000111110",
  21084=>"111000000",
  21085=>"000001001",
  21086=>"111111000",
  21087=>"110110110",
  21088=>"000000111",
  21089=>"111110101",
  21090=>"111000000",
  21091=>"110111110",
  21092=>"000100110",
  21093=>"010000000",
  21094=>"010111110",
  21095=>"101110010",
  21096=>"010000001",
  21097=>"011000111",
  21098=>"111111011",
  21099=>"000000000",
  21100=>"111111000",
  21101=>"111100111",
  21102=>"011010000",
  21103=>"000000000",
  21104=>"000001111",
  21105=>"000000010",
  21106=>"000100111",
  21107=>"000000010",
  21108=>"100101000",
  21109=>"000000000",
  21110=>"111010001",
  21111=>"111001100",
  21112=>"000111000",
  21113=>"000010011",
  21114=>"100111110",
  21115=>"000000000",
  21116=>"110110101",
  21117=>"100100000",
  21118=>"000100000",
  21119=>"111101000",
  21120=>"000000000",
  21121=>"000000110",
  21122=>"010010000",
  21123=>"000000000",
  21124=>"110111111",
  21125=>"011011000",
  21126=>"110110100",
  21127=>"011110110",
  21128=>"110110110",
  21129=>"100000010",
  21130=>"000100111",
  21131=>"011000000",
  21132=>"111000000",
  21133=>"000000010",
  21134=>"000101100",
  21135=>"001011100",
  21136=>"000111010",
  21137=>"000000111",
  21138=>"000000001",
  21139=>"111001000",
  21140=>"100110111",
  21141=>"000010000",
  21142=>"111110010",
  21143=>"000001100",
  21144=>"010110000",
  21145=>"111101001",
  21146=>"110000110",
  21147=>"111101010",
  21148=>"111001110",
  21149=>"000100100",
  21150=>"111000000",
  21151=>"100000000",
  21152=>"001010010",
  21153=>"010010000",
  21154=>"101111111",
  21155=>"100000000",
  21156=>"111010100",
  21157=>"000111111",
  21158=>"100111110",
  21159=>"011111000",
  21160=>"001110111",
  21161=>"100100000",
  21162=>"111000000",
  21163=>"111100000",
  21164=>"101001000",
  21165=>"101100100",
  21166=>"100000000",
  21167=>"111110111",
  21168=>"000000000",
  21169=>"001111101",
  21170=>"001111111",
  21171=>"000000100",
  21172=>"000010110",
  21173=>"011111000",
  21174=>"011100100",
  21175=>"000100101",
  21176=>"100100011",
  21177=>"101111011",
  21178=>"000011000",
  21179=>"111000010",
  21180=>"110000000",
  21181=>"111110000",
  21182=>"100100100",
  21183=>"000000011",
  21184=>"101100001",
  21185=>"010010000",
  21186=>"000000101",
  21187=>"000111111",
  21188=>"011010000",
  21189=>"111001011",
  21190=>"000110111",
  21191=>"110111111",
  21192=>"101100010",
  21193=>"001100000",
  21194=>"011000000",
  21195=>"111000000",
  21196=>"011011001",
  21197=>"111101000",
  21198=>"100010000",
  21199=>"110000101",
  21200=>"000010111",
  21201=>"010110111",
  21202=>"111010100",
  21203=>"111000000",
  21204=>"000111000",
  21205=>"100100000",
  21206=>"000011010",
  21207=>"111111111",
  21208=>"011000001",
  21209=>"100000110",
  21210=>"101010011",
  21211=>"111000000",
  21212=>"110100111",
  21213=>"000000000",
  21214=>"010111111",
  21215=>"011000000",
  21216=>"111010000",
  21217=>"101100110",
  21218=>"010111110",
  21219=>"011001111",
  21220=>"101000000",
  21221=>"001111111",
  21222=>"000010111",
  21223=>"010011111",
  21224=>"000010111",
  21225=>"101110111",
  21226=>"000111100",
  21227=>"111101100",
  21228=>"000000000",
  21229=>"000010111",
  21230=>"011000010",
  21231=>"000000000",
  21232=>"011011010",
  21233=>"011100110",
  21234=>"001000010",
  21235=>"000110101",
  21236=>"100100111",
  21237=>"111111111",
  21238=>"000000010",
  21239=>"000010001",
  21240=>"111011000",
  21241=>"001010011",
  21242=>"000001101",
  21243=>"100111111",
  21244=>"111000000",
  21245=>"111100000",
  21246=>"111001000",
  21247=>"111011001",
  21248=>"011011000",
  21249=>"111000001",
  21250=>"101000001",
  21251=>"110000111",
  21252=>"100111111",
  21253=>"000000110",
  21254=>"000111110",
  21255=>"001101101",
  21256=>"000001000",
  21257=>"111000100",
  21258=>"000010000",
  21259=>"111101101",
  21260=>"101000000",
  21261=>"000000001",
  21262=>"000000011",
  21263=>"000001101",
  21264=>"011010111",
  21265=>"111100000",
  21266=>"010110111",
  21267=>"000001010",
  21268=>"110111111",
  21269=>"111111111",
  21270=>"110000101",
  21271=>"000111111",
  21272=>"000001100",
  21273=>"111111111",
  21274=>"000101000",
  21275=>"101000001",
  21276=>"110110101",
  21277=>"000000111",
  21278=>"000111011",
  21279=>"000000111",
  21280=>"111000000",
  21281=>"110100110",
  21282=>"000000000",
  21283=>"111111000",
  21284=>"010111100",
  21285=>"100111111",
  21286=>"101000000",
  21287=>"010010000",
  21288=>"110100101",
  21289=>"000001111",
  21290=>"001111000",
  21291=>"101000000",
  21292=>"111111111",
  21293=>"101011000",
  21294=>"111001001",
  21295=>"010000100",
  21296=>"010101000",
  21297=>"100100110",
  21298=>"111100110",
  21299=>"111101111",
  21300=>"000010111",
  21301=>"111000000",
  21302=>"111111011",
  21303=>"101000011",
  21304=>"001000000",
  21305=>"100100010",
  21306=>"000001111",
  21307=>"111101101",
  21308=>"010011011",
  21309=>"111111001",
  21310=>"100000000",
  21311=>"001100110",
  21312=>"111100101",
  21313=>"000111111",
  21314=>"111111000",
  21315=>"000110011",
  21316=>"111101111",
  21317=>"111000010",
  21318=>"010010111",
  21319=>"010110110",
  21320=>"111101100",
  21321=>"001000001",
  21322=>"110001001",
  21323=>"000011111",
  21324=>"000000000",
  21325=>"101101101",
  21326=>"010111011",
  21327=>"000000000",
  21328=>"000000111",
  21329=>"111000000",
  21330=>"011000111",
  21331=>"000011100",
  21332=>"101000000",
  21333=>"111101100",
  21334=>"100111111",
  21335=>"101111111",
  21336=>"111000001",
  21337=>"100100111",
  21338=>"100101101",
  21339=>"010011111",
  21340=>"111000000",
  21341=>"001001001",
  21342=>"111101111",
  21343=>"101110110",
  21344=>"000111110",
  21345=>"000011011",
  21346=>"101000101",
  21347=>"100101001",
  21348=>"100110000",
  21349=>"011000001",
  21350=>"111110010",
  21351=>"000011100",
  21352=>"000000010",
  21353=>"010100001",
  21354=>"111000010",
  21355=>"010000001",
  21356=>"101000001",
  21357=>"010111111",
  21358=>"000010111",
  21359=>"001000001",
  21360=>"100100111",
  21361=>"111111001",
  21362=>"111011110",
  21363=>"000000000",
  21364=>"111101101",
  21365=>"101001111",
  21366=>"000011010",
  21367=>"001000000",
  21368=>"111000000",
  21369=>"110111111",
  21370=>"000000111",
  21371=>"001001111",
  21372=>"100110010",
  21373=>"000100000",
  21374=>"000000000",
  21375=>"001000001",
  21376=>"111010000",
  21377=>"100101000",
  21378=>"010000000",
  21379=>"000000000",
  21380=>"001000000",
  21381=>"000010000",
  21382=>"001011111",
  21383=>"001010001",
  21384=>"011111011",
  21385=>"111111010",
  21386=>"000101000",
  21387=>"110000111",
  21388=>"000000000",
  21389=>"111111111",
  21390=>"011101000",
  21391=>"000000101",
  21392=>"100100100",
  21393=>"101001101",
  21394=>"011010000",
  21395=>"101000111",
  21396=>"111000000",
  21397=>"000010011",
  21398=>"110110000",
  21399=>"110100100",
  21400=>"101110010",
  21401=>"111111110",
  21402=>"111010110",
  21403=>"000000000",
  21404=>"011111011",
  21405=>"111010000",
  21406=>"111010010",
  21407=>"000000000",
  21408=>"010100001",
  21409=>"101000000",
  21410=>"111101000",
  21411=>"110000001",
  21412=>"000000111",
  21413=>"110110010",
  21414=>"111001101",
  21415=>"011101000",
  21416=>"111110111",
  21417=>"111011000",
  21418=>"010000101",
  21419=>"000001101",
  21420=>"010001111",
  21421=>"000000000",
  21422=>"111111111",
  21423=>"110111111",
  21424=>"000000101",
  21425=>"001100110",
  21426=>"000000000",
  21427=>"000000010",
  21428=>"000000101",
  21429=>"000000000",
  21430=>"110000100",
  21431=>"001000010",
  21432=>"011110010",
  21433=>"110010000",
  21434=>"011001101",
  21435=>"000000011",
  21436=>"110101100",
  21437=>"110101111",
  21438=>"100000000",
  21439=>"111000000",
  21440=>"011111010",
  21441=>"000111010",
  21442=>"000010111",
  21443=>"001001001",
  21444=>"011000000",
  21445=>"100010001",
  21446=>"011000000",
  21447=>"111111110",
  21448=>"011010000",
  21449=>"101101111",
  21450=>"111000010",
  21451=>"100110000",
  21452=>"000011111",
  21453=>"000110010",
  21454=>"000111111",
  21455=>"000000000",
  21456=>"000000000",
  21457=>"001011011",
  21458=>"010111111",
  21459=>"000100001",
  21460=>"000010110",
  21461=>"110100101",
  21462=>"110100000",
  21463=>"000000000",
  21464=>"111111000",
  21465=>"000101101",
  21466=>"111011000",
  21467=>"000000100",
  21468=>"001000001",
  21469=>"100111100",
  21470=>"111111111",
  21471=>"010110111",
  21472=>"100000000",
  21473=>"010000000",
  21474=>"000000100",
  21475=>"001111111",
  21476=>"000011111",
  21477=>"010000111",
  21478=>"111101111",
  21479=>"011000101",
  21480=>"101100111",
  21481=>"111000010",
  21482=>"000111011",
  21483=>"111101000",
  21484=>"000000000",
  21485=>"101101000",
  21486=>"000000000",
  21487=>"111000000",
  21488=>"111101101",
  21489=>"000000100",
  21490=>"000000010",
  21491=>"000000111",
  21492=>"111111001",
  21493=>"100111011",
  21494=>"110101100",
  21495=>"000000000",
  21496=>"000111000",
  21497=>"101000010",
  21498=>"010111000",
  21499=>"111111101",
  21500=>"111010001",
  21501=>"000011011",
  21502=>"010000000",
  21503=>"000010000",
  21504=>"100110010",
  21505=>"000101000",
  21506=>"011001000",
  21507=>"101000001",
  21508=>"111110001",
  21509=>"111001001",
  21510=>"101101111",
  21511=>"111111000",
  21512=>"010001001",
  21513=>"110000000",
  21514=>"011111110",
  21515=>"111110110",
  21516=>"000000010",
  21517=>"000010010",
  21518=>"001110110",
  21519=>"000000010",
  21520=>"111110110",
  21521=>"000000110",
  21522=>"000000000",
  21523=>"110100110",
  21524=>"000111111",
  21525=>"111110000",
  21526=>"111110111",
  21527=>"111000101",
  21528=>"111000000",
  21529=>"111000001",
  21530=>"010000010",
  21531=>"000000000",
  21532=>"001000110",
  21533=>"100000010",
  21534=>"000001000",
  21535=>"101101111",
  21536=>"111111111",
  21537=>"111111111",
  21538=>"000010000",
  21539=>"001000011",
  21540=>"100010000",
  21541=>"100000110",
  21542=>"010000000",
  21543=>"001000000",
  21544=>"000001000",
  21545=>"111111111",
  21546=>"101000111",
  21547=>"000000000",
  21548=>"000001001",
  21549=>"000000000",
  21550=>"110110111",
  21551=>"111111010",
  21552=>"111111111",
  21553=>"111110011",
  21554=>"001000000",
  21555=>"000011010",
  21556=>"111111111",
  21557=>"001011010",
  21558=>"100001010",
  21559=>"100101101",
  21560=>"010111000",
  21561=>"000000111",
  21562=>"111111010",
  21563=>"101000001",
  21564=>"000001100",
  21565=>"101111111",
  21566=>"100001111",
  21567=>"100100001",
  21568=>"001111110",
  21569=>"110000000",
  21570=>"111000001",
  21571=>"011011001",
  21572=>"001111111",
  21573=>"111111010",
  21574=>"000000000",
  21575=>"010010111",
  21576=>"000000000",
  21577=>"000000111",
  21578=>"000111110",
  21579=>"110111111",
  21580=>"111001000",
  21581=>"011110001",
  21582=>"110110001",
  21583=>"011111111",
  21584=>"101000001",
  21585=>"111111111",
  21586=>"011101111",
  21587=>"111110001",
  21588=>"101000101",
  21589=>"100111001",
  21590=>"011000100",
  21591=>"111000000",
  21592=>"111010111",
  21593=>"000110111",
  21594=>"101001101",
  21595=>"111111111",
  21596=>"000110010",
  21597=>"000111000",
  21598=>"000000000",
  21599=>"110101001",
  21600=>"000000000",
  21601=>"111000000",
  21602=>"000110011",
  21603=>"101101001",
  21604=>"100110111",
  21605=>"000000101",
  21606=>"101000101",
  21607=>"110000000",
  21608=>"110111001",
  21609=>"000000000",
  21610=>"000000100",
  21611=>"110000101",
  21612=>"111111010",
  21613=>"000111110",
  21614=>"101001000",
  21615=>"000010000",
  21616=>"011110110",
  21617=>"000000001",
  21618=>"110100100",
  21619=>"000000000",
  21620=>"000000000",
  21621=>"110000000",
  21622=>"000000000",
  21623=>"110100000",
  21624=>"001010000",
  21625=>"110000000",
  21626=>"000101110",
  21627=>"000000010",
  21628=>"000000100",
  21629=>"101011110",
  21630=>"111010000",
  21631=>"001010100",
  21632=>"111000001",
  21633=>"101110111",
  21634=>"000011111",
  21635=>"000111100",
  21636=>"000111111",
  21637=>"000000000",
  21638=>"011100111",
  21639=>"001001111",
  21640=>"011011011",
  21641=>"010010110",
  21642=>"011111011",
  21643=>"111000111",
  21644=>"111111000",
  21645=>"000011000",
  21646=>"000110110",
  21647=>"101110110",
  21648=>"001000100",
  21649=>"111111111",
  21650=>"111110000",
  21651=>"000011111",
  21652=>"000011111",
  21653=>"111111111",
  21654=>"000110110",
  21655=>"110111110",
  21656=>"110000101",
  21657=>"111111101",
  21658=>"101000100",
  21659=>"000000001",
  21660=>"010011010",
  21661=>"000100000",
  21662=>"000000000",
  21663=>"001101111",
  21664=>"100110000",
  21665=>"000000000",
  21666=>"111000000",
  21667=>"010001101",
  21668=>"000001111",
  21669=>"100111111",
  21670=>"011111001",
  21671=>"001001111",
  21672=>"111100111",
  21673=>"000010000",
  21674=>"000011011",
  21675=>"001000111",
  21676=>"111111101",
  21677=>"000100111",
  21678=>"000011011",
  21679=>"110111000",
  21680=>"001000000",
  21681=>"100100100",
  21682=>"111111111",
  21683=>"100010000",
  21684=>"001000000",
  21685=>"000000011",
  21686=>"110110000",
  21687=>"100000000",
  21688=>"000100001",
  21689=>"000110101",
  21690=>"010010110",
  21691=>"000110111",
  21692=>"110000000",
  21693=>"111101100",
  21694=>"011101110",
  21695=>"110111000",
  21696=>"000000101",
  21697=>"101000000",
  21698=>"000010101",
  21699=>"110010011",
  21700=>"000000000",
  21701=>"100100000",
  21702=>"000001111",
  21703=>"111000010",
  21704=>"000011100",
  21705=>"111111101",
  21706=>"111111111",
  21707=>"100000000",
  21708=>"101000000",
  21709=>"000001001",
  21710=>"100101101",
  21711=>"111111110",
  21712=>"011000001",
  21713=>"111100000",
  21714=>"110101111",
  21715=>"001101101",
  21716=>"111000001",
  21717=>"010111011",
  21718=>"010000000",
  21719=>"110000000",
  21720=>"001000000",
  21721=>"001000101",
  21722=>"000100111",
  21723=>"000111111",
  21724=>"011111000",
  21725=>"010010111",
  21726=>"111001000",
  21727=>"010010111",
  21728=>"111100110",
  21729=>"000001111",
  21730=>"010100010",
  21731=>"111111110",
  21732=>"110110000",
  21733=>"111011000",
  21734=>"000000000",
  21735=>"100000000",
  21736=>"001011010",
  21737=>"000110110",
  21738=>"111011101",
  21739=>"001000101",
  21740=>"111111111",
  21741=>"101111010",
  21742=>"010000011",
  21743=>"010010000",
  21744=>"011000100",
  21745=>"011000010",
  21746=>"000000000",
  21747=>"000100000",
  21748=>"000001011",
  21749=>"101101101",
  21750=>"000001101",
  21751=>"010000000",
  21752=>"111111000",
  21753=>"100000000",
  21754=>"011000001",
  21755=>"110101101",
  21756=>"000000101",
  21757=>"111111111",
  21758=>"000000001",
  21759=>"001000111",
  21760=>"111101101",
  21761=>"110111111",
  21762=>"001000001",
  21763=>"100001001",
  21764=>"000000000",
  21765=>"100010010",
  21766=>"100000000",
  21767=>"000111101",
  21768=>"000000000",
  21769=>"110010110",
  21770=>"101101000",
  21771=>"000100110",
  21772=>"001001001",
  21773=>"100000100",
  21774=>"111010111",
  21775=>"110110101",
  21776=>"101000000",
  21777=>"110010110",
  21778=>"000000100",
  21779=>"000000110",
  21780=>"001101001",
  21781=>"111001111",
  21782=>"111101111",
  21783=>"000000000",
  21784=>"110110000",
  21785=>"101000111",
  21786=>"000000000",
  21787=>"100110101",
  21788=>"000101111",
  21789=>"100000011",
  21790=>"000011111",
  21791=>"110100001",
  21792=>"101101100",
  21793=>"000000000",
  21794=>"110110010",
  21795=>"000110000",
  21796=>"111111111",
  21797=>"000010000",
  21798=>"100000001",
  21799=>"100110100",
  21800=>"111101111",
  21801=>"001001010",
  21802=>"000010110",
  21803=>"011011001",
  21804=>"110100001",
  21805=>"110011011",
  21806=>"000011011",
  21807=>"011110111",
  21808=>"000000110",
  21809=>"100100001",
  21810=>"010001100",
  21811=>"001111110",
  21812=>"001000100",
  21813=>"000010011",
  21814=>"000100111",
  21815=>"110111100",
  21816=>"001001100",
  21817=>"100100110",
  21818=>"000000000",
  21819=>"100010001",
  21820=>"001001001",
  21821=>"000000000",
  21822=>"011011011",
  21823=>"100001000",
  21824=>"111001011",
  21825=>"000001101",
  21826=>"011000000",
  21827=>"011011001",
  21828=>"000010110",
  21829=>"000010010",
  21830=>"000100100",
  21831=>"000000011",
  21832=>"100111101",
  21833=>"000100000",
  21834=>"111111111",
  21835=>"100000001",
  21836=>"001001011",
  21837=>"111100111",
  21838=>"111011111",
  21839=>"001011001",
  21840=>"011001001",
  21841=>"000000000",
  21842=>"111110001",
  21843=>"101100100",
  21844=>"001000000",
  21845=>"011010011",
  21846=>"111101100",
  21847=>"010011110",
  21848=>"111110110",
  21849=>"000100100",
  21850=>"010000100",
  21851=>"001101000",
  21852=>"110110100",
  21853=>"000100100",
  21854=>"101001011",
  21855=>"001001101",
  21856=>"100110110",
  21857=>"101111101",
  21858=>"101001011",
  21859=>"110110110",
  21860=>"000100100",
  21861=>"111111111",
  21862=>"000100000",
  21863=>"000000000",
  21864=>"101111101",
  21865=>"000111111",
  21866=>"101011000",
  21867=>"011101011",
  21868=>"000001001",
  21869=>"101000101",
  21870=>"001000100",
  21871=>"100101110",
  21872=>"011010011",
  21873=>"000001000",
  21874=>"111011011",
  21875=>"011111001",
  21876=>"011111101",
  21877=>"011011010",
  21878=>"100100000",
  21879=>"000000011",
  21880=>"001011001",
  21881=>"100100100",
  21882=>"111111111",
  21883=>"011000011",
  21884=>"000000000",
  21885=>"000000000",
  21886=>"000000001",
  21887=>"111000001",
  21888=>"101011011",
  21889=>"101001101",
  21890=>"100101000",
  21891=>"000011001",
  21892=>"011001100",
  21893=>"101111111",
  21894=>"001101111",
  21895=>"110110001",
  21896=>"111111111",
  21897=>"100000000",
  21898=>"111001001",
  21899=>"001000001",
  21900=>"101101011",
  21901=>"001101001",
  21902=>"000000000",
  21903=>"000010000",
  21904=>"111111111",
  21905=>"111101101",
  21906=>"100100100",
  21907=>"011001000",
  21908=>"100000000",
  21909=>"101011011",
  21910=>"001001101",
  21911=>"100100100",
  21912=>"001000000",
  21913=>"000011000",
  21914=>"001001001",
  21915=>"111011011",
  21916=>"000100000",
  21917=>"100000111",
  21918=>"101111001",
  21919=>"011011011",
  21920=>"111101101",
  21921=>"111000111",
  21922=>"000000001",
  21923=>"011001101",
  21924=>"101001101",
  21925=>"000000100",
  21926=>"100110000",
  21927=>"100101100",
  21928=>"000110011",
  21929=>"110100001",
  21930=>"011001011",
  21931=>"101000001",
  21932=>"000000011",
  21933=>"001001001",
  21934=>"001001001",
  21935=>"000000000",
  21936=>"010100011",
  21937=>"111011110",
  21938=>"000000001",
  21939=>"000001000",
  21940=>"111100110",
  21941=>"011001100",
  21942=>"100110111",
  21943=>"000101011",
  21944=>"110100100",
  21945=>"110010000",
  21946=>"100110100",
  21947=>"001001001",
  21948=>"001101101",
  21949=>"001001001",
  21950=>"111000111",
  21951=>"000011100",
  21952=>"000011011",
  21953=>"100100100",
  21954=>"001000011",
  21955=>"111000001",
  21956=>"000000000",
  21957=>"000001011",
  21958=>"101101100",
  21959=>"100111111",
  21960=>"000100100",
  21961=>"101010011",
  21962=>"011101001",
  21963=>"100011111",
  21964=>"111111000",
  21965=>"111100100",
  21966=>"110100100",
  21967=>"111101000",
  21968=>"101001101",
  21969=>"001010001",
  21970=>"100101001",
  21971=>"000000000",
  21972=>"001101111",
  21973=>"000000011",
  21974=>"001001001",
  21975=>"101111101",
  21976=>"110000100",
  21977=>"100100100",
  21978=>"001001000",
  21979=>"001000000",
  21980=>"101001001",
  21981=>"111000000",
  21982=>"100100000",
  21983=>"001000000",
  21984=>"011001000",
  21985=>"011000000",
  21986=>"101011001",
  21987=>"111100000",
  21988=>"001000000",
  21989=>"101100001",
  21990=>"100000110",
  21991=>"100001111",
  21992=>"110011111",
  21993=>"000111110",
  21994=>"100000011",
  21995=>"000010011",
  21996=>"100010011",
  21997=>"100100110",
  21998=>"000000000",
  21999=>"000000000",
  22000=>"010011101",
  22001=>"110111011",
  22002=>"100111111",
  22003=>"000000000",
  22004=>"010110110",
  22005=>"001011011",
  22006=>"011101100",
  22007=>"110000000",
  22008=>"000001011",
  22009=>"100111100",
  22010=>"000001001",
  22011=>"101111101",
  22012=>"001001101",
  22013=>"000001001",
  22014=>"001010110",
  22015=>"101111001",
  22016=>"110011100",
  22017=>"010000010",
  22018=>"101000111",
  22019=>"000000111",
  22020=>"000000100",
  22021=>"010001111",
  22022=>"000110011",
  22023=>"010111110",
  22024=>"111001000",
  22025=>"101000101",
  22026=>"110011000",
  22027=>"000011111",
  22028=>"000000001",
  22029=>"000110010",
  22030=>"000101000",
  22031=>"111110010",
  22032=>"010110000",
  22033=>"010111011",
  22034=>"110000001",
  22035=>"000000101",
  22036=>"100100101",
  22037=>"000000111",
  22038=>"111111100",
  22039=>"010010111",
  22040=>"101000000",
  22041=>"001111001",
  22042=>"000000000",
  22043=>"111111000",
  22044=>"011010110",
  22045=>"111001000",
  22046=>"111111000",
  22047=>"101111110",
  22048=>"101101101",
  22049=>"000101111",
  22050=>"100000110",
  22051=>"000000111",
  22052=>"110100100",
  22053=>"011010101",
  22054=>"100110010",
  22055=>"000111010",
  22056=>"000010011",
  22057=>"000111110",
  22058=>"000010000",
  22059=>"100111110",
  22060=>"000111111",
  22061=>"111110111",
  22062=>"010000011",
  22063=>"001001000",
  22064=>"110111111",
  22065=>"110111100",
  22066=>"111001101",
  22067=>"001101000",
  22068=>"111111000",
  22069=>"111100000",
  22070=>"011010010",
  22071=>"101000000",
  22072=>"000000011",
  22073=>"111000000",
  22074=>"101000100",
  22075=>"000000000",
  22076=>"100110110",
  22077=>"010000000",
  22078=>"000000000",
  22079=>"001011101",
  22080=>"011001101",
  22081=>"001111000",
  22082=>"100001101",
  22083=>"110011111",
  22084=>"000000000",
  22085=>"100001000",
  22086=>"011001000",
  22087=>"111111111",
  22088=>"110100011",
  22089=>"000001000",
  22090=>"111101000",
  22091=>"000010000",
  22092=>"100010010",
  22093=>"011011010",
  22094=>"000111011",
  22095=>"000110111",
  22096=>"001010010",
  22097=>"010010101",
  22098=>"011111000",
  22099=>"000001000",
  22100=>"000100111",
  22101=>"111100000",
  22102=>"011011010",
  22103=>"111101111",
  22104=>"101000110",
  22105=>"010000001",
  22106=>"100100011",
  22107=>"110111110",
  22108=>"110000000",
  22109=>"000001000",
  22110=>"011000101",
  22111=>"010100000",
  22112=>"000111111",
  22113=>"011000111",
  22114=>"101111111",
  22115=>"010000100",
  22116=>"000111100",
  22117=>"110000100",
  22118=>"100000111",
  22119=>"100000000",
  22120=>"000101110",
  22121=>"111100000",
  22122=>"010000111",
  22123=>"011010111",
  22124=>"011000000",
  22125=>"101110101",
  22126=>"011101111",
  22127=>"111110111",
  22128=>"000011011",
  22129=>"000000000",
  22130=>"110011000",
  22131=>"111011010",
  22132=>"000111111",
  22133=>"111000000",
  22134=>"000000100",
  22135=>"010111010",
  22136=>"111000001",
  22137=>"000010000",
  22138=>"100010111",
  22139=>"000000000",
  22140=>"000100110",
  22141=>"000100000",
  22142=>"101101111",
  22143=>"100001111",
  22144=>"010000000",
  22145=>"010000000",
  22146=>"010000001",
  22147=>"010001101",
  22148=>"110010001",
  22149=>"111101101",
  22150=>"100011001",
  22151=>"000000110",
  22152=>"000110100",
  22153=>"000111010",
  22154=>"111000100",
  22155=>"000110001",
  22156=>"000000101",
  22157=>"000010000",
  22158=>"110000000",
  22159=>"000000000",
  22160=>"101000000",
  22161=>"111000111",
  22162=>"000000000",
  22163=>"011000000",
  22164=>"010011111",
  22165=>"000101100",
  22166=>"010111110",
  22167=>"000010011",
  22168=>"111111000",
  22169=>"111011111",
  22170=>"010111111",
  22171=>"001001111",
  22172=>"011000000",
  22173=>"110000111",
  22174=>"101000000",
  22175=>"000111000",
  22176=>"101011010",
  22177=>"111101111",
  22178=>"111001111",
  22179=>"111000111",
  22180=>"111111000",
  22181=>"100011011",
  22182=>"001010110",
  22183=>"110000000",
  22184=>"110111100",
  22185=>"000000110",
  22186=>"101000111",
  22187=>"110110000",
  22188=>"000110000",
  22189=>"000000000",
  22190=>"111001100",
  22191=>"111111111",
  22192=>"000000000",
  22193=>"000000001",
  22194=>"000001000",
  22195=>"011001000",
  22196=>"110111101",
  22197=>"010000000",
  22198=>"000111100",
  22199=>"000000100",
  22200=>"001011111",
  22201=>"011110011",
  22202=>"110110111",
  22203=>"111000000",
  22204=>"011110111",
  22205=>"101101011",
  22206=>"100100100",
  22207=>"111011011",
  22208=>"000000100",
  22209=>"000000000",
  22210=>"000100000",
  22211=>"100000000",
  22212=>"111111111",
  22213=>"110110000",
  22214=>"111111000",
  22215=>"000000000",
  22216=>"000011110",
  22217=>"000000000",
  22218=>"010000000",
  22219=>"000111111",
  22220=>"011010000",
  22221=>"000011010",
  22222=>"110100111",
  22223=>"101101000",
  22224=>"000110111",
  22225=>"000111011",
  22226=>"010000110",
  22227=>"011111111",
  22228=>"000000000",
  22229=>"011000000",
  22230=>"000010111",
  22231=>"001000001",
  22232=>"001101101",
  22233=>"010100000",
  22234=>"000101101",
  22235=>"101000000",
  22236=>"110011001",
  22237=>"000010111",
  22238=>"111011000",
  22239=>"001011000",
  22240=>"011100001",
  22241=>"111111011",
  22242=>"111000101",
  22243=>"010001001",
  22244=>"101100100",
  22245=>"000000001",
  22246=>"010111111",
  22247=>"010011111",
  22248=>"110100111",
  22249=>"000100111",
  22250=>"001010000",
  22251=>"010000000",
  22252=>"000000101",
  22253=>"000000000",
  22254=>"000000010",
  22255=>"010000010",
  22256=>"111000000",
  22257=>"011011000",
  22258=>"010111010",
  22259=>"111111000",
  22260=>"010010101",
  22261=>"011001011",
  22262=>"000000010",
  22263=>"101110000",
  22264=>"000000000",
  22265=>"001001101",
  22266=>"111101100",
  22267=>"000000011",
  22268=>"000111011",
  22269=>"000000000",
  22270=>"010100001",
  22271=>"000111000",
  22272=>"101011001",
  22273=>"010101111",
  22274=>"100000000",
  22275=>"000000001",
  22276=>"000100100",
  22277=>"000000001",
  22278=>"000000000",
  22279=>"000111011",
  22280=>"000000010",
  22281=>"000100111",
  22282=>"001000000",
  22283=>"000000001",
  22284=>"000000101",
  22285=>"100111001",
  22286=>"100000110",
  22287=>"000000000",
  22288=>"111001010",
  22289=>"000000010",
  22290=>"000111010",
  22291=>"110111110",
  22292=>"100101111",
  22293=>"000100000",
  22294=>"111011100",
  22295=>"111111111",
  22296=>"100100000",
  22297=>"111001000",
  22298=>"110000000",
  22299=>"000001111",
  22300=>"011101111",
  22301=>"000000000",
  22302=>"110111001",
  22303=>"000010011",
  22304=>"111101101",
  22305=>"010001111",
  22306=>"000000000",
  22307=>"111101110",
  22308=>"100100100",
  22309=>"111110111",
  22310=>"001000000",
  22311=>"000000101",
  22312=>"111001111",
  22313=>"011001000",
  22314=>"110000001",
  22315=>"000000010",
  22316=>"110100010",
  22317=>"111010111",
  22318=>"100000001",
  22319=>"111110110",
  22320=>"111000000",
  22321=>"010100110",
  22322=>"111110111",
  22323=>"100101000",
  22324=>"000000001",
  22325=>"000000001",
  22326=>"100110100",
  22327=>"100110010",
  22328=>"111010000",
  22329=>"000000000",
  22330=>"000000111",
  22331=>"101111111",
  22332=>"001001011",
  22333=>"111111111",
  22334=>"000000000",
  22335=>"110111011",
  22336=>"110100000",
  22337=>"111001111",
  22338=>"101000000",
  22339=>"011011111",
  22340=>"111110010",
  22341=>"000000000",
  22342=>"011001001",
  22343=>"111111010",
  22344=>"101011110",
  22345=>"010000011",
  22346=>"000001001",
  22347=>"000000000",
  22348=>"111111011",
  22349=>"001001011",
  22350=>"000000001",
  22351=>"111110100",
  22352=>"101101111",
  22353=>"110111111",
  22354=>"001110111",
  22355=>"011000001",
  22356=>"000000000",
  22357=>"001001110",
  22358=>"000000101",
  22359=>"001111111",
  22360=>"101101111",
  22361=>"001101111",
  22362=>"011011111",
  22363=>"100000101",
  22364=>"111111010",
  22365=>"010001011",
  22366=>"110111110",
  22367=>"100100101",
  22368=>"111000000",
  22369=>"010000100",
  22370=>"000000001",
  22371=>"110010100",
  22372=>"110110110",
  22373=>"000001000",
  22374=>"010111010",
  22375=>"111110010",
  22376=>"000010011",
  22377=>"110101000",
  22378=>"011100010",
  22379=>"011001111",
  22380=>"100000000",
  22381=>"000001001",
  22382=>"000000000",
  22383=>"000000111",
  22384=>"000100100",
  22385=>"001000111",
  22386=>"111111000",
  22387=>"100000000",
  22388=>"000111010",
  22389=>"100000000",
  22390=>"011111111",
  22391=>"101001001",
  22392=>"011000010",
  22393=>"000011011",
  22394=>"110110111",
  22395=>"100110111",
  22396=>"100110101",
  22397=>"110000000",
  22398=>"000000001",
  22399=>"000000111",
  22400=>"111001000",
  22401=>"000101110",
  22402=>"000011111",
  22403=>"001110010",
  22404=>"010100000",
  22405=>"000000001",
  22406=>"100110011",
  22407=>"110010010",
  22408=>"110111111",
  22409=>"111000000",
  22410=>"000000000",
  22411=>"101101111",
  22412=>"101010000",
  22413=>"101000001",
  22414=>"000000000",
  22415=>"001000000",
  22416=>"111001001",
  22417=>"111110110",
  22418=>"000011000",
  22419=>"000000000",
  22420=>"000000110",
  22421=>"001000111",
  22422=>"011111010",
  22423=>"010100001",
  22424=>"011000010",
  22425=>"000110111",
  22426=>"000011010",
  22427=>"101100100",
  22428=>"111100000",
  22429=>"000110111",
  22430=>"101001111",
  22431=>"111001111",
  22432=>"101111111",
  22433=>"010111111",
  22434=>"100110100",
  22435=>"111000101",
  22436=>"000100111",
  22437=>"101001000",
  22438=>"001001001",
  22439=>"110111111",
  22440=>"010001000",
  22441=>"000011111",
  22442=>"111000000",
  22443=>"111000000",
  22444=>"111110000",
  22445=>"000000101",
  22446=>"011111110",
  22447=>"000000000",
  22448=>"111111111",
  22449=>"011001000",
  22450=>"010000000",
  22451=>"000000000",
  22452=>"011011101",
  22453=>"001000101",
  22454=>"000000100",
  22455=>"111100011",
  22456=>"000000100",
  22457=>"000110111",
  22458=>"000010111",
  22459=>"111010010",
  22460=>"111011110",
  22461=>"000010111",
  22462=>"000111000",
  22463=>"010111011",
  22464=>"001000000",
  22465=>"000000111",
  22466=>"111001010",
  22467=>"001001001",
  22468=>"000000000",
  22469=>"111000101",
  22470=>"110111100",
  22471=>"111111111",
  22472=>"000010111",
  22473=>"000001000",
  22474=>"110011111",
  22475=>"000000000",
  22476=>"000011011",
  22477=>"111111101",
  22478=>"011000000",
  22479=>"011110001",
  22480=>"000111111",
  22481=>"001001000",
  22482=>"000001001",
  22483=>"010101111",
  22484=>"001000101",
  22485=>"110110000",
  22486=>"101111111",
  22487=>"000000010",
  22488=>"000111111",
  22489=>"000111010",
  22490=>"101101110",
  22491=>"101000001",
  22492=>"110000000",
  22493=>"100010011",
  22494=>"000000000",
  22495=>"000001111",
  22496=>"111000000",
  22497=>"111101001",
  22498=>"000000000",
  22499=>"011010110",
  22500=>"111000000",
  22501=>"111001000",
  22502=>"000111111",
  22503=>"100111000",
  22504=>"100000101",
  22505=>"010111000",
  22506=>"000000000",
  22507=>"111000000",
  22508=>"000000011",
  22509=>"101001101",
  22510=>"101001001",
  22511=>"000000110",
  22512=>"100110101",
  22513=>"111100110",
  22514=>"011011011",
  22515=>"100000011",
  22516=>"001111110",
  22517=>"000000000",
  22518=>"000000110",
  22519=>"100010000",
  22520=>"001111111",
  22521=>"000000011",
  22522=>"111100111",
  22523=>"000000010",
  22524=>"111111010",
  22525=>"111101100",
  22526=>"001011001",
  22527=>"100000000",
  22528=>"001000111",
  22529=>"110100111",
  22530=>"001000111",
  22531=>"010101100",
  22532=>"110100100",
  22533=>"111111111",
  22534=>"000101001",
  22535=>"011001111",
  22536=>"000101101",
  22537=>"000011011",
  22538=>"111110001",
  22539=>"001011001",
  22540=>"111111010",
  22541=>"000000101",
  22542=>"101111000",
  22543=>"000001111",
  22544=>"111011110",
  22545=>"010010010",
  22546=>"010111010",
  22547=>"111110101",
  22548=>"100101101",
  22549=>"011011111",
  22550=>"010111010",
  22551=>"010111011",
  22552=>"110100100",
  22553=>"001111110",
  22554=>"100100111",
  22555=>"000011111",
  22556=>"010011100",
  22557=>"100101001",
  22558=>"111101111",
  22559=>"010111000",
  22560=>"011100111",
  22561=>"001011011",
  22562=>"011000011",
  22563=>"101101100",
  22564=>"111111010",
  22565=>"100111111",
  22566=>"100000000",
  22567=>"000011000",
  22568=>"100100101",
  22569=>"000101000",
  22570=>"100110011",
  22571=>"010000000",
  22572=>"110111110",
  22573=>"111111010",
  22574=>"000001100",
  22575=>"111101101",
  22576=>"000110010",
  22577=>"011011110",
  22578=>"000000010",
  22579=>"011000010",
  22580=>"011000010",
  22581=>"100010000",
  22582=>"100000001",
  22583=>"010111001",
  22584=>"011000000",
  22585=>"010000000",
  22586=>"010001000",
  22587=>"000000000",
  22588=>"100011100",
  22589=>"111111011",
  22590=>"000010000",
  22591=>"010111001",
  22592=>"000000111",
  22593=>"101011000",
  22594=>"111111000",
  22595=>"110111000",
  22596=>"101100000",
  22597=>"000000000",
  22598=>"000000000",
  22599=>"111010111",
  22600=>"100000100",
  22601=>"011010100",
  22602=>"000000000",
  22603=>"111101100",
  22604=>"111111010",
  22605=>"111100011",
  22606=>"011011001",
  22607=>"111010111",
  22608=>"011001000",
  22609=>"111111100",
  22610=>"011000110",
  22611=>"011011000",
  22612=>"101101101",
  22613=>"110100111",
  22614=>"011000000",
  22615=>"000111000",
  22616=>"100111100",
  22617=>"111111110",
  22618=>"110110000",
  22619=>"011111001",
  22620=>"010010000",
  22621=>"000000001",
  22622=>"000111000",
  22623=>"011111011",
  22624=>"000100000",
  22625=>"010110010",
  22626=>"101100101",
  22627=>"000110100",
  22628=>"010011110",
  22629=>"111010111",
  22630=>"001011000",
  22631=>"101111010",
  22632=>"010010011",
  22633=>"011000100",
  22634=>"000011011",
  22635=>"111000111",
  22636=>"011111001",
  22637=>"011011000",
  22638=>"000011000",
  22639=>"110000000",
  22640=>"001001000",
  22641=>"010101100",
  22642=>"011000110",
  22643=>"111101111",
  22644=>"101100110",
  22645=>"000000010",
  22646=>"100101000",
  22647=>"001100000",
  22648=>"000001001",
  22649=>"010110000",
  22650=>"000010111",
  22651=>"001001000",
  22652=>"111111111",
  22653=>"000110010",
  22654=>"010011010",
  22655=>"010111010",
  22656=>"100000110",
  22657=>"111111011",
  22658=>"000001010",
  22659=>"000000001",
  22660=>"000000111",
  22661=>"000010000",
  22662=>"000010011",
  22663=>"011001000",
  22664=>"000011000",
  22665=>"010000100",
  22666=>"010000000",
  22667=>"011111111",
  22668=>"000001000",
  22669=>"000010000",
  22670=>"101111111",
  22671=>"000001011",
  22672=>"110110111",
  22673=>"000100000",
  22674=>"110011011",
  22675=>"111100101",
  22676=>"000000000",
  22677=>"000000000",
  22678=>"111101000",
  22679=>"010100011",
  22680=>"011011000",
  22681=>"000101111",
  22682=>"101100100",
  22683=>"000111111",
  22684=>"000011011",
  22685=>"100100110",
  22686=>"101000010",
  22687=>"101000000",
  22688=>"000011001",
  22689=>"101001010",
  22690=>"000011011",
  22691=>"100010011",
  22692=>"100000000",
  22693=>"100100100",
  22694=>"010111011",
  22695=>"000000000",
  22696=>"000011000",
  22697=>"100101111",
  22698=>"111011010",
  22699=>"000010000",
  22700=>"010010011",
  22701=>"101100111",
  22702=>"111110100",
  22703=>"000111001",
  22704=>"000010111",
  22705=>"110001110",
  22706=>"111100100",
  22707=>"000100010",
  22708=>"000011010",
  22709=>"000010010",
  22710=>"110100000",
  22711=>"000010100",
  22712=>"000010001",
  22713=>"001000011",
  22714=>"111011000",
  22715=>"111111011",
  22716=>"000011011",
  22717=>"111111110",
  22718=>"001011111",
  22719=>"010000000",
  22720=>"000000000",
  22721=>"010111011",
  22722=>"001111111",
  22723=>"100100111",
  22724=>"000000101",
  22725=>"110110110",
  22726=>"000101111",
  22727=>"000000100",
  22728=>"101000000",
  22729=>"100000000",
  22730=>"000000010",
  22731=>"000011011",
  22732=>"010000000",
  22733=>"100111011",
  22734=>"111010011",
  22735=>"000011010",
  22736=>"000100000",
  22737=>"011000000",
  22738=>"000101000",
  22739=>"111011000",
  22740=>"000111111",
  22741=>"110110110",
  22742=>"000000000",
  22743=>"011010000",
  22744=>"001101111",
  22745=>"000010111",
  22746=>"000110010",
  22747=>"000000000",
  22748=>"001100011",
  22749=>"101101011",
  22750=>"000000011",
  22751=>"111110000",
  22752=>"111111111",
  22753=>"101010101",
  22754=>"000100101",
  22755=>"001011011",
  22756=>"000100000",
  22757=>"111100111",
  22758=>"011000000",
  22759=>"011010010",
  22760=>"101100100",
  22761=>"000100110",
  22762=>"111001000",
  22763=>"000000000",
  22764=>"000000110",
  22765=>"111010000",
  22766=>"111111010",
  22767=>"010000111",
  22768=>"000100100",
  22769=>"111001001",
  22770=>"100000000",
  22771=>"010011000",
  22772=>"000000000",
  22773=>"000110100",
  22774=>"000111110",
  22775=>"010100000",
  22776=>"000010010",
  22777=>"000100000",
  22778=>"000111011",
  22779=>"111001111",
  22780=>"111101111",
  22781=>"100100111",
  22782=>"001000001",
  22783=>"000011011",
  22784=>"001100101",
  22785=>"000000000",
  22786=>"101000001",
  22787=>"101000000",
  22788=>"000100001",
  22789=>"010000100",
  22790=>"010001111",
  22791=>"001011000",
  22792=>"101111000",
  22793=>"111000111",
  22794=>"000111111",
  22795=>"111000000",
  22796=>"111111011",
  22797=>"000000010",
  22798=>"000100100",
  22799=>"001111000",
  22800=>"100100111",
  22801=>"000111111",
  22802=>"101000000",
  22803=>"111110000",
  22804=>"000000000",
  22805=>"010010000",
  22806=>"100110100",
  22807=>"100111111",
  22808=>"000000101",
  22809=>"110111111",
  22810=>"010111111",
  22811=>"000010000",
  22812=>"000111111",
  22813=>"000010111",
  22814=>"100110011",
  22815=>"011011000",
  22816=>"111101100",
  22817=>"101000101",
  22818=>"000000000",
  22819=>"101100000",
  22820=>"001010011",
  22821=>"111011110",
  22822=>"011111001",
  22823=>"101000100",
  22824=>"000001101",
  22825=>"101001100",
  22826=>"111111100",
  22827=>"111101101",
  22828=>"111110110",
  22829=>"110000111",
  22830=>"000000111",
  22831=>"010111000",
  22832=>"000000101",
  22833=>"100111011",
  22834=>"000010111",
  22835=>"111010001",
  22836=>"000011000",
  22837=>"111111110",
  22838=>"110011011",
  22839=>"110011010",
  22840=>"010011010",
  22841=>"000000000",
  22842=>"000000000",
  22843=>"000000000",
  22844=>"111111001",
  22845=>"111111111",
  22846=>"101000000",
  22847=>"010011001",
  22848=>"111111001",
  22849=>"011111111",
  22850=>"000101000",
  22851=>"001000110",
  22852=>"010000000",
  22853=>"000010000",
  22854=>"111111001",
  22855=>"000010111",
  22856=>"001010000",
  22857=>"000000000",
  22858=>"000000000",
  22859=>"000000111",
  22860=>"100011011",
  22861=>"110111111",
  22862=>"001111001",
  22863=>"000001000",
  22864=>"011011011",
  22865=>"010111111",
  22866=>"111111100",
  22867=>"000000100",
  22868=>"011111000",
  22869=>"101111111",
  22870=>"000011011",
  22871=>"111100111",
  22872=>"011111011",
  22873=>"100011010",
  22874=>"101111001",
  22875=>"111111011",
  22876=>"111111010",
  22877=>"000010110",
  22878=>"101000100",
  22879=>"101001011",
  22880=>"011111001",
  22881=>"100000000",
  22882=>"111101111",
  22883=>"110111001",
  22884=>"001000001",
  22885=>"111010000",
  22886=>"000000000",
  22887=>"100101101",
  22888=>"000000000",
  22889=>"000110111",
  22890=>"111011011",
  22891=>"111111101",
  22892=>"000000001",
  22893=>"000100000",
  22894=>"000011010",
  22895=>"000010111",
  22896=>"011011011",
  22897=>"111111110",
  22898=>"011110110",
  22899=>"000001011",
  22900=>"000010010",
  22901=>"001000000",
  22902=>"000010001",
  22903=>"000111000",
  22904=>"000000000",
  22905=>"101000100",
  22906=>"000001111",
  22907=>"001000000",
  22908=>"111111000",
  22909=>"000000000",
  22910=>"101000101",
  22911=>"010010000",
  22912=>"111110101",
  22913=>"000011011",
  22914=>"000010000",
  22915=>"000000111",
  22916=>"011111111",
  22917=>"111111111",
  22918=>"111111101",
  22919=>"111101111",
  22920=>"110110110",
  22921=>"101101101",
  22922=>"000100111",
  22923=>"100011100",
  22924=>"000000000",
  22925=>"111000000",
  22926=>"111011100",
  22927=>"001000010",
  22928=>"010111110",
  22929=>"101010000",
  22930=>"001100110",
  22931=>"001011001",
  22932=>"111011011",
  22933=>"100100000",
  22934=>"111111000",
  22935=>"111000001",
  22936=>"000000101",
  22937=>"000000000",
  22938=>"010111010",
  22939=>"111000100",
  22940=>"010011111",
  22941=>"111000000",
  22942=>"110111101",
  22943=>"010111011",
  22944=>"100010010",
  22945=>"111111000",
  22946=>"000000000",
  22947=>"101111111",
  22948=>"111111011",
  22949=>"110111110",
  22950=>"110111110",
  22951=>"101100000",
  22952=>"110001111",
  22953=>"010000000",
  22954=>"000011000",
  22955=>"000010011",
  22956=>"101000100",
  22957=>"011101100",
  22958=>"101111110",
  22959=>"101100100",
  22960=>"101010000",
  22961=>"111010000",
  22962=>"000100100",
  22963=>"001010011",
  22964=>"001011001",
  22965=>"000011000",
  22966=>"000000000",
  22967=>"100101100",
  22968=>"111111011",
  22969=>"001010011",
  22970=>"001011111",
  22971=>"111111111",
  22972=>"011001111",
  22973=>"000010011",
  22974=>"000110100",
  22975=>"000011011",
  22976=>"101100000",
  22977=>"100100000",
  22978=>"010010011",
  22979=>"110111011",
  22980=>"010100111",
  22981=>"000001101",
  22982=>"011111001",
  22983=>"111101111",
  22984=>"000010000",
  22985=>"010111111",
  22986=>"000000010",
  22987=>"001001011",
  22988=>"100000000",
  22989=>"011101011",
  22990=>"110000111",
  22991=>"100010111",
  22992=>"100010000",
  22993=>"100100100",
  22994=>"111111101",
  22995=>"111111111",
  22996=>"000001001",
  22997=>"100010000",
  22998=>"000000000",
  22999=>"000010010",
  23000=>"111111000",
  23001=>"011000000",
  23002=>"001001000",
  23003=>"001100101",
  23004=>"001111100",
  23005=>"010010110",
  23006=>"010001011",
  23007=>"111111111",
  23008=>"000111111",
  23009=>"000101011",
  23010=>"111111100",
  23011=>"001011011",
  23012=>"000000000",
  23013=>"111111000",
  23014=>"111111010",
  23015=>"111011011",
  23016=>"011110010",
  23017=>"000110111",
  23018=>"111011000",
  23019=>"010110010",
  23020=>"110111111",
  23021=>"101101010",
  23022=>"111101101",
  23023=>"011000000",
  23024=>"000011000",
  23025=>"100100111",
  23026=>"000000100",
  23027=>"001000000",
  23028=>"110000110",
  23029=>"010010111",
  23030=>"111010100",
  23031=>"100100111",
  23032=>"111001010",
  23033=>"001000000",
  23034=>"000010010",
  23035=>"010010000",
  23036=>"000000000",
  23037=>"000100000",
  23038=>"101111111",
  23039=>"101011001",
  23040=>"100101100",
  23041=>"000000000",
  23042=>"111001000",
  23043=>"011110101",
  23044=>"000101011",
  23045=>"101100010",
  23046=>"000010110",
  23047=>"001011111",
  23048=>"000001111",
  23049=>"000000010",
  23050=>"000110111",
  23051=>"000111011",
  23052=>"100100000",
  23053=>"110110000",
  23054=>"110101101",
  23055=>"001100000",
  23056=>"110111011",
  23057=>"111000000",
  23058=>"000100000",
  23059=>"101001000",
  23060=>"000010000",
  23061=>"110111011",
  23062=>"000100000",
  23063=>"111000100",
  23064=>"010000000",
  23065=>"000110010",
  23066=>"000111111",
  23067=>"000000111",
  23068=>"101101001",
  23069=>"011111000",
  23070=>"000000011",
  23071=>"111000000",
  23072=>"111000000",
  23073=>"000000101",
  23074=>"000000000",
  23075=>"001101100",
  23076=>"001101111",
  23077=>"000100111",
  23078=>"111000111",
  23079=>"000000110",
  23080=>"111010110",
  23081=>"000000111",
  23082=>"100000111",
  23083=>"100110000",
  23084=>"010110101",
  23085=>"010111101",
  23086=>"110011010",
  23087=>"010111100",
  23088=>"011111001",
  23089=>"000100101",
  23090=>"000010001",
  23091=>"000000111",
  23092=>"001101110",
  23093=>"000000101",
  23094=>"001000000",
  23095=>"000000111",
  23096=>"001110111",
  23097=>"101000011",
  23098=>"111101100",
  23099=>"000000000",
  23100=>"001001111",
  23101=>"000010111",
  23102=>"000000000",
  23103=>"000010011",
  23104=>"000000110",
  23105=>"000100111",
  23106=>"111101101",
  23107=>"100110110",
  23108=>"010111000",
  23109=>"000000000",
  23110=>"000110000",
  23111=>"010101101",
  23112=>"001110111",
  23113=>"000111010",
  23114=>"011011111",
  23115=>"111100000",
  23116=>"101000010",
  23117=>"110111011",
  23118=>"000000100",
  23119=>"101111111",
  23120=>"111001001",
  23121=>"111111111",
  23122=>"101111111",
  23123=>"000101000",
  23124=>"111000000",
  23125=>"011001110",
  23126=>"000100100",
  23127=>"000000010",
  23128=>"010001000",
  23129=>"010011110",
  23130=>"011000100",
  23131=>"100110101",
  23132=>"101000111",
  23133=>"010000000",
  23134=>"111111110",
  23135=>"011011011",
  23136=>"000000000",
  23137=>"110111010",
  23138=>"111100000",
  23139=>"111000000",
  23140=>"011011101",
  23141=>"000011011",
  23142=>"111111110",
  23143=>"000011111",
  23144=>"000010011",
  23145=>"111110000",
  23146=>"000111111",
  23147=>"111111111",
  23148=>"010011111",
  23149=>"111000000",
  23150=>"000000000",
  23151=>"000101100",
  23152=>"111111101",
  23153=>"000010111",
  23154=>"110000000",
  23155=>"110100000",
  23156=>"000111101",
  23157=>"000000001",
  23158=>"110000000",
  23159=>"000000010",
  23160=>"111000010",
  23161=>"111111010",
  23162=>"101011001",
  23163=>"000101001",
  23164=>"010110000",
  23165=>"110101000",
  23166=>"111110000",
  23167=>"111101111",
  23168=>"000000000",
  23169=>"000111000",
  23170=>"000011011",
  23171=>"000011111",
  23172=>"000011110",
  23173=>"000000001",
  23174=>"000001111",
  23175=>"000000011",
  23176=>"110110100",
  23177=>"000011111",
  23178=>"000011100",
  23179=>"100100000",
  23180=>"110000000",
  23181=>"100000100",
  23182=>"000100111",
  23183=>"000000000",
  23184=>"010011111",
  23185=>"000100000",
  23186=>"111110010",
  23187=>"111111111",
  23188=>"000010001",
  23189=>"111110010",
  23190=>"111111111",
  23191=>"000001011",
  23192=>"101001101",
  23193=>"110111011",
  23194=>"000001000",
  23195=>"111101000",
  23196=>"000110111",
  23197=>"000101011",
  23198=>"000111011",
  23199=>"010101011",
  23200=>"110110110",
  23201=>"000000101",
  23202=>"110111111",
  23203=>"110010000",
  23204=>"111010011",
  23205=>"000100100",
  23206=>"100101001",
  23207=>"010111011",
  23208=>"100001000",
  23209=>"000000100",
  23210=>"010101000",
  23211=>"101000000",
  23212=>"001101101",
  23213=>"000100010",
  23214=>"011011000",
  23215=>"111101000",
  23216=>"001111111",
  23217=>"011010100",
  23218=>"100001000",
  23219=>"000000110",
  23220=>"010011101",
  23221=>"100100100",
  23222=>"000000000",
  23223=>"100100000",
  23224=>"000110011",
  23225=>"000010111",
  23226=>"000111111",
  23227=>"010111111",
  23228=>"011110010",
  23229=>"111100000",
  23230=>"000100110",
  23231=>"000000010",
  23232=>"110110010",
  23233=>"100000010",
  23234=>"101011001",
  23235=>"111111011",
  23236=>"000000111",
  23237=>"111100101",
  23238=>"000000110",
  23239=>"000111011",
  23240=>"111110110",
  23241=>"101000110",
  23242=>"111000000",
  23243=>"111001011",
  23244=>"000111111",
  23245=>"000001011",
  23246=>"010000000",
  23247=>"100000111",
  23248=>"101001010",
  23249=>"000011000",
  23250=>"000000011",
  23251=>"000010100",
  23252=>"000010000",
  23253=>"111001001",
  23254=>"001111111",
  23255=>"000110010",
  23256=>"111010110",
  23257=>"000001000",
  23258=>"000001000",
  23259=>"111101000",
  23260=>"001001011",
  23261=>"100100001",
  23262=>"000000000",
  23263=>"001110111",
  23264=>"001001011",
  23265=>"011111100",
  23266=>"111011000",
  23267=>"011111000",
  23268=>"111110110",
  23269=>"000110111",
  23270=>"101100111",
  23271=>"000000000",
  23272=>"000110011",
  23273=>"010010001",
  23274=>"000011111",
  23275=>"111101100",
  23276=>"000000011",
  23277=>"000001011",
  23278=>"000001000",
  23279=>"001111111",
  23280=>"000101111",
  23281=>"000001101",
  23282=>"000111010",
  23283=>"000101001",
  23284=>"000001110",
  23285=>"111000100",
  23286=>"110100000",
  23287=>"000111000",
  23288=>"000000000",
  23289=>"011111000",
  23290=>"000010010",
  23291=>"110100101",
  23292=>"101111111",
  23293=>"110000111",
  23294=>"000110111",
  23295=>"010100001",
  23296=>"111011011",
  23297=>"111111101",
  23298=>"101000101",
  23299=>"110000101",
  23300=>"011111001",
  23301=>"110110101",
  23302=>"000101010",
  23303=>"000110000",
  23304=>"000100111",
  23305=>"111000101",
  23306=>"100000000",
  23307=>"000000111",
  23308=>"011111111",
  23309=>"000000000",
  23310=>"111001100",
  23311=>"000100000",
  23312=>"010000000",
  23313=>"000000000",
  23314=>"000000111",
  23315=>"011010000",
  23316=>"111111110",
  23317=>"000000010",
  23318=>"110111111",
  23319=>"100101101",
  23320=>"001010000",
  23321=>"111111111",
  23322=>"011010100",
  23323=>"110101101",
  23324=>"101101101",
  23325=>"001001010",
  23326=>"000000011",
  23327=>"001000001",
  23328=>"111010101",
  23329=>"110101111",
  23330=>"101000111",
  23331=>"010010000",
  23332=>"000011011",
  23333=>"111110110",
  23334=>"000000000",
  23335=>"001101111",
  23336=>"111001101",
  23337=>"001100010",
  23338=>"000000000",
  23339=>"010101111",
  23340=>"111111011",
  23341=>"101101100",
  23342=>"110010101",
  23343=>"000101110",
  23344=>"110101001",
  23345=>"011011101",
  23346=>"000110000",
  23347=>"110000010",
  23348=>"000000010",
  23349=>"010111011",
  23350=>"001000000",
  23351=>"000000111",
  23352=>"101000100",
  23353=>"000011011",
  23354=>"011001010",
  23355=>"111000100",
  23356=>"110100101",
  23357=>"111111000",
  23358=>"000000001",
  23359=>"100100100",
  23360=>"000001111",
  23361=>"111111101",
  23362=>"101000111",
  23363=>"011000001",
  23364=>"000001000",
  23365=>"001011010",
  23366=>"100110010",
  23367=>"001000101",
  23368=>"110100010",
  23369=>"010111111",
  23370=>"000001101",
  23371=>"001111110",
  23372=>"000010010",
  23373=>"010010111",
  23374=>"000111010",
  23375=>"001100100",
  23376=>"000000000",
  23377=>"111000110",
  23378=>"010001000",
  23379=>"011001000",
  23380=>"100110101",
  23381=>"101001101",
  23382=>"111101000",
  23383=>"111000000",
  23384=>"100110111",
  23385=>"000111111",
  23386=>"111000000",
  23387=>"001100110",
  23388=>"010000000",
  23389=>"010000000",
  23390=>"010110010",
  23391=>"100000100",
  23392=>"100111111",
  23393=>"000111011",
  23394=>"000000001",
  23395=>"111101010",
  23396=>"101000000",
  23397=>"111100111",
  23398=>"110110010",
  23399=>"000000111",
  23400=>"111001011",
  23401=>"000000010",
  23402=>"000111111",
  23403=>"010011101",
  23404=>"111111001",
  23405=>"000010010",
  23406=>"001000100",
  23407=>"000011111",
  23408=>"101001011",
  23409=>"000000110",
  23410=>"100000000",
  23411=>"000010000",
  23412=>"010100100",
  23413=>"101000001",
  23414=>"111101010",
  23415=>"000000111",
  23416=>"101101101",
  23417=>"111111111",
  23418=>"011111110",
  23419=>"010111110",
  23420=>"010010100",
  23421=>"110100100",
  23422=>"001010111",
  23423=>"101001001",
  23424=>"010110000",
  23425=>"111111111",
  23426=>"101100000",
  23427=>"000111111",
  23428=>"010111111",
  23429=>"111101001",
  23430=>"110011001",
  23431=>"000100011",
  23432=>"001110110",
  23433=>"111010000",
  23434=>"000111101",
  23435=>"000000000",
  23436=>"000110110",
  23437=>"001000001",
  23438=>"101000101",
  23439=>"000000000",
  23440=>"001110110",
  23441=>"111101101",
  23442=>"000110000",
  23443=>"000111111",
  23444=>"111111000",
  23445=>"110110000",
  23446=>"010011111",
  23447=>"000100110",
  23448=>"101111000",
  23449=>"000111101",
  23450=>"010100111",
  23451=>"000101111",
  23452=>"110111011",
  23453=>"010101101",
  23454=>"000001100",
  23455=>"000111011",
  23456=>"000000111",
  23457=>"101000101",
  23458=>"000001000",
  23459=>"000100000",
  23460=>"000101100",
  23461=>"000110010",
  23462=>"001010110",
  23463=>"000000000",
  23464=>"111111100",
  23465=>"000001101",
  23466=>"111000001",
  23467=>"111101000",
  23468=>"000010111",
  23469=>"101001101",
  23470=>"110011111",
  23471=>"000101111",
  23472=>"011011101",
  23473=>"001111110",
  23474=>"010001000",
  23475=>"000001000",
  23476=>"000001011",
  23477=>"101111111",
  23478=>"000111011",
  23479=>"111111010",
  23480=>"011001100",
  23481=>"001011110",
  23482=>"000000101",
  23483=>"010010111",
  23484=>"111010000",
  23485=>"111111111",
  23486=>"000010100",
  23487=>"000100111",
  23488=>"000000000",
  23489=>"011000100",
  23490=>"111101101",
  23491=>"000010011",
  23492=>"111010000",
  23493=>"001110100",
  23494=>"010110111",
  23495=>"111001000",
  23496=>"000000000",
  23497=>"000011110",
  23498=>"110000011",
  23499=>"100100111",
  23500=>"000000100",
  23501=>"001001011",
  23502=>"010000000",
  23503=>"111111110",
  23504=>"001000000",
  23505=>"011111110",
  23506=>"000111111",
  23507=>"001101010",
  23508=>"010000000",
  23509=>"000000111",
  23510=>"110000100",
  23511=>"000101101",
  23512=>"011101000",
  23513=>"001111101",
  23514=>"100000001",
  23515=>"100000000",
  23516=>"110111001",
  23517=>"101000101",
  23518=>"100111111",
  23519=>"111000111",
  23520=>"111100100",
  23521=>"111001000",
  23522=>"111111110",
  23523=>"111111011",
  23524=>"000000000",
  23525=>"110111000",
  23526=>"111101101",
  23527=>"100100111",
  23528=>"010101010",
  23529=>"000000001",
  23530=>"111110000",
  23531=>"001000000",
  23532=>"000010011",
  23533=>"101111010",
  23534=>"000000011",
  23535=>"000000000",
  23536=>"110111100",
  23537=>"111111100",
  23538=>"010001111",
  23539=>"000100010",
  23540=>"110110110",
  23541=>"101000000",
  23542=>"000000000",
  23543=>"111101111",
  23544=>"010000000",
  23545=>"100101101",
  23546=>"000000000",
  23547=>"000111111",
  23548=>"101100111",
  23549=>"110100100",
  23550=>"010000110",
  23551=>"111000000",
  23552=>"100001001",
  23553=>"111000000",
  23554=>"000000000",
  23555=>"110111011",
  23556=>"100110111",
  23557=>"001000111",
  23558=>"100111111",
  23559=>"101001011",
  23560=>"001101101",
  23561=>"000111111",
  23562=>"000110110",
  23563=>"101101000",
  23564=>"000000001",
  23565=>"100100000",
  23566=>"111011110",
  23567=>"001001000",
  23568=>"100111110",
  23569=>"000001000",
  23570=>"000110000",
  23571=>"000011111",
  23572=>"111111101",
  23573=>"101101000",
  23574=>"111111111",
  23575=>"000000010",
  23576=>"110101000",
  23577=>"111111111",
  23578=>"100101001",
  23579=>"100111011",
  23580=>"101101000",
  23581=>"010000010",
  23582=>"001011111",
  23583=>"001001001",
  23584=>"000000101",
  23585=>"000110011",
  23586=>"111011000",
  23587=>"101001111",
  23588=>"110110000",
  23589=>"011111111",
  23590=>"111111111",
  23591=>"011111000",
  23592=>"011000000",
  23593=>"100111010",
  23594=>"000111111",
  23595=>"111111000",
  23596=>"011010110",
  23597=>"110111100",
  23598=>"110110111",
  23599=>"000000111",
  23600=>"111000000",
  23601=>"110110011",
  23602=>"000001010",
  23603=>"101011110",
  23604=>"001000000",
  23605=>"110000110",
  23606=>"111110110",
  23607=>"101000000",
  23608=>"111000000",
  23609=>"000000100",
  23610=>"000011111",
  23611=>"110000010",
  23612=>"001000100",
  23613=>"011011111",
  23614=>"000000100",
  23615=>"110110111",
  23616=>"101101000",
  23617=>"001111100",
  23618=>"111111110",
  23619=>"000000100",
  23620=>"000000000",
  23621=>"000000111",
  23622=>"001011001",
  23623=>"111111110",
  23624=>"011011010",
  23625=>"001111111",
  23626=>"100000000",
  23627=>"100000011",
  23628=>"100001001",
  23629=>"110011011",
  23630=>"011000010",
  23631=>"011111111",
  23632=>"000010010",
  23633=>"010111011",
  23634=>"011001000",
  23635=>"011001111",
  23636=>"000101101",
  23637=>"001001111",
  23638=>"010011001",
  23639=>"001001001",
  23640=>"000110110",
  23641=>"111110001",
  23642=>"100001000",
  23643=>"110111110",
  23644=>"001001101",
  23645=>"010011000",
  23646=>"100101101",
  23647=>"000001011",
  23648=>"000000000",
  23649=>"000000100",
  23650=>"101101100",
  23651=>"101111110",
  23652=>"111111110",
  23653=>"110010100",
  23654=>"101101000",
  23655=>"101000000",
  23656=>"001011001",
  23657=>"111111111",
  23658=>"101111111",
  23659=>"101001001",
  23660=>"001000000",
  23661=>"101101000",
  23662=>"001000101",
  23663=>"100000010",
  23664=>"011001111",
  23665=>"101111000",
  23666=>"111001011",
  23667=>"011000000",
  23668=>"000000000",
  23669=>"000000100",
  23670=>"111111111",
  23671=>"000000000",
  23672=>"000111101",
  23673=>"111111101",
  23674=>"101100001",
  23675=>"011000111",
  23676=>"001000011",
  23677=>"010100100",
  23678=>"000010000",
  23679=>"000111111",
  23680=>"111101000",
  23681=>"000111111",
  23682=>"100100100",
  23683=>"111010010",
  23684=>"010000101",
  23685=>"111111110",
  23686=>"100111111",
  23687=>"100000110",
  23688=>"110000000",
  23689=>"111011010",
  23690=>"011101000",
  23691=>"101101000",
  23692=>"101101111",
  23693=>"101101101",
  23694=>"010111111",
  23695=>"000100101",
  23696=>"011010100",
  23697=>"000101101",
  23698=>"101101111",
  23699=>"001001100",
  23700=>"111110100",
  23701=>"000101001",
  23702=>"000010010",
  23703=>"110101001",
  23704=>"010101111",
  23705=>"101001001",
  23706=>"000000010",
  23707=>"001111111",
  23708=>"100011000",
  23709=>"000100000",
  23710=>"111111100",
  23711=>"000101001",
  23712=>"110100010",
  23713=>"001101100",
  23714=>"001010011",
  23715=>"101000000",
  23716=>"010010111",
  23717=>"111011010",
  23718=>"111001000",
  23719=>"000010111",
  23720=>"010100111",
  23721=>"000001011",
  23722=>"101000011",
  23723=>"001111001",
  23724=>"000100000",
  23725=>"000000000",
  23726=>"000000000",
  23727=>"101100100",
  23728=>"001001101",
  23729=>"001001011",
  23730=>"111000110",
  23731=>"011010010",
  23732=>"100111100",
  23733=>"111110001",
  23734=>"100000100",
  23735=>"001101101",
  23736=>"100000101",
  23737=>"001001011",
  23738=>"111101111",
  23739=>"001100100",
  23740=>"111110111",
  23741=>"101111111",
  23742=>"111001111",
  23743=>"001100000",
  23744=>"000000100",
  23745=>"010011100",
  23746=>"000000001",
  23747=>"010010010",
  23748=>"111111110",
  23749=>"011111100",
  23750=>"000100101",
  23751=>"010010010",
  23752=>"101100111",
  23753=>"011001000",
  23754=>"000101011",
  23755=>"101100110",
  23756=>"000001111",
  23757=>"000100111",
  23758=>"000000101",
  23759=>"000000101",
  23760=>"110010110",
  23761=>"010111001",
  23762=>"100010001",
  23763=>"101111000",
  23764=>"000000111",
  23765=>"001000000",
  23766=>"000101101",
  23767=>"010011111",
  23768=>"101001111",
  23769=>"111101001",
  23770=>"011001100",
  23771=>"110110010",
  23772=>"111111111",
  23773=>"110001100",
  23774=>"111111110",
  23775=>"111110111",
  23776=>"000001111",
  23777=>"000111100",
  23778=>"110011111",
  23779=>"010110110",
  23780=>"100001101",
  23781=>"101001010",
  23782=>"101000100",
  23783=>"000000000",
  23784=>"100101111",
  23785=>"000110101",
  23786=>"000001000",
  23787=>"001000000",
  23788=>"000000001",
  23789=>"101000111",
  23790=>"111111000",
  23791=>"111001101",
  23792=>"011011011",
  23793=>"111010001",
  23794=>"001000000",
  23795=>"000001001",
  23796=>"011110110",
  23797=>"111111111",
  23798=>"010001101",
  23799=>"000000010",
  23800=>"100101111",
  23801=>"110110010",
  23802=>"111111111",
  23803=>"111111111",
  23804=>"000010010",
  23805=>"111011111",
  23806=>"110111011",
  23807=>"010010110",
  23808=>"011001100",
  23809=>"000000101",
  23810=>"000000101",
  23811=>"000000001",
  23812=>"101111000",
  23813=>"001100000",
  23814=>"000000001",
  23815=>"000000010",
  23816=>"001001101",
  23817=>"000001000",
  23818=>"000110001",
  23819=>"111111111",
  23820=>"001000000",
  23821=>"000111110",
  23822=>"101001001",
  23823=>"001110010",
  23824=>"101111110",
  23825=>"000000001",
  23826=>"000101111",
  23827=>"000000000",
  23828=>"000000111",
  23829=>"110010010",
  23830=>"110101011",
  23831=>"000101011",
  23832=>"000101111",
  23833=>"001100111",
  23834=>"000101111",
  23835=>"111111000",
  23836=>"000100101",
  23837=>"110110111",
  23838=>"111111000",
  23839=>"111000010",
  23840=>"000000101",
  23841=>"111110110",
  23842=>"000000000",
  23843=>"000000000",
  23844=>"110000000",
  23845=>"100110111",
  23846=>"111101000",
  23847=>"001111111",
  23848=>"010110100",
  23849=>"111111111",
  23850=>"001011111",
  23851=>"010000010",
  23852=>"111111110",
  23853=>"000101111",
  23854=>"000111111",
  23855=>"001000001",
  23856=>"000000111",
  23857=>"010011011",
  23858=>"111011101",
  23859=>"111111111",
  23860=>"111111011",
  23861=>"110010000",
  23862=>"011011000",
  23863=>"101000111",
  23864=>"111000000",
  23865=>"111000000",
  23866=>"000000000",
  23867=>"000000100",
  23868=>"010111000",
  23869=>"011011000",
  23870=>"100000000",
  23871=>"000000000",
  23872=>"111111000",
  23873=>"100111101",
  23874=>"111101011",
  23875=>"100100100",
  23876=>"010000000",
  23877=>"000111111",
  23878=>"101001001",
  23879=>"111110010",
  23880=>"011111111",
  23881=>"001111110",
  23882=>"101000110",
  23883=>"000000111",
  23884=>"001000001",
  23885=>"100100000",
  23886=>"000111100",
  23887=>"111011000",
  23888=>"111000000",
  23889=>"000111011",
  23890=>"000000000",
  23891=>"001001000",
  23892=>"000000000",
  23893=>"111111111",
  23894=>"011001001",
  23895=>"000010111",
  23896=>"010001110",
  23897=>"011011000",
  23898=>"111000001",
  23899=>"100010100",
  23900=>"111000000",
  23901=>"001001001",
  23902=>"111111011",
  23903=>"011011001",
  23904=>"101000000",
  23905=>"001010000",
  23906=>"000000101",
  23907=>"101100101",
  23908=>"111111110",
  23909=>"110100111",
  23910=>"000110101",
  23911=>"010000111",
  23912=>"111101000",
  23913=>"000000000",
  23914=>"111011000",
  23915=>"111111001",
  23916=>"000010011",
  23917=>"011010110",
  23918=>"000000000",
  23919=>"100101111",
  23920=>"111111011",
  23921=>"010110111",
  23922=>"110110000",
  23923=>"000000011",
  23924=>"000010000",
  23925=>"000101000",
  23926=>"111111111",
  23927=>"000000000",
  23928=>"010010000",
  23929=>"010000001",
  23930=>"101111111",
  23931=>"000000001",
  23932=>"100110011",
  23933=>"100100000",
  23934=>"010111100",
  23935=>"010010111",
  23936=>"000001011",
  23937=>"000100000",
  23938=>"100010111",
  23939=>"111100100",
  23940=>"000100000",
  23941=>"101001100",
  23942=>"100011001",
  23943=>"001000000",
  23944=>"101111101",
  23945=>"010010111",
  23946=>"101100111",
  23947=>"110101101",
  23948=>"111000000",
  23949=>"111011111",
  23950=>"100001111",
  23951=>"000000000",
  23952=>"111011111",
  23953=>"111011000",
  23954=>"001000010",
  23955=>"101010000",
  23956=>"101101000",
  23957=>"001111011",
  23958=>"111111111",
  23959=>"001011111",
  23960=>"111110011",
  23961=>"010010111",
  23962=>"101000000",
  23963=>"101100011",
  23964=>"000000000",
  23965=>"111101111",
  23966=>"101111111",
  23967=>"000001000",
  23968=>"110111111",
  23969=>"111101111",
  23970=>"110111111",
  23971=>"000000010",
  23972=>"100001000",
  23973=>"110000000",
  23974=>"010110010",
  23975=>"111111111",
  23976=>"000110111",
  23977=>"010110111",
  23978=>"111001000",
  23979=>"111110010",
  23980=>"010000010",
  23981=>"010000000",
  23982=>"111111110",
  23983=>"011000001",
  23984=>"000000000",
  23985=>"110001111",
  23986=>"111111000",
  23987=>"101110110",
  23988=>"011011110",
  23989=>"100100101",
  23990=>"101000000",
  23991=>"110110101",
  23992=>"001001001",
  23993=>"111101001",
  23994=>"000110111",
  23995=>"000011111",
  23996=>"010010010",
  23997=>"111111011",
  23998=>"000001001",
  23999=>"000000010",
  24000=>"000000001",
  24001=>"000000000",
  24002=>"110100010",
  24003=>"111001001",
  24004=>"000000111",
  24005=>"100100101",
  24006=>"000001111",
  24007=>"111000000",
  24008=>"011101100",
  24009=>"010000000",
  24010=>"000000000",
  24011=>"000000110",
  24012=>"111111110",
  24013=>"011011111",
  24014=>"000000000",
  24015=>"000000000",
  24016=>"101000111",
  24017=>"100111111",
  24018=>"000011010",
  24019=>"111110110",
  24020=>"101001111",
  24021=>"100100110",
  24022=>"110110000",
  24023=>"001000111",
  24024=>"000010110",
  24025=>"000111111",
  24026=>"111111100",
  24027=>"000101101",
  24028=>"111110110",
  24029=>"000001001",
  24030=>"111110010",
  24031=>"000111010",
  24032=>"000000000",
  24033=>"100000011",
  24034=>"110110010",
  24035=>"000100110",
  24036=>"001000000",
  24037=>"000110110",
  24038=>"101101111",
  24039=>"101101101",
  24040=>"111111000",
  24041=>"000001111",
  24042=>"000011001",
  24043=>"101000000",
  24044=>"110111000",
  24045=>"000000000",
  24046=>"000010000",
  24047=>"111100000",
  24048=>"111111110",
  24049=>"100001001",
  24050=>"000001000",
  24051=>"100100100",
  24052=>"110101001",
  24053=>"010010111",
  24054=>"000000000",
  24055=>"101000000",
  24056=>"010110111",
  24057=>"111000010",
  24058=>"110010000",
  24059=>"000000000",
  24060=>"111101000",
  24061=>"000000000",
  24062=>"011101000",
  24063=>"000000000",
  24064=>"010000111",
  24065=>"110110111",
  24066=>"100100101",
  24067=>"111000111",
  24068=>"100000100",
  24069=>"001101100",
  24070=>"101100101",
  24071=>"000000111",
  24072=>"111010000",
  24073=>"000000100",
  24074=>"110110111",
  24075=>"111100000",
  24076=>"001000111",
  24077=>"010010000",
  24078=>"000000000",
  24079=>"000000000",
  24080=>"000000000",
  24081=>"110100000",
  24082=>"011000000",
  24083=>"100001000",
  24084=>"011111111",
  24085=>"011111111",
  24086=>"001111011",
  24087=>"000111111",
  24088=>"101100111",
  24089=>"111111101",
  24090=>"111011000",
  24091=>"100101000",
  24092=>"010011010",
  24093=>"011010000",
  24094=>"110111111",
  24095=>"011111000",
  24096=>"111101111",
  24097=>"100011110",
  24098=>"000111111",
  24099=>"001011011",
  24100=>"011100000",
  24101=>"110010010",
  24102=>"011011010",
  24103=>"000000111",
  24104=>"110000011",
  24105=>"000000001",
  24106=>"110101100",
  24107=>"000000000",
  24108=>"111111011",
  24109=>"011000000",
  24110=>"010001111",
  24111=>"011100100",
  24112=>"001111000",
  24113=>"000000100",
  24114=>"000000010",
  24115=>"111000011",
  24116=>"000010000",
  24117=>"111110000",
  24118=>"001010000",
  24119=>"000000101",
  24120=>"000000111",
  24121=>"111101000",
  24122=>"010111010",
  24123=>"111111011",
  24124=>"011011111",
  24125=>"000011011",
  24126=>"000000000",
  24127=>"000000000",
  24128=>"101001000",
  24129=>"000111101",
  24130=>"000111010",
  24131=>"000100000",
  24132=>"111111001",
  24133=>"000100100",
  24134=>"111101011",
  24135=>"100111011",
  24136=>"010010110",
  24137=>"011101101",
  24138=>"100100001",
  24139=>"101100000",
  24140=>"000000000",
  24141=>"011000000",
  24142=>"110100001",
  24143=>"010110011",
  24144=>"000010000",
  24145=>"111111111",
  24146=>"011111000",
  24147=>"001001001",
  24148=>"011010000",
  24149=>"011011110",
  24150=>"001100011",
  24151=>"001010011",
  24152=>"111111111",
  24153=>"010011111",
  24154=>"101001000",
  24155=>"000000000",
  24156=>"000000000",
  24157=>"011001010",
  24158=>"111000101",
  24159=>"001001101",
  24160=>"111101000",
  24161=>"001000011",
  24162=>"111000011",
  24163=>"100110100",
  24164=>"111000000",
  24165=>"100011111",
  24166=>"100011001",
  24167=>"011000101",
  24168=>"101011111",
  24169=>"101111111",
  24170=>"001000111",
  24171=>"111101000",
  24172=>"111000001",
  24173=>"111101000",
  24174=>"100110110",
  24175=>"000101101",
  24176=>"101000100",
  24177=>"100100101",
  24178=>"111011000",
  24179=>"101000000",
  24180=>"101101000",
  24181=>"111000010",
  24182=>"111100000",
  24183=>"010010010",
  24184=>"001111010",
  24185=>"000011111",
  24186=>"111101110",
  24187=>"010000111",
  24188=>"100100010",
  24189=>"011110110",
  24190=>"100000111",
  24191=>"100110000",
  24192=>"111000000",
  24193=>"100100110",
  24194=>"000000110",
  24195=>"001000111",
  24196=>"011101001",
  24197=>"100000010",
  24198=>"000011001",
  24199=>"010010000",
  24200=>"100000100",
  24201=>"000010000",
  24202=>"111111000",
  24203=>"111100111",
  24204=>"101101100",
  24205=>"111101101",
  24206=>"000101111",
  24207=>"111000000",
  24208=>"010000000",
  24209=>"100100000",
  24210=>"100000010",
  24211=>"111111000",
  24212=>"011010000",
  24213=>"100100000",
  24214=>"111110101",
  24215=>"011000000",
  24216=>"111101000",
  24217=>"000011010",
  24218=>"110111111",
  24219=>"000000100",
  24220=>"000000000",
  24221=>"111101111",
  24222=>"000000000",
  24223=>"000100000",
  24224=>"000011101",
  24225=>"001111111",
  24226=>"011000000",
  24227=>"000111111",
  24228=>"101011110",
  24229=>"100001000",
  24230=>"010001011",
  24231=>"000000000",
  24232=>"010000110",
  24233=>"111010000",
  24234=>"110101001",
  24235=>"010111101",
  24236=>"000110110",
  24237=>"100000100",
  24238=>"010110101",
  24239=>"000000001",
  24240=>"010000000",
  24241=>"111111001",
  24242=>"111100000",
  24243=>"001000001",
  24244=>"000101000",
  24245=>"010111011",
  24246=>"111011100",
  24247=>"000111111",
  24248=>"001011011",
  24249=>"100010011",
  24250=>"111011111",
  24251=>"100101110",
  24252=>"111000010",
  24253=>"111100111",
  24254=>"110100010",
  24255=>"000000000",
  24256=>"011011000",
  24257=>"110101000",
  24258=>"100000000",
  24259=>"111000100",
  24260=>"101111101",
  24261=>"001100111",
  24262=>"111101101",
  24263=>"000011110",
  24264=>"010000101",
  24265=>"000011111",
  24266=>"000101111",
  24267=>"101101111",
  24268=>"010000000",
  24269=>"110010000",
  24270=>"110111111",
  24271=>"111000101",
  24272=>"111011001",
  24273=>"010100101",
  24274=>"111000011",
  24275=>"000101000",
  24276=>"101101101",
  24277=>"011110000",
  24278=>"111111000",
  24279=>"111111000",
  24280=>"000011000",
  24281=>"010000000",
  24282=>"000111110",
  24283=>"101100100",
  24284=>"110111110",
  24285=>"110010010",
  24286=>"111100000",
  24287=>"000101100",
  24288=>"000111001",
  24289=>"111101111",
  24290=>"011010111",
  24291=>"011001100",
  24292=>"100000000",
  24293=>"111101101",
  24294=>"110000000",
  24295=>"000010101",
  24296=>"111100000",
  24297=>"000000000",
  24298=>"001111110",
  24299=>"011111111",
  24300=>"000000111",
  24301=>"011000000",
  24302=>"000000010",
  24303=>"110111010",
  24304=>"111111010",
  24305=>"000110001",
  24306=>"100101111",
  24307=>"010110110",
  24308=>"011101110",
  24309=>"001111101",
  24310=>"100000000",
  24311=>"000000000",
  24312=>"000100011",
  24313=>"000001010",
  24314=>"000011111",
  24315=>"101111010",
  24316=>"101101000",
  24317=>"010110010",
  24318=>"100000000",
  24319=>"111100111",
  24320=>"011001011",
  24321=>"111110011",
  24322=>"000100100",
  24323=>"000000011",
  24324=>"100011001",
  24325=>"010110100",
  24326=>"111011011",
  24327=>"111001011",
  24328=>"100110100",
  24329=>"000000000",
  24330=>"000111111",
  24331=>"011101110",
  24332=>"000000000",
  24333=>"000000000",
  24334=>"100100111",
  24335=>"110010010",
  24336=>"100000001",
  24337=>"101111100",
  24338=>"010000000",
  24339=>"100110011",
  24340=>"101111000",
  24341=>"101111101",
  24342=>"000101111",
  24343=>"100000111",
  24344=>"000000000",
  24345=>"011111011",
  24346=>"000011010",
  24347=>"111100100",
  24348=>"101100011",
  24349=>"111010001",
  24350=>"111111010",
  24351=>"000111110",
  24352=>"000100101",
  24353=>"110110111",
  24354=>"000001000",
  24355=>"000000000",
  24356=>"001000000",
  24357=>"100000011",
  24358=>"111011011",
  24359=>"000100000",
  24360=>"100111101",
  24361=>"001010111",
  24362=>"000000011",
  24363=>"001000010",
  24364=>"110001011",
  24365=>"011110111",
  24366=>"110110100",
  24367=>"000101100",
  24368=>"000001011",
  24369=>"011010110",
  24370=>"111100000",
  24371=>"000111011",
  24372=>"101111111",
  24373=>"000011011",
  24374=>"111011111",
  24375=>"000001000",
  24376=>"010010000",
  24377=>"111100110",
  24378=>"011000000",
  24379=>"000011000",
  24380=>"111001000",
  24381=>"111111110",
  24382=>"101100100",
  24383=>"110111111",
  24384=>"111111011",
  24385=>"000100110",
  24386=>"110000001",
  24387=>"001111011",
  24388=>"000000001",
  24389=>"011000000",
  24390=>"001011011",
  24391=>"011011111",
  24392=>"111110100",
  24393=>"100000011",
  24394=>"000100100",
  24395=>"000100000",
  24396=>"100100100",
  24397=>"111111101",
  24398=>"001111111",
  24399=>"000011111",
  24400=>"000000000",
  24401=>"111100100",
  24402=>"000101011",
  24403=>"000001011",
  24404=>"100100100",
  24405=>"111110010",
  24406=>"000100110",
  24407=>"101000000",
  24408=>"000000000",
  24409=>"000000001",
  24410=>"000000011",
  24411=>"110110111",
  24412=>"000000000",
  24413=>"011000010",
  24414=>"000011111",
  24415=>"110110001",
  24416=>"000011011",
  24417=>"000000001",
  24418=>"000000100",
  24419=>"001000001",
  24420=>"110110011",
  24421=>"110110111",
  24422=>"100100010",
  24423=>"110100000",
  24424=>"011111011",
  24425=>"011011111",
  24426=>"011010000",
  24427=>"100101111",
  24428=>"100100110",
  24429=>"001011101",
  24430=>"110110100",
  24431=>"000000000",
  24432=>"000000000",
  24433=>"111000000",
  24434=>"011111111",
  24435=>"111100100",
  24436=>"000000000",
  24437=>"100100100",
  24438=>"001011000",
  24439=>"000011011",
  24440=>"000010001",
  24441=>"100000011",
  24442=>"011100110",
  24443=>"000000001",
  24444=>"001100000",
  24445=>"000000000",
  24446=>"111100111",
  24447=>"111100100",
  24448=>"100000011",
  24449=>"011011100",
  24450=>"000001000",
  24451=>"000001010",
  24452=>"100110111",
  24453=>"100111111",
  24454=>"010110110",
  24455=>"010000000",
  24456=>"110111101",
  24457=>"000001000",
  24458=>"110000010",
  24459=>"011000000",
  24460=>"000000000",
  24461=>"100111000",
  24462=>"000001011",
  24463=>"000000000",
  24464=>"000000000",
  24465=>"000100111",
  24466=>"001100100",
  24467=>"111100101",
  24468=>"110111100",
  24469=>"111101000",
  24470=>"000011110",
  24471=>"110011011",
  24472=>"000111011",
  24473=>"111100001",
  24474=>"100100101",
  24475=>"000010011",
  24476=>"000000000",
  24477=>"110111011",
  24478=>"000001011",
  24479=>"100100111",
  24480=>"000100000",
  24481=>"100110000",
  24482=>"010011001",
  24483=>"100011011",
  24484=>"101100100",
  24485=>"100010011",
  24486=>"110010011",
  24487=>"010011011",
  24488=>"011100000",
  24489=>"001011111",
  24490=>"000110111",
  24491=>"100110111",
  24492=>"010011100",
  24493=>"010100001",
  24494=>"100100100",
  24495=>"011011011",
  24496=>"010100100",
  24497=>"001100100",
  24498=>"100010111",
  24499=>"001100000",
  24500=>"000001001",
  24501=>"011011000",
  24502=>"000001011",
  24503=>"000000000",
  24504=>"010010000",
  24505=>"010010111",
  24506=>"001001111",
  24507=>"000001011",
  24508=>"111001000",
  24509=>"011111110",
  24510=>"000001000",
  24511=>"011001000",
  24512=>"011111111",
  24513=>"000011011",
  24514=>"000011011",
  24515=>"100100110",
  24516=>"010100000",
  24517=>"011010110",
  24518=>"000000010",
  24519=>"111111000",
  24520=>"100000011",
  24521=>"110001010",
  24522=>"000011011",
  24523=>"111111111",
  24524=>"100011010",
  24525=>"100111110",
  24526=>"011011000",
  24527=>"100110110",
  24528=>"000100110",
  24529=>"001111111",
  24530=>"001000100",
  24531=>"000111011",
  24532=>"000100100",
  24533=>"011010000",
  24534=>"011100110",
  24535=>"110010111",
  24536=>"011000101",
  24537=>"010000000",
  24538=>"100111111",
  24539=>"110100000",
  24540=>"101111111",
  24541=>"011011110",
  24542=>"000011011",
  24543=>"100110011",
  24544=>"000000000",
  24545=>"111110000",
  24546=>"101111110",
  24547=>"000000101",
  24548=>"111100100",
  24549=>"000111101",
  24550=>"111110000",
  24551=>"011111000",
  24552=>"111100100",
  24553=>"011100100",
  24554=>"111001101",
  24555=>"000011011",
  24556=>"000000000",
  24557=>"011100100",
  24558=>"011000000",
  24559=>"100100000",
  24560=>"111100100",
  24561=>"101001100",
  24562=>"011000000",
  24563=>"101110111",
  24564=>"010011010",
  24565=>"010000100",
  24566=>"001000001",
  24567=>"110110100",
  24568=>"000001111",
  24569=>"110010011",
  24570=>"001001001",
  24571=>"011011111",
  24572=>"111000111",
  24573=>"110100100",
  24574=>"000011011",
  24575=>"100111011",
  24576=>"001000000",
  24577=>"000001101",
  24578=>"101000101",
  24579=>"011000011",
  24580=>"000011111",
  24581=>"111101101",
  24582=>"111000101",
  24583=>"111011101",
  24584=>"011000000",
  24585=>"100000100",
  24586=>"100111001",
  24587=>"110010010",
  24588=>"011001011",
  24589=>"111111000",
  24590=>"100111100",
  24591=>"011010000",
  24592=>"000100111",
  24593=>"101101001",
  24594=>"000001110",
  24595=>"101000001",
  24596=>"111111111",
  24597=>"000111000",
  24598=>"110000111",
  24599=>"111111110",
  24600=>"000000100",
  24601=>"001000100",
  24602=>"110111011",
  24603=>"000111111",
  24604=>"000000101",
  24605=>"000000101",
  24606=>"111100111",
  24607=>"000000000",
  24608=>"001000011",
  24609=>"101111010",
  24610=>"100101001",
  24611=>"101000101",
  24612=>"001111111",
  24613=>"100001000",
  24614=>"010000000",
  24615=>"000111101",
  24616=>"100010100",
  24617=>"001001001",
  24618=>"010111011",
  24619=>"001000111",
  24620=>"000111110",
  24621=>"111110011",
  24622=>"111001100",
  24623=>"001000000",
  24624=>"000101000",
  24625=>"111010000",
  24626=>"000000000",
  24627=>"100000100",
  24628=>"111011000",
  24629=>"101111001",
  24630=>"101101100",
  24631=>"111111000",
  24632=>"111010010",
  24633=>"101111111",
  24634=>"000010010",
  24635=>"000111000",
  24636=>"011111011",
  24637=>"000000001",
  24638=>"000000101",
  24639=>"011111011",
  24640=>"101101101",
  24641=>"000000101",
  24642=>"000000000",
  24643=>"011011001",
  24644=>"111111010",
  24645=>"001000000",
  24646=>"011010000",
  24647=>"000010011",
  24648=>"111111111",
  24649=>"010111010",
  24650=>"010001001",
  24651=>"010001000",
  24652=>"111000000",
  24653=>"111111011",
  24654=>"001000111",
  24655=>"000111111",
  24656=>"000000000",
  24657=>"111111111",
  24658=>"111111000",
  24659=>"011001000",
  24660=>"101101000",
  24661=>"001011110",
  24662=>"001100011",
  24663=>"111101101",
  24664=>"000000011",
  24665=>"000011010",
  24666=>"100011010",
  24667=>"000100100",
  24668=>"000101101",
  24669=>"000100110",
  24670=>"011000010",
  24671=>"110110101",
  24672=>"000000100",
  24673=>"001010000",
  24674=>"111001111",
  24675=>"000111010",
  24676=>"000001010",
  24677=>"011010000",
  24678=>"010110111",
  24679=>"111111010",
  24680=>"010011001",
  24681=>"010010110",
  24682=>"110000110",
  24683=>"111111111",
  24684=>"000000111",
  24685=>"001111110",
  24686=>"001001000",
  24687=>"010101110",
  24688=>"001110000",
  24689=>"000010110",
  24690=>"101101001",
  24691=>"000000000",
  24692=>"111100000",
  24693=>"010000000",
  24694=>"000011111",
  24695=>"111000100",
  24696=>"000000111",
  24697=>"000111011",
  24698=>"100111000",
  24699=>"010111111",
  24700=>"001001101",
  24701=>"010100000",
  24702=>"000111000",
  24703=>"000111000",
  24704=>"110111001",
  24705=>"010000010",
  24706=>"000111101",
  24707=>"000000100",
  24708=>"111111111",
  24709=>"111110001",
  24710=>"001000011",
  24711=>"000001100",
  24712=>"100011010",
  24713=>"001000000",
  24714=>"011111010",
  24715=>"000010111",
  24716=>"100001101",
  24717=>"001101101",
  24718=>"101010111",
  24719=>"000000000",
  24720=>"111111000",
  24721=>"001111000",
  24722=>"111110000",
  24723=>"100000111",
  24724=>"101000011",
  24725=>"101000101",
  24726=>"000010111",
  24727=>"010000100",
  24728=>"000011000",
  24729=>"100000001",
  24730=>"111111000",
  24731=>"000000111",
  24732=>"111111110",
  24733=>"100000110",
  24734=>"110010011",
  24735=>"101000110",
  24736=>"100010001",
  24737=>"111101101",
  24738=>"000000010",
  24739=>"010111010",
  24740=>"010110011",
  24741=>"101000000",
  24742=>"010001100",
  24743=>"101111101",
  24744=>"100100100",
  24745=>"110111001",
  24746=>"111000001",
  24747=>"111101101",
  24748=>"001101011",
  24749=>"110000000",
  24750=>"000000000",
  24751=>"111000010",
  24752=>"100000101",
  24753=>"001000111",
  24754=>"000010000",
  24755=>"001001011",
  24756=>"111111011",
  24757=>"000001001",
  24758=>"000000000",
  24759=>"101110010",
  24760=>"100111110",
  24761=>"000000110",
  24762=>"111000000",
  24763=>"011000111",
  24764=>"000000000",
  24765=>"111111100",
  24766=>"110011000",
  24767=>"000000000",
  24768=>"111000000",
  24769=>"000001001",
  24770=>"111110001",
  24771=>"111010000",
  24772=>"001111000",
  24773=>"111001101",
  24774=>"011000010",
  24775=>"001001101",
  24776=>"110110000",
  24777=>"010100000",
  24778=>"000000001",
  24779=>"001000000",
  24780=>"000001000",
  24781=>"000100101",
  24782=>"000000101",
  24783=>"000001111",
  24784=>"000110000",
  24785=>"111110100",
  24786=>"100110111",
  24787=>"010011000",
  24788=>"101001111",
  24789=>"100000011",
  24790=>"010011111",
  24791=>"010010111",
  24792=>"001011001",
  24793=>"000000010",
  24794=>"000000000",
  24795=>"000010000",
  24796=>"010101011",
  24797=>"110111110",
  24798=>"000000010",
  24799=>"101110010",
  24800=>"111000000",
  24801=>"111100001",
  24802=>"100110001",
  24803=>"001111111",
  24804=>"000000000",
  24805=>"111111001",
  24806=>"001011111",
  24807=>"001001000",
  24808=>"000010111",
  24809=>"101011111",
  24810=>"001111100",
  24811=>"000000001",
  24812=>"000000000",
  24813=>"000010010",
  24814=>"000000000",
  24815=>"010101111",
  24816=>"111110000",
  24817=>"111110000",
  24818=>"111101111",
  24819=>"111110110",
  24820=>"000111011",
  24821=>"000000000",
  24822=>"000000100",
  24823=>"100111001",
  24824=>"011001011",
  24825=>"011011000",
  24826=>"000011000",
  24827=>"000101101",
  24828=>"010000101",
  24829=>"000001000",
  24830=>"101111110",
  24831=>"011010001",
  24832=>"011101111",
  24833=>"001000000",
  24834=>"000000000",
  24835=>"000100110",
  24836=>"111011001",
  24837=>"000001111",
  24838=>"101100000",
  24839=>"111111010",
  24840=>"001001111",
  24841=>"000001000",
  24842=>"011100100",
  24843=>"000000000",
  24844=>"000000111",
  24845=>"000000100",
  24846=>"110111111",
  24847=>"101111101",
  24848=>"100111111",
  24849=>"000000111",
  24850=>"111111000",
  24851=>"000000000",
  24852=>"110110000",
  24853=>"100000010",
  24854=>"101111111",
  24855=>"111111011",
  24856=>"000001001",
  24857=>"000000111",
  24858=>"000000111",
  24859=>"000000001",
  24860=>"101111101",
  24861=>"000011111",
  24862=>"111111111",
  24863=>"000110110",
  24864=>"000000010",
  24865=>"000000000",
  24866=>"111011100",
  24867=>"000000000",
  24868=>"111001001",
  24869=>"101001001",
  24870=>"000000001",
  24871=>"111011100",
  24872=>"111010000",
  24873=>"000001010",
  24874=>"111001111",
  24875=>"111111111",
  24876=>"001101111",
  24877=>"011000000",
  24878=>"111111101",
  24879=>"110111111",
  24880=>"000000000",
  24881=>"111111011",
  24882=>"000000001",
  24883=>"101111100",
  24884=>"000111110",
  24885=>"111110111",
  24886=>"000000010",
  24887=>"011011111",
  24888=>"111111001",
  24889=>"010001000",
  24890=>"000000111",
  24891=>"100000010",
  24892=>"001001001",
  24893=>"111111111",
  24894=>"000000111",
  24895=>"111001001",
  24896=>"010001000",
  24897=>"010000000",
  24898=>"000111111",
  24899=>"111110110",
  24900=>"110000000",
  24901=>"101111100",
  24902=>"111110110",
  24903=>"010100100",
  24904=>"010101101",
  24905=>"111101101",
  24906=>"111101111",
  24907=>"000101111",
  24908=>"000001000",
  24909=>"111111010",
  24910=>"100110110",
  24911=>"100000110",
  24912=>"000100111",
  24913=>"111111000",
  24914=>"000000111",
  24915=>"001000000",
  24916=>"111000000",
  24917=>"000100100",
  24918=>"001011110",
  24919=>"000000010",
  24920=>"011000111",
  24921=>"001001001",
  24922=>"110000011",
  24923=>"000100111",
  24924=>"001001111",
  24925=>"101000001",
  24926=>"111111000",
  24927=>"111101110",
  24928=>"111111111",
  24929=>"000100110",
  24930=>"000000000",
  24931=>"111010000",
  24932=>"100000100",
  24933=>"000000000",
  24934=>"000101001",
  24935=>"111011010",
  24936=>"010000000",
  24937=>"100001101",
  24938=>"111000000",
  24939=>"000000000",
  24940=>"000111011",
  24941=>"000000000",
  24942=>"000000000",
  24943=>"000000101",
  24944=>"100000110",
  24945=>"000000111",
  24946=>"010000000",
  24947=>"000101111",
  24948=>"100101101",
  24949=>"000101101",
  24950=>"000000000",
  24951=>"110101100",
  24952=>"111100000",
  24953=>"000001111",
  24954=>"011000001",
  24955=>"111110000",
  24956=>"110110100",
  24957=>"100000001",
  24958=>"111111010",
  24959=>"000000111",
  24960=>"000001000",
  24961=>"111111111",
  24962=>"110111111",
  24963=>"001011100",
  24964=>"100110110",
  24965=>"101100011",
  24966=>"000000100",
  24967=>"000000000",
  24968=>"011001011",
  24969=>"110111111",
  24970=>"111111011",
  24971=>"000000100",
  24972=>"000000000",
  24973=>"001101110",
  24974=>"011110000",
  24975=>"000000000",
  24976=>"011011001",
  24977=>"111000100",
  24978=>"000001000",
  24979=>"111110010",
  24980=>"000111111",
  24981=>"000000100",
  24982=>"111111111",
  24983=>"001001011",
  24984=>"000001110",
  24985=>"111111100",
  24986=>"011111000",
  24987=>"000110000",
  24988=>"100000000",
  24989=>"000000001",
  24990=>"101110110",
  24991=>"101111111",
  24992=>"001000001",
  24993=>"101110111",
  24994=>"111001111",
  24995=>"000100000",
  24996=>"101111011",
  24997=>"001001101",
  24998=>"100100111",
  24999=>"111111111",
  25000=>"000111111",
  25001=>"011110000",
  25002=>"000000000",
  25003=>"001000000",
  25004=>"011010001",
  25005=>"000000001",
  25006=>"011010110",
  25007=>"011010000",
  25008=>"111000000",
  25009=>"101000101",
  25010=>"000100110",
  25011=>"000000100",
  25012=>"011111101",
  25013=>"111111111",
  25014=>"010000000",
  25015=>"000000000",
  25016=>"110000101",
  25017=>"001010010",
  25018=>"001000101",
  25019=>"011010100",
  25020=>"000010000",
  25021=>"000101000",
  25022=>"101100100",
  25023=>"000101111",
  25024=>"111010010",
  25025=>"011001111",
  25026=>"000111010",
  25027=>"001001001",
  25028=>"000111000",
  25029=>"000000000",
  25030=>"011101111",
  25031=>"110111111",
  25032=>"111110000",
  25033=>"010001001",
  25034=>"110000000",
  25035=>"000000000",
  25036=>"011111010",
  25037=>"111011011",
  25038=>"000000000",
  25039=>"000001011",
  25040=>"000111111",
  25041=>"110111111",
  25042=>"000000000",
  25043=>"101111111",
  25044=>"000000000",
  25045=>"001001001",
  25046=>"101000001",
  25047=>"000111011",
  25048=>"111111110",
  25049=>"011111010",
  25050=>"100000110",
  25051=>"000001000",
  25052=>"010111101",
  25053=>"000000100",
  25054=>"000010110",
  25055=>"001101111",
  25056=>"000000000",
  25057=>"000000000",
  25058=>"111000000",
  25059=>"100111111",
  25060=>"001001011",
  25061=>"100001100",
  25062=>"000000000",
  25063=>"111100100",
  25064=>"000000111",
  25065=>"000000010",
  25066=>"110001001",
  25067=>"000000100",
  25068=>"000000000",
  25069=>"000000000",
  25070=>"000000001",
  25071=>"001000000",
  25072=>"000100111",
  25073=>"000000100",
  25074=>"001101100",
  25075=>"111111111",
  25076=>"100101001",
  25077=>"110111101",
  25078=>"000000100",
  25079=>"000001011",
  25080=>"111110010",
  25081=>"000110100",
  25082=>"111111111",
  25083=>"000010010",
  25084=>"111111010",
  25085=>"000000000",
  25086=>"110110110",
  25087=>"111111111",
  25088=>"110010111",
  25089=>"011110110",
  25090=>"001001111",
  25091=>"000010111",
  25092=>"010011110",
  25093=>"000011011",
  25094=>"100110100",
  25095=>"100110001",
  25096=>"010000001",
  25097=>"011000011",
  25098=>"110101001",
  25099=>"111111011",
  25100=>"011001011",
  25101=>"001001001",
  25102=>"100010000",
  25103=>"101100000",
  25104=>"100100001",
  25105=>"000100100",
  25106=>"001001000",
  25107=>"001100100",
  25108=>"110110100",
  25109=>"011011011",
  25110=>"110000110",
  25111=>"001100101",
  25112=>"100000001",
  25113=>"101001001",
  25114=>"001000110",
  25115=>"000100110",
  25116=>"111101110",
  25117=>"011011011",
  25118=>"100000011",
  25119=>"001001000",
  25120=>"001001101",
  25121=>"100101101",
  25122=>"111001011",
  25123=>"001011001",
  25124=>"010000000",
  25125=>"111101100",
  25126=>"111110010",
  25127=>"000100001",
  25128=>"010111111",
  25129=>"100110001",
  25130=>"110100100",
  25131=>"000001111",
  25132=>"111111110",
  25133=>"110110101",
  25134=>"010000110",
  25135=>"001001000",
  25136=>"100100000",
  25137=>"010011110",
  25138=>"000000000",
  25139=>"101101000",
  25140=>"000000001",
  25141=>"110111110",
  25142=>"011011000",
  25143=>"110011000",
  25144=>"000111011",
  25145=>"110000011",
  25146=>"001001110",
  25147=>"000100100",
  25148=>"011010010",
  25149=>"111011111",
  25150=>"001001001",
  25151=>"000110000",
  25152=>"101101011",
  25153=>"001010111",
  25154=>"011001000",
  25155=>"001011101",
  25156=>"010011010",
  25157=>"000000100",
  25158=>"000000100",
  25159=>"011111011",
  25160=>"111111011",
  25161=>"110100110",
  25162=>"100100000",
  25163=>"011000001",
  25164=>"001000100",
  25165=>"111011001",
  25166=>"111000101",
  25167=>"101111100",
  25168=>"010000100",
  25169=>"000011011",
  25170=>"001100101",
  25171=>"101111000",
  25172=>"100100010",
  25173=>"000000000",
  25174=>"100000010",
  25175=>"101001111",
  25176=>"110110111",
  25177=>"110111001",
  25178=>"100101111",
  25179=>"011001000",
  25180=>"101101101",
  25181=>"010011100",
  25182=>"001111111",
  25183=>"010000011",
  25184=>"011011011",
  25185=>"010001000",
  25186=>"001001001",
  25187=>"000010000",
  25188=>"000001010",
  25189=>"011011001",
  25190=>"111110101",
  25191=>"111011011",
  25192=>"100101011",
  25193=>"101101111",
  25194=>"100000100",
  25195=>"110011001",
  25196=>"011001110",
  25197=>"110100100",
  25198=>"101000011",
  25199=>"001111100",
  25200=>"010000001",
  25201=>"100000000",
  25202=>"000001001",
  25203=>"000011000",
  25204=>"001001001",
  25205=>"000001010",
  25206=>"001001010",
  25207=>"000011000",
  25208=>"110111110",
  25209=>"000000110",
  25210=>"100100101",
  25211=>"000010000",
  25212=>"101011011",
  25213=>"001001000",
  25214=>"000100011",
  25215=>"011011001",
  25216=>"001101100",
  25217=>"010010001",
  25218=>"011001101",
  25219=>"010011111",
  25220=>"101101101",
  25221=>"011011111",
  25222=>"100111110",
  25223=>"100111001",
  25224=>"000000001",
  25225=>"011000000",
  25226=>"001100000",
  25227=>"000000100",
  25228=>"001110001",
  25229=>"010011111",
  25230=>"000110100",
  25231=>"111001000",
  25232=>"110011011",
  25233=>"100011110",
  25234=>"001100000",
  25235=>"111011001",
  25236=>"111110100",
  25237=>"001000100",
  25238=>"110110100",
  25239=>"000010000",
  25240=>"111111011",
  25241=>"011100110",
  25242=>"011011001",
  25243=>"001011011",
  25244=>"111111001",
  25245=>"000000001",
  25246=>"100100111",
  25247=>"011101111",
  25248=>"111100001",
  25249=>"100100001",
  25250=>"000010110",
  25251=>"001011010",
  25252=>"100100101",
  25253=>"100000000",
  25254=>"100001001",
  25255=>"111110111",
  25256=>"011100100",
  25257=>"100100000",
  25258=>"001001111",
  25259=>"001001001",
  25260=>"001001100",
  25261=>"000001001",
  25262=>"111111000",
  25263=>"101011001",
  25264=>"001000000",
  25265=>"110100011",
  25266=>"101011110",
  25267=>"101001001",
  25268=>"010110110",
  25269=>"011110110",
  25270=>"101001011",
  25271=>"100111110",
  25272=>"000000000",
  25273=>"000000000",
  25274=>"000011011",
  25275=>"110111100",
  25276=>"101001111",
  25277=>"001001011",
  25278=>"001000000",
  25279=>"010010000",
  25280=>"011001100",
  25281=>"000100001",
  25282=>"100011100",
  25283=>"011010000",
  25284=>"100100100",
  25285=>"010001000",
  25286=>"001101100",
  25287=>"011011110",
  25288=>"100110000",
  25289=>"011000000",
  25290=>"011111011",
  25291=>"111110011",
  25292=>"110111001",
  25293=>"110010000",
  25294=>"000001011",
  25295=>"001111001",
  25296=>"101111001",
  25297=>"010111011",
  25298=>"111011001",
  25299=>"001000000",
  25300=>"001001001",
  25301=>"110110110",
  25302=>"100001001",
  25303=>"100100100",
  25304=>"100110100",
  25305=>"100001000",
  25306=>"011000000",
  25307=>"100101100",
  25308=>"000110000",
  25309=>"000010000",
  25310=>"110010000",
  25311=>"000001111",
  25312=>"110001000",
  25313=>"100001010",
  25314=>"100100110",
  25315=>"001000001",
  25316=>"011000100",
  25317=>"011111011",
  25318=>"111011011",
  25319=>"000111110",
  25320=>"111011111",
  25321=>"000110110",
  25322=>"000100110",
  25323=>"111100110",
  25324=>"011011001",
  25325=>"101101110",
  25326=>"000001110",
  25327=>"110000100",
  25328=>"110000100",
  25329=>"111111111",
  25330=>"100000100",
  25331=>"110110000",
  25332=>"011010001",
  25333=>"100111110",
  25334=>"000000100",
  25335=>"110010110",
  25336=>"100100001",
  25337=>"100011000",
  25338=>"011011111",
  25339=>"100010100",
  25340=>"011110100",
  25341=>"001010011",
  25342=>"110011111",
  25343=>"000001110",
  25344=>"000111000",
  25345=>"010000011",
  25346=>"101100001",
  25347=>"111111010",
  25348=>"100110100",
  25349=>"100000111",
  25350=>"111000100",
  25351=>"010000000",
  25352=>"110010000",
  25353=>"010000001",
  25354=>"111101100",
  25355=>"000111000",
  25356=>"101000101",
  25357=>"111111011",
  25358=>"000000000",
  25359=>"000000000",
  25360=>"011111111",
  25361=>"111110110",
  25362=>"101100111",
  25363=>"001000000",
  25364=>"100000111",
  25365=>"111101100",
  25366=>"111111100",
  25367=>"110110111",
  25368=>"000001111",
  25369=>"000001100",
  25370=>"000000000",
  25371=>"110111001",
  25372=>"111111011",
  25373=>"010000010",
  25374=>"101011000",
  25375=>"111111111",
  25376=>"111111000",
  25377=>"001000000",
  25378=>"000000110",
  25379=>"000000000",
  25380=>"000000000",
  25381=>"110100000",
  25382=>"000000000",
  25383=>"111111111",
  25384=>"111000111",
  25385=>"000010010",
  25386=>"111111111",
  25387=>"000111110",
  25388=>"111110111",
  25389=>"000000000",
  25390=>"000111111",
  25391=>"000100000",
  25392=>"000110000",
  25393=>"000111110",
  25394=>"000001111",
  25395=>"111110010",
  25396=>"101100111",
  25397=>"010111010",
  25398=>"011001110",
  25399=>"001001011",
  25400=>"111000000",
  25401=>"000000000",
  25402=>"100110111",
  25403=>"000000011",
  25404=>"100110110",
  25405=>"111111111",
  25406=>"000000000",
  25407=>"111111101",
  25408=>"011000001",
  25409=>"010110000",
  25410=>"000000000",
  25411=>"110101100",
  25412=>"000010000",
  25413=>"001001100",
  25414=>"101001000",
  25415=>"001000111",
  25416=>"000000000",
  25417=>"110111010",
  25418=>"001000000",
  25419=>"111110111",
  25420=>"000000000",
  25421=>"111001110",
  25422=>"000001001",
  25423=>"011010111",
  25424=>"111111111",
  25425=>"110110111",
  25426=>"000000000",
  25427=>"001001000",
  25428=>"111110110",
  25429=>"100011011",
  25430=>"001001000",
  25431=>"111111111",
  25432=>"000000111",
  25433=>"000001110",
  25434=>"001001000",
  25435=>"111111111",
  25436=>"000000000",
  25437=>"001100010",
  25438=>"001001000",
  25439=>"111111111",
  25440=>"111110110",
  25441=>"111010010",
  25442=>"101000000",
  25443=>"000111100",
  25444=>"100000110",
  25445=>"000111111",
  25446=>"111111110",
  25447=>"000000000",
  25448=>"111111000",
  25449=>"000000000",
  25450=>"100000111",
  25451=>"010000000",
  25452=>"000000000",
  25453=>"110110000",
  25454=>"111111000",
  25455=>"110000000",
  25456=>"111111011",
  25457=>"000000010",
  25458=>"000110010",
  25459=>"000001101",
  25460=>"000001001",
  25461=>"001001001",
  25462=>"011111111",
  25463=>"011111111",
  25464=>"111111111",
  25465=>"110010010",
  25466=>"000111001",
  25467=>"000000100",
  25468=>"111110000",
  25469=>"110110000",
  25470=>"111111001",
  25471=>"111111110",
  25472=>"001101000",
  25473=>"111111100",
  25474=>"000110000",
  25475=>"000000000",
  25476=>"111101000",
  25477=>"000011111",
  25478=>"011011001",
  25479=>"010010110",
  25480=>"011111011",
  25481=>"000000001",
  25482=>"010011111",
  25483=>"001000000",
  25484=>"000001000",
  25485=>"111111111",
  25486=>"000111100",
  25487=>"101001001",
  25488=>"000001011",
  25489=>"111000000",
  25490=>"111111000",
  25491=>"111111000",
  25492=>"011111111",
  25493=>"111111011",
  25494=>"011111001",
  25495=>"010011010",
  25496=>"111111111",
  25497=>"101000000",
  25498=>"111111001",
  25499=>"110111111",
  25500=>"010010000",
  25501=>"010111000",
  25502=>"011111111",
  25503=>"000111111",
  25504=>"000000000",
  25505=>"010110010",
  25506=>"111111000",
  25507=>"000000001",
  25508=>"100010111",
  25509=>"100010010",
  25510=>"000000000",
  25511=>"000100100",
  25512=>"010000010",
  25513=>"000100101",
  25514=>"000000000",
  25515=>"110110110",
  25516=>"101101111",
  25517=>"101000000",
  25518=>"111111110",
  25519=>"000000001",
  25520=>"000000101",
  25521=>"000000111",
  25522=>"000110100",
  25523=>"100000001",
  25524=>"000010011",
  25525=>"011001111",
  25526=>"000000110",
  25527=>"000001101",
  25528=>"000011111",
  25529=>"110110010",
  25530=>"000010111",
  25531=>"110111010",
  25532=>"101010011",
  25533=>"111111110",
  25534=>"100110111",
  25535=>"000000111",
  25536=>"111000101",
  25537=>"010011011",
  25538=>"011010000",
  25539=>"111010111",
  25540=>"000000000",
  25541=>"110000000",
  25542=>"010000000",
  25543=>"110100000",
  25544=>"000101111",
  25545=>"000111010",
  25546=>"000101000",
  25547=>"111111001",
  25548=>"011011011",
  25549=>"111001000",
  25550=>"000000000",
  25551=>"010110000",
  25552=>"111111000",
  25553=>"110110010",
  25554=>"010001000",
  25555=>"000000000",
  25556=>"010001100",
  25557=>"000000000",
  25558=>"101101101",
  25559=>"111111111",
  25560=>"000000001",
  25561=>"110010101",
  25562=>"000010001",
  25563=>"111111101",
  25564=>"001111110",
  25565=>"000000100",
  25566=>"000000000",
  25567=>"100001000",
  25568=>"000000000",
  25569=>"000000001",
  25570=>"000000000",
  25571=>"011111011",
  25572=>"000011101",
  25573=>"000000000",
  25574=>"001111101",
  25575=>"011011010",
  25576=>"110000000",
  25577=>"111110100",
  25578=>"111001001",
  25579=>"000111111",
  25580=>"000111111",
  25581=>"111101000",
  25582=>"110110000",
  25583=>"000000110",
  25584=>"000000001",
  25585=>"011001000",
  25586=>"000000011",
  25587=>"000110000",
  25588=>"000111011",
  25589=>"111111001",
  25590=>"111000010",
  25591=>"000000000",
  25592=>"110111001",
  25593=>"000000000",
  25594=>"000110000",
  25595=>"000000010",
  25596=>"111111000",
  25597=>"000000000",
  25598=>"001100011",
  25599=>"001111111",
  25600=>"100001001",
  25601=>"100100111",
  25602=>"100000100",
  25603=>"010001100",
  25604=>"111111011",
  25605=>"110101110",
  25606=>"111010011",
  25607=>"000000000",
  25608=>"010011011",
  25609=>"100100110",
  25610=>"000100000",
  25611=>"100100100",
  25612=>"110000110",
  25613=>"110100000",
  25614=>"100110111",
  25615=>"000001000",
  25616=>"111000001",
  25617=>"000000111",
  25618=>"010110111",
  25619=>"100110000",
  25620=>"110000110",
  25621=>"000100111",
  25622=>"101000111",
  25623=>"111100101",
  25624=>"100000110",
  25625=>"100100111",
  25626=>"110100100",
  25627=>"011001000",
  25628=>"100001111",
  25629=>"010010000",
  25630=>"101100100",
  25631=>"011011011",
  25632=>"111001000",
  25633=>"111100011",
  25634=>"000000001",
  25635=>"000000000",
  25636=>"001001001",
  25637=>"000000000",
  25638=>"000011011",
  25639=>"011010000",
  25640=>"110100000",
  25641=>"000000011",
  25642=>"100100100",
  25643=>"111110110",
  25644=>"111010111",
  25645=>"100011011",
  25646=>"001100110",
  25647=>"101111010",
  25648=>"001011010",
  25649=>"100110111",
  25650=>"001011011",
  25651=>"011111110",
  25652=>"110100110",
  25653=>"000010011",
  25654=>"000110111",
  25655=>"011011011",
  25656=>"011111000",
  25657=>"100100100",
  25658=>"010110110",
  25659=>"000000100",
  25660=>"000010010",
  25661=>"011011010",
  25662=>"010000100",
  25663=>"101001000",
  25664=>"110100100",
  25665=>"000000000",
  25666=>"000001011",
  25667=>"110110111",
  25668=>"011111000",
  25669=>"000000000",
  25670=>"101101111",
  25671=>"101111000",
  25672=>"000011011",
  25673=>"000000110",
  25674=>"010000000",
  25675=>"100100110",
  25676=>"001000100",
  25677=>"111011111",
  25678=>"011000000",
  25679=>"001011011",
  25680=>"000000001",
  25681=>"100000000",
  25682=>"100110111",
  25683=>"101000000",
  25684=>"100100000",
  25685=>"000000011",
  25686=>"110001001",
  25687=>"000100100",
  25688=>"110100000",
  25689=>"001111111",
  25690=>"001000000",
  25691=>"111110110",
  25692=>"000011011",
  25693=>"000101100",
  25694=>"000001011",
  25695=>"100000001",
  25696=>"001011011",
  25697=>"011011000",
  25698=>"100100100",
  25699=>"111111111",
  25700=>"010010010",
  25701=>"111111100",
  25702=>"100100110",
  25703=>"011000000",
  25704=>"011011000",
  25705=>"001010100",
  25706=>"000000111",
  25707=>"110110100",
  25708=>"011011011",
  25709=>"100100111",
  25710=>"001000000",
  25711=>"000100110",
  25712=>"001001001",
  25713=>"011110110",
  25714=>"111011011",
  25715=>"011111001",
  25716=>"100110011",
  25717=>"100100010",
  25718=>"111100100",
  25719=>"000000001",
  25720=>"111100111",
  25721=>"011011011",
  25722=>"000110111",
  25723=>"110100110",
  25724=>"011100100",
  25725=>"010010000",
  25726=>"111011000",
  25727=>"000100111",
  25728=>"000110000",
  25729=>"000000000",
  25730=>"010000011",
  25731=>"011011001",
  25732=>"100100100",
  25733=>"010011011",
  25734=>"100100011",
  25735=>"011100101",
  25736=>"100011110",
  25737=>"001000010",
  25738=>"101100111",
  25739=>"011011010",
  25740=>"000011011",
  25741=>"100111111",
  25742=>"011011011",
  25743=>"100000010",
  25744=>"000000000",
  25745=>"010110110",
  25746=>"111110110",
  25747=>"011110111",
  25748=>"011011000",
  25749=>"110100100",
  25750=>"000001001",
  25751=>"000000001",
  25752=>"000000000",
  25753=>"000101011",
  25754=>"011011110",
  25755=>"000000000",
  25756=>"001110110",
  25757=>"101001101",
  25758=>"111110010",
  25759=>"001000100",
  25760=>"010100101",
  25761=>"100100110",
  25762=>"010001011",
  25763=>"010111000",
  25764=>"100100100",
  25765=>"011000110",
  25766=>"111111000",
  25767=>"011111011",
  25768=>"101011111",
  25769=>"000011011",
  25770=>"000110100",
  25771=>"110100000",
  25772=>"011011000",
  25773=>"111001001",
  25774=>"110110111",
  25775=>"111011011",
  25776=>"001100010",
  25777=>"001001001",
  25778=>"111111100",
  25779=>"110010110",
  25780=>"010001001",
  25781=>"000000000",
  25782=>"011011100",
  25783=>"001100100",
  25784=>"110100100",
  25785=>"001011000",
  25786=>"110100000",
  25787=>"011001000",
  25788=>"000100001",
  25789=>"000011011",
  25790=>"011011001",
  25791=>"000000000",
  25792=>"100100100",
  25793=>"000100000",
  25794=>"000000011",
  25795=>"001101011",
  25796=>"011111111",
  25797=>"001011010",
  25798=>"011011001",
  25799=>"111100100",
  25800=>"011001010",
  25801=>"111011001",
  25802=>"011011101",
  25803=>"000000111",
  25804=>"111000011",
  25805=>"001000110",
  25806=>"011111101",
  25807=>"011011010",
  25808=>"110100100",
  25809=>"100111111",
  25810=>"010100100",
  25811=>"111000011",
  25812=>"011100000",
  25813=>"111111111",
  25814=>"000000110",
  25815=>"110000000",
  25816=>"110000000",
  25817=>"011000000",
  25818=>"000010110",
  25819=>"100100100",
  25820=>"011010100",
  25821=>"011111001",
  25822=>"010000010",
  25823=>"000000000",
  25824=>"010110100",
  25825=>"100110100",
  25826=>"100100100",
  25827=>"011001010",
  25828=>"100100100",
  25829=>"011000000",
  25830=>"111100100",
  25831=>"001011011",
  25832=>"110100100",
  25833=>"011000100",
  25834=>"100100110",
  25835=>"101100101",
  25836=>"010010010",
  25837=>"111100100",
  25838=>"000000000",
  25839=>"011101011",
  25840=>"001000000",
  25841=>"111111001",
  25842=>"111000000",
  25843=>"001110100",
  25844=>"010010010",
  25845=>"000000001",
  25846=>"110100000",
  25847=>"000001000",
  25848=>"100100100",
  25849=>"111100011",
  25850=>"010010110",
  25851=>"111011011",
  25852=>"011011011",
  25853=>"001011010",
  25854=>"000000000",
  25855=>"000000100",
  25856=>"011101000",
  25857=>"000000000",
  25858=>"000101111",
  25859=>"110110111",
  25860=>"000011100",
  25861=>"000001000",
  25862=>"011010100",
  25863=>"110110000",
  25864=>"010111111",
  25865=>"011111111",
  25866=>"011111110",
  25867=>"000000000",
  25868=>"111111111",
  25869=>"010000001",
  25870=>"001111011",
  25871=>"111101111",
  25872=>"001011111",
  25873=>"111101101",
  25874=>"100010010",
  25875=>"111011000",
  25876=>"010000000",
  25877=>"111001000",
  25878=>"011100111",
  25879=>"000111111",
  25880=>"001000001",
  25881=>"000101111",
  25882=>"101111111",
  25883=>"000100000",
  25884=>"100001001",
  25885=>"011111111",
  25886=>"111010010",
  25887=>"000010100",
  25888=>"000100000",
  25889=>"000000000",
  25890=>"111111101",
  25891=>"100101111",
  25892=>"001111001",
  25893=>"110100100",
  25894=>"111111000",
  25895=>"001011111",
  25896=>"000111000",
  25897=>"100010000",
  25898=>"111001011",
  25899=>"011111011",
  25900=>"111111111",
  25901=>"011111111",
  25902=>"111100000",
  25903=>"010001001",
  25904=>"001011000",
  25905=>"100100000",
  25906=>"110001111",
  25907=>"110110110",
  25908=>"000011001",
  25909=>"110000000",
  25910=>"000001001",
  25911=>"000000001",
  25912=>"100111110",
  25913=>"101000001",
  25914=>"101111111",
  25915=>"111111111",
  25916=>"000000001",
  25917=>"111111111",
  25918=>"111001000",
  25919=>"000101110",
  25920=>"100000000",
  25921=>"000000010",
  25922=>"000000000",
  25923=>"000000100",
  25924=>"111010000",
  25925=>"111011000",
  25926=>"110000000",
  25927=>"111111111",
  25928=>"111111001",
  25929=>"101101101",
  25930=>"101000000",
  25931=>"101000000",
  25932=>"001000101",
  25933=>"110100100",
  25934=>"000011011",
  25935=>"111111110",
  25936=>"000000000",
  25937=>"000111000",
  25938=>"111011111",
  25939=>"111111001",
  25940=>"010001011",
  25941=>"000100001",
  25942=>"110111101",
  25943=>"000111111",
  25944=>"111111101",
  25945=>"001110010",
  25946=>"001000001",
  25947=>"100111001",
  25948=>"010010111",
  25949=>"011011001",
  25950=>"000000000",
  25951=>"000001001",
  25952=>"000110110",
  25953=>"000011111",
  25954=>"101001000",
  25955=>"100100110",
  25956=>"111111111",
  25957=>"011111111",
  25958=>"110010000",
  25959=>"111111111",
  25960=>"101000001",
  25961=>"101010000",
  25962=>"001000000",
  25963=>"111101000",
  25964=>"000000000",
  25965=>"001000000",
  25966=>"001001101",
  25967=>"010000000",
  25968=>"000001000",
  25969=>"010011111",
  25970=>"000100100",
  25971=>"011111111",
  25972=>"010000111",
  25973=>"001000111",
  25974=>"110000000",
  25975=>"010000000",
  25976=>"000111001",
  25977=>"000000111",
  25978=>"000000101",
  25979=>"110010011",
  25980=>"110110110",
  25981=>"111110100",
  25982=>"110111111",
  25983=>"110110101",
  25984=>"111001000",
  25985=>"000000000",
  25986=>"000000000",
  25987=>"000000011",
  25988=>"100011111",
  25989=>"101010000",
  25990=>"011001000",
  25991=>"011011011",
  25992=>"100000001",
  25993=>"101010000",
  25994=>"010110100",
  25995=>"111111000",
  25996=>"000000010",
  25997=>"000100000",
  25998=>"000000101",
  25999=>"111001101",
  26000=>"111111110",
  26001=>"101000000",
  26002=>"011101111",
  26003=>"111011111",
  26004=>"110011111",
  26005=>"000000000",
  26006=>"111111111",
  26007=>"011001000",
  26008=>"000000000",
  26009=>"000111111",
  26010=>"111111111",
  26011=>"000111111",
  26012=>"000000000",
  26013=>"000000000",
  26014=>"011111000",
  26015=>"010000000",
  26016=>"001001000",
  26017=>"011111100",
  26018=>"011001100",
  26019=>"101111111",
  26020=>"011000001",
  26021=>"110111111",
  26022=>"111111111",
  26023=>"000001001",
  26024=>"011111010",
  26025=>"100110110",
  26026=>"101101101",
  26027=>"010000000",
  26028=>"110010010",
  26029=>"110000000",
  26030=>"111111000",
  26031=>"111110000",
  26032=>"000000000",
  26033=>"011101100",
  26034=>"100110000",
  26035=>"100000000",
  26036=>"011110010",
  26037=>"011111011",
  26038=>"111111110",
  26039=>"110100001",
  26040=>"001000000",
  26041=>"010110110",
  26042=>"111001111",
  26043=>"000001101",
  26044=>"111111111",
  26045=>"000000000",
  26046=>"000111111",
  26047=>"011011011",
  26048=>"111111111",
  26049=>"111111001",
  26050=>"111000000",
  26051=>"011111101",
  26052=>"010011010",
  26053=>"100101000",
  26054=>"111011110",
  26055=>"000000001",
  26056=>"111110000",
  26057=>"110000011",
  26058=>"111111001",
  26059=>"111111111",
  26060=>"111100000",
  26061=>"011111111",
  26062=>"000100111",
  26063=>"101000000",
  26064=>"110100000",
  26065=>"001011011",
  26066=>"111111111",
  26067=>"011111111",
  26068=>"110111111",
  26069=>"100100100",
  26070=>"100110111",
  26071=>"010011110",
  26072=>"110111111",
  26073=>"000000011",
  26074=>"100100000",
  26075=>"000000111",
  26076=>"010001100",
  26077=>"000000011",
  26078=>"111111011",
  26079=>"111111111",
  26080=>"110011011",
  26081=>"110110100",
  26082=>"010111011",
  26083=>"010111110",
  26084=>"111100110",
  26085=>"000000000",
  26086=>"000000000",
  26087=>"100100100",
  26088=>"000000101",
  26089=>"111101111",
  26090=>"110111111",
  26091=>"111101111",
  26092=>"000010010",
  26093=>"110111111",
  26094=>"111110000",
  26095=>"111101111",
  26096=>"000001111",
  26097=>"001010000",
  26098=>"111100111",
  26099=>"111111111",
  26100=>"010011011",
  26101=>"001110111",
  26102=>"101101111",
  26103=>"010100100",
  26104=>"000000000",
  26105=>"111111110",
  26106=>"000001001",
  26107=>"010100100",
  26108=>"000111111",
  26109=>"001000000",
  26110=>"001001001",
  26111=>"000100000",
  26112=>"110110111",
  26113=>"000000101",
  26114=>"111011001",
  26115=>"101101111",
  26116=>"111000101",
  26117=>"000001001",
  26118=>"000001010",
  26119=>"111111101",
  26120=>"111101111",
  26121=>"010000011",
  26122=>"000010000",
  26123=>"100011110",
  26124=>"101000101",
  26125=>"111111111",
  26126=>"100010010",
  26127=>"111111110",
  26128=>"111111111",
  26129=>"111111111",
  26130=>"010110000",
  26131=>"000001111",
  26132=>"111101111",
  26133=>"110000111",
  26134=>"000000000",
  26135=>"000111000",
  26136=>"110000000",
  26137=>"000011000",
  26138=>"100000000",
  26139=>"101100100",
  26140=>"000100110",
  26141=>"101111111",
  26142=>"011111101",
  26143=>"101000111",
  26144=>"101110111",
  26145=>"010111011",
  26146=>"000000000",
  26147=>"010001111",
  26148=>"000111111",
  26149=>"011101110",
  26150=>"100111000",
  26151=>"000000011",
  26152=>"101111000",
  26153=>"111111001",
  26154=>"000101000",
  26155=>"011000111",
  26156=>"000111011",
  26157=>"110111001",
  26158=>"000111000",
  26159=>"110000110",
  26160=>"111110000",
  26161=>"001110000",
  26162=>"010000000",
  26163=>"011111111",
  26164=>"000010000",
  26165=>"010011111",
  26166=>"100000000",
  26167=>"111010111",
  26168=>"101000111",
  26169=>"001000110",
  26170=>"000000000",
  26171=>"000010011",
  26172=>"001111110",
  26173=>"001000000",
  26174=>"111111110",
  26175=>"000001010",
  26176=>"111111100",
  26177=>"001000011",
  26178=>"010100010",
  26179=>"010100100",
  26180=>"101001110",
  26181=>"111000101",
  26182=>"000001011",
  26183=>"101110111",
  26184=>"001111010",
  26185=>"100011101",
  26186=>"111001000",
  26187=>"111001000",
  26188=>"110010110",
  26189=>"001111111",
  26190=>"010111010",
  26191=>"000101101",
  26192=>"111110111",
  26193=>"101111101",
  26194=>"001101111",
  26195=>"101111000",
  26196=>"001000010",
  26197=>"100000000",
  26198=>"000000010",
  26199=>"111101100",
  26200=>"011011110",
  26201=>"110100000",
  26202=>"000000110",
  26203=>"111011000",
  26204=>"101101110",
  26205=>"100100001",
  26206=>"101101111",
  26207=>"010000001",
  26208=>"000000000",
  26209=>"011000100",
  26210=>"011000110",
  26211=>"000001001",
  26212=>"011001100",
  26213=>"000111010",
  26214=>"000000001",
  26215=>"000001111",
  26216=>"000100111",
  26217=>"000000000",
  26218=>"000100001",
  26219=>"001000101",
  26220=>"000111000",
  26221=>"111111011",
  26222=>"110000111",
  26223=>"000111001",
  26224=>"110000000",
  26225=>"111000000",
  26226=>"010010000",
  26227=>"000100001",
  26228=>"100000010",
  26229=>"101000000",
  26230=>"001000001",
  26231=>"111001101",
  26232=>"101111001",
  26233=>"011111000",
  26234=>"000001011",
  26235=>"110111000",
  26236=>"011011110",
  26237=>"000001000",
  26238=>"111111011",
  26239=>"000000011",
  26240=>"111111000",
  26241=>"000011001",
  26242=>"000000110",
  26243=>"101100010",
  26244=>"001101000",
  26245=>"000010000",
  26246=>"111001011",
  26247=>"000001110",
  26248=>"011000000",
  26249=>"000000000",
  26250=>"111111111",
  26251=>"000010011",
  26252=>"011001111",
  26253=>"110010110",
  26254=>"111000000",
  26255=>"000000000",
  26256=>"000101100",
  26257=>"010000000",
  26258=>"011111000",
  26259=>"100101001",
  26260=>"101000101",
  26261=>"110111111",
  26262=>"000111011",
  26263=>"111100000",
  26264=>"011111101",
  26265=>"111100011",
  26266=>"110111111",
  26267=>"111001000",
  26268=>"101101101",
  26269=>"111110000",
  26270=>"000110111",
  26271=>"000111110",
  26272=>"000000000",
  26273=>"111111111",
  26274=>"101111110",
  26275=>"011110111",
  26276=>"000111000",
  26277=>"011011000",
  26278=>"111001001",
  26279=>"010000100",
  26280=>"111111111",
  26281=>"111001001",
  26282=>"111100001",
  26283=>"000010111",
  26284=>"111100001",
  26285=>"111100100",
  26286=>"111111111",
  26287=>"100101000",
  26288=>"111000100",
  26289=>"001011011",
  26290=>"000111010",
  26291=>"000000000",
  26292=>"010111000",
  26293=>"101010101",
  26294=>"011001000",
  26295=>"001000010",
  26296=>"100111011",
  26297=>"001001011",
  26298=>"000000000",
  26299=>"011000000",
  26300=>"100000011",
  26301=>"000001100",
  26302=>"011000110",
  26303=>"010010000",
  26304=>"000101101",
  26305=>"000000000",
  26306=>"110100111",
  26307=>"000000000",
  26308=>"110000000",
  26309=>"000111111",
  26310=>"010111000",
  26311=>"000011101",
  26312=>"010010011",
  26313=>"001000000",
  26314=>"111010111",
  26315=>"101001000",
  26316=>"001000010",
  26317=>"111110111",
  26318=>"010010110",
  26319=>"110000101",
  26320=>"111101000",
  26321=>"010011001",
  26322=>"111111111",
  26323=>"101001110",
  26324=>"111000111",
  26325=>"000000011",
  26326=>"101001111",
  26327=>"001111110",
  26328=>"001111011",
  26329=>"111001110",
  26330=>"000000000",
  26331=>"011110000",
  26332=>"000000000",
  26333=>"110000111",
  26334=>"000110000",
  26335=>"001100001",
  26336=>"101000001",
  26337=>"001111111",
  26338=>"000001011",
  26339=>"111101001",
  26340=>"101000000",
  26341=>"111010011",
  26342=>"101100111",
  26343=>"111110111",
  26344=>"001000010",
  26345=>"101000101",
  26346=>"010010110",
  26347=>"001000111",
  26348=>"111000100",
  26349=>"000000000",
  26350=>"111000000",
  26351=>"110000110",
  26352=>"000000000",
  26353=>"001100111",
  26354=>"000101101",
  26355=>"101111110",
  26356=>"000100101",
  26357=>"000000000",
  26358=>"110000110",
  26359=>"001011011",
  26360=>"011111111",
  26361=>"000010001",
  26362=>"111111000",
  26363=>"100000000",
  26364=>"010111111",
  26365=>"101101010",
  26366=>"000001011",
  26367=>"111111110",
  26368=>"001101001",
  26369=>"010000010",
  26370=>"111100100",
  26371=>"000100111",
  26372=>"111011001",
  26373=>"111001010",
  26374=>"100101100",
  26375=>"101101010",
  26376=>"100110111",
  26377=>"000111000",
  26378=>"111100001",
  26379=>"000000000",
  26380=>"101000000",
  26381=>"111101101",
  26382=>"000111111",
  26383=>"101011100",
  26384=>"011000110",
  26385=>"000010011",
  26386=>"101000111",
  26387=>"000000010",
  26388=>"111101111",
  26389=>"000000000",
  26390=>"100100100",
  26391=>"110011010",
  26392=>"111100001",
  26393=>"000111011",
  26394=>"000000100",
  26395=>"100100101",
  26396=>"000010011",
  26397=>"000000100",
  26398=>"001000000",
  26399=>"100100101",
  26400=>"010010000",
  26401=>"010011000",
  26402=>"000000100",
  26403=>"100011011",
  26404=>"010000010",
  26405=>"110111111",
  26406=>"010000000",
  26407=>"101010111",
  26408=>"011011011",
  26409=>"010111010",
  26410=>"000011000",
  26411=>"111000101",
  26412=>"000100000",
  26413=>"101000011",
  26414=>"110100100",
  26415=>"010110010",
  26416=>"111100000",
  26417=>"101111111",
  26418=>"000011100",
  26419=>"011011010",
  26420=>"111000000",
  26421=>"111111110",
  26422=>"100110000",
  26423=>"010111011",
  26424=>"111111110",
  26425=>"000000000",
  26426=>"011101111",
  26427=>"000010011",
  26428=>"000111110",
  26429=>"111111001",
  26430=>"100000100",
  26431=>"110011000",
  26432=>"001010011",
  26433=>"010011000",
  26434=>"010111110",
  26435=>"010110100",
  26436=>"000010000",
  26437=>"000000000",
  26438=>"000111000",
  26439=>"111101100",
  26440=>"100000100",
  26441=>"100100111",
  26442=>"101101101",
  26443=>"011001100",
  26444=>"000111111",
  26445=>"101111111",
  26446=>"000111111",
  26447=>"111001011",
  26448=>"000000101",
  26449=>"110111100",
  26450=>"111110100",
  26451=>"011001000",
  26452=>"011000000",
  26453=>"010110100",
  26454=>"000111011",
  26455=>"000000000",
  26456=>"101110101",
  26457=>"100100000",
  26458=>"100110100",
  26459=>"011100111",
  26460=>"000000010",
  26461=>"110101101",
  26462=>"111111100",
  26463=>"011011000",
  26464=>"000110010",
  26465=>"100100110",
  26466=>"100000110",
  26467=>"011001000",
  26468=>"000111010",
  26469=>"000100000",
  26470=>"110000100",
  26471=>"000111011",
  26472=>"111000000",
  26473=>"111101111",
  26474=>"111000001",
  26475=>"111011011",
  26476=>"111000000",
  26477=>"111000111",
  26478=>"000011011",
  26479=>"111000011",
  26480=>"101110010",
  26481=>"011000011",
  26482=>"001000000",
  26483=>"100100000",
  26484=>"000010011",
  26485=>"010000000",
  26486=>"000010010",
  26487=>"011111011",
  26488=>"011000000",
  26489=>"100100100",
  26490=>"100000100",
  26491=>"111111111",
  26492=>"000110110",
  26493=>"011000000",
  26494=>"111101100",
  26495=>"100000000",
  26496=>"011000000",
  26497=>"100100000",
  26498=>"010011011",
  26499=>"111100111",
  26500=>"111001000",
  26501=>"000100000",
  26502=>"011111110",
  26503=>"000011011",
  26504=>"100001110",
  26505=>"000000000",
  26506=>"111101100",
  26507=>"111111010",
  26508=>"000111010",
  26509=>"100011111",
  26510=>"000010000",
  26511=>"111101001",
  26512=>"111111010",
  26513=>"000000010",
  26514=>"010010011",
  26515=>"001000000",
  26516=>"000001011",
  26517=>"011010010",
  26518=>"110110000",
  26519=>"100011011",
  26520=>"011011001",
  26521=>"000100100",
  26522=>"011011000",
  26523=>"111100100",
  26524=>"000100100",
  26525=>"011011110",
  26526=>"001000000",
  26527=>"100100100",
  26528=>"111001100",
  26529=>"011101100",
  26530=>"111101010",
  26531=>"111000100",
  26532=>"011000011",
  26533=>"100011111",
  26534=>"000011011",
  26535=>"010011111",
  26536=>"011010001",
  26537=>"101000111",
  26538=>"011011000",
  26539=>"110000111",
  26540=>"011001000",
  26541=>"100110111",
  26542=>"010000000",
  26543=>"000100000",
  26544=>"011001010",
  26545=>"010000000",
  26546=>"101100110",
  26547=>"000110011",
  26548=>"001100111",
  26549=>"101111001",
  26550=>"011011011",
  26551=>"000011011",
  26552=>"000011011",
  26553=>"000011011",
  26554=>"100011011",
  26555=>"111111000",
  26556=>"111111111",
  26557=>"011011011",
  26558=>"011011000",
  26559=>"010000100",
  26560=>"011000111",
  26561=>"000011111",
  26562=>"000000000",
  26563=>"101101101",
  26564=>"011011111",
  26565=>"110000000",
  26566=>"010001111",
  26567=>"100011001",
  26568=>"000101111",
  26569=>"011000000",
  26570=>"111111111",
  26571=>"111001000",
  26572=>"000011011",
  26573=>"000001010",
  26574=>"000010000",
  26575=>"011000011",
  26576=>"100111011",
  26577=>"010110110",
  26578=>"000010010",
  26579=>"010111011",
  26580=>"111111010",
  26581=>"000000011",
  26582=>"100000100",
  26583=>"100100000",
  26584=>"111101000",
  26585=>"111100111",
  26586=>"111100010",
  26587=>"111101111",
  26588=>"100100100",
  26589=>"000000101",
  26590=>"011111111",
  26591=>"011001001",
  26592=>"100100100",
  26593=>"101100100",
  26594=>"011101111",
  26595=>"111100000",
  26596=>"111100000",
  26597=>"010000010",
  26598=>"011000111",
  26599=>"011000000",
  26600=>"111101110",
  26601=>"010000100",
  26602=>"100100100",
  26603=>"110000111",
  26604=>"001001000",
  26605=>"000011011",
  26606=>"000000000",
  26607=>"000000010",
  26608=>"000000000",
  26609=>"000000100",
  26610=>"010001101",
  26611=>"101111111",
  26612=>"000100100",
  26613=>"111100000",
  26614=>"000001011",
  26615=>"100101100",
  26616=>"011000000",
  26617=>"111011110",
  26618=>"111100100",
  26619=>"000000101",
  26620=>"000000000",
  26621=>"011000000",
  26622=>"011111100",
  26623=>"101100100",
  26624=>"000010001",
  26625=>"000000010",
  26626=>"010011100",
  26627=>"010001001",
  26628=>"101100000",
  26629=>"000001001",
  26630=>"011001100",
  26631=>"011010011",
  26632=>"010000000",
  26633=>"000010010",
  26634=>"010000000",
  26635=>"010001000",
  26636=>"001001001",
  26637=>"101101001",
  26638=>"100001000",
  26639=>"111011001",
  26640=>"010010000",
  26641=>"011011000",
  26642=>"000100110",
  26643=>"000000011",
  26644=>"011001001",
  26645=>"000001111",
  26646=>"010011101",
  26647=>"001111011",
  26648=>"001100100",
  26649=>"111111100",
  26650=>"011001001",
  26651=>"111001001",
  26652=>"011101111",
  26653=>"000100000",
  26654=>"011101001",
  26655=>"010010000",
  26656=>"011001001",
  26657=>"000100101",
  26658=>"111001000",
  26659=>"110011011",
  26660=>"100110100",
  26661=>"010000101",
  26662=>"010110010",
  26663=>"101101000",
  26664=>"110110011",
  26665=>"010010000",
  26666=>"100111011",
  26667=>"000000001",
  26668=>"111111110",
  26669=>"001001100",
  26670=>"011111100",
  26671=>"100100010",
  26672=>"111001000",
  26673=>"110100000",
  26674=>"011000000",
  26675=>"111110011",
  26676=>"011001000",
  26677=>"010001010",
  26678=>"100000100",
  26679=>"001101000",
  26680=>"000100100",
  26681=>"001100100",
  26682=>"000100100",
  26683=>"001010000",
  26684=>"000000011",
  26685=>"110110010",
  26686=>"011001001",
  26687=>"000100110",
  26688=>"001001101",
  26689=>"011000100",
  26690=>"110110011",
  26691=>"000001001",
  26692=>"000111001",
  26693=>"001001000",
  26694=>"110110010",
  26695=>"111111111",
  26696=>"000100011",
  26697=>"111010010",
  26698=>"011001001",
  26699=>"001110110",
  26700=>"000000100",
  26701=>"101110010",
  26702=>"000000110",
  26703=>"111010011",
  26704=>"000001000",
  26705=>"110110110",
  26706=>"011001001",
  26707=>"000011010",
  26708=>"010111111",
  26709=>"111000000",
  26710=>"000100111",
  26711=>"010010111",
  26712=>"011111111",
  26713=>"000110000",
  26714=>"101000010",
  26715=>"110100110",
  26716=>"011001000",
  26717=>"000000100",
  26718=>"111111011",
  26719=>"011010000",
  26720=>"100100000",
  26721=>"011001001",
  26722=>"100011111",
  26723=>"000101101",
  26724=>"110110110",
  26725=>"100100000",
  26726=>"111111000",
  26727=>"110110010",
  26728=>"110010101",
  26729=>"100100111",
  26730=>"000111011",
  26731=>"111111011",
  26732=>"110011111",
  26733=>"101101111",
  26734=>"000000000",
  26735=>"010100100",
  26736=>"101110010",
  26737=>"010100100",
  26738=>"110011010",
  26739=>"011000000",
  26740=>"110100110",
  26741=>"000101001",
  26742=>"111110011",
  26743=>"000110110",
  26744=>"011001001",
  26745=>"011000110",
  26746=>"100101011",
  26747=>"001001111",
  26748=>"101100110",
  26749=>"111001001",
  26750=>"010000111",
  26751=>"000011000",
  26752=>"010110001",
  26753=>"100100101",
  26754=>"001001001",
  26755=>"000100000",
  26756=>"000110101",
  26757=>"110111000",
  26758=>"001000100",
  26759=>"010010000",
  26760=>"110100101",
  26761=>"001010000",
  26762=>"001111000",
  26763=>"111001000",
  26764=>"100000011",
  26765=>"100011011",
  26766=>"011011110",
  26767=>"001000001",
  26768=>"000110110",
  26769=>"000010011",
  26770=>"000110000",
  26771=>"100000000",
  26772=>"000110010",
  26773=>"011000001",
  26774=>"010110111",
  26775=>"000000000",
  26776=>"111000010",
  26777=>"110000010",
  26778=>"110100000",
  26779=>"110100000",
  26780=>"001001001",
  26781=>"000001010",
  26782=>"011001110",
  26783=>"100101111",
  26784=>"000100000",
  26785=>"011000001",
  26786=>"110100100",
  26787=>"010011001",
  26788=>"110111111",
  26789=>"101011001",
  26790=>"111000000",
  26791=>"110111001",
  26792=>"011011011",
  26793=>"001100100",
  26794=>"100000000",
  26795=>"000000001",
  26796=>"001011111",
  26797=>"110100010",
  26798=>"011000000",
  26799=>"111011001",
  26800=>"000000111",
  26801=>"011001110",
  26802=>"000101100",
  26803=>"000100110",
  26804=>"100110011",
  26805=>"111100010",
  26806=>"000100110",
  26807=>"010000000",
  26808=>"000100000",
  26809=>"111000110",
  26810=>"011011001",
  26811=>"000100011",
  26812=>"100100000",
  26813=>"110110011",
  26814=>"101110011",
  26815=>"011011100",
  26816=>"011001000",
  26817=>"011011000",
  26818=>"011100110",
  26819=>"010110000",
  26820=>"001100100",
  26821=>"111111100",
  26822=>"010100111",
  26823=>"011010001",
  26824=>"000000001",
  26825=>"000100000",
  26826=>"100110110",
  26827=>"011011010",
  26828=>"000011011",
  26829=>"110000101",
  26830=>"001000000",
  26831=>"010100000",
  26832=>"100110111",
  26833=>"001000010",
  26834=>"000010000",
  26835=>"111011011",
  26836=>"100000101",
  26837=>"011101000",
  26838=>"001000100",
  26839=>"010001000",
  26840=>"101110010",
  26841=>"111000111",
  26842=>"101001110",
  26843=>"101001001",
  26844=>"111100100",
  26845=>"000110111",
  26846=>"001111111",
  26847=>"011000001",
  26848=>"011011001",
  26849=>"101001001",
  26850=>"100111011",
  26851=>"100110110",
  26852=>"010000001",
  26853=>"110110100",
  26854=>"111000111",
  26855=>"100100111",
  26856=>"111101111",
  26857=>"011100000",
  26858=>"111100010",
  26859=>"100110011",
  26860=>"011001001",
  26861=>"000000000",
  26862=>"000001001",
  26863=>"000000100",
  26864=>"100011011",
  26865=>"000000100",
  26866=>"011001001",
  26867=>"110101110",
  26868=>"111001001",
  26869=>"100110011",
  26870=>"000001000",
  26871=>"100100110",
  26872=>"001001001",
  26873=>"100000000",
  26874=>"011001000",
  26875=>"100110110",
  26876=>"011010110",
  26877=>"110100011",
  26878=>"100100111",
  26879=>"011110111",
  26880=>"000000011",
  26881=>"001000111",
  26882=>"000010111",
  26883=>"000000100",
  26884=>"000111111",
  26885=>"101001100",
  26886=>"110100010",
  26887=>"000111010",
  26888=>"010000000",
  26889=>"010011001",
  26890=>"111111110",
  26891=>"000000000",
  26892=>"001000000",
  26893=>"000000110",
  26894=>"011100100",
  26895=>"110110101",
  26896=>"000111011",
  26897=>"010110110",
  26898=>"000000101",
  26899=>"111111111",
  26900=>"000000111",
  26901=>"000000000",
  26902=>"100000100",
  26903=>"011111111",
  26904=>"000000011",
  26905=>"000000001",
  26906=>"011000000",
  26907=>"000000111",
  26908=>"110010010",
  26909=>"010101111",
  26910=>"000010010",
  26911=>"001000000",
  26912=>"000010000",
  26913=>"001111111",
  26914=>"000000111",
  26915=>"111101111",
  26916=>"111100100",
  26917=>"000101000",
  26918=>"000111011",
  26919=>"000111111",
  26920=>"000111111",
  26921=>"011100000",
  26922=>"000000000",
  26923=>"100000101",
  26924=>"100110111",
  26925=>"111010110",
  26926=>"000110111",
  26927=>"001001000",
  26928=>"110111111",
  26929=>"101111011",
  26930=>"000101000",
  26931=>"010010000",
  26932=>"001111111",
  26933=>"011111101",
  26934=>"000100011",
  26935=>"000001101",
  26936=>"111111001",
  26937=>"001000111",
  26938=>"111000000",
  26939=>"010011000",
  26940=>"011011111",
  26941=>"101100101",
  26942=>"110000000",
  26943=>"100011111",
  26944=>"111111000",
  26945=>"000110000",
  26946=>"111000000",
  26947=>"110011011",
  26948=>"111000000",
  26949=>"001010011",
  26950=>"111011110",
  26951=>"001000000",
  26952=>"001001011",
  26953=>"000111111",
  26954=>"001100111",
  26955=>"010011000",
  26956=>"111000000",
  26957=>"011111111",
  26958=>"001111110",
  26959=>"111101100",
  26960=>"000000111",
  26961=>"111000000",
  26962=>"010000001",
  26963=>"010101100",
  26964=>"000010110",
  26965=>"100110111",
  26966=>"111011011",
  26967=>"000111111",
  26968=>"111000000",
  26969=>"010000000",
  26970=>"111000000",
  26971=>"010000000",
  26972=>"111111111",
  26973=>"110110000",
  26974=>"111111000",
  26975=>"011110111",
  26976=>"111001000",
  26977=>"011000010",
  26978=>"001000000",
  26979=>"111011000",
  26980=>"111101000",
  26981=>"101100000",
  26982=>"000111011",
  26983=>"000000000",
  26984=>"001111101",
  26985=>"111111000",
  26986=>"111111000",
  26987=>"000000000",
  26988=>"111111001",
  26989=>"110111111",
  26990=>"111101111",
  26991=>"000000001",
  26992=>"001100110",
  26993=>"111000000",
  26994=>"001001001",
  26995=>"000101000",
  26996=>"001101111",
  26997=>"000000000",
  26998=>"111101000",
  26999=>"000011000",
  27000=>"000000111",
  27001=>"000000101",
  27002=>"111101000",
  27003=>"010111111",
  27004=>"111100111",
  27005=>"010100000",
  27006=>"000101000",
  27007=>"000000110",
  27008=>"010001000",
  27009=>"010011111",
  27010=>"000001111",
  27011=>"001000101",
  27012=>"010110111",
  27013=>"111000001",
  27014=>"000110000",
  27015=>"111100000",
  27016=>"101001011",
  27017=>"110011000",
  27018=>"000100011",
  27019=>"000000010",
  27020=>"111000000",
  27021=>"110000000",
  27022=>"111000000",
  27023=>"110110000",
  27024=>"011101111",
  27025=>"001001000",
  27026=>"100000000",
  27027=>"001000110",
  27028=>"000001111",
  27029=>"111110000",
  27030=>"011000000",
  27031=>"111110100",
  27032=>"010000000",
  27033=>"000000010",
  27034=>"010011011",
  27035=>"000100010",
  27036=>"111000000",
  27037=>"101110111",
  27038=>"100000000",
  27039=>"000000101",
  27040=>"001101111",
  27041=>"111010101",
  27042=>"111101001",
  27043=>"111000000",
  27044=>"111111101",
  27045=>"000000011",
  27046=>"111100100",
  27047=>"110000000",
  27048=>"111110111",
  27049=>"111111001",
  27050=>"111000000",
  27051=>"000000101",
  27052=>"011000111",
  27053=>"000111111",
  27054=>"011011111",
  27055=>"011000000",
  27056=>"101001001",
  27057=>"111100000",
  27058=>"101111110",
  27059=>"001000101",
  27060=>"011111110",
  27061=>"111001000",
  27062=>"000100111",
  27063=>"000110000",
  27064=>"100110100",
  27065=>"000010111",
  27066=>"000000000",
  27067=>"000011111",
  27068=>"100011000",
  27069=>"111111111",
  27070=>"110100111",
  27071=>"100000000",
  27072=>"000010111",
  27073=>"111000000",
  27074=>"001101111",
  27075=>"000100100",
  27076=>"000111101",
  27077=>"111000001",
  27078=>"101111111",
  27079=>"100000000",
  27080=>"000000110",
  27081=>"111001111",
  27082=>"111001001",
  27083=>"000010000",
  27084=>"000010000",
  27085=>"110011111",
  27086=>"000000111",
  27087=>"000000111",
  27088=>"000111111",
  27089=>"111011000",
  27090=>"001001011",
  27091=>"101000001",
  27092=>"110000000",
  27093=>"011011011",
  27094=>"111100000",
  27095=>"000000001",
  27096=>"000111000",
  27097=>"010111101",
  27098=>"000000101",
  27099=>"100000000",
  27100=>"001011001",
  27101=>"000100000",
  27102=>"111000000",
  27103=>"001110111",
  27104=>"000000111",
  27105=>"011000111",
  27106=>"000111111",
  27107=>"000101110",
  27108=>"100000000",
  27109=>"011000001",
  27110=>"111010111",
  27111=>"110110011",
  27112=>"111111000",
  27113=>"011000101",
  27114=>"110110111",
  27115=>"111100000",
  27116=>"001111111",
  27117=>"000111111",
  27118=>"010010110",
  27119=>"111101000",
  27120=>"000001000",
  27121=>"111000100",
  27122=>"111001000",
  27123=>"111001000",
  27124=>"000000110",
  27125=>"111000000",
  27126=>"111000000",
  27127=>"000000000",
  27128=>"000111111",
  27129=>"111111101",
  27130=>"100000111",
  27131=>"111110000",
  27132=>"110000010",
  27133=>"001000000",
  27134=>"111011111",
  27135=>"111111100",
  27136=>"010101100",
  27137=>"010011010",
  27138=>"001000000",
  27139=>"010001001",
  27140=>"010110011",
  27141=>"000101111",
  27142=>"000010011",
  27143=>"111101000",
  27144=>"101000000",
  27145=>"011011010",
  27146=>"010111111",
  27147=>"111001001",
  27148=>"111001001",
  27149=>"100000001",
  27150=>"111111111",
  27151=>"111111111",
  27152=>"010010000",
  27153=>"110010000",
  27154=>"110100111",
  27155=>"000000000",
  27156=>"100001000",
  27157=>"101000000",
  27158=>"000000011",
  27159=>"111100111",
  27160=>"010100010",
  27161=>"100111011",
  27162=>"100100000",
  27163=>"000001001",
  27164=>"000101000",
  27165=>"111111000",
  27166=>"000001111",
  27167=>"000000000",
  27168=>"000000000",
  27169=>"010110010",
  27170=>"110000000",
  27171=>"100000000",
  27172=>"000000000",
  27173=>"110111001",
  27174=>"101000000",
  27175=>"100111110",
  27176=>"000001000",
  27177=>"101001000",
  27178=>"011001000",
  27179=>"000000100",
  27180=>"111110010",
  27181=>"111101101",
  27182=>"000000111",
  27183=>"000110110",
  27184=>"000000000",
  27185=>"001011000",
  27186=>"000001111",
  27187=>"100010110",
  27188=>"000111111",
  27189=>"011000000",
  27190=>"111010001",
  27191=>"101101100",
  27192=>"111111101",
  27193=>"101000111",
  27194=>"001000000",
  27195=>"000111001",
  27196=>"111001011",
  27197=>"010111011",
  27198=>"000000000",
  27199=>"111111111",
  27200=>"000000111",
  27201=>"100110110",
  27202=>"010000111",
  27203=>"111111110",
  27204=>"111100000",
  27205=>"000100001",
  27206=>"000000000",
  27207=>"000000000",
  27208=>"001101001",
  27209=>"000111011",
  27210=>"101000101",
  27211=>"111111001",
  27212=>"111000000",
  27213=>"000000000",
  27214=>"100011100",
  27215=>"101000000",
  27216=>"001001000",
  27217=>"110111111",
  27218=>"000000001",
  27219=>"001001000",
  27220=>"000111010",
  27221=>"001000100",
  27222=>"110110110",
  27223=>"111000110",
  27224=>"101101011",
  27225=>"011111110",
  27226=>"110010000",
  27227=>"111111111",
  27228=>"000010111",
  27229=>"000000100",
  27230=>"000111110",
  27231=>"111111011",
  27232=>"111101000",
  27233=>"110111111",
  27234=>"000111011",
  27235=>"111111010",
  27236=>"011001011",
  27237=>"011111111",
  27238=>"110111000",
  27239=>"001111011",
  27240=>"111001000",
  27241=>"111111010",
  27242=>"000110111",
  27243=>"100101001",
  27244=>"110000001",
  27245=>"011111111",
  27246=>"000000000",
  27247=>"111000110",
  27248=>"010110110",
  27249=>"111111111",
  27250=>"010000000",
  27251=>"010110110",
  27252=>"100001000",
  27253=>"101101101",
  27254=>"111111111",
  27255=>"111111011",
  27256=>"000000000",
  27257=>"000000010",
  27258=>"000111111",
  27259=>"101000111",
  27260=>"111011101",
  27261=>"100000010",
  27262=>"000000000",
  27263=>"101111111",
  27264=>"111000010",
  27265=>"111110000",
  27266=>"010010011",
  27267=>"000000000",
  27268=>"101111111",
  27269=>"100000000",
  27270=>"011011100",
  27271=>"110010011",
  27272=>"100011000",
  27273=>"111011000",
  27274=>"000000000",
  27275=>"001000000",
  27276=>"000111111",
  27277=>"001010010",
  27278=>"111001011",
  27279=>"101000000",
  27280=>"000110110",
  27281=>"001101111",
  27282=>"111111001",
  27283=>"000010000",
  27284=>"111001001",
  27285=>"010010010",
  27286=>"111111010",
  27287=>"110100100",
  27288=>"001101001",
  27289=>"111011000",
  27290=>"000000000",
  27291=>"000000000",
  27292=>"000000000",
  27293=>"101000000",
  27294=>"111101000",
  27295=>"111000111",
  27296=>"001001001",
  27297=>"110011110",
  27298=>"000000000",
  27299=>"000000111",
  27300=>"000000110",
  27301=>"000000110",
  27302=>"111001000",
  27303=>"100000000",
  27304=>"010111011",
  27305=>"111100100",
  27306=>"000000000",
  27307=>"111110110",
  27308=>"110110100",
  27309=>"010100101",
  27310=>"111111111",
  27311=>"000000010",
  27312=>"000000101",
  27313=>"000110110",
  27314=>"000011011",
  27315=>"000100111",
  27316=>"000101111",
  27317=>"100000000",
  27318=>"001000000",
  27319=>"010110000",
  27320=>"010011111",
  27321=>"111011011",
  27322=>"000111111",
  27323=>"000000000",
  27324=>"000011111",
  27325=>"111111111",
  27326=>"100101111",
  27327=>"111110110",
  27328=>"010010111",
  27329=>"000000100",
  27330=>"001001001",
  27331=>"001000000",
  27332=>"000000001",
  27333=>"111100000",
  27334=>"000000001",
  27335=>"000000111",
  27336=>"101100010",
  27337=>"111000000",
  27338=>"000000101",
  27339=>"101000000",
  27340=>"010111111",
  27341=>"110110100",
  27342=>"000010010",
  27343=>"000101111",
  27344=>"010110000",
  27345=>"011011011",
  27346=>"000010101",
  27347=>"011111111",
  27348=>"001111111",
  27349=>"000000000",
  27350=>"101000101",
  27351=>"111010000",
  27352=>"000000001",
  27353=>"000110010",
  27354=>"011000010",
  27355=>"101000110",
  27356=>"000000010",
  27357=>"001100111",
  27358=>"010111110",
  27359=>"010111011",
  27360=>"000010010",
  27361=>"100110111",
  27362=>"000111111",
  27363=>"011111110",
  27364=>"011111110",
  27365=>"000111000",
  27366=>"101001011",
  27367=>"000111111",
  27368=>"101011011",
  27369=>"000100000",
  27370=>"011111111",
  27371=>"111111111",
  27372=>"111101001",
  27373=>"100001000",
  27374=>"000000100",
  27375=>"000001111",
  27376=>"111101111",
  27377=>"101001000",
  27378=>"001000111",
  27379=>"110001111",
  27380=>"000010111",
  27381=>"000010000",
  27382=>"010111000",
  27383=>"001000111",
  27384=>"000110111",
  27385=>"111000000",
  27386=>"111101111",
  27387=>"111110100",
  27388=>"001000001",
  27389=>"010111111",
  27390=>"000000000",
  27391=>"111000000",
  27392=>"000110111",
  27393=>"000000000",
  27394=>"111000001",
  27395=>"111011111",
  27396=>"111011110",
  27397=>"100000111",
  27398=>"000000000",
  27399=>"010111010",
  27400=>"111111000",
  27401=>"000000001",
  27402=>"100101111",
  27403=>"100101000",
  27404=>"001101111",
  27405=>"010100101",
  27406=>"000010111",
  27407=>"000000111",
  27408=>"010111111",
  27409=>"100100001",
  27410=>"100010111",
  27411=>"110000000",
  27412=>"010111110",
  27413=>"110010110",
  27414=>"101101001",
  27415=>"001111101",
  27416=>"101110011",
  27417=>"011100110",
  27418=>"000001011",
  27419=>"111000101",
  27420=>"000011110",
  27421=>"000100000",
  27422=>"101101111",
  27423=>"000000000",
  27424=>"101100100",
  27425=>"011101110",
  27426=>"000000101",
  27427=>"000111111",
  27428=>"110110011",
  27429=>"101101001",
  27430=>"100101111",
  27431=>"000100000",
  27432=>"101111111",
  27433=>"000101000",
  27434=>"001100001",
  27435=>"000010101",
  27436=>"111111010",
  27437=>"101010111",
  27438=>"000101111",
  27439=>"110110000",
  27440=>"011110011",
  27441=>"111000100",
  27442=>"000001000",
  27443=>"000111110",
  27444=>"000000101",
  27445=>"001101011",
  27446=>"000110100",
  27447=>"000110000",
  27448=>"111111000",
  27449=>"000001111",
  27450=>"000000000",
  27451=>"101000010",
  27452=>"000000101",
  27453=>"111010010",
  27454=>"000000101",
  27455=>"110100101",
  27456=>"100000000",
  27457=>"100101011",
  27458=>"000000000",
  27459=>"111111111",
  27460=>"100101111",
  27461=>"000000101",
  27462=>"001111000",
  27463=>"010000000",
  27464=>"000100010",
  27465=>"010111010",
  27466=>"000101000",
  27467=>"001110101",
  27468=>"100000111",
  27469=>"001100110",
  27470=>"110100011",
  27471=>"010000111",
  27472=>"100110100",
  27473=>"111010110",
  27474=>"100010001",
  27475=>"000000011",
  27476=>"000000100",
  27477=>"001000000",
  27478=>"000010011",
  27479=>"010110111",
  27480=>"101111110",
  27481=>"001000001",
  27482=>"011001011",
  27483=>"001010010",
  27484=>"100111110",
  27485=>"101000101",
  27486=>"111000111",
  27487=>"101101111",
  27488=>"000000000",
  27489=>"000100000",
  27490=>"000000001",
  27491=>"111110111",
  27492=>"000010010",
  27493=>"000100000",
  27494=>"110110000",
  27495=>"111101011",
  27496=>"010011011",
  27497=>"100111010",
  27498=>"100101010",
  27499=>"101100111",
  27500=>"001100111",
  27501=>"101111111",
  27502=>"000000000",
  27503=>"111111111",
  27504=>"110100100",
  27505=>"101001011",
  27506=>"000111110",
  27507=>"101000000",
  27508=>"111010010",
  27509=>"000100100",
  27510=>"010000000",
  27511=>"010110100",
  27512=>"100100111",
  27513=>"111100110",
  27514=>"000000101",
  27515=>"111111101",
  27516=>"000000001",
  27517=>"001001111",
  27518=>"000000011",
  27519=>"000000011",
  27520=>"000000010",
  27521=>"101001111",
  27522=>"010011000",
  27523=>"111000000",
  27524=>"111111111",
  27525=>"000001001",
  27526=>"100011100",
  27527=>"000100001",
  27528=>"001110010",
  27529=>"011010010",
  27530=>"100111110",
  27531=>"100100000",
  27532=>"100000000",
  27533=>"000100100",
  27534=>"100000010",
  27535=>"000000000",
  27536=>"110001000",
  27537=>"111100100",
  27538=>"000101111",
  27539=>"001010101",
  27540=>"111111010",
  27541=>"011000101",
  27542=>"101011001",
  27543=>"000100100",
  27544=>"000000010",
  27545=>"100100100",
  27546=>"011000000",
  27547=>"010000000",
  27548=>"000000100",
  27549=>"011010000",
  27550=>"111100111",
  27551=>"100000010",
  27552=>"111101011",
  27553=>"111111111",
  27554=>"010101111",
  27555=>"011111111",
  27556=>"011010101",
  27557=>"000010111",
  27558=>"100111000",
  27559=>"111000000",
  27560=>"000000001",
  27561=>"000000000",
  27562=>"011100100",
  27563=>"000101101",
  27564=>"110110111",
  27565=>"000010001",
  27566=>"000111011",
  27567=>"001111111",
  27568=>"011010100",
  27569=>"000000000",
  27570=>"100000000",
  27571=>"101010011",
  27572=>"011011111",
  27573=>"001000000",
  27574=>"000000100",
  27575=>"000000000",
  27576=>"000100101",
  27577=>"000010110",
  27578=>"010000011",
  27579=>"010010111",
  27580=>"101011111",
  27581=>"111000000",
  27582=>"000000000",
  27583=>"010111000",
  27584=>"100100000",
  27585=>"100000010",
  27586=>"010010000",
  27587=>"011001000",
  27588=>"000011001",
  27589=>"001111010",
  27590=>"010111000",
  27591=>"110100011",
  27592=>"000101011",
  27593=>"001101101",
  27594=>"010010010",
  27595=>"100111111",
  27596=>"011011000",
  27597=>"000000100",
  27598=>"100111000",
  27599=>"011111111",
  27600=>"111110010",
  27601=>"001101111",
  27602=>"101111011",
  27603=>"100110111",
  27604=>"111100101",
  27605=>"000100100",
  27606=>"100000101",
  27607=>"100000000",
  27608=>"111110000",
  27609=>"001011011",
  27610=>"111110011",
  27611=>"101000000",
  27612=>"001100100",
  27613=>"001101101",
  27614=>"100000100",
  27615=>"000001111",
  27616=>"111110111",
  27617=>"000100000",
  27618=>"111111111",
  27619=>"100010011",
  27620=>"101000010",
  27621=>"011011000",
  27622=>"101011111",
  27623=>"110100110",
  27624=>"100100111",
  27625=>"110001000",
  27626=>"100110111",
  27627=>"000111111",
  27628=>"111000000",
  27629=>"000101111",
  27630=>"100000000",
  27631=>"111011100",
  27632=>"101111111",
  27633=>"101101111",
  27634=>"000000001",
  27635=>"110010100",
  27636=>"000000111",
  27637=>"101101010",
  27638=>"100000111",
  27639=>"111010100",
  27640=>"111000000",
  27641=>"010001011",
  27642=>"001101111",
  27643=>"000001000",
  27644=>"000011111",
  27645=>"000110000",
  27646=>"110111011",
  27647=>"111111010",
  27648=>"001000111",
  27649=>"111000000",
  27650=>"100110111",
  27651=>"110110111",
  27652=>"101101000",
  27653=>"110110110",
  27654=>"100110111",
  27655=>"010111001",
  27656=>"100000100",
  27657=>"100100110",
  27658=>"010010101",
  27659=>"011011001",
  27660=>"100000100",
  27661=>"111000000",
  27662=>"111101100",
  27663=>"011001001",
  27664=>"000001001",
  27665=>"001111011",
  27666=>"000100011",
  27667=>"011001001",
  27668=>"110110110",
  27669=>"111110110",
  27670=>"100100110",
  27671=>"000111011",
  27672=>"110000010",
  27673=>"011011000",
  27674=>"011001001",
  27675=>"100110111",
  27676=>"000000000",
  27677=>"001011001",
  27678=>"100110100",
  27679=>"011001001",
  27680=>"100110111",
  27681=>"100110100",
  27682=>"001000011",
  27683=>"011011000",
  27684=>"101111001",
  27685=>"011001000",
  27686=>"001001001",
  27687=>"101011000",
  27688=>"001011011",
  27689=>"111000001",
  27690=>"011000010",
  27691=>"000000001",
  27692=>"101110001",
  27693=>"110001011",
  27694=>"111011111",
  27695=>"000110011",
  27696=>"001100000",
  27697=>"000100001",
  27698=>"001001011",
  27699=>"100100001",
  27700=>"011000011",
  27701=>"011011010",
  27702=>"110001110",
  27703=>"111011010",
  27704=>"110100111",
  27705=>"110110111",
  27706=>"100011000",
  27707=>"000010000",
  27708=>"111111001",
  27709=>"010011010",
  27710=>"110100100",
  27711=>"101100100",
  27712=>"000011101",
  27713=>"001010001",
  27714=>"100100111",
  27715=>"101110000",
  27716=>"000000010",
  27717=>"110110110",
  27718=>"001011000",
  27719=>"000001000",
  27720=>"110111011",
  27721=>"010110111",
  27722=>"110000011",
  27723=>"011100010",
  27724=>"010000000",
  27725=>"101111111",
  27726=>"000111111",
  27727=>"011011100",
  27728=>"111110110",
  27729=>"001111111",
  27730=>"110100111",
  27731=>"001000000",
  27732=>"000000100",
  27733=>"000000010",
  27734=>"001001001",
  27735=>"100100110",
  27736=>"000111001",
  27737=>"000000000",
  27738=>"100000000",
  27739=>"001011010",
  27740=>"100100011",
  27741=>"000000011",
  27742=>"001001100",
  27743=>"110100111",
  27744=>"110110111",
  27745=>"001000000",
  27746=>"100100111",
  27747=>"000100000",
  27748=>"110101000",
  27749=>"001001010",
  27750=>"010001000",
  27751=>"011001001",
  27752=>"100100101",
  27753=>"000011101",
  27754=>"001000011",
  27755=>"001011000",
  27756=>"100101111",
  27757=>"011001000",
  27758=>"000110011",
  27759=>"000010011",
  27760=>"110111001",
  27761=>"010011000",
  27762=>"101001100",
  27763=>"001001000",
  27764=>"001001000",
  27765=>"011011010",
  27766=>"100011001",
  27767=>"001100110",
  27768=>"110110010",
  27769=>"000001010",
  27770=>"000011111",
  27771=>"111110111",
  27772=>"101111011",
  27773=>"001001001",
  27774=>"100100110",
  27775=>"110110110",
  27776=>"011001010",
  27777=>"011000100",
  27778=>"011110110",
  27779=>"101111001",
  27780=>"111100000",
  27781=>"111111000",
  27782=>"001100000",
  27783=>"000001000",
  27784=>"100101111",
  27785=>"000100110",
  27786=>"111110011",
  27787=>"011001100",
  27788=>"110100110",
  27789=>"110100010",
  27790=>"110110011",
  27791=>"001000001",
  27792=>"000001100",
  27793=>"110000100",
  27794=>"011000000",
  27795=>"100000111",
  27796=>"000001001",
  27797=>"100100100",
  27798=>"100100101",
  27799=>"011010001",
  27800=>"011011000",
  27801=>"000000010",
  27802=>"111111000",
  27803=>"110110110",
  27804=>"011010101",
  27805=>"110111100",
  27806=>"000000100",
  27807=>"100110100",
  27808=>"011000001",
  27809=>"111000010",
  27810=>"010000100",
  27811=>"110100000",
  27812=>"111110000",
  27813=>"011011001",
  27814=>"000001000",
  27815=>"011000010",
  27816=>"111110011",
  27817=>"110011011",
  27818=>"110110110",
  27819=>"100100110",
  27820=>"111000100",
  27821=>"100100100",
  27822=>"110110001",
  27823=>"010001000",
  27824=>"111000100",
  27825=>"000010111",
  27826=>"111110111",
  27827=>"000000000",
  27828=>"011001001",
  27829=>"001000111",
  27830=>"001001001",
  27831=>"001111010",
  27832=>"000000010",
  27833=>"001011011",
  27834=>"001011001",
  27835=>"111110110",
  27836=>"011000000",
  27837=>"110111010",
  27838=>"110110111",
  27839=>"011011000",
  27840=>"000000011",
  27841=>"110010011",
  27842=>"100001100",
  27843=>"001001001",
  27844=>"001000000",
  27845=>"101100100",
  27846=>"001001000",
  27847=>"100100111",
  27848=>"001111011",
  27849=>"011111000",
  27850=>"011011001",
  27851=>"111111111",
  27852=>"011000001",
  27853=>"110101110",
  27854=>"111111110",
  27855=>"111001100",
  27856=>"111110110",
  27857=>"011011000",
  27858=>"001001001",
  27859=>"100110000",
  27860=>"000000100",
  27861=>"111100000",
  27862=>"110100110",
  27863=>"111111111",
  27864=>"001011000",
  27865=>"011011011",
  27866=>"111100110",
  27867=>"110100111",
  27868=>"110110110",
  27869=>"011001111",
  27870=>"011011010",
  27871=>"101000000",
  27872=>"110110111",
  27873=>"110110111",
  27874=>"111111110",
  27875=>"000000001",
  27876=>"110100110",
  27877=>"101101000",
  27878=>"011101100",
  27879=>"001100110",
  27880=>"001000111",
  27881=>"111111000",
  27882=>"010110110",
  27883=>"100000000",
  27884=>"110110110",
  27885=>"011011000",
  27886=>"000100000",
  27887=>"011010000",
  27888=>"001001000",
  27889=>"001100110",
  27890=>"000100110",
  27891=>"011011000",
  27892=>"110110101",
  27893=>"110100110",
  27894=>"000001000",
  27895=>"000001000",
  27896=>"000111011",
  27897=>"100101111",
  27898=>"011010001",
  27899=>"010110001",
  27900=>"001000000",
  27901=>"101000110",
  27902=>"010000001",
  27903=>"110110110",
  27904=>"011011100",
  27905=>"000110111",
  27906=>"000000110",
  27907=>"000000000",
  27908=>"000101000",
  27909=>"001100100",
  27910=>"010100100",
  27911=>"010010010",
  27912=>"001001111",
  27913=>"000000000",
  27914=>"001011110",
  27915=>"100111101",
  27916=>"111001001",
  27917=>"100000011",
  27918=>"100000001",
  27919=>"000110010",
  27920=>"001000001",
  27921=>"001000110",
  27922=>"101001110",
  27923=>"001111000",
  27924=>"010110111",
  27925=>"101101111",
  27926=>"011111011",
  27927=>"110001000",
  27928=>"100100000",
  27929=>"110001001",
  27930=>"000000111",
  27931=>"100000010",
  27932=>"100000000",
  27933=>"011010011",
  27934=>"101100011",
  27935=>"010110101",
  27936=>"000000101",
  27937=>"100110110",
  27938=>"000010010",
  27939=>"000111011",
  27940=>"001000100",
  27941=>"101001000",
  27942=>"000001111",
  27943=>"100001010",
  27944=>"011111111",
  27945=>"110101100",
  27946=>"000000000",
  27947=>"000111000",
  27948=>"110000110",
  27949=>"111101111",
  27950=>"111111101",
  27951=>"100000111",
  27952=>"111111100",
  27953=>"111100100",
  27954=>"001000001",
  27955=>"101011000",
  27956=>"000010000",
  27957=>"111010110",
  27958=>"100001011",
  27959=>"000101111",
  27960=>"010101111",
  27961=>"000001011",
  27962=>"000001001",
  27963=>"001000000",
  27964=>"000100101",
  27965=>"111111010",
  27966=>"000000010",
  27967=>"111111111",
  27968=>"110000000",
  27969=>"010000010",
  27970=>"010111001",
  27971=>"100000001",
  27972=>"000010010",
  27973=>"110100000",
  27974=>"000111111",
  27975=>"101111111",
  27976=>"010000100",
  27977=>"111111111",
  27978=>"000001110",
  27979=>"111010000",
  27980=>"000101101",
  27981=>"100000010",
  27982=>"110001001",
  27983=>"001000010",
  27984=>"000111111",
  27985=>"101100000",
  27986=>"111111010",
  27987=>"011001000",
  27988=>"000111110",
  27989=>"001000000",
  27990=>"000101001",
  27991=>"000000010",
  27992=>"001001111",
  27993=>"011001011",
  27994=>"000000100",
  27995=>"010100111",
  27996=>"000000100",
  27997=>"000011010",
  27998=>"010101011",
  27999=>"100100101",
  28000=>"000000000",
  28001=>"010111111",
  28002=>"101000010",
  28003=>"011001011",
  28004=>"110000000",
  28005=>"001011000",
  28006=>"101111100",
  28007=>"000010000",
  28008=>"010001000",
  28009=>"111001000",
  28010=>"101111101",
  28011=>"110000000",
  28012=>"111011000",
  28013=>"111000111",
  28014=>"000000000",
  28015=>"011111111",
  28016=>"000101111",
  28017=>"100101110",
  28018=>"000111110",
  28019=>"111000000",
  28020=>"110001111",
  28021=>"100000000",
  28022=>"111111000",
  28023=>"000000000",
  28024=>"000001000",
  28025=>"000000000",
  28026=>"111000000",
  28027=>"111001101",
  28028=>"101100000",
  28029=>"111000000",
  28030=>"010010111",
  28031=>"111001111",
  28032=>"100010010",
  28033=>"110110111",
  28034=>"101111011",
  28035=>"110111111",
  28036=>"010001011",
  28037=>"010111000",
  28038=>"111011010",
  28039=>"100000000",
  28040=>"100001011",
  28041=>"010000000",
  28042=>"101101001",
  28043=>"000100111",
  28044=>"000100100",
  28045=>"111101010",
  28046=>"000101111",
  28047=>"001100100",
  28048=>"111111001",
  28049=>"000010111",
  28050=>"010001111",
  28051=>"100100011",
  28052=>"000100010",
  28053=>"001000000",
  28054=>"111110010",
  28055=>"111000001",
  28056=>"111111000",
  28057=>"011011000",
  28058=>"000111111",
  28059=>"000000100",
  28060=>"000111000",
  28061=>"001000000",
  28062=>"010100110",
  28063=>"101101110",
  28064=>"001100111",
  28065=>"000010111",
  28066=>"000000111",
  28067=>"000110111",
  28068=>"101110010",
  28069=>"001111111",
  28070=>"111000110",
  28071=>"000110111",
  28072=>"101000010",
  28073=>"110110000",
  28074=>"101100110",
  28075=>"100011110",
  28076=>"100000000",
  28077=>"000101111",
  28078=>"001011110",
  28079=>"001011111",
  28080=>"000111111",
  28081=>"001000101",
  28082=>"001010000",
  28083=>"011011111",
  28084=>"011111101",
  28085=>"000111000",
  28086=>"100000011",
  28087=>"110000011",
  28088=>"010001101",
  28089=>"001101010",
  28090=>"001101000",
  28091=>"000000000",
  28092=>"111000111",
  28093=>"111000110",
  28094=>"100001101",
  28095=>"000111111",
  28096=>"000111011",
  28097=>"100000000",
  28098=>"000101110",
  28099=>"000010111",
  28100=>"000000000",
  28101=>"001111100",
  28102=>"111010010",
  28103=>"000000110",
  28104=>"111100101",
  28105=>"000000111",
  28106=>"000000001",
  28107=>"011010011",
  28108=>"000101010",
  28109=>"101000100",
  28110=>"000010011",
  28111=>"111001000",
  28112=>"000000111",
  28113=>"110001101",
  28114=>"010100000",
  28115=>"001101110",
  28116=>"111000000",
  28117=>"000000000",
  28118=>"000101000",
  28119=>"000101000",
  28120=>"010011001",
  28121=>"001110111",
  28122=>"111011110",
  28123=>"101000000",
  28124=>"111111111",
  28125=>"100000101",
  28126=>"110111110",
  28127=>"101110000",
  28128=>"011000100",
  28129=>"001011111",
  28130=>"000000001",
  28131=>"001000111",
  28132=>"000110000",
  28133=>"111100100",
  28134=>"101101111",
  28135=>"000101101",
  28136=>"111101111",
  28137=>"111001010",
  28138=>"100100011",
  28139=>"101011010",
  28140=>"000000000",
  28141=>"001001101",
  28142=>"001000100",
  28143=>"001011000",
  28144=>"100000000",
  28145=>"100101011",
  28146=>"001101100",
  28147=>"100110110",
  28148=>"111110001",
  28149=>"101101111",
  28150=>"001001000",
  28151=>"000010000",
  28152=>"000000000",
  28153=>"110011011",
  28154=>"111111111",
  28155=>"111000000",
  28156=>"101111000",
  28157=>"001010011",
  28158=>"101011010",
  28159=>"001001000",
  28160=>"000000000",
  28161=>"000100101",
  28162=>"000111111",
  28163=>"111111111",
  28164=>"001110111",
  28165=>"111001000",
  28166=>"001000000",
  28167=>"011010000",
  28168=>"011111110",
  28169=>"010110101",
  28170=>"011001001",
  28171=>"000000001",
  28172=>"101000111",
  28173=>"000011000",
  28174=>"110110011",
  28175=>"101111111",
  28176=>"111101000",
  28177=>"111111111",
  28178=>"110111010",
  28179=>"001000001",
  28180=>"000010100",
  28181=>"010000010",
  28182=>"100000100",
  28183=>"000000000",
  28184=>"000000000",
  28185=>"000001101",
  28186=>"111011000",
  28187=>"000010011",
  28188=>"000101101",
  28189=>"000000000",
  28190=>"111000000",
  28191=>"011000001",
  28192=>"010110100",
  28193=>"010000000",
  28194=>"010000100",
  28195=>"000000110",
  28196=>"011111110",
  28197=>"000000000",
  28198=>"111000000",
  28199=>"110111111",
  28200=>"111110000",
  28201=>"101101101",
  28202=>"101101111",
  28203=>"111111111",
  28204=>"001001001",
  28205=>"010000000",
  28206=>"111000001",
  28207=>"000000000",
  28208=>"000000000",
  28209=>"111111111",
  28210=>"111011100",
  28211=>"000011011",
  28212=>"001000100",
  28213=>"111111111",
  28214=>"111001000",
  28215=>"000000110",
  28216=>"111100000",
  28217=>"000000100",
  28218=>"000101101",
  28219=>"000010111",
  28220=>"001011111",
  28221=>"000001001",
  28222=>"011111101",
  28223=>"111111011",
  28224=>"111000000",
  28225=>"100000000",
  28226=>"111111001",
  28227=>"111111111",
  28228=>"000010000",
  28229=>"000000111",
  28230=>"111010010",
  28231=>"011011111",
  28232=>"000000000",
  28233=>"111111010",
  28234=>"000011101",
  28235=>"010111000",
  28236=>"000001111",
  28237=>"111111111",
  28238=>"111111010",
  28239=>"000000000",
  28240=>"111111001",
  28241=>"110111111",
  28242=>"111111110",
  28243=>"001000000",
  28244=>"111111111",
  28245=>"000001011",
  28246=>"000001000",
  28247=>"101101111",
  28248=>"011001101",
  28249=>"101111001",
  28250=>"000000100",
  28251=>"000010011",
  28252=>"111111000",
  28253=>"001001001",
  28254=>"000111111",
  28255=>"111111111",
  28256=>"110010000",
  28257=>"111100000",
  28258=>"000010000",
  28259=>"000000000",
  28260=>"000110100",
  28261=>"000000001",
  28262=>"110000000",
  28263=>"000111111",
  28264=>"111111100",
  28265=>"000000001",
  28266=>"111001000",
  28267=>"000111001",
  28268=>"101011000",
  28269=>"000000000",
  28270=>"011000000",
  28271=>"000000000",
  28272=>"110110100",
  28273=>"000000101",
  28274=>"011000110",
  28275=>"111111111",
  28276=>"101110110",
  28277=>"000000000",
  28278=>"111111111",
  28279=>"101111111",
  28280=>"000000001",
  28281=>"000000101",
  28282=>"000000111",
  28283=>"101111000",
  28284=>"100110110",
  28285=>"100001001",
  28286=>"111111110",
  28287=>"111111110",
  28288=>"000101010",
  28289=>"111000000",
  28290=>"111111111",
  28291=>"101001101",
  28292=>"110000110",
  28293=>"001011000",
  28294=>"001011001",
  28295=>"100001011",
  28296=>"011011011",
  28297=>"111110100",
  28298=>"011011000",
  28299=>"001111111",
  28300=>"111111001",
  28301=>"011010010",
  28302=>"000000000",
  28303=>"111111100",
  28304=>"011111111",
  28305=>"110101000",
  28306=>"111111111",
  28307=>"000000000",
  28308=>"000011111",
  28309=>"101100111",
  28310=>"111001000",
  28311=>"110000000",
  28312=>"100000000",
  28313=>"000001111",
  28314=>"010111111",
  28315=>"000010000",
  28316=>"010011001",
  28317=>"000100000",
  28318=>"111000000",
  28319=>"000000000",
  28320=>"000100000",
  28321=>"000111111",
  28322=>"111111111",
  28323=>"010100001",
  28324=>"010101101",
  28325=>"001000000",
  28326=>"001001111",
  28327=>"001001000",
  28328=>"111000001",
  28329=>"001000010",
  28330=>"000010000",
  28331=>"111110101",
  28332=>"101000101",
  28333=>"111110111",
  28334=>"011001000",
  28335=>"011111101",
  28336=>"111110000",
  28337=>"011001000",
  28338=>"001000000",
  28339=>"000010110",
  28340=>"100000111",
  28341=>"100011111",
  28342=>"100100000",
  28343=>"100000111",
  28344=>"000100011",
  28345=>"001100111",
  28346=>"111101000",
  28347=>"001111111",
  28348=>"000110111",
  28349=>"111111111",
  28350=>"111111110",
  28351=>"010101000",
  28352=>"001001111",
  28353=>"011010000",
  28354=>"100100111",
  28355=>"000110110",
  28356=>"000000000",
  28357=>"000000001",
  28358=>"110111000",
  28359=>"010111011",
  28360=>"001001110",
  28361=>"000000000",
  28362=>"001111010",
  28363=>"000000111",
  28364=>"111111011",
  28365=>"000011011",
  28366=>"000000000",
  28367=>"011110010",
  28368=>"000011111",
  28369=>"011011001",
  28370=>"111000000",
  28371=>"011011111",
  28372=>"111110010",
  28373=>"111100001",
  28374=>"101000000",
  28375=>"001000111",
  28376=>"010111111",
  28377=>"000111111",
  28378=>"000000000",
  28379=>"000011011",
  28380=>"011000110",
  28381=>"000011111",
  28382=>"010001111",
  28383=>"011110110",
  28384=>"111111000",
  28385=>"011000001",
  28386=>"110110110",
  28387=>"111110110",
  28388=>"111000000",
  28389=>"101101111",
  28390=>"000000001",
  28391=>"011101000",
  28392=>"111111011",
  28393=>"110100111",
  28394=>"110100000",
  28395=>"000001111",
  28396=>"111001000",
  28397=>"001001111",
  28398=>"010000000",
  28399=>"000010010",
  28400=>"000000100",
  28401=>"000000001",
  28402=>"000000101",
  28403=>"001011100",
  28404=>"110001000",
  28405=>"111111111",
  28406=>"111111011",
  28407=>"000000011",
  28408=>"000000001",
  28409=>"000000000",
  28410=>"000001100",
  28411=>"000000010",
  28412=>"011111010",
  28413=>"101111011",
  28414=>"100100000",
  28415=>"000000100",
  28416=>"101111011",
  28417=>"000000000",
  28418=>"010110110",
  28419=>"111000000",
  28420=>"001111111",
  28421=>"000000110",
  28422=>"000000001",
  28423=>"011110111",
  28424=>"000000000",
  28425=>"001000111",
  28426=>"011000100",
  28427=>"111111111",
  28428=>"010010000",
  28429=>"111111001",
  28430=>"111101111",
  28431=>"000111110",
  28432=>"111011000",
  28433=>"101000110",
  28434=>"000000110",
  28435=>"000000001",
  28436=>"111101111",
  28437=>"000010010",
  28438=>"000000111",
  28439=>"111110110",
  28440=>"000000111",
  28441=>"000010000",
  28442=>"101111111",
  28443=>"110111111",
  28444=>"100111011",
  28445=>"101101000",
  28446=>"101111011",
  28447=>"000000000",
  28448=>"101000111",
  28449=>"111111011",
  28450=>"110000000",
  28451=>"000000000",
  28452=>"111100101",
  28453=>"111011111",
  28454=>"110010010",
  28455=>"110111111",
  28456=>"101010010",
  28457=>"100010111",
  28458=>"111111111",
  28459=>"000000000",
  28460=>"100101111",
  28461=>"000000000",
  28462=>"110010111",
  28463=>"011111111",
  28464=>"111100110",
  28465=>"101001001",
  28466=>"000111000",
  28467=>"101000000",
  28468=>"101101101",
  28469=>"000111101",
  28470=>"000001001",
  28471=>"111001001",
  28472=>"111000010",
  28473=>"000110111",
  28474=>"101000000",
  28475=>"000000000",
  28476=>"111011001",
  28477=>"111111111",
  28478=>"000000100",
  28479=>"100110101",
  28480=>"000011111",
  28481=>"101101111",
  28482=>"100001010",
  28483=>"011111111",
  28484=>"000001000",
  28485=>"000001000",
  28486=>"110011101",
  28487=>"001000000",
  28488=>"111001111",
  28489=>"111111000",
  28490=>"111001001",
  28491=>"000000000",
  28492=>"101100100",
  28493=>"001111111",
  28494=>"111101001",
  28495=>"111010101",
  28496=>"100111111",
  28497=>"111111111",
  28498=>"000000001",
  28499=>"100000101",
  28500=>"000000110",
  28501=>"000011111",
  28502=>"000000010",
  28503=>"110111101",
  28504=>"001110000",
  28505=>"001010000",
  28506=>"111111111",
  28507=>"001001001",
  28508=>"111001000",
  28509=>"100100100",
  28510=>"101000000",
  28511=>"110000011",
  28512=>"000000011",
  28513=>"001011001",
  28514=>"000001101",
  28515=>"011010011",
  28516=>"011111111",
  28517=>"000011101",
  28518=>"110011101",
  28519=>"111110110",
  28520=>"001000000",
  28521=>"111101110",
  28522=>"111000110",
  28523=>"111111111",
  28524=>"111110000",
  28525=>"111011010",
  28526=>"011001000",
  28527=>"001111000",
  28528=>"001001001",
  28529=>"111111111",
  28530=>"011110100",
  28531=>"000000000",
  28532=>"111000000",
  28533=>"000000000",
  28534=>"010110000",
  28535=>"000101111",
  28536=>"000010111",
  28537=>"000000000",
  28538=>"000000000",
  28539=>"111010000",
  28540=>"101101101",
  28541=>"111000101",
  28542=>"111011000",
  28543=>"101101000",
  28544=>"010000000",
  28545=>"000000000",
  28546=>"111101111",
  28547=>"100000010",
  28548=>"111000000",
  28549=>"000010111",
  28550=>"100101111",
  28551=>"100000000",
  28552=>"110011001",
  28553=>"001000000",
  28554=>"111000101",
  28555=>"111111010",
  28556=>"101000100",
  28557=>"100001110",
  28558=>"000100111",
  28559=>"011010000",
  28560=>"100100100",
  28561=>"010111111",
  28562=>"110010000",
  28563=>"111111000",
  28564=>"110100101",
  28565=>"001000111",
  28566=>"011111111",
  28567=>"000100100",
  28568=>"010111111",
  28569=>"010000101",
  28570=>"010110110",
  28571=>"000001111",
  28572=>"001011111",
  28573=>"001101111",
  28574=>"111110001",
  28575=>"011111110",
  28576=>"110110110",
  28577=>"000111111",
  28578=>"111111000",
  28579=>"110100111",
  28580=>"000000111",
  28581=>"000001100",
  28582=>"001110110",
  28583=>"000111111",
  28584=>"001000000",
  28585=>"000000000",
  28586=>"110111111",
  28587=>"011010010",
  28588=>"000000000",
  28589=>"111000000",
  28590=>"111011000",
  28591=>"111000000",
  28592=>"011011000",
  28593=>"101011100",
  28594=>"101101100",
  28595=>"101001101",
  28596=>"001110110",
  28597=>"101001000",
  28598=>"000000001",
  28599=>"111010001",
  28600=>"010110000",
  28601=>"001001100",
  28602=>"010111101",
  28603=>"000010000",
  28604=>"101100010",
  28605=>"111101101",
  28606=>"000100000",
  28607=>"100101110",
  28608=>"111000000",
  28609=>"110101111",
  28610=>"111111111",
  28611=>"101110001",
  28612=>"100111110",
  28613=>"111100001",
  28614=>"111110000",
  28615=>"101101101",
  28616=>"101000001",
  28617=>"000000000",
  28618=>"110010011",
  28619=>"000000000",
  28620=>"000010111",
  28621=>"101000001",
  28622=>"000000100",
  28623=>"000000000",
  28624=>"010110111",
  28625=>"100111110",
  28626=>"000000000",
  28627=>"011001000",
  28628=>"101111111",
  28629=>"000000110",
  28630=>"111111111",
  28631=>"111000001",
  28632=>"111100001",
  28633=>"000000001",
  28634=>"000000011",
  28635=>"111000000",
  28636=>"011011111",
  28637=>"011010010",
  28638=>"000010000",
  28639=>"111010000",
  28640=>"000111011",
  28641=>"100111001",
  28642=>"111110100",
  28643=>"111111000",
  28644=>"101000010",
  28645=>"111101000",
  28646=>"100111111",
  28647=>"100101000",
  28648=>"000000111",
  28649=>"000000000",
  28650=>"111100100",
  28651=>"001001000",
  28652=>"000111010",
  28653=>"001111000",
  28654=>"000110100",
  28655=>"111000100",
  28656=>"111101000",
  28657=>"111001110",
  28658=>"111000000",
  28659=>"101111111",
  28660=>"101101100",
  28661=>"101000000",
  28662=>"000000000",
  28663=>"111101111",
  28664=>"000111111",
  28665=>"111000000",
  28666=>"101101101",
  28667=>"101111111",
  28668=>"010111111",
  28669=>"101000000",
  28670=>"000000110",
  28671=>"111110111",
  28672=>"011011000",
  28673=>"000111110",
  28674=>"101000110",
  28675=>"000000100",
  28676=>"110110000",
  28677=>"100110000",
  28678=>"111101110",
  28679=>"000000100",
  28680=>"110010000",
  28681=>"001000101",
  28682=>"001110111",
  28683=>"010110111",
  28684=>"000000001",
  28685=>"000000001",
  28686=>"100001010",
  28687=>"111111111",
  28688=>"110110010",
  28689=>"100111111",
  28690=>"000000010",
  28691=>"100101000",
  28692=>"111111111",
  28693=>"111110000",
  28694=>"100100110",
  28695=>"000011110",
  28696=>"110101111",
  28697=>"111111010",
  28698=>"000000001",
  28699=>"100111111",
  28700=>"000001111",
  28701=>"011101111",
  28702=>"111000000",
  28703=>"000101100",
  28704=>"000000010",
  28705=>"000000101",
  28706=>"111111101",
  28707=>"101000000",
  28708=>"000100100",
  28709=>"010001011",
  28710=>"000010111",
  28711=>"111000000",
  28712=>"010010110",
  28713=>"110110110",
  28714=>"111000011",
  28715=>"110110110",
  28716=>"011011111",
  28717=>"101000000",
  28718=>"011110000",
  28719=>"010001000",
  28720=>"010000000",
  28721=>"000101001",
  28722=>"010000000",
  28723=>"111111011",
  28724=>"001000100",
  28725=>"010111111",
  28726=>"111011011",
  28727=>"011011001",
  28728=>"111111110",
  28729=>"011000110",
  28730=>"100110000",
  28731=>"111111000",
  28732=>"011011001",
  28733=>"101101111",
  28734=>"000001101",
  28735=>"111111111",
  28736=>"000110111",
  28737=>"101001010",
  28738=>"000100000",
  28739=>"011011000",
  28740=>"000001111",
  28741=>"000000000",
  28742=>"000000000",
  28743=>"000011101",
  28744=>"001101111",
  28745=>"011110010",
  28746=>"000000000",
  28747=>"111111000",
  28748=>"111101101",
  28749=>"011011000",
  28750=>"000100100",
  28751=>"111111111",
  28752=>"101101101",
  28753=>"101111111",
  28754=>"000000111",
  28755=>"001101010",
  28756=>"010110010",
  28757=>"101111111",
  28758=>"000011001",
  28759=>"001000111",
  28760=>"010101111",
  28761=>"001101011",
  28762=>"101111111",
  28763=>"110110111",
  28764=>"001000101",
  28765=>"001001111",
  28766=>"111111000",
  28767=>"010010000",
  28768=>"111111111",
  28769=>"001111000",
  28770=>"111011000",
  28771=>"111111100",
  28772=>"110111111",
  28773=>"000100100",
  28774=>"010000000",
  28775=>"110001000",
  28776=>"111111110",
  28777=>"000000011",
  28778=>"111010110",
  28779=>"110011111",
  28780=>"111111111",
  28781=>"111111010",
  28782=>"001000100",
  28783=>"011101111",
  28784=>"011001000",
  28785=>"000000111",
  28786=>"111100110",
  28787=>"111010110",
  28788=>"100101010",
  28789=>"100000000",
  28790=>"111101110",
  28791=>"110010001",
  28792=>"010111111",
  28793=>"110000000",
  28794=>"010110111",
  28795=>"100000000",
  28796=>"111101111",
  28797=>"110100000",
  28798=>"011010000",
  28799=>"101101000",
  28800=>"010010010",
  28801=>"000001000",
  28802=>"111011011",
  28803=>"000011011",
  28804=>"001001000",
  28805=>"011110101",
  28806=>"101100100",
  28807=>"010110010",
  28808=>"000111001",
  28809=>"111111111",
  28810=>"111001000",
  28811=>"010011000",
  28812=>"100111011",
  28813=>"110000000",
  28814=>"000111001",
  28815=>"101001011",
  28816=>"110101000",
  28817=>"000010111",
  28818=>"001000111",
  28819=>"000000111",
  28820=>"000111111",
  28821=>"000000001",
  28822=>"111011010",
  28823=>"001011011",
  28824=>"111111111",
  28825=>"111111111",
  28826=>"101000000",
  28827=>"110100000",
  28828=>"111001000",
  28829=>"111111010",
  28830=>"000010100",
  28831=>"010000001",
  28832=>"001001111",
  28833=>"111111111",
  28834=>"000000111",
  28835=>"111011111",
  28836=>"111111000",
  28837=>"010111110",
  28838=>"011101111",
  28839=>"000000001",
  28840=>"111000010",
  28841=>"000110111",
  28842=>"000000000",
  28843=>"000101110",
  28844=>"111111101",
  28845=>"101000000",
  28846=>"111001011",
  28847=>"010010000",
  28848=>"000001101",
  28849=>"011101111",
  28850=>"001000111",
  28851=>"000101110",
  28852=>"100111111",
  28853=>"000111110",
  28854=>"010110100",
  28855=>"000000000",
  28856=>"111110001",
  28857=>"000110111",
  28858=>"110000111",
  28859=>"000111111",
  28860=>"010111100",
  28861=>"100111111",
  28862=>"111010000",
  28863=>"010000100",
  28864=>"110000110",
  28865=>"000000011",
  28866=>"000110111",
  28867=>"100101010",
  28868=>"110111001",
  28869=>"110100101",
  28870=>"000000111",
  28871=>"001000001",
  28872=>"110000000",
  28873=>"000111001",
  28874=>"000000001",
  28875=>"110111110",
  28876=>"111111010",
  28877=>"010111110",
  28878=>"111110010",
  28879=>"000000000",
  28880=>"111110000",
  28881=>"111110011",
  28882=>"111100110",
  28883=>"000000101",
  28884=>"101000000",
  28885=>"100100110",
  28886=>"000000000",
  28887=>"000001111",
  28888=>"000000111",
  28889=>"000000000",
  28890=>"000000101",
  28891=>"101100000",
  28892=>"011011101",
  28893=>"010110010",
  28894=>"110110010",
  28895=>"011000000",
  28896=>"001101101",
  28897=>"001000000",
  28898=>"000000100",
  28899=>"101010000",
  28900=>"000000000",
  28901=>"000111101",
  28902=>"010011000",
  28903=>"010011000",
  28904=>"000000010",
  28905=>"000000001",
  28906=>"100111110",
  28907=>"000110111",
  28908=>"000000111",
  28909=>"000100101",
  28910=>"000000000",
  28911=>"001111000",
  28912=>"000010010",
  28913=>"011100111",
  28914=>"111110011",
  28915=>"111111111",
  28916=>"100100100",
  28917=>"111111101",
  28918=>"000011011",
  28919=>"111111111",
  28920=>"010011111",
  28921=>"101000110",
  28922=>"111111111",
  28923=>"000001001",
  28924=>"000000000",
  28925=>"000111110",
  28926=>"100010000",
  28927=>"000000101",
  28928=>"111001001",
  28929=>"110111000",
  28930=>"001110000",
  28931=>"001001000",
  28932=>"000011010",
  28933=>"011111000",
  28934=>"111100110",
  28935=>"100000011",
  28936=>"011010000",
  28937=>"000000001",
  28938=>"111000000",
  28939=>"000000000",
  28940=>"001011000",
  28941=>"001111010",
  28942=>"101100001",
  28943=>"001100000",
  28944=>"111111011",
  28945=>"000000111",
  28946=>"110110100",
  28947=>"000100010",
  28948=>"100011111",
  28949=>"010111010",
  28950=>"110110111",
  28951=>"111101111",
  28952=>"101100101",
  28953=>"101100100",
  28954=>"011111011",
  28955=>"111111100",
  28956=>"101110110",
  28957=>"100100110",
  28958=>"111111101",
  28959=>"000110011",
  28960=>"000000000",
  28961=>"011011000",
  28962=>"101001000",
  28963=>"110000100",
  28964=>"011011011",
  28965=>"011001000",
  28966=>"010111010",
  28967=>"111101000",
  28968=>"010000000",
  28969=>"110111100",
  28970=>"000010000",
  28971=>"000000000",
  28972=>"111111011",
  28973=>"101001011",
  28974=>"101011001",
  28975=>"000000000",
  28976=>"000000111",
  28977=>"100100000",
  28978=>"111010001",
  28979=>"010111111",
  28980=>"011111111",
  28981=>"000000000",
  28982=>"100011011",
  28983=>"001000001",
  28984=>"001011110",
  28985=>"000111010",
  28986=>"000010000",
  28987=>"010011011",
  28988=>"011101100",
  28989=>"110111111",
  28990=>"000000001",
  28991=>"100000110",
  28992=>"011101111",
  28993=>"111111111",
  28994=>"010010000",
  28995=>"001000010",
  28996=>"111111111",
  28997=>"000000100",
  28998=>"111111010",
  28999=>"000111011",
  29000=>"000100000",
  29001=>"000000000",
  29002=>"000000001",
  29003=>"111000000",
  29004=>"111111111",
  29005=>"101111111",
  29006=>"011111101",
  29007=>"111011000",
  29008=>"001111111",
  29009=>"110111111",
  29010=>"111111111",
  29011=>"111111111",
  29012=>"111111101",
  29013=>"101110111",
  29014=>"111011101",
  29015=>"001000000",
  29016=>"000000000",
  29017=>"011110110",
  29018=>"100100101",
  29019=>"010110010",
  29020=>"000000100",
  29021=>"111001001",
  29022=>"111111111",
  29023=>"101000011",
  29024=>"111111111",
  29025=>"111000000",
  29026=>"010010010",
  29027=>"111011101",
  29028=>"111111111",
  29029=>"111100001",
  29030=>"000001000",
  29031=>"110100111",
  29032=>"000000000",
  29033=>"111011000",
  29034=>"010010110",
  29035=>"111111000",
  29036=>"111111111",
  29037=>"100001000",
  29038=>"011001000",
  29039=>"111111111",
  29040=>"101001001",
  29041=>"100011000",
  29042=>"000100110",
  29043=>"100000111",
  29044=>"000000011",
  29045=>"000000001",
  29046=>"000111100",
  29047=>"001100001",
  29048=>"010000000",
  29049=>"111111000",
  29050=>"011000111",
  29051=>"000000110",
  29052=>"011101111",
  29053=>"001000000",
  29054=>"000001111",
  29055=>"101000111",
  29056=>"111111101",
  29057=>"000000000",
  29058=>"111101000",
  29059=>"111110000",
  29060=>"111111011",
  29061=>"011011111",
  29062=>"110111000",
  29063=>"111100110",
  29064=>"100100100",
  29065=>"111011111",
  29066=>"100111100",
  29067=>"001000000",
  29068=>"000000011",
  29069=>"000000100",
  29070=>"100000110",
  29071=>"011000001",
  29072=>"000011110",
  29073=>"000010010",
  29074=>"111000011",
  29075=>"001000011",
  29076=>"111101001",
  29077=>"000111011",
  29078=>"011111011",
  29079=>"000011011",
  29080=>"000000000",
  29081=>"111111000",
  29082=>"000101001",
  29083=>"101000000",
  29084=>"000111111",
  29085=>"111001011",
  29086=>"000001111",
  29087=>"010010000",
  29088=>"000000000",
  29089=>"000111101",
  29090=>"110000101",
  29091=>"111111000",
  29092=>"011110101",
  29093=>"010011011",
  29094=>"100000100",
  29095=>"111111101",
  29096=>"111011011",
  29097=>"000111010",
  29098=>"000000000",
  29099=>"000000000",
  29100=>"100100110",
  29101=>"011111111",
  29102=>"101001001",
  29103=>"111111110",
  29104=>"000010000",
  29105=>"000000000",
  29106=>"110110100",
  29107=>"111011011",
  29108=>"100101000",
  29109=>"000000000",
  29110=>"011000000",
  29111=>"100000000",
  29112=>"100110101",
  29113=>"111000001",
  29114=>"001111011",
  29115=>"111000000",
  29116=>"100000001",
  29117=>"010010010",
  29118=>"111001001",
  29119=>"000000000",
  29120=>"101100100",
  29121=>"101000011",
  29122=>"111000011",
  29123=>"110110111",
  29124=>"011001001",
  29125=>"111100000",
  29126=>"011011000",
  29127=>"100100000",
  29128=>"110000100",
  29129=>"000011011",
  29130=>"010100000",
  29131=>"111011000",
  29132=>"101100000",
  29133=>"111111111",
  29134=>"000101111",
  29135=>"000000000",
  29136=>"111100111",
  29137=>"010110110",
  29138=>"000010101",
  29139=>"010010000",
  29140=>"101001111",
  29141=>"100100110",
  29142=>"010111111",
  29143=>"101011111",
  29144=>"000000000",
  29145=>"010000010",
  29146=>"100000000",
  29147=>"000000000",
  29148=>"111111110",
  29149=>"100000000",
  29150=>"000001001",
  29151=>"001111101",
  29152=>"100000100",
  29153=>"000100101",
  29154=>"000000101",
  29155=>"110101001",
  29156=>"111101000",
  29157=>"100100110",
  29158=>"001000000",
  29159=>"101101100",
  29160=>"110111101",
  29161=>"111100111",
  29162=>"110000000",
  29163=>"000000010",
  29164=>"000000001",
  29165=>"000101101",
  29166=>"111010110",
  29167=>"001000101",
  29168=>"000000000",
  29169=>"101001011",
  29170=>"111111000",
  29171=>"011011011",
  29172=>"111101101",
  29173=>"000000011",
  29174=>"111011010",
  29175=>"111111101",
  29176=>"011001000",
  29177=>"000001011",
  29178=>"000010000",
  29179=>"101101101",
  29180=>"000111111",
  29181=>"111001111",
  29182=>"110110010",
  29183=>"110000000",
  29184=>"011101100",
  29185=>"100000011",
  29186=>"000101111",
  29187=>"000000110",
  29188=>"011011111",
  29189=>"110111011",
  29190=>"111011010",
  29191=>"110011111",
  29192=>"010000101",
  29193=>"111000001",
  29194=>"011000000",
  29195=>"011001111",
  29196=>"110001111",
  29197=>"011001000",
  29198=>"011000010",
  29199=>"110000110",
  29200=>"111101000",
  29201=>"101100000",
  29202=>"000000000",
  29203=>"111111000",
  29204=>"010110111",
  29205=>"001111110",
  29206=>"000110110",
  29207=>"111110100",
  29208=>"000110000",
  29209=>"111110010",
  29210=>"000111111",
  29211=>"001101011",
  29212=>"110011010",
  29213=>"000001100",
  29214=>"000011011",
  29215=>"010000000",
  29216=>"000000000",
  29217=>"000001110",
  29218=>"010000000",
  29219=>"110011000",
  29220=>"100001000",
  29221=>"100101110",
  29222=>"000010110",
  29223=>"110110000",
  29224=>"111111111",
  29225=>"001001011",
  29226=>"010000000",
  29227=>"000111000",
  29228=>"010100011",
  29229=>"110111111",
  29230=>"111110111",
  29231=>"100000111",
  29232=>"000000000",
  29233=>"111111111",
  29234=>"000001001",
  29235=>"111111000",
  29236=>"001000000",
  29237=>"111010110",
  29238=>"100000101",
  29239=>"111111000",
  29240=>"100111111",
  29241=>"110010000",
  29242=>"111000000",
  29243=>"111011011",
  29244=>"110010110",
  29245=>"111010010",
  29246=>"001000000",
  29247=>"001110110",
  29248=>"111000011",
  29249=>"100100110",
  29250=>"000001000",
  29251=>"001100111",
  29252=>"010000000",
  29253=>"011010000",
  29254=>"110010000",
  29255=>"010010101",
  29256=>"010011110",
  29257=>"010000010",
  29258=>"101000000",
  29259=>"111100000",
  29260=>"000000001",
  29261=>"001111111",
  29262=>"111111110",
  29263=>"000001100",
  29264=>"001000111",
  29265=>"101001000",
  29266=>"011101000",
  29267=>"001100000",
  29268=>"010010001",
  29269=>"100001011",
  29270=>"100100100",
  29271=>"110001011",
  29272=>"101100111",
  29273=>"011011011",
  29274=>"001001110",
  29275=>"110100100",
  29276=>"000001111",
  29277=>"001001001",
  29278=>"000111111",
  29279=>"100001111",
  29280=>"000000111",
  29281=>"000000100",
  29282=>"000000111",
  29283=>"100110110",
  29284=>"111110100",
  29285=>"000011001",
  29286=>"001111110",
  29287=>"010010000",
  29288=>"011110011",
  29289=>"010010010",
  29290=>"100100111",
  29291=>"110000001",
  29292=>"000100111",
  29293=>"111111000",
  29294=>"001001000",
  29295=>"010010000",
  29296=>"011001011",
  29297=>"111001000",
  29298=>"111101001",
  29299=>"110011000",
  29300=>"000010010",
  29301=>"101001000",
  29302=>"110000100",
  29303=>"000000001",
  29304=>"000010110",
  29305=>"111010000",
  29306=>"111001001",
  29307=>"001111101",
  29308=>"110011011",
  29309=>"100000000",
  29310=>"101111111",
  29311=>"111000101",
  29312=>"000000000",
  29313=>"101100111",
  29314=>"010011111",
  29315=>"000111111",
  29316=>"011111111",
  29317=>"000000100",
  29318=>"101111010",
  29319=>"000000000",
  29320=>"111101100",
  29321=>"000000000",
  29322=>"111000000",
  29323=>"000000110",
  29324=>"111111111",
  29325=>"000000000",
  29326=>"001111000",
  29327=>"001000000",
  29328=>"011100110",
  29329=>"111000110",
  29330=>"111011011",
  29331=>"010111101",
  29332=>"101010100",
  29333=>"101000000",
  29334=>"111000111",
  29335=>"100000001",
  29336=>"011001000",
  29337=>"000010111",
  29338=>"001000111",
  29339=>"001001111",
  29340=>"010011011",
  29341=>"001101101",
  29342=>"010000010",
  29343=>"111010000",
  29344=>"110100111",
  29345=>"101101000",
  29346=>"101000000",
  29347=>"101101110",
  29348=>"001111000",
  29349=>"110010000",
  29350=>"110111010",
  29351=>"000001001",
  29352=>"111111111",
  29353=>"000000110",
  29354=>"001111111",
  29355=>"001000000",
  29356=>"000001000",
  29357=>"000110000",
  29358=>"101011011",
  29359=>"111000000",
  29360=>"001000101",
  29361=>"111111011",
  29362=>"000100000",
  29363=>"000000010",
  29364=>"110111011",
  29365=>"111011010",
  29366=>"111000000",
  29367=>"110111000",
  29368=>"011000001",
  29369=>"010110000",
  29370=>"000000111",
  29371=>"111000010",
  29372=>"101000010",
  29373=>"101000111",
  29374=>"000001111",
  29375=>"000011000",
  29376=>"010000000",
  29377=>"111010000",
  29378=>"000101010",
  29379=>"011000100",
  29380=>"000010000",
  29381=>"100001111",
  29382=>"011111011",
  29383=>"111000001",
  29384=>"111010011",
  29385=>"111101100",
  29386=>"100000000",
  29387=>"000100111",
  29388=>"011000010",
  29389=>"011110110",
  29390=>"111010000",
  29391=>"110001111",
  29392=>"010000000",
  29393=>"011001011",
  29394=>"011010010",
  29395=>"011010000",
  29396=>"010000111",
  29397=>"101100110",
  29398=>"001000111",
  29399=>"000000000",
  29400=>"110010000",
  29401=>"001111001",
  29402=>"001001000",
  29403=>"101100001",
  29404=>"000110110",
  29405=>"000010111",
  29406=>"111010000",
  29407=>"101110101",
  29408=>"000001101",
  29409=>"100111110",
  29410=>"000111111",
  29411=>"100101010",
  29412=>"110100000",
  29413=>"011000000",
  29414=>"010010000",
  29415=>"101101001",
  29416=>"000000000",
  29417=>"010010101",
  29418=>"000000001",
  29419=>"101000000",
  29420=>"000001111",
  29421=>"000110000",
  29422=>"011000001",
  29423=>"111111000",
  29424=>"111000000",
  29425=>"000001111",
  29426=>"010111111",
  29427=>"111000000",
  29428=>"110001011",
  29429=>"011011111",
  29430=>"111000000",
  29431=>"110101111",
  29432=>"000000000",
  29433=>"000010000",
  29434=>"001101000",
  29435=>"011111110",
  29436=>"011000000",
  29437=>"001101111",
  29438=>"110111101",
  29439=>"100001000",
  29440=>"100011010",
  29441=>"000010110",
  29442=>"011001001",
  29443=>"111111001",
  29444=>"101000011",
  29445=>"000001110",
  29446=>"111001011",
  29447=>"000110110",
  29448=>"000001110",
  29449=>"011001011",
  29450=>"100001000",
  29451=>"000000100",
  29452=>"000000100",
  29453=>"000000000",
  29454=>"100000111",
  29455=>"011001000",
  29456=>"000110110",
  29457=>"011001001",
  29458=>"110011000",
  29459=>"011000000",
  29460=>"001111100",
  29461=>"111101100",
  29462=>"011011010",
  29463=>"111001110",
  29464=>"010001001",
  29465=>"011111100",
  29466=>"100001001",
  29467=>"100100100",
  29468=>"011111001",
  29469=>"010000001",
  29470=>"100110110",
  29471=>"100100000",
  29472=>"100001000",
  29473=>"001100110",
  29474=>"111011001",
  29475=>"001110100",
  29476=>"100010101",
  29477=>"010111001",
  29478=>"000000000",
  29479=>"100110000",
  29480=>"011001111",
  29481=>"010110110",
  29482=>"011000010",
  29483=>"111001001",
  29484=>"100100101",
  29485=>"100110101",
  29486=>"110111000",
  29487=>"011001000",
  29488=>"111011010",
  29489=>"000011011",
  29490=>"011100000",
  29491=>"110100001",
  29492=>"011011001",
  29493=>"111111101",
  29494=>"000000000",
  29495=>"100110100",
  29496=>"100100000",
  29497=>"000000110",
  29498=>"000001000",
  29499=>"001011111",
  29500=>"011011111",
  29501=>"000110001",
  29502=>"000001001",
  29503=>"101110110",
  29504=>"011001100",
  29505=>"000100110",
  29506=>"010000100",
  29507=>"010110110",
  29508=>"000011000",
  29509=>"000000011",
  29510=>"111001001",
  29511=>"011110100",
  29512=>"111111110",
  29513=>"100010000",
  29514=>"000110110",
  29515=>"111000111",
  29516=>"110110100",
  29517=>"000000000",
  29518=>"000000000",
  29519=>"111111101",
  29520=>"110010011",
  29521=>"100111111",
  29522=>"001001100",
  29523=>"010011000",
  29524=>"000011001",
  29525=>"111001111",
  29526=>"010011100",
  29527=>"000001011",
  29528=>"111011100",
  29529=>"001001110",
  29530=>"110000000",
  29531=>"100110110",
  29532=>"100100000",
  29533=>"100010000",
  29534=>"111100001",
  29535=>"110111111",
  29536=>"000000000",
  29537=>"110001011",
  29538=>"111001001",
  29539=>"101111011",
  29540=>"000100110",
  29541=>"001001000",
  29542=>"100110000",
  29543=>"111001001",
  29544=>"100011000",
  29545=>"110001000",
  29546=>"001001100",
  29547=>"110110000",
  29548=>"110110000",
  29549=>"011001011",
  29550=>"110001001",
  29551=>"000000100",
  29552=>"100111111",
  29553=>"100000100",
  29554=>"000000110",
  29555=>"000000011",
  29556=>"110110000",
  29557=>"010001000",
  29558=>"010000100",
  29559=>"001001000",
  29560=>"111001001",
  29561=>"110111110",
  29562=>"111001001",
  29563=>"000001111",
  29564=>"011001100",
  29565=>"100000100",
  29566=>"101111011",
  29567=>"100110001",
  29568=>"110111001",
  29569=>"000110110",
  29570=>"111111100",
  29571=>"010011110",
  29572=>"100101100",
  29573=>"000000111",
  29574=>"000100010",
  29575=>"000010110",
  29576=>"000100000",
  29577=>"110100000",
  29578=>"011001001",
  29579=>"011111011",
  29580=>"111001001",
  29581=>"011001001",
  29582=>"111101101",
  29583=>"011001011",
  29584=>"100111101",
  29585=>"100110010",
  29586=>"011001011",
  29587=>"110110000",
  29588=>"110010100",
  29589=>"111000010",
  29590=>"100100100",
  29591=>"000111100",
  29592=>"111100100",
  29593=>"000100110",
  29594=>"011001001",
  29595=>"011001001",
  29596=>"110100000",
  29597=>"111000001",
  29598=>"110110010",
  29599=>"000100110",
  29600=>"011011111",
  29601=>"001001011",
  29602=>"000110110",
  29603=>"000011110",
  29604=>"100100000",
  29605=>"101101100",
  29606=>"010110000",
  29607=>"010110000",
  29608=>"011001000",
  29609=>"010100111",
  29610=>"011001001",
  29611=>"000001000",
  29612=>"111101001",
  29613=>"110000000",
  29614=>"001000000",
  29615=>"101001011",
  29616=>"101000000",
  29617=>"110110001",
  29618=>"110000111",
  29619=>"010001101",
  29620=>"100110101",
  29621=>"001001011",
  29622=>"000001001",
  29623=>"010001001",
  29624=>"100000011",
  29625=>"011100101",
  29626=>"111011011",
  29627=>"110110100",
  29628=>"110100001",
  29629=>"011011111",
  29630=>"001001000",
  29631=>"101011000",
  29632=>"111001001",
  29633=>"111001000",
  29634=>"110110100",
  29635=>"010000000",
  29636=>"010011111",
  29637=>"011011001",
  29638=>"000100110",
  29639=>"001001011",
  29640=>"011110001",
  29641=>"001110110",
  29642=>"011010000",
  29643=>"000100000",
  29644=>"010001000",
  29645=>"011111111",
  29646=>"001000000",
  29647=>"111000000",
  29648=>"100001000",
  29649=>"010000100",
  29650=>"000110100",
  29651=>"100110000",
  29652=>"000010011",
  29653=>"100000000",
  29654=>"000110100",
  29655=>"001000111",
  29656=>"110100000",
  29657=>"000101000",
  29658=>"001001001",
  29659=>"011001001",
  29660=>"100001000",
  29661=>"111101001",
  29662=>"001001000",
  29663=>"000101111",
  29664=>"101111111",
  29665=>"110001001",
  29666=>"111011010",
  29667=>"011110110",
  29668=>"011000011",
  29669=>"100110110",
  29670=>"110000001",
  29671=>"000001011",
  29672=>"101001110",
  29673=>"011001011",
  29674=>"111001001",
  29675=>"011001001",
  29676=>"000110110",
  29677=>"110011000",
  29678=>"000000110",
  29679=>"000111111",
  29680=>"000000001",
  29681=>"011000001",
  29682=>"010110110",
  29683=>"000000100",
  29684=>"110001011",
  29685=>"100001001",
  29686=>"010001010",
  29687=>"101001000",
  29688=>"100001111",
  29689=>"110110111",
  29690=>"110111111",
  29691=>"010111101",
  29692=>"111011101",
  29693=>"001001000",
  29694=>"000011110",
  29695=>"111011101",
  29696=>"111011111",
  29697=>"000111111",
  29698=>"000010000",
  29699=>"110000000",
  29700=>"010100001",
  29701=>"011000000",
  29702=>"010010101",
  29703=>"111101001",
  29704=>"000000101",
  29705=>"111111000",
  29706=>"110010100",
  29707=>"101111010",
  29708=>"001000000",
  29709=>"010000000",
  29710=>"001001011",
  29711=>"000110110",
  29712=>"101111111",
  29713=>"000000000",
  29714=>"000000111",
  29715=>"111100111",
  29716=>"110101001",
  29717=>"000000000",
  29718=>"111111111",
  29719=>"010110111",
  29720=>"100000010",
  29721=>"010001101",
  29722=>"111111111",
  29723=>"111111000",
  29724=>"100000100",
  29725=>"010000000",
  29726=>"111100010",
  29727=>"011111010",
  29728=>"000000000",
  29729=>"000011001",
  29730=>"001101000",
  29731=>"011100000",
  29732=>"000000100",
  29733=>"101001111",
  29734=>"000010110",
  29735=>"111111111",
  29736=>"110111111",
  29737=>"100000001",
  29738=>"101100010",
  29739=>"000000000",
  29740=>"111110000",
  29741=>"110111111",
  29742=>"111111101",
  29743=>"000000000",
  29744=>"111111111",
  29745=>"011001110",
  29746=>"000000101",
  29747=>"101000000",
  29748=>"000001001",
  29749=>"000000000",
  29750=>"100001001",
  29751=>"111111110",
  29752=>"101111001",
  29753=>"000000110",
  29754=>"000000100",
  29755=>"010110000",
  29756=>"011010011",
  29757=>"111111111",
  29758=>"000001111",
  29759=>"011111011",
  29760=>"111011011",
  29761=>"100100111",
  29762=>"111111110",
  29763=>"001000101",
  29764=>"111111111",
  29765=>"111101000",
  29766=>"100000111",
  29767=>"101101101",
  29768=>"011111110",
  29769=>"000000000",
  29770=>"000000000",
  29771=>"001000101",
  29772=>"101000100",
  29773=>"000000000",
  29774=>"000000000",
  29775=>"111111111",
  29776=>"011111011",
  29777=>"000000000",
  29778=>"001101110",
  29779=>"111110110",
  29780=>"000001001",
  29781=>"110000111",
  29782=>"110110001",
  29783=>"010010000",
  29784=>"110000000",
  29785=>"100111110",
  29786=>"001011111",
  29787=>"110111111",
  29788=>"101111111",
  29789=>"000000011",
  29790=>"000000000",
  29791=>"110010111",
  29792=>"111111111",
  29793=>"111111011",
  29794=>"001001000",
  29795=>"010110110",
  29796=>"000000111",
  29797=>"101111111",
  29798=>"111110100",
  29799=>"000100100",
  29800=>"111000010",
  29801=>"000010010",
  29802=>"111001011",
  29803=>"111111101",
  29804=>"000101011",
  29805=>"000000000",
  29806=>"111000000",
  29807=>"110110100",
  29808=>"110110111",
  29809=>"000010011",
  29810=>"001101100",
  29811=>"111110000",
  29812=>"101001111",
  29813=>"000000000",
  29814=>"011000000",
  29815=>"011111000",
  29816=>"110100000",
  29817=>"100001100",
  29818=>"010111011",
  29819=>"000000000",
  29820=>"000111011",
  29821=>"100000000",
  29822=>"000101001",
  29823=>"000100111",
  29824=>"101111011",
  29825=>"010110000",
  29826=>"111110110",
  29827=>"100100111",
  29828=>"100101111",
  29829=>"000001110",
  29830=>"101100100",
  29831=>"100110000",
  29832=>"001001110",
  29833=>"001011010",
  29834=>"000001100",
  29835=>"001111101",
  29836=>"000101010",
  29837=>"011000000",
  29838=>"000000111",
  29839=>"111001011",
  29840=>"000000011",
  29841=>"000111111",
  29842=>"000000111",
  29843=>"000000000",
  29844=>"010111010",
  29845=>"001000000",
  29846=>"000000110",
  29847=>"000101110",
  29848=>"011000000",
  29849=>"101000000",
  29850=>"000111101",
  29851=>"000001000",
  29852=>"111101000",
  29853=>"110111010",
  29854=>"100101001",
  29855=>"000000001",
  29856=>"010011111",
  29857=>"000111010",
  29858=>"000001110",
  29859=>"010000111",
  29860=>"111000010",
  29861=>"011111111",
  29862=>"111000110",
  29863=>"110010100",
  29864=>"111111000",
  29865=>"000111100",
  29866=>"111111111",
  29867=>"000000000",
  29868=>"000000000",
  29869=>"010111111",
  29870=>"011111011",
  29871=>"100110001",
  29872=>"000000111",
  29873=>"000000000",
  29874=>"000000000",
  29875=>"000111111",
  29876=>"110110100",
  29877=>"000000000",
  29878=>"110000011",
  29879=>"000110111",
  29880=>"111010000",
  29881=>"111000000",
  29882=>"111101111",
  29883=>"111011101",
  29884=>"000011101",
  29885=>"000001010",
  29886=>"110110110",
  29887=>"000000001",
  29888=>"010000000",
  29889=>"011000010",
  29890=>"111101111",
  29891=>"101000101",
  29892=>"000110111",
  29893=>"111000000",
  29894=>"100101000",
  29895=>"111110010",
  29896=>"111000001",
  29897=>"100100111",
  29898=>"100101111",
  29899=>"000001101",
  29900=>"000000000",
  29901=>"101011111",
  29902=>"101001001",
  29903=>"111111011",
  29904=>"111000000",
  29905=>"011111111",
  29906=>"111111101",
  29907=>"111111000",
  29908=>"000000101",
  29909=>"001000111",
  29910=>"111101111",
  29911=>"000001010",
  29912=>"000001111",
  29913=>"000001011",
  29914=>"000110011",
  29915=>"000111000",
  29916=>"111011011",
  29917=>"110110010",
  29918=>"000010011",
  29919=>"110111011",
  29920=>"001111100",
  29921=>"001000111",
  29922=>"111111101",
  29923=>"001011111",
  29924=>"101000001",
  29925=>"111000011",
  29926=>"000001000",
  29927=>"010011001",
  29928=>"010001000",
  29929=>"000000000",
  29930=>"010011000",
  29931=>"011110000",
  29932=>"111101001",
  29933=>"000101111",
  29934=>"010010000",
  29935=>"000100010",
  29936=>"000000000",
  29937=>"110000111",
  29938=>"111111001",
  29939=>"000000001",
  29940=>"111100100",
  29941=>"000000010",
  29942=>"011100001",
  29943=>"111111111",
  29944=>"101001111",
  29945=>"100001011",
  29946=>"010001111",
  29947=>"111011000",
  29948=>"101111111",
  29949=>"000001011",
  29950=>"110001101",
  29951=>"011011111",
  29952=>"000010001",
  29953=>"110010010",
  29954=>"000100000",
  29955=>"000000000",
  29956=>"111111111",
  29957=>"110110000",
  29958=>"011111111",
  29959=>"000011111",
  29960=>"000000110",
  29961=>"000101101",
  29962=>"001001110",
  29963=>"000111111",
  29964=>"100010011",
  29965=>"001111011",
  29966=>"001010010",
  29967=>"001101001",
  29968=>"000111111",
  29969=>"111111110",
  29970=>"111001111",
  29971=>"000000100",
  29972=>"001111111",
  29973=>"110101111",
  29974=>"100100011",
  29975=>"000000000",
  29976=>"000000110",
  29977=>"010111111",
  29978=>"011001011",
  29979=>"000001100",
  29980=>"001111111",
  29981=>"000100111",
  29982=>"001011100",
  29983=>"001101001",
  29984=>"000000000",
  29985=>"000111111",
  29986=>"111111000",
  29987=>"111011000",
  29988=>"000111110",
  29989=>"110100100",
  29990=>"010111001",
  29991=>"000000001",
  29992=>"010110000",
  29993=>"110111111",
  29994=>"011000111",
  29995=>"001101101",
  29996=>"000000001",
  29997=>"010111111",
  29998=>"110111010",
  29999=>"010110111",
  30000=>"011010000",
  30001=>"010001101",
  30002=>"100111100",
  30003=>"000000101",
  30004=>"010000101",
  30005=>"101001110",
  30006=>"110100000",
  30007=>"000000110",
  30008=>"111101101",
  30009=>"111001011",
  30010=>"010011010",
  30011=>"111000000",
  30012=>"100110110",
  30013=>"111101111",
  30014=>"000000000",
  30015=>"110111011",
  30016=>"111000010",
  30017=>"111111000",
  30018=>"000000111",
  30019=>"011111100",
  30020=>"000000000",
  30021=>"111111011",
  30022=>"110001001",
  30023=>"111100111",
  30024=>"010110101",
  30025=>"111000000",
  30026=>"000000001",
  30027=>"001000001",
  30028=>"111111111",
  30029=>"111111011",
  30030=>"001100110",
  30031=>"000000111",
  30032=>"000011001",
  30033=>"100111111",
  30034=>"000000001",
  30035=>"010010001",
  30036=>"111110010",
  30037=>"000001111",
  30038=>"110110011",
  30039=>"000111011",
  30040=>"101001000",
  30041=>"000000001",
  30042=>"111100000",
  30043=>"100100111",
  30044=>"000000111",
  30045=>"001000010",
  30046=>"011101111",
  30047=>"000001001",
  30048=>"011010000",
  30049=>"001111100",
  30050=>"100101101",
  30051=>"111000100",
  30052=>"110000010",
  30053=>"000000011",
  30054=>"011010111",
  30055=>"001101000",
  30056=>"010010001",
  30057=>"000011111",
  30058=>"010111000",
  30059=>"010001001",
  30060=>"000110011",
  30061=>"110111011",
  30062=>"011011010",
  30063=>"001111000",
  30064=>"111100101",
  30065=>"100000101",
  30066=>"001000000",
  30067=>"111111111",
  30068=>"100111100",
  30069=>"000000101",
  30070=>"111010000",
  30071=>"111111000",
  30072=>"010000000",
  30073=>"010010111",
  30074=>"000001000",
  30075=>"100110111",
  30076=>"100100010",
  30077=>"011011100",
  30078=>"000000011",
  30079=>"001111000",
  30080=>"000000010",
  30081=>"111111100",
  30082=>"000110111",
  30083=>"101100111",
  30084=>"111111011",
  30085=>"001001011",
  30086=>"111011101",
  30087=>"000001001",
  30088=>"100110001",
  30089=>"101101001",
  30090=>"101110111",
  30091=>"101001111",
  30092=>"010010000",
  30093=>"111000000",
  30094=>"001101111",
  30095=>"001000000",
  30096=>"110111110",
  30097=>"111110000",
  30098=>"000000000",
  30099=>"000000111",
  30100=>"000000000",
  30101=>"010000011",
  30102=>"010010011",
  30103=>"011010000",
  30104=>"011111111",
  30105=>"000000000",
  30106=>"111111000",
  30107=>"001000000",
  30108=>"101000000",
  30109=>"010111011",
  30110=>"000010111",
  30111=>"110010000",
  30112=>"000010010",
  30113=>"111010000",
  30114=>"000010000",
  30115=>"111101000",
  30116=>"000000000",
  30117=>"000110010",
  30118=>"110010001",
  30119=>"000010011",
  30120=>"000000011",
  30121=>"100000000",
  30122=>"110010110",
  30123=>"000111000",
  30124=>"110000101",
  30125=>"000100000",
  30126=>"010010000",
  30127=>"000000111",
  30128=>"111111111",
  30129=>"011111110",
  30130=>"000111111",
  30131=>"000101000",
  30132=>"101010000",
  30133=>"011000000",
  30134=>"111011011",
  30135=>"110111000",
  30136=>"001011001",
  30137=>"010110110",
  30138=>"001000101",
  30139=>"000110110",
  30140=>"001001111",
  30141=>"010111100",
  30142=>"001010011",
  30143=>"111100010",
  30144=>"111101001",
  30145=>"011011111",
  30146=>"110111010",
  30147=>"011011101",
  30148=>"011101000",
  30149=>"000110001",
  30150=>"010000110",
  30151=>"111001000",
  30152=>"000111111",
  30153=>"111000111",
  30154=>"111110111",
  30155=>"000101111",
  30156=>"000111000",
  30157=>"010001110",
  30158=>"111111111",
  30159=>"000100100",
  30160=>"001111101",
  30161=>"011010100",
  30162=>"000000111",
  30163=>"000010010",
  30164=>"111010111",
  30165=>"111111111",
  30166=>"111101001",
  30167=>"000000000",
  30168=>"010000111",
  30169=>"100100110",
  30170=>"001000011",
  30171=>"110011001",
  30172=>"001100101",
  30173=>"111000001",
  30174=>"111000011",
  30175=>"111101110",
  30176=>"101101100",
  30177=>"100000101",
  30178=>"001000010",
  30179=>"100000110",
  30180=>"011000000",
  30181=>"011111000",
  30182=>"100110110",
  30183=>"111001000",
  30184=>"101111011",
  30185=>"111111111",
  30186=>"100100000",
  30187=>"110110010",
  30188=>"000101001",
  30189=>"111110110",
  30190=>"000011011",
  30191=>"110010000",
  30192=>"000000000",
  30193=>"000110110",
  30194=>"001000111",
  30195=>"001000100",
  30196=>"000011110",
  30197=>"111111111",
  30198=>"000100110",
  30199=>"001101101",
  30200=>"000000011",
  30201=>"000010111",
  30202=>"100111111",
  30203=>"000001101",
  30204=>"101000111",
  30205=>"011111100",
  30206=>"011111100",
  30207=>"111010010",
  30208=>"111011011",
  30209=>"000000001",
  30210=>"101100010",
  30211=>"101001000",
  30212=>"100100001",
  30213=>"111001011",
  30214=>"101101100",
  30215=>"111100001",
  30216=>"011000111",
  30217=>"000000111",
  30218=>"011001100",
  30219=>"101011111",
  30220=>"000001011",
  30221=>"000000000",
  30222=>"100100101",
  30223=>"011111111",
  30224=>"000000010",
  30225=>"000000111",
  30226=>"111111000",
  30227=>"000000111",
  30228=>"111110101",
  30229=>"111111111",
  30230=>"111101101",
  30231=>"000010111",
  30232=>"000000001",
  30233=>"010111111",
  30234=>"111000011",
  30235=>"000000011",
  30236=>"000000010",
  30237=>"101011000",
  30238=>"111110000",
  30239=>"000000101",
  30240=>"001010101",
  30241=>"111011001",
  30242=>"000110110",
  30243=>"000010010",
  30244=>"000111110",
  30245=>"010011001",
  30246=>"110010010",
  30247=>"000110110",
  30248=>"000011001",
  30249=>"111111000",
  30250=>"000000110",
  30251=>"011111111",
  30252=>"010000000",
  30253=>"111100000",
  30254=>"111101101",
  30255=>"001101101",
  30256=>"101001000",
  30257=>"000101111",
  30258=>"010000010",
  30259=>"010000111",
  30260=>"010011011",
  30261=>"101000101",
  30262=>"000000011",
  30263=>"000000000",
  30264=>"111101000",
  30265=>"000000000",
  30266=>"000000000",
  30267=>"010000010",
  30268=>"010000001",
  30269=>"010111001",
  30270=>"000000100",
  30271=>"000111111",
  30272=>"000111111",
  30273=>"101000000",
  30274=>"010000000",
  30275=>"110001110",
  30276=>"000000001",
  30277=>"000100101",
  30278=>"000001001",
  30279=>"101111110",
  30280=>"001000000",
  30281=>"111000000",
  30282=>"111111000",
  30283=>"000011001",
  30284=>"000000111",
  30285=>"010000000",
  30286=>"001001101",
  30287=>"101000010",
  30288=>"000000000",
  30289=>"100101011",
  30290=>"111001101",
  30291=>"000000110",
  30292=>"110100111",
  30293=>"001111111",
  30294=>"011011010",
  30295=>"101010111",
  30296=>"010000100",
  30297=>"100000111",
  30298=>"011001101",
  30299=>"110011000",
  30300=>"000111000",
  30301=>"001000000",
  30302=>"000111010",
  30303=>"110100000",
  30304=>"000111111",
  30305=>"001000000",
  30306=>"111000000",
  30307=>"111111110",
  30308=>"000001011",
  30309=>"100111111",
  30310=>"110000011",
  30311=>"111000000",
  30312=>"111111000",
  30313=>"111111001",
  30314=>"111000010",
  30315=>"111000000",
  30316=>"111000000",
  30317=>"101000001",
  30318=>"101001111",
  30319=>"000000001",
  30320=>"111111001",
  30321=>"111101000",
  30322=>"000000110",
  30323=>"000000000",
  30324=>"111100001",
  30325=>"111000100",
  30326=>"001000000",
  30327=>"000110000",
  30328=>"000001000",
  30329=>"111111111",
  30330=>"111111111",
  30331=>"111110010",
  30332=>"010001011",
  30333=>"000100000",
  30334=>"001011011",
  30335=>"000001111",
  30336=>"111111010",
  30337=>"100111000",
  30338=>"000010000",
  30339=>"110111101",
  30340=>"111111011",
  30341=>"100110001",
  30342=>"110100100",
  30343=>"000010111",
  30344=>"110111101",
  30345=>"111111111",
  30346=>"101000111",
  30347=>"110010110",
  30348=>"000110000",
  30349=>"000000111",
  30350=>"100000111",
  30351=>"000000011",
  30352=>"011001011",
  30353=>"100000010",
  30354=>"000010000",
  30355=>"000010111",
  30356=>"000010111",
  30357=>"000000111",
  30358=>"000011110",
  30359=>"000100000",
  30360=>"000001011",
  30361=>"000000010",
  30362=>"000010010",
  30363=>"000100111",
  30364=>"111100000",
  30365=>"010110101",
  30366=>"110111010",
  30367=>"111101111",
  30368=>"110101011",
  30369=>"111001010",
  30370=>"111010000",
  30371=>"001001011",
  30372=>"111101101",
  30373=>"000110110",
  30374=>"011010101",
  30375=>"000000000",
  30376=>"001000111",
  30377=>"000001111",
  30378=>"001101001",
  30379=>"111101011",
  30380=>"101111110",
  30381=>"101000100",
  30382=>"000001101",
  30383=>"111111111",
  30384=>"101110100",
  30385=>"000000111",
  30386=>"001100000",
  30387=>"011011011",
  30388=>"010000000",
  30389=>"000000000",
  30390=>"000111111",
  30391=>"111010101",
  30392=>"010100000",
  30393=>"000110111",
  30394=>"010000000",
  30395=>"111010111",
  30396=>"000111111",
  30397=>"011111111",
  30398=>"110111011",
  30399=>"111000000",
  30400=>"011111111",
  30401=>"000000000",
  30402=>"011100010",
  30403=>"100111110",
  30404=>"111111111",
  30405=>"001111100",
  30406=>"100010011",
  30407=>"000111111",
  30408=>"110111111",
  30409=>"010110000",
  30410=>"111111001",
  30411=>"010111111",
  30412=>"000000000",
  30413=>"010100111",
  30414=>"011101111",
  30415=>"010111110",
  30416=>"001000100",
  30417=>"000001001",
  30418=>"000000101",
  30419=>"011100111",
  30420=>"000010111",
  30421=>"000000000",
  30422=>"111000000",
  30423=>"111100010",
  30424=>"111001000",
  30425=>"000010111",
  30426=>"010111100",
  30427=>"000010010",
  30428=>"111011111",
  30429=>"000001101",
  30430=>"010000000",
  30431=>"101000111",
  30432=>"010000000",
  30433=>"111000111",
  30434=>"101011101",
  30435=>"010111111",
  30436=>"110000000",
  30437=>"000111001",
  30438=>"000000111",
  30439=>"110011010",
  30440=>"000000110",
  30441=>"000000000",
  30442=>"110100000",
  30443=>"000111101",
  30444=>"111110111",
  30445=>"000011111",
  30446=>"000010000",
  30447=>"101000111",
  30448=>"000000111",
  30449=>"100101101",
  30450=>"111011000",
  30451=>"000001001",
  30452=>"111100110",
  30453=>"111110111",
  30454=>"100000110",
  30455=>"111111111",
  30456=>"001111010",
  30457=>"110111101",
  30458=>"111010010",
  30459=>"000011111",
  30460=>"011111111",
  30461=>"111110000",
  30462=>"000111011",
  30463=>"111111110",
  30464=>"000100111",
  30465=>"011011011",
  30466=>"000100000",
  30467=>"000000001",
  30468=>"000010110",
  30469=>"011111111",
  30470=>"100111111",
  30471=>"100011001",
  30472=>"000000111",
  30473=>"000011111",
  30474=>"011110100",
  30475=>"000010111",
  30476=>"111110000",
  30477=>"000011011",
  30478=>"100101001",
  30479=>"111001001",
  30480=>"010000100",
  30481=>"111010000",
  30482=>"000000100",
  30483=>"111111111",
  30484=>"100101000",
  30485=>"000000111",
  30486=>"111100110",
  30487=>"111111011",
  30488=>"111011000",
  30489=>"111000101",
  30490=>"000000010",
  30491=>"110100100",
  30492=>"011011000",
  30493=>"001001101",
  30494=>"000111011",
  30495=>"101000011",
  30496=>"000111111",
  30497=>"111000110",
  30498=>"101000111",
  30499=>"000010011",
  30500=>"111110110",
  30501=>"110111110",
  30502=>"000010111",
  30503=>"001000100",
  30504=>"000000111",
  30505=>"010000111",
  30506=>"101000000",
  30507=>"111000000",
  30508=>"011000100",
  30509=>"101000000",
  30510=>"111111100",
  30511=>"000000101",
  30512=>"000110111",
  30513=>"011001000",
  30514=>"111111111",
  30515=>"111111101",
  30516=>"111111100",
  30517=>"111100111",
  30518=>"000110110",
  30519=>"101000000",
  30520=>"011000001",
  30521=>"111111000",
  30522=>"100000000",
  30523=>"111110100",
  30524=>"111011010",
  30525=>"110100010",
  30526=>"100001101",
  30527=>"001010110",
  30528=>"001101100",
  30529=>"111111111",
  30530=>"010000000",
  30531=>"001011011",
  30532=>"000000000",
  30533=>"100000000",
  30534=>"000111100",
  30535=>"001011001",
  30536=>"011101011",
  30537=>"100111111",
  30538=>"111101101",
  30539=>"010100000",
  30540=>"000011111",
  30541=>"001001011",
  30542=>"000000100",
  30543=>"111101101",
  30544=>"101101111",
  30545=>"011000000",
  30546=>"000011011",
  30547=>"100100111",
  30548=>"001000000",
  30549=>"110011100",
  30550=>"001011011",
  30551=>"111111011",
  30552=>"000000110",
  30553=>"000000000",
  30554=>"110110001",
  30555=>"010100111",
  30556=>"010000000",
  30557=>"111100100",
  30558=>"111101000",
  30559=>"000110010",
  30560=>"000010010",
  30561=>"010001110",
  30562=>"110110000",
  30563=>"011001000",
  30564=>"111101001",
  30565=>"111111100",
  30566=>"111100110",
  30567=>"001001010",
  30568=>"000101101",
  30569=>"011001101",
  30570=>"111111111",
  30571=>"000011111",
  30572=>"111011111",
  30573=>"111101000",
  30574=>"000000000",
  30575=>"001001000",
  30576=>"000001110",
  30577=>"000000000",
  30578=>"011011101",
  30579=>"111101110",
  30580=>"000000001",
  30581=>"000000100",
  30582=>"001000000",
  30583=>"100000111",
  30584=>"000111101",
  30585=>"111010000",
  30586=>"001101111",
  30587=>"000000000",
  30588=>"010000000",
  30589=>"000001111",
  30590=>"100001000",
  30591=>"100011011",
  30592=>"000010010",
  30593=>"000010011",
  30594=>"111010110",
  30595=>"111000000",
  30596=>"000001111",
  30597=>"101101111",
  30598=>"111111111",
  30599=>"000100100",
  30600=>"010110111",
  30601=>"100100101",
  30602=>"111100100",
  30603=>"000000000",
  30604=>"000000011",
  30605=>"000000000",
  30606=>"111111000",
  30607=>"000000001",
  30608=>"101111000",
  30609=>"100000111",
  30610=>"010011111",
  30611=>"000000011",
  30612=>"000000101",
  30613=>"011010000",
  30614=>"111011000",
  30615=>"000100011",
  30616=>"010011101",
  30617=>"000000000",
  30618=>"000010011",
  30619=>"111111101",
  30620=>"111111001",
  30621=>"101100110",
  30622=>"111011101",
  30623=>"100110111",
  30624=>"010011011",
  30625=>"111000000",
  30626=>"000001010",
  30627=>"101000000",
  30628=>"010111111",
  30629=>"000001111",
  30630=>"000000111",
  30631=>"111111111",
  30632=>"111100000",
  30633=>"000001000",
  30634=>"000010110",
  30635=>"010110111",
  30636=>"000000111",
  30637=>"101000000",
  30638=>"011111110",
  30639=>"111101101",
  30640=>"000111101",
  30641=>"001001101",
  30642=>"111011000",
  30643=>"001000000",
  30644=>"110110100",
  30645=>"111111011",
  30646=>"000110110",
  30647=>"100100111",
  30648=>"001100000",
  30649=>"000000100",
  30650=>"111111011",
  30651=>"111011011",
  30652=>"110110101",
  30653=>"000111111",
  30654=>"000000011",
  30655=>"000000011",
  30656=>"111101100",
  30657=>"110000000",
  30658=>"111111111",
  30659=>"010000100",
  30660=>"001000100",
  30661=>"011000000",
  30662=>"000011111",
  30663=>"010000000",
  30664=>"100111000",
  30665=>"111000100",
  30666=>"111011111",
  30667=>"011011110",
  30668=>"100100110",
  30669=>"011000000",
  30670=>"000000000",
  30671=>"000110100",
  30672=>"100010010",
  30673=>"000010110",
  30674=>"101101111",
  30675=>"111100000",
  30676=>"000000100",
  30677=>"011001111",
  30678=>"111011011",
  30679=>"111000100",
  30680=>"101100100",
  30681=>"011011111",
  30682=>"011100000",
  30683=>"000000101",
  30684=>"111000001",
  30685=>"010011011",
  30686=>"100101100",
  30687=>"000011111",
  30688=>"101100100",
  30689=>"100101000",
  30690=>"111000000",
  30691=>"000000001",
  30692=>"000000111",
  30693=>"010110010",
  30694=>"101011111",
  30695=>"100000000",
  30696=>"111111101",
  30697=>"000000000",
  30698=>"110111101",
  30699=>"111111111",
  30700=>"000000100",
  30701=>"001010110",
  30702=>"000000000",
  30703=>"000000010",
  30704=>"000010111",
  30705=>"011101110",
  30706=>"011010001",
  30707=>"111001000",
  30708=>"011010010",
  30709=>"001101101",
  30710=>"100000010",
  30711=>"101110100",
  30712=>"111111000",
  30713=>"110101101",
  30714=>"111100010",
  30715=>"001001100",
  30716=>"111010000",
  30717=>"000000100",
  30718=>"000110000",
  30719=>"111111000",
  30720=>"011011100",
  30721=>"000100111",
  30722=>"111000000",
  30723=>"000000010",
  30724=>"110110011",
  30725=>"000000000",
  30726=>"110101111",
  30727=>"000000110",
  30728=>"001101001",
  30729=>"111011110",
  30730=>"011111111",
  30731=>"011001000",
  30732=>"000000000",
  30733=>"111111111",
  30734=>"110110010",
  30735=>"000000001",
  30736=>"000111001",
  30737=>"010111111",
  30738=>"110110000",
  30739=>"000011111",
  30740=>"111110011",
  30741=>"110000111",
  30742=>"110111110",
  30743=>"110111111",
  30744=>"111001111",
  30745=>"111001001",
  30746=>"000000110",
  30747=>"111111110",
  30748=>"111111010",
  30749=>"101000000",
  30750=>"110000000",
  30751=>"010110000",
  30752=>"110110010",
  30753=>"111111100",
  30754=>"000101001",
  30755=>"000111111",
  30756=>"111111010",
  30757=>"110010110",
  30758=>"000111101",
  30759=>"001111111",
  30760=>"000001111",
  30761=>"000000110",
  30762=>"010111001",
  30763=>"111111111",
  30764=>"110111111",
  30765=>"000000001",
  30766=>"101000111",
  30767=>"000000000",
  30768=>"000000000",
  30769=>"111111001",
  30770=>"000010000",
  30771=>"111110000",
  30772=>"101111000",
  30773=>"000000000",
  30774=>"111111011",
  30775=>"001000000",
  30776=>"111110010",
  30777=>"101111111",
  30778=>"010000000",
  30779=>"110110010",
  30780=>"011001001",
  30781=>"100111101",
  30782=>"000000000",
  30783=>"001000110",
  30784=>"111111000",
  30785=>"000100000",
  30786=>"000100111",
  30787=>"010000110",
  30788=>"110111111",
  30789=>"000001011",
  30790=>"010011010",
  30791=>"000000001",
  30792=>"001010001",
  30793=>"000000111",
  30794=>"001001111",
  30795=>"000000000",
  30796=>"000000000",
  30797=>"010110000",
  30798=>"110110110",
  30799=>"010000110",
  30800=>"001100101",
  30801=>"110111110",
  30802=>"011011111",
  30803=>"011000000",
  30804=>"000000010",
  30805=>"100000100",
  30806=>"110110100",
  30807=>"101000111",
  30808=>"111111111",
  30809=>"000000011",
  30810=>"111111111",
  30811=>"000000000",
  30812=>"001101101",
  30813=>"111100110",
  30814=>"110111111",
  30815=>"111111111",
  30816=>"111111111",
  30817=>"110011111",
  30818=>"111111000",
  30819=>"110110001",
  30820=>"001011011",
  30821=>"001000000",
  30822=>"110111100",
  30823=>"001000000",
  30824=>"011000001",
  30825=>"011000000",
  30826=>"011111110",
  30827=>"000000010",
  30828=>"110000111",
  30829=>"110111110",
  30830=>"011010000",
  30831=>"111111110",
  30832=>"110100100",
  30833=>"110000000",
  30834=>"111111100",
  30835=>"000110000",
  30836=>"111111001",
  30837=>"000000001",
  30838=>"000101000",
  30839=>"101001010",
  30840=>"000101101",
  30841=>"110111111",
  30842=>"011111111",
  30843=>"000000000",
  30844=>"110111110",
  30845=>"000000000",
  30846=>"000001111",
  30847=>"111001000",
  30848=>"000111000",
  30849=>"111100000",
  30850=>"111000001",
  30851=>"000000000",
  30852=>"111011110",
  30853=>"000001001",
  30854=>"111111110",
  30855=>"011111000",
  30856=>"111010010",
  30857=>"000000001",
  30858=>"000111011",
  30859=>"001000000",
  30860=>"110101101",
  30861=>"111110111",
  30862=>"000000000",
  30863=>"000001001",
  30864=>"100000000",
  30865=>"000101111",
  30866=>"000000011",
  30867=>"000011001",
  30868=>"110010100",
  30869=>"111101010",
  30870=>"000000000",
  30871=>"000100000",
  30872=>"110111100",
  30873=>"000000000",
  30874=>"000000010",
  30875=>"000000000",
  30876=>"110110110",
  30877=>"111000110",
  30878=>"111001001",
  30879=>"000000000",
  30880=>"001001001",
  30881=>"111110000",
  30882=>"000000000",
  30883=>"000000001",
  30884=>"011011111",
  30885=>"000000000",
  30886=>"000100000",
  30887=>"000000000",
  30888=>"000111111",
  30889=>"000000100",
  30890=>"111110111",
  30891=>"111110111",
  30892=>"000001111",
  30893=>"101000100",
  30894=>"111110110",
  30895=>"000011001",
  30896=>"000000111",
  30897=>"110110100",
  30898=>"110100000",
  30899=>"111010000",
  30900=>"000000000",
  30901=>"000000000",
  30902=>"001000000",
  30903=>"111111111",
  30904=>"010100100",
  30905=>"100111001",
  30906=>"111111111",
  30907=>"000001111",
  30908=>"000000000",
  30909=>"111110100",
  30910=>"100000000",
  30911=>"000000111",
  30912=>"101001000",
  30913=>"011000000",
  30914=>"001000000",
  30915=>"001000001",
  30916=>"000001111",
  30917=>"110100110",
  30918=>"000000111",
  30919=>"000110110",
  30920=>"011000000",
  30921=>"000000000",
  30922=>"000000111",
  30923=>"000000000",
  30924=>"111011000",
  30925=>"111111111",
  30926=>"001101000",
  30927=>"100001001",
  30928=>"111110000",
  30929=>"110110000",
  30930=>"100011000",
  30931=>"000000000",
  30932=>"001001111",
  30933=>"010111011",
  30934=>"111111000",
  30935=>"000000000",
  30936=>"000000001",
  30937=>"010111111",
  30938=>"100000000",
  30939=>"000000000",
  30940=>"011111110",
  30941=>"111010000",
  30942=>"000010000",
  30943=>"111101111",
  30944=>"000000000",
  30945=>"110101101",
  30946=>"000111111",
  30947=>"000001100",
  30948=>"000000001",
  30949=>"111111100",
  30950=>"111111111",
  30951=>"111111011",
  30952=>"000111111",
  30953=>"010111111",
  30954=>"111111111",
  30955=>"000010111",
  30956=>"011111111",
  30957=>"000111111",
  30958=>"110110000",
  30959=>"111000111",
  30960=>"111010001",
  30961=>"111011011",
  30962=>"110000001",
  30963=>"110110100",
  30964=>"100100000",
  30965=>"110110111",
  30966=>"000000000",
  30967=>"000000000",
  30968=>"011000000",
  30969=>"000000000",
  30970=>"000000000",
  30971=>"111001000",
  30972=>"100101101",
  30973=>"000010000",
  30974=>"100011000",
  30975=>"001000000",
  30976=>"100000001",
  30977=>"111011000",
  30978=>"111000000",
  30979=>"101111000",
  30980=>"111100100",
  30981=>"001110001",
  30982=>"111111111",
  30983=>"111101101",
  30984=>"000001110",
  30985=>"000101111",
  30986=>"110111000",
  30987=>"111111000",
  30988=>"000100111",
  30989=>"110110000",
  30990=>"000001000",
  30991=>"111111100",
  30992=>"000111111",
  30993=>"000111111",
  30994=>"111001101",
  30995=>"001000000",
  30996=>"101111111",
  30997=>"111000000",
  30998=>"111000100",
  30999=>"111111000",
  31000=>"111000000",
  31001=>"111011111",
  31002=>"111101001",
  31003=>"100111111",
  31004=>"100000010",
  31005=>"111000000",
  31006=>"111000000",
  31007=>"001000000",
  31008=>"110110000",
  31009=>"111101000",
  31010=>"011111001",
  31011=>"000000101",
  31012=>"100111011",
  31013=>"111001000",
  31014=>"111001000",
  31015=>"000001111",
  31016=>"111001000",
  31017=>"110100000",
  31018=>"110000000",
  31019=>"110000111",
  31020=>"011111001",
  31021=>"111101010",
  31022=>"111000000",
  31023=>"111011111",
  31024=>"000100000",
  31025=>"101111100",
  31026=>"111101000",
  31027=>"111011000",
  31028=>"001000100",
  31029=>"000000100",
  31030=>"001110000",
  31031=>"111111111",
  31032=>"111111111",
  31033=>"110110000",
  31034=>"011111000",
  31035=>"111111000",
  31036=>"000010100",
  31037=>"111011010",
  31038=>"001000100",
  31039=>"011011000",
  31040=>"010000111",
  31041=>"000000101",
  31042=>"100001111",
  31043=>"100101111",
  31044=>"011011011",
  31045=>"010000001",
  31046=>"111111000",
  31047=>"110111111",
  31048=>"111011011",
  31049=>"000000111",
  31050=>"111000111",
  31051=>"000110111",
  31052=>"000001101",
  31053=>"000011110",
  31054=>"100110011",
  31055=>"111010111",
  31056=>"111101000",
  31057=>"111010010",
  31058=>"000000000",
  31059=>"000111011",
  31060=>"101101111",
  31061=>"011100101",
  31062=>"011000000",
  31063=>"000101101",
  31064=>"101101000",
  31065=>"000111110",
  31066=>"111101000",
  31067=>"000111111",
  31068=>"000001111",
  31069=>"000000000",
  31070=>"111000011",
  31071=>"001000001",
  31072=>"000000000",
  31073=>"001101000",
  31074=>"011101111",
  31075=>"111101000",
  31076=>"000010010",
  31077=>"000100011",
  31078=>"001001110",
  31079=>"000000110",
  31080=>"111000000",
  31081=>"101001001",
  31082=>"000000101",
  31083=>"010000000",
  31084=>"010000001",
  31085=>"000011010",
  31086=>"000000111",
  31087=>"111111001",
  31088=>"110100010",
  31089=>"100111111",
  31090=>"111011001",
  31091=>"000000000",
  31092=>"111111111",
  31093=>"000100000",
  31094=>"111010000",
  31095=>"000000010",
  31096=>"000001000",
  31097=>"000101000",
  31098=>"110010111",
  31099=>"001000010",
  31100=>"111111001",
  31101=>"000001000",
  31102=>"111111110",
  31103=>"000000111",
  31104=>"000000011",
  31105=>"111100110",
  31106=>"000010111",
  31107=>"100000000",
  31108=>"000000000",
  31109=>"000011111",
  31110=>"011000000",
  31111=>"010011001",
  31112=>"000001111",
  31113=>"101000111",
  31114=>"111100000",
  31115=>"000110111",
  31116=>"011000111",
  31117=>"000111110",
  31118=>"000000111",
  31119=>"000100111",
  31120=>"011110111",
  31121=>"111101101",
  31122=>"010000000",
  31123=>"010000101",
  31124=>"001110110",
  31125=>"000000010",
  31126=>"111110100",
  31127=>"001100110",
  31128=>"000111111",
  31129=>"110000000",
  31130=>"111000000",
  31131=>"011000000",
  31132=>"100001111",
  31133=>"010000100",
  31134=>"111111111",
  31135=>"000100010",
  31136=>"001111110",
  31137=>"111101000",
  31138=>"000000000",
  31139=>"100111101",
  31140=>"001000000",
  31141=>"000100110",
  31142=>"000010111",
  31143=>"001101000",
  31144=>"000011111",
  31145=>"000101011",
  31146=>"111111111",
  31147=>"001000110",
  31148=>"111011111",
  31149=>"000101111",
  31150=>"011111000",
  31151=>"000101111",
  31152=>"001001011",
  31153=>"110110000",
  31154=>"001101010",
  31155=>"100000001",
  31156=>"001100111",
  31157=>"011011000",
  31158=>"011000000",
  31159=>"011010000",
  31160=>"000001001",
  31161=>"100110110",
  31162=>"011000000",
  31163=>"111111101",
  31164=>"000111101",
  31165=>"111111000",
  31166=>"000100001",
  31167=>"101111110",
  31168=>"100001010",
  31169=>"000000111",
  31170=>"000010100",
  31171=>"110110110",
  31172=>"000000100",
  31173=>"100011001",
  31174=>"000000000",
  31175=>"000000111",
  31176=>"110111111",
  31177=>"000000111",
  31178=>"100001101",
  31179=>"000000001",
  31180=>"111100000",
  31181=>"111000110",
  31182=>"111001000",
  31183=>"111111100",
  31184=>"111111000",
  31185=>"110011001",
  31186=>"000010111",
  31187=>"000111111",
  31188=>"000001111",
  31189=>"111101100",
  31190=>"111100100",
  31191=>"111111111",
  31192=>"000011111",
  31193=>"000000010",
  31194=>"101111001",
  31195=>"000011010",
  31196=>"110000011",
  31197=>"001100010",
  31198=>"000111111",
  31199=>"101111111",
  31200=>"100000000",
  31201=>"100000111",
  31202=>"001001111",
  31203=>"001110110",
  31204=>"000000110",
  31205=>"000000000",
  31206=>"000100000",
  31207=>"010011010",
  31208=>"000000111",
  31209=>"010000011",
  31210=>"111110000",
  31211=>"010000001",
  31212=>"110000111",
  31213=>"111111001",
  31214=>"000000000",
  31215=>"000100110",
  31216=>"110100000",
  31217=>"101100100",
  31218=>"000010100",
  31219=>"000111001",
  31220=>"001111110",
  31221=>"111001000",
  31222=>"100000100",
  31223=>"000000111",
  31224=>"100100111",
  31225=>"101111000",
  31226=>"110100010",
  31227=>"000010111",
  31228=>"111010000",
  31229=>"000000101",
  31230=>"000000000",
  31231=>"001000111",
  31232=>"111111000",
  31233=>"000111011",
  31234=>"000110110",
  31235=>"000000011",
  31236=>"011111110",
  31237=>"000000000",
  31238=>"111001011",
  31239=>"010000001",
  31240=>"100111111",
  31241=>"111101111",
  31242=>"010100100",
  31243=>"111000010",
  31244=>"101000000",
  31245=>"111110000",
  31246=>"000001001",
  31247=>"000000100",
  31248=>"000000001",
  31249=>"001001001",
  31250=>"010100101",
  31251=>"001100000",
  31252=>"101000111",
  31253=>"010111110",
  31254=>"011110000",
  31255=>"011111101",
  31256=>"100100100",
  31257=>"101100111",
  31258=>"010000100",
  31259=>"000000000",
  31260=>"101111111",
  31261=>"101111110",
  31262=>"000110111",
  31263=>"001001011",
  31264=>"010111011",
  31265=>"000000000",
  31266=>"000111111",
  31267=>"111011111",
  31268=>"000100110",
  31269=>"100100010",
  31270=>"010111000",
  31271=>"101111001",
  31272=>"111111111",
  31273=>"000000000",
  31274=>"111010010",
  31275=>"000000000",
  31276=>"000100100",
  31277=>"010000000",
  31278=>"010000000",
  31279=>"001000000",
  31280=>"110000001",
  31281=>"000000000",
  31282=>"000110111",
  31283=>"100000001",
  31284=>"000000010",
  31285=>"111111000",
  31286=>"000100010",
  31287=>"011111111",
  31288=>"010111111",
  31289=>"000000000",
  31290=>"000000101",
  31291=>"000000000",
  31292=>"011011111",
  31293=>"111111011",
  31294=>"000000000",
  31295=>"101110000",
  31296=>"111101101",
  31297=>"111100001",
  31298=>"000000000",
  31299=>"011001100",
  31300=>"000000111",
  31301=>"101000001",
  31302=>"110011011",
  31303=>"111110111",
  31304=>"000000000",
  31305=>"011010010",
  31306=>"101000000",
  31307=>"011001011",
  31308=>"000100111",
  31309=>"001111111",
  31310=>"100000000",
  31311=>"000000000",
  31312=>"100100100",
  31313=>"000111111",
  31314=>"000000101",
  31315=>"001000000",
  31316=>"111111010",
  31317=>"001100100",
  31318=>"001001101",
  31319=>"000110101",
  31320=>"111000110",
  31321=>"000000001",
  31322=>"011100000",
  31323=>"011001100",
  31324=>"011111110",
  31325=>"001001011",
  31326=>"010111011",
  31327=>"111111011",
  31328=>"000000100",
  31329=>"000101001",
  31330=>"000000101",
  31331=>"100110000",
  31332=>"100100111",
  31333=>"100000000",
  31334=>"100000001",
  31335=>"110110111",
  31336=>"111111010",
  31337=>"000100111",
  31338=>"110100100",
  31339=>"010000010",
  31340=>"101101101",
  31341=>"101111000",
  31342=>"000000000",
  31343=>"000000111",
  31344=>"001000011",
  31345=>"000000000",
  31346=>"000000000",
  31347=>"010010011",
  31348=>"000000011",
  31349=>"000000111",
  31350=>"111110111",
  31351=>"100100011",
  31352=>"000111111",
  31353=>"001001111",
  31354=>"000000111",
  31355=>"101101101",
  31356=>"100110111",
  31357=>"100100000",
  31358=>"011010000",
  31359=>"010011111",
  31360=>"111101011",
  31361=>"111011010",
  31362=>"100000101",
  31363=>"000001101",
  31364=>"100000000",
  31365=>"111101001",
  31366=>"011001110",
  31367=>"000100000",
  31368=>"100011011",
  31369=>"101000000",
  31370=>"011011000",
  31371=>"100010000",
  31372=>"011111010",
  31373=>"011111111",
  31374=>"001011011",
  31375=>"100000001",
  31376=>"001001001",
  31377=>"111000010",
  31378=>"011011000",
  31379=>"000000001",
  31380=>"101111111",
  31381=>"000000100",
  31382=>"111111111",
  31383=>"000000000",
  31384=>"101010110",
  31385=>"001111111",
  31386=>"000111010",
  31387=>"000000000",
  31388=>"101111000",
  31389=>"101000000",
  31390=>"000000111",
  31391=>"111101000",
  31392=>"100011101",
  31393=>"010011010",
  31394=>"000011000",
  31395=>"000010000",
  31396=>"011101000",
  31397=>"111101111",
  31398=>"000110000",
  31399=>"100111111",
  31400=>"111110111",
  31401=>"011000100",
  31402=>"000000000",
  31403=>"000000000",
  31404=>"000001000",
  31405=>"000000001",
  31406=>"111111110",
  31407=>"111111110",
  31408=>"111110000",
  31409=>"111011000",
  31410=>"000000100",
  31411=>"100100100",
  31412=>"001111000",
  31413=>"111111010",
  31414=>"100100100",
  31415=>"000000000",
  31416=>"100111111",
  31417=>"100110100",
  31418=>"000000100",
  31419=>"011111111",
  31420=>"000000111",
  31421=>"001001111",
  31422=>"110011111",
  31423=>"111111111",
  31424=>"000111111",
  31425=>"111011010",
  31426=>"001110010",
  31427=>"000000000",
  31428=>"001000000",
  31429=>"001100010",
  31430=>"111110111",
  31431=>"100000011",
  31432=>"001111001",
  31433=>"111100111",
  31434=>"111111111",
  31435=>"010111000",
  31436=>"001000011",
  31437=>"001001011",
  31438=>"000000000",
  31439=>"000101001",
  31440=>"011111110",
  31441=>"001001000",
  31442=>"011000110",
  31443=>"001000111",
  31444=>"011011010",
  31445=>"100111111",
  31446=>"000000100",
  31447=>"000001011",
  31448=>"011111000",
  31449=>"111101101",
  31450=>"001101101",
  31451=>"001000000",
  31452=>"110011110",
  31453=>"011010111",
  31454=>"010000111",
  31455=>"110111111",
  31456=>"000000101",
  31457=>"100000001",
  31458=>"101101000",
  31459=>"100000000",
  31460=>"010000000",
  31461=>"010010011",
  31462=>"101000000",
  31463=>"111111011",
  31464=>"101000000",
  31465=>"110111101",
  31466=>"110011001",
  31467=>"000010101",
  31468=>"000000000",
  31469=>"101101111",
  31470=>"000000000",
  31471=>"100000010",
  31472=>"101000000",
  31473=>"010001000",
  31474=>"000000101",
  31475=>"000000000",
  31476=>"101000101",
  31477=>"010111001",
  31478=>"000000111",
  31479=>"000000000",
  31480=>"000100111",
  31481=>"000000100",
  31482=>"010111110",
  31483=>"001101101",
  31484=>"010110100",
  31485=>"000000000",
  31486=>"100100111",
  31487=>"110100001",
  31488=>"011110000",
  31489=>"010000010",
  31490=>"000010110",
  31491=>"000000001",
  31492=>"000011001",
  31493=>"010000000",
  31494=>"000000101",
  31495=>"111000100",
  31496=>"111011100",
  31497=>"011010010",
  31498=>"110111001",
  31499=>"000000000",
  31500=>"111111111",
  31501=>"111111000",
  31502=>"100011111",
  31503=>"110001111",
  31504=>"010000010",
  31505=>"111111010",
  31506=>"000001101",
  31507=>"011010110",
  31508=>"010000111",
  31509=>"100000000",
  31510=>"111000000",
  31511=>"100100111",
  31512=>"101100101",
  31513=>"111111110",
  31514=>"011101000",
  31515=>"000010000",
  31516=>"010000011",
  31517=>"100000111",
  31518=>"011110010",
  31519=>"001111011",
  31520=>"000000000",
  31521=>"000000010",
  31522=>"100000011",
  31523=>"000000000",
  31524=>"100110110",
  31525=>"110101000",
  31526=>"000000101",
  31527=>"111111011",
  31528=>"010100000",
  31529=>"011000000",
  31530=>"010000010",
  31531=>"011000000",
  31532=>"111000100",
  31533=>"111000110",
  31534=>"111101101",
  31535=>"110100111",
  31536=>"111111011",
  31537=>"100100001",
  31538=>"100000001",
  31539=>"111011010",
  31540=>"011011010",
  31541=>"001110110",
  31542=>"110000001",
  31543=>"000000001",
  31544=>"000000000",
  31545=>"001001111",
  31546=>"000000101",
  31547=>"000010000",
  31548=>"100000001",
  31549=>"111101111",
  31550=>"000010000",
  31551=>"100000100",
  31552=>"000111011",
  31553=>"111001111",
  31554=>"000000000",
  31555=>"000000101",
  31556=>"111110110",
  31557=>"010000101",
  31558=>"111111000",
  31559=>"000010100",
  31560=>"101001101",
  31561=>"011111000",
  31562=>"101101111",
  31563=>"111111111",
  31564=>"000001101",
  31565=>"011011011",
  31566=>"011011100",
  31567=>"100000000",
  31568=>"000001101",
  31569=>"010000010",
  31570=>"111000111",
  31571=>"001110110",
  31572=>"010010000",
  31573=>"100100010",
  31574=>"000000000",
  31575=>"010110000",
  31576=>"110111111",
  31577=>"111111011",
  31578=>"110110110",
  31579=>"000100100",
  31580=>"001000000",
  31581=>"001000001",
  31582=>"111111110",
  31583=>"000000001",
  31584=>"101000101",
  31585=>"001000000",
  31586=>"000000101",
  31587=>"000001000",
  31588=>"101001101",
  31589=>"001100100",
  31590=>"000001011",
  31591=>"001101101",
  31592=>"000000111",
  31593=>"111100000",
  31594=>"111001000",
  31595=>"111000111",
  31596=>"100000000",
  31597=>"111111101",
  31598=>"111000000",
  31599=>"111111111",
  31600=>"011110101",
  31601=>"000000110",
  31602=>"011000010",
  31603=>"000111101",
  31604=>"101111111",
  31605=>"000000111",
  31606=>"001110111",
  31607=>"110000100",
  31608=>"010010010",
  31609=>"111000000",
  31610=>"000000010",
  31611=>"111001101",
  31612=>"000110100",
  31613=>"100101101",
  31614=>"011000000",
  31615=>"000001101",
  31616=>"011000000",
  31617=>"000000010",
  31618=>"111000000",
  31619=>"111100011",
  31620=>"111101111",
  31621=>"101101101",
  31622=>"011001100",
  31623=>"000001101",
  31624=>"100101100",
  31625=>"111001101",
  31626=>"001000000",
  31627=>"000011111",
  31628=>"000000000",
  31629=>"011110110",
  31630=>"101101101",
  31631=>"000000100",
  31632=>"100100110",
  31633=>"111000100",
  31634=>"111000000",
  31635=>"000010010",
  31636=>"000010100",
  31637=>"010010110",
  31638=>"010010010",
  31639=>"000000010",
  31640=>"010000010",
  31641=>"111010010",
  31642=>"010011010",
  31643=>"001010000",
  31644=>"000001001",
  31645=>"000111111",
  31646=>"000111111",
  31647=>"001000001",
  31648=>"001101001",
  31649=>"000011010",
  31650=>"111111101",
  31651=>"000000010",
  31652=>"000000011",
  31653=>"100001001",
  31654=>"110010111",
  31655=>"010111010",
  31656=>"011010110",
  31657=>"000000000",
  31658=>"110111110",
  31659=>"000011010",
  31660=>"111000100",
  31661=>"010011000",
  31662=>"100100101",
  31663=>"010100101",
  31664=>"111100111",
  31665=>"001110111",
  31666=>"000000101",
  31667=>"000110000",
  31668=>"001101101",
  31669=>"100111111",
  31670=>"111000100",
  31671=>"011111110",
  31672=>"000000000",
  31673=>"000100101",
  31674=>"111000010",
  31675=>"001010010",
  31676=>"011100000",
  31677=>"110111111",
  31678=>"001100001",
  31679=>"011000000",
  31680=>"010000010",
  31681=>"101101111",
  31682=>"000110111",
  31683=>"001001000",
  31684=>"000000111",
  31685=>"110010010",
  31686=>"111111000",
  31687=>"010111111",
  31688=>"000000000",
  31689=>"111101011",
  31690=>"000000110",
  31691=>"101000111",
  31692=>"111100000",
  31693=>"000010000",
  31694=>"001111000",
  31695=>"000000011",
  31696=>"000010100",
  31697=>"101000101",
  31698=>"000111110",
  31699=>"111111101",
  31700=>"000000111",
  31701=>"111111101",
  31702=>"110010000",
  31703=>"100101101",
  31704=>"000000001",
  31705=>"111000000",
  31706=>"100101101",
  31707=>"000001111",
  31708=>"000000010",
  31709=>"010000111",
  31710=>"010110111",
  31711=>"000000010",
  31712=>"010010000",
  31713=>"111111111",
  31714=>"000001000",
  31715=>"010001110",
  31716=>"010111010",
  31717=>"110000000",
  31718=>"001000001",
  31719=>"011001000",
  31720=>"000000000",
  31721=>"111101100",
  31722=>"011111110",
  31723=>"111111111",
  31724=>"111111000",
  31725=>"000111011",
  31726=>"000010000",
  31727=>"000000111",
  31728=>"000000010",
  31729=>"011011100",
  31730=>"111000000",
  31731=>"101101101",
  31732=>"111101001",
  31733=>"101101100",
  31734=>"100000000",
  31735=>"000000000",
  31736=>"000000011",
  31737=>"000000111",
  31738=>"010000110",
  31739=>"000110101",
  31740=>"100000010",
  31741=>"101100100",
  31742=>"110110111",
  31743=>"001000000",
  31744=>"100100100",
  31745=>"101111010",
  31746=>"111000000",
  31747=>"110111111",
  31748=>"000101101",
  31749=>"110101000",
  31750=>"000111011",
  31751=>"000111111",
  31752=>"111000000",
  31753=>"011000101",
  31754=>"000000000",
  31755=>"000001110",
  31756=>"001101001",
  31757=>"110010010",
  31758=>"100011001",
  31759=>"101000001",
  31760=>"100010100",
  31761=>"000000000",
  31762=>"110000010",
  31763=>"101111011",
  31764=>"111111000",
  31765=>"011111001",
  31766=>"000101011",
  31767=>"111111111",
  31768=>"000000111",
  31769=>"010000110",
  31770=>"000000000",
  31771=>"000101111",
  31772=>"111000010",
  31773=>"001001010",
  31774=>"010100101",
  31775=>"000000000",
  31776=>"000000000",
  31777=>"010001101",
  31778=>"010010010",
  31779=>"111111111",
  31780=>"101100000",
  31781=>"001011001",
  31782=>"000111010",
  31783=>"011011001",
  31784=>"000101111",
  31785=>"100111000",
  31786=>"000000010",
  31787=>"010111010",
  31788=>"000111101",
  31789=>"101100011",
  31790=>"110000000",
  31791=>"111001000",
  31792=>"011011000",
  31793=>"100000000",
  31794=>"000001111",
  31795=>"000111111",
  31796=>"001001000",
  31797=>"110010100",
  31798=>"001001001",
  31799=>"110110000",
  31800=>"101110000",
  31801=>"000111111",
  31802=>"000000100",
  31803=>"000111111",
  31804=>"001011011",
  31805=>"111000011",
  31806=>"000000101",
  31807=>"001001000",
  31808=>"111111111",
  31809=>"010101010",
  31810=>"011110011",
  31811=>"111100001",
  31812=>"111111111",
  31813=>"010010000",
  31814=>"000000111",
  31815=>"100010010",
  31816=>"001101011",
  31817=>"001101111",
  31818=>"001001001",
  31819=>"011000001",
  31820=>"111011111",
  31821=>"100101101",
  31822=>"010000000",
  31823=>"101111111",
  31824=>"000000000",
  31825=>"101111111",
  31826=>"111101010",
  31827=>"110110100",
  31828=>"110100101",
  31829=>"100001000",
  31830=>"101101001",
  31831=>"111001101",
  31832=>"001011101",
  31833=>"001101001",
  31834=>"001101101",
  31835=>"111000000",
  31836=>"001010000",
  31837=>"000001111",
  31838=>"111111000",
  31839=>"101001000",
  31840=>"111110000",
  31841=>"000000011",
  31842=>"111000000",
  31843=>"100111111",
  31844=>"000100101",
  31845=>"000000101",
  31846=>"000101011",
  31847=>"000000010",
  31848=>"110111001",
  31849=>"000100010",
  31850=>"001001000",
  31851=>"111000011",
  31852=>"001010000",
  31853=>"010000100",
  31854=>"011000000",
  31855=>"000101111",
  31856=>"001001100",
  31857=>"011101111",
  31858=>"100100100",
  31859=>"011000001",
  31860=>"101101010",
  31861=>"000000110",
  31862=>"010100101",
  31863=>"011000000",
  31864=>"000010000",
  31865=>"000100010",
  31866=>"000000101",
  31867=>"000000000",
  31868=>"000000101",
  31869=>"011001001",
  31870=>"111101000",
  31871=>"111000000",
  31872=>"111101101",
  31873=>"110011000",
  31874=>"101100000",
  31875=>"100101110",
  31876=>"111011111",
  31877=>"101111111",
  31878=>"100100110",
  31879=>"000001001",
  31880=>"100101011",
  31881=>"011111111",
  31882=>"010100011",
  31883=>"001001001",
  31884=>"010101111",
  31885=>"011011000",
  31886=>"001111010",
  31887=>"011000111",
  31888=>"001101101",
  31889=>"110111111",
  31890=>"000001111",
  31891=>"110111101",
  31892=>"111011101",
  31893=>"111001000",
  31894=>"110001001",
  31895=>"001011000",
  31896=>"000100000",
  31897=>"111111111",
  31898=>"111111111",
  31899=>"111111000",
  31900=>"011111111",
  31901=>"110010010",
  31902=>"000001111",
  31903=>"000000101",
  31904=>"000000000",
  31905=>"001001111",
  31906=>"111111011",
  31907=>"111111111",
  31908=>"010001100",
  31909=>"001001001",
  31910=>"000100111",
  31911=>"000000000",
  31912=>"010000010",
  31913=>"111110000",
  31914=>"111000000",
  31915=>"011000000",
  31916=>"010000111",
  31917=>"000000000",
  31918=>"001011001",
  31919=>"001001010",
  31920=>"101010010",
  31921=>"000100100",
  31922=>"001101111",
  31923=>"000100101",
  31924=>"100101011",
  31925=>"000001010",
  31926=>"010000101",
  31927=>"000101111",
  31928=>"100100101",
  31929=>"111100111",
  31930=>"111111100",
  31931=>"101111101",
  31932=>"000000000",
  31933=>"111010010",
  31934=>"111000000",
  31935=>"000000000",
  31936=>"000101101",
  31937=>"000111001",
  31938=>"011111111",
  31939=>"100100100",
  31940=>"011000000",
  31941=>"101001011",
  31942=>"111011111",
  31943=>"111010000",
  31944=>"011000000",
  31945=>"010001000",
  31946=>"010000110",
  31947=>"011111100",
  31948=>"100111000",
  31949=>"000001101",
  31950=>"110000000",
  31951=>"111001011",
  31952=>"001101111",
  31953=>"000000000",
  31954=>"110110111",
  31955=>"110101000",
  31956=>"000000000",
  31957=>"000101011",
  31958=>"000100000",
  31959=>"101001000",
  31960=>"101111011",
  31961=>"000011011",
  31962=>"000001001",
  31963=>"011000000",
  31964=>"001101100",
  31965=>"101111011",
  31966=>"011010010",
  31967=>"001110110",
  31968=>"111000000",
  31969=>"000000111",
  31970=>"101111010",
  31971=>"011101100",
  31972=>"010000101",
  31973=>"000001001",
  31974=>"111000000",
  31975=>"000101111",
  31976=>"011111011",
  31977=>"000111111",
  31978=>"100000000",
  31979=>"000001001",
  31980=>"000000000",
  31981=>"110101110",
  31982=>"100000000",
  31983=>"011000000",
  31984=>"101000100",
  31985=>"010000100",
  31986=>"000101000",
  31987=>"001111000",
  31988=>"001001111",
  31989=>"000000001",
  31990=>"100000101",
  31991=>"000011010",
  31992=>"111111000",
  31993=>"001111011",
  31994=>"000111111",
  31995=>"000000111",
  31996=>"111111010",
  31997=>"000110000",
  31998=>"000001001",
  31999=>"110111000",
  32000=>"000011110",
  32001=>"100111001",
  32002=>"100000000",
  32003=>"100000111",
  32004=>"000011010",
  32005=>"101001111",
  32006=>"000000000",
  32007=>"000010000",
  32008=>"000000101",
  32009=>"000010000",
  32010=>"000011000",
  32011=>"100000101",
  32012=>"101010010",
  32013=>"000000000",
  32014=>"101011001",
  32015=>"111111000",
  32016=>"100010010",
  32017=>"000000010",
  32018=>"101100101",
  32019=>"000010011",
  32020=>"111111010",
  32021=>"101000100",
  32022=>"001000100",
  32023=>"111111010",
  32024=>"000101001",
  32025=>"000111101",
  32026=>"000000110",
  32027=>"000000101",
  32028=>"101100111",
  32029=>"100001110",
  32030=>"011000000",
  32031=>"101101111",
  32032=>"010000001",
  32033=>"001111000",
  32034=>"000010000",
  32035=>"101001111",
  32036=>"011001001",
  32037=>"011101111",
  32038=>"101000111",
  32039=>"000010010",
  32040=>"100100111",
  32041=>"101100111",
  32042=>"010111000",
  32043=>"011011000",
  32044=>"110111011",
  32045=>"000000110",
  32046=>"110110110",
  32047=>"111001111",
  32048=>"100100111",
  32049=>"001001100",
  32050=>"100000000",
  32051=>"101000011",
  32052=>"011011011",
  32053=>"101111100",
  32054=>"011011100",
  32055=>"000111000",
  32056=>"100000111",
  32057=>"111100110",
  32058=>"000101111",
  32059=>"000000111",
  32060=>"111010111",
  32061=>"010011110",
  32062=>"000000000",
  32063=>"101001001",
  32064=>"001011111",
  32065=>"010110010",
  32066=>"100000111",
  32067=>"100000110",
  32068=>"000000000",
  32069=>"000100000",
  32070=>"000111000",
  32071=>"101000101",
  32072=>"000001101",
  32073=>"011011010",
  32074=>"111100111",
  32075=>"011100001",
  32076=>"111101111",
  32077=>"100111111",
  32078=>"000110110",
  32079=>"111111111",
  32080=>"011010111",
  32081=>"010000010",
  32082=>"101000100",
  32083=>"011001000",
  32084=>"011000000",
  32085=>"001100100",
  32086=>"100110110",
  32087=>"000011111",
  32088=>"001101101",
  32089=>"100001110",
  32090=>"110110110",
  32091=>"000001000",
  32092=>"000000001",
  32093=>"000001001",
  32094=>"101101101",
  32095=>"110110001",
  32096=>"011001111",
  32097=>"000000010",
  32098=>"101100101",
  32099=>"011001010",
  32100=>"101000110",
  32101=>"001001000",
  32102=>"011110111",
  32103=>"110110111",
  32104=>"000100110",
  32105=>"000100100",
  32106=>"111111111",
  32107=>"101111111",
  32108=>"000000000",
  32109=>"011111001",
  32110=>"000000000",
  32111=>"011100011",
  32112=>"011001000",
  32113=>"000000010",
  32114=>"111111000",
  32115=>"010011111",
  32116=>"111111000",
  32117=>"000000001",
  32118=>"001100111",
  32119=>"111011100",
  32120=>"001011010",
  32121=>"100101010",
  32122=>"101010111",
  32123=>"111101111",
  32124=>"110110010",
  32125=>"110100000",
  32126=>"010111000",
  32127=>"111101100",
  32128=>"001011000",
  32129=>"000110110",
  32130=>"111000111",
  32131=>"100101110",
  32132=>"111111111",
  32133=>"000000001",
  32134=>"011111001",
  32135=>"001011000",
  32136=>"101101000",
  32137=>"001010000",
  32138=>"000111010",
  32139=>"010000000",
  32140=>"110100100",
  32141=>"000111000",
  32142=>"000111001",
  32143=>"100000000",
  32144=>"100100011",
  32145=>"111000011",
  32146=>"010011110",
  32147=>"011111000",
  32148=>"000001000",
  32149=>"100000111",
  32150=>"111111010",
  32151=>"110000000",
  32152=>"001111111",
  32153=>"000011110",
  32154=>"101100111",
  32155=>"110100110",
  32156=>"000000100",
  32157=>"000000111",
  32158=>"010011010",
  32159=>"001001111",
  32160=>"101100101",
  32161=>"000101001",
  32162=>"111100110",
  32163=>"111101000",
  32164=>"100000000",
  32165=>"100111000",
  32166=>"111010000",
  32167=>"000100100",
  32168=>"001000111",
  32169=>"111010010",
  32170=>"101100111",
  32171=>"000000000",
  32172=>"100100011",
  32173=>"101000000",
  32174=>"010010010",
  32175=>"111010000",
  32176=>"100000000",
  32177=>"010010001",
  32178=>"011010000",
  32179=>"100010100",
  32180=>"000111111",
  32181=>"111011000",
  32182=>"010010010",
  32183=>"010111101",
  32184=>"101111111",
  32185=>"100011000",
  32186=>"000111011",
  32187=>"010111011",
  32188=>"110010011",
  32189=>"011111111",
  32190=>"001000110",
  32191=>"010010011",
  32192=>"000000000",
  32193=>"010011000",
  32194=>"000111010",
  32195=>"100100100",
  32196=>"010010000",
  32197=>"110100101",
  32198=>"000011011",
  32199=>"000000001",
  32200=>"010100101",
  32201=>"110011000",
  32202=>"111111111",
  32203=>"011000000",
  32204=>"000001001",
  32205=>"000011000",
  32206=>"001001000",
  32207=>"111000000",
  32208=>"001000000",
  32209=>"001001011",
  32210=>"110010111",
  32211=>"001001000",
  32212=>"001000000",
  32213=>"110110111",
  32214=>"101000100",
  32215=>"110000000",
  32216=>"010000000",
  32217=>"111111111",
  32218=>"010010011",
  32219=>"111010000",
  32220=>"100100100",
  32221=>"110000000",
  32222=>"100000000",
  32223=>"011001000",
  32224=>"111000011",
  32225=>"111000111",
  32226=>"111111000",
  32227=>"111110110",
  32228=>"000000111",
  32229=>"000010111",
  32230=>"000000000",
  32231=>"011001110",
  32232=>"001111111",
  32233=>"000110100",
  32234=>"011111100",
  32235=>"000011010",
  32236=>"101101111",
  32237=>"111000011",
  32238=>"000000000",
  32239=>"101100111",
  32240=>"100100101",
  32241=>"011001001",
  32242=>"010000011",
  32243=>"100110000",
  32244=>"110110000",
  32245=>"001101100",
  32246=>"000000011",
  32247=>"000000000",
  32248=>"010010000",
  32249=>"010010101",
  32250=>"011100001",
  32251=>"001011110",
  32252=>"001000000",
  32253=>"100000100",
  32254=>"000000001",
  32255=>"110101111",
  32256=>"001011011",
  32257=>"111110000",
  32258=>"001000000",
  32259=>"111000000",
  32260=>"001111011",
  32261=>"101011011",
  32262=>"001111100",
  32263=>"000111111",
  32264=>"000001001",
  32265=>"100101101",
  32266=>"110100100",
  32267=>"000000000",
  32268=>"001000000",
  32269=>"000011000",
  32270=>"100100000",
  32271=>"111010011",
  32272=>"101000111",
  32273=>"000000010",
  32274=>"111001000",
  32275=>"111110000",
  32276=>"111010010",
  32277=>"010000000",
  32278=>"001001000",
  32279=>"000000111",
  32280=>"101111110",
  32281=>"010100111",
  32282=>"000100010",
  32283=>"000000000",
  32284=>"100110011",
  32285=>"110111100",
  32286=>"011000000",
  32287=>"010001101",
  32288=>"000111111",
  32289=>"101001100",
  32290=>"010001001",
  32291=>"000011111",
  32292=>"000001111",
  32293=>"100000110",
  32294=>"100111010",
  32295=>"000010110",
  32296=>"000010010",
  32297=>"111111110",
  32298=>"111101101",
  32299=>"111100000",
  32300=>"111100000",
  32301=>"001001001",
  32302=>"000000000",
  32303=>"001000100",
  32304=>"001101111",
  32305=>"000000000",
  32306=>"111111000",
  32307=>"111111110",
  32308=>"000000000",
  32309=>"111111101",
  32310=>"110000000",
  32311=>"110101101",
  32312=>"101000000",
  32313=>"000111000",
  32314=>"010011001",
  32315=>"010110111",
  32316=>"000000000",
  32317=>"111111001",
  32318=>"000010000",
  32319=>"001001011",
  32320=>"001000000",
  32321=>"111011110",
  32322=>"111010111",
  32323=>"001001111",
  32324=>"111001001",
  32325=>"001001100",
  32326=>"010010001",
  32327=>"000111011",
  32328=>"000001100",
  32329=>"000001101",
  32330=>"000100101",
  32331=>"010000000",
  32332=>"000001101",
  32333=>"000100101",
  32334=>"000110100",
  32335=>"111000010",
  32336=>"111001101",
  32337=>"010111111",
  32338=>"000011000",
  32339=>"001011011",
  32340=>"110111000",
  32341=>"000000000",
  32342=>"100101010",
  32343=>"101001111",
  32344=>"011010101",
  32345=>"011101011",
  32346=>"111101100",
  32347=>"001110010",
  32348=>"000000011",
  32349=>"010111001",
  32350=>"001000010",
  32351=>"100100100",
  32352=>"111001101",
  32353=>"111100000",
  32354=>"001001000",
  32355=>"110100100",
  32356=>"000110111",
  32357=>"010010110",
  32358=>"000000001",
  32359=>"100111010",
  32360=>"001010100",
  32361=>"000001000",
  32362=>"110111000",
  32363=>"100000000",
  32364=>"111111000",
  32365=>"111111110",
  32366=>"011111111",
  32367=>"010000000",
  32368=>"000010111",
  32369=>"011111111",
  32370=>"011001001",
  32371=>"101101110",
  32372=>"100100010",
  32373=>"000000000",
  32374=>"111000000",
  32375=>"000000101",
  32376=>"110101111",
  32377=>"010000000",
  32378=>"111101001",
  32379=>"000000011",
  32380=>"011001000",
  32381=>"100100100",
  32382=>"111111111",
  32383=>"111110010",
  32384=>"110100111",
  32385=>"100111000",
  32386=>"010000000",
  32387=>"111100100",
  32388=>"101111110",
  32389=>"111110010",
  32390=>"011000011",
  32391=>"011111011",
  32392=>"100101011",
  32393=>"000000010",
  32394=>"011111111",
  32395=>"000000001",
  32396=>"000011111",
  32397=>"111100101",
  32398=>"000011111",
  32399=>"110000000",
  32400=>"001011001",
  32401=>"000000000",
  32402=>"001001011",
  32403=>"111111000",
  32404=>"000000010",
  32405=>"000101101",
  32406=>"111011000",
  32407=>"000000001",
  32408=>"010011111",
  32409=>"000000000",
  32410=>"111111010",
  32411=>"111111001",
  32412=>"010111000",
  32413=>"100111000",
  32414=>"001111101",
  32415=>"110110000",
  32416=>"001011001",
  32417=>"110111111",
  32418=>"111101101",
  32419=>"010000111",
  32420=>"000111111",
  32421=>"100111011",
  32422=>"011011110",
  32423=>"110111111",
  32424=>"011000110",
  32425=>"001000110",
  32426=>"101100000",
  32427=>"111111111",
  32428=>"111010100",
  32429=>"101001100",
  32430=>"110110100",
  32431=>"101010011",
  32432=>"001001111",
  32433=>"011111001",
  32434=>"001111101",
  32435=>"000001000",
  32436=>"011101111",
  32437=>"111111111",
  32438=>"000000101",
  32439=>"000001000",
  32440=>"000000100",
  32441=>"010010110",
  32442=>"000000010",
  32443=>"001000001",
  32444=>"111000000",
  32445=>"111111111",
  32446=>"100100100",
  32447=>"111100001",
  32448=>"111010011",
  32449=>"000000010",
  32450=>"110000100",
  32451=>"001001000",
  32452=>"000000011",
  32453=>"100100001",
  32454=>"001000000",
  32455=>"000000000",
  32456=>"111111110",
  32457=>"000000010",
  32458=>"000110101",
  32459=>"100100110",
  32460=>"000100111",
  32461=>"110100001",
  32462=>"111111000",
  32463=>"000001111",
  32464=>"000000000",
  32465=>"001000011",
  32466=>"011111110",
  32467=>"111100101",
  32468=>"011000110",
  32469=>"111111100",
  32470=>"111111000",
  32471=>"010111010",
  32472=>"001111111",
  32473=>"000000000",
  32474=>"100101000",
  32475=>"001000110",
  32476=>"011000000",
  32477=>"100000000",
  32478=>"010110000",
  32479=>"000000101",
  32480=>"010111111",
  32481=>"110000000",
  32482=>"010010111",
  32483=>"011011111",
  32484=>"000110000",
  32485=>"000000000",
  32486=>"000000100",
  32487=>"111111011",
  32488=>"000101111",
  32489=>"111010000",
  32490=>"011011011",
  32491=>"101011111",
  32492=>"000000000",
  32493=>"000011011",
  32494=>"101111000",
  32495=>"001000101",
  32496=>"000110011",
  32497=>"001001101",
  32498=>"010000000",
  32499=>"110000000",
  32500=>"100110110",
  32501=>"011010110",
  32502=>"010000010",
  32503=>"010000100",
  32504=>"000000111",
  32505=>"111111011",
  32506=>"101111001",
  32507=>"110111001",
  32508=>"110000000",
  32509=>"111101000",
  32510=>"000111100",
  32511=>"000010100",
  32512=>"111101000",
  32513=>"110001110",
  32514=>"000000111",
  32515=>"101001111",
  32516=>"111101010",
  32517=>"100000000",
  32518=>"000000000",
  32519=>"000001000",
  32520=>"000110000",
  32521=>"000010110",
  32522=>"000000110",
  32523=>"000000000",
  32524=>"011000000",
  32525=>"111011010",
  32526=>"100111010",
  32527=>"000000000",
  32528=>"001111000",
  32529=>"000110110",
  32530=>"111111000",
  32531=>"000000000",
  32532=>"011111000",
  32533=>"111111111",
  32534=>"100100001",
  32535=>"111011111",
  32536=>"001000011",
  32537=>"110111111",
  32538=>"111111010",
  32539=>"000000011",
  32540=>"101111011",
  32541=>"111010110",
  32542=>"001111000",
  32543=>"011101000",
  32544=>"010000000",
  32545=>"111110000",
  32546=>"001000000",
  32547=>"000000000",
  32548=>"001001000",
  32549=>"001101100",
  32550=>"110110100",
  32551=>"001001000",
  32552=>"000000111",
  32553=>"001000101",
  32554=>"001110110",
  32555=>"000111111",
  32556=>"010011011",
  32557=>"000110010",
  32558=>"111111111",
  32559=>"101000101",
  32560=>"000011111",
  32561=>"000000001",
  32562=>"111111000",
  32563=>"000010111",
  32564=>"000000111",
  32565=>"000000000",
  32566=>"000111011",
  32567=>"001000000",
  32568=>"111111000",
  32569=>"111101001",
  32570=>"000111100",
  32571=>"000000001",
  32572=>"111111111",
  32573=>"101111001",
  32574=>"000000000",
  32575=>"101110110",
  32576=>"111111111",
  32577=>"101111110",
  32578=>"111000000",
  32579=>"011111111",
  32580=>"000000000",
  32581=>"111100011",
  32582=>"011000000",
  32583=>"000000101",
  32584=>"010111001",
  32585=>"111111111",
  32586=>"111001001",
  32587=>"110110000",
  32588=>"111111000",
  32589=>"000010110",
  32590=>"010001000",
  32591=>"111111111",
  32592=>"111111111",
  32593=>"110110010",
  32594=>"001000111",
  32595=>"001010000",
  32596=>"000000011",
  32597=>"110111110",
  32598=>"001001000",
  32599=>"111111111",
  32600=>"000000100",
  32601=>"001000001",
  32602=>"111001000",
  32603=>"011010000",
  32604=>"111111000",
  32605=>"111101001",
  32606=>"001000001",
  32607=>"010011011",
  32608=>"010110010",
  32609=>"010111011",
  32610=>"110100110",
  32611=>"001100100",
  32612=>"111101000",
  32613=>"111111001",
  32614=>"111111000",
  32615=>"000011111",
  32616=>"101101000",
  32617=>"011000010",
  32618=>"010000101",
  32619=>"111111000",
  32620=>"111111111",
  32621=>"000000000",
  32622=>"111001111",
  32623=>"110010000",
  32624=>"110100000",
  32625=>"100111111",
  32626=>"000111110",
  32627=>"000000011",
  32628=>"111000000",
  32629=>"000000000",
  32630=>"110111110",
  32631=>"111010000",
  32632=>"000000111",
  32633=>"111000000",
  32634=>"100000000",
  32635=>"000000000",
  32636=>"111111111",
  32637=>"110100000",
  32638=>"111111111",
  32639=>"011110110",
  32640=>"101111010",
  32641=>"110100000",
  32642=>"011011010",
  32643=>"011001000",
  32644=>"000000000",
  32645=>"101010000",
  32646=>"000111000",
  32647=>"110110110",
  32648=>"111111111",
  32649=>"111101000",
  32650=>"101011011",
  32651=>"101100101",
  32652=>"000000000",
  32653=>"111111110",
  32654=>"001111110",
  32655=>"000000011",
  32656=>"101111001",
  32657=>"111011000",
  32658=>"000000000",
  32659=>"100110000",
  32660=>"110111110",
  32661=>"100111111",
  32662=>"100001000",
  32663=>"010000000",
  32664=>"000000010",
  32665=>"010111010",
  32666=>"100111111",
  32667=>"000000000",
  32668=>"110100001",
  32669=>"000000111",
  32670=>"111000000",
  32671=>"000000010",
  32672=>"111111101",
  32673=>"111111111",
  32674=>"111111111",
  32675=>"001000111",
  32676=>"010110011",
  32677=>"110110010",
  32678=>"000000000",
  32679=>"011111111",
  32680=>"000000111",
  32681=>"110000111",
  32682=>"001000101",
  32683=>"000000110",
  32684=>"111111111",
  32685=>"111010110",
  32686=>"111101001",
  32687=>"000000001",
  32688=>"111000000",
  32689=>"111001001",
  32690=>"011011011",
  32691=>"101011000",
  32692=>"111011110",
  32693=>"111111111",
  32694=>"111101001",
  32695=>"001110101",
  32696=>"011111101",
  32697=>"111111111",
  32698=>"110100111",
  32699=>"010010111",
  32700=>"000000000",
  32701=>"111111110",
  32702=>"011001100",
  32703=>"110001111",
  32704=>"000011111",
  32705=>"111011011",
  32706=>"111110101",
  32707=>"111011110",
  32708=>"011000000",
  32709=>"111000100",
  32710=>"000000100",
  32711=>"011011000",
  32712=>"000000100",
  32713=>"111001000",
  32714=>"101001111",
  32715=>"111111011",
  32716=>"001111011",
  32717=>"011011101",
  32718=>"000000110",
  32719=>"000011000",
  32720=>"000000010",
  32721=>"100110000",
  32722=>"100000111",
  32723=>"001100000",
  32724=>"000000001",
  32725=>"100000000",
  32726=>"000000000",
  32727=>"010000000",
  32728=>"000000000",
  32729=>"100010000",
  32730=>"000011010",
  32731=>"001000110",
  32732=>"001010000",
  32733=>"011011011",
  32734=>"000000111",
  32735=>"101000010",
  32736=>"110111111",
  32737=>"000000111",
  32738=>"000000000",
  32739=>"111111000",
  32740=>"000000000",
  32741=>"000000000",
  32742=>"000000000",
  32743=>"011111010",
  32744=>"101000001",
  32745=>"000000000",
  32746=>"000001111",
  32747=>"111001000",
  32748=>"111000000",
  32749=>"001000010",
  32750=>"000010000",
  32751=>"010000000",
  32752=>"000000000",
  32753=>"111001001",
  32754=>"110111111",
  32755=>"010100000",
  32756=>"100011000",
  32757=>"101101111",
  32758=>"010110010",
  32759=>"000000111",
  32760=>"010110000",
  32761=>"111000000",
  32762=>"000001111",
  32763=>"111011000",
  32764=>"110010000",
  32765=>"101101111",
  32766=>"111100000",
  32767=>"001111111",
  32768=>"000100100",
  32769=>"100111110",
  32770=>"100100111",
  32771=>"000000011",
  32772=>"011111100",
  32773=>"000001000",
  32774=>"100100000",
  32775=>"001011011",
  32776=>"011011001",
  32777=>"000011011",
  32778=>"000000000",
  32779=>"000100011",
  32780=>"001011100",
  32781=>"100100111",
  32782=>"100001011",
  32783=>"110001011",
  32784=>"111010000",
  32785=>"000000000",
  32786=>"110110010",
  32787=>"111000000",
  32788=>"100100011",
  32789=>"000000000",
  32790=>"110111111",
  32791=>"111011010",
  32792=>"001111001",
  32793=>"111101100",
  32794=>"001011000",
  32795=>"000100110",
  32796=>"000010001",
  32797=>"100110110",
  32798=>"100000000",
  32799=>"111110100",
  32800=>"011011010",
  32801=>"011001101",
  32802=>"110000000",
  32803=>"001011000",
  32804=>"001111111",
  32805=>"011111110",
  32806=>"010011011",
  32807=>"000001000",
  32808=>"100100111",
  32809=>"010100110",
  32810=>"110000100",
  32811=>"110100111",
  32812=>"000001001",
  32813=>"100011001",
  32814=>"100110011",
  32815=>"111011011",
  32816=>"011010010",
  32817=>"100111011",
  32818=>"011011011",
  32819=>"110100000",
  32820=>"100100110",
  32821=>"101111010",
  32822=>"110100011",
  32823=>"011000011",
  32824=>"011110011",
  32825=>"000000011",
  32826=>"000000000",
  32827=>"100110000",
  32828=>"011111111",
  32829=>"011111100",
  32830=>"100000111",
  32831=>"001011001",
  32832=>"011000000",
  32833=>"011010000",
  32834=>"011011001",
  32835=>"011100100",
  32836=>"110101101",
  32837=>"100000000",
  32838=>"000011010",
  32839=>"001011111",
  32840=>"010010011",
  32841=>"001011010",
  32842=>"011100111",
  32843=>"000011110",
  32844=>"100000000",
  32845=>"110110011",
  32846=>"111100011",
  32847=>"111011011",
  32848=>"010000111",
  32849=>"110110111",
  32850=>"110111011",
  32851=>"001000010",
  32852=>"100100110",
  32853=>"100000000",
  32854=>"001001001",
  32855=>"110100011",
  32856=>"011100111",
  32857=>"010011011",
  32858=>"111001010",
  32859=>"010101111",
  32860=>"011011000",
  32861=>"001000001",
  32862=>"110100110",
  32863=>"000100000",
  32864=>"011011000",
  32865=>"011001011",
  32866=>"000111111",
  32867=>"011100111",
  32868=>"110110111",
  32869=>"011111011",
  32870=>"010000000",
  32871=>"111111011",
  32872=>"010011011",
  32873=>"001100000",
  32874=>"011011011",
  32875=>"000110100",
  32876=>"001111000",
  32877=>"100100111",
  32878=>"000010010",
  32879=>"001011011",
  32880=>"000001010",
  32881=>"011011011",
  32882=>"000000110",
  32883=>"100011000",
  32884=>"000001011",
  32885=>"010000000",
  32886=>"000010011",
  32887=>"000100100",
  32888=>"101000011",
  32889=>"111110110",
  32890=>"111100100",
  32891=>"100101101",
  32892=>"011011011",
  32893=>"110110000",
  32894=>"000100011",
  32895=>"000000110",
  32896=>"011000000",
  32897=>"110100110",
  32898=>"011011010",
  32899=>"000100011",
  32900=>"011011011",
  32901=>"101010000",
  32902=>"010001001",
  32903=>"111101000",
  32904=>"111011000",
  32905=>"000000000",
  32906=>"100100000",
  32907=>"001100000",
  32908=>"100100110",
  32909=>"000100101",
  32910=>"011000000",
  32911=>"111000010",
  32912=>"101111000",
  32913=>"000110100",
  32914=>"000001011",
  32915=>"011010000",
  32916=>"001011001",
  32917=>"100100100",
  32918=>"011011000",
  32919=>"010001001",
  32920=>"011011000",
  32921=>"000011011",
  32922=>"011011101",
  32923=>"011011011",
  32924=>"001110000",
  32925=>"011010111",
  32926=>"011011000",
  32927=>"101011001",
  32928=>"000000000",
  32929=>"000100111",
  32930=>"010111000",
  32931=>"111110111",
  32932=>"011111100",
  32933=>"001011000",
  32934=>"111001000",
  32935=>"001011000",
  32936=>"100011011",
  32937=>"000011011",
  32938=>"001000110",
  32939=>"001000100",
  32940=>"111000100",
  32941=>"011001011",
  32942=>"010110111",
  32943=>"011111011",
  32944=>"011011010",
  32945=>"101100100",
  32946=>"111100111",
  32947=>"100110111",
  32948=>"010011110",
  32949=>"110000100",
  32950=>"011010001",
  32951=>"111101110",
  32952=>"011011011",
  32953=>"001011000",
  32954=>"001000000",
  32955=>"000001010",
  32956=>"101010000",
  32957=>"110111111",
  32958=>"011011010",
  32959=>"100100001",
  32960=>"100100111",
  32961=>"100100110",
  32962=>"011010001",
  32963=>"100111100",
  32964=>"000000000",
  32965=>"101110000",
  32966=>"111110100",
  32967=>"010111111",
  32968=>"001001011",
  32969=>"100100100",
  32970=>"111111111",
  32971=>"000100111",
  32972=>"000001010",
  32973=>"000100011",
  32974=>"100000110",
  32975=>"011111011",
  32976=>"000000011",
  32977=>"111011001",
  32978=>"011011001",
  32979=>"100001011",
  32980=>"011011000",
  32981=>"111010101",
  32982=>"010000011",
  32983=>"001011011",
  32984=>"111110000",
  32985=>"100100000",
  32986=>"100110110",
  32987=>"100100100",
  32988=>"111101011",
  32989=>"110100100",
  32990=>"110001000",
  32991=>"100100110",
  32992=>"100000010",
  32993=>"100100111",
  32994=>"000000010",
  32995=>"101111001",
  32996=>"111100111",
  32997=>"100100100",
  32998=>"001000001",
  32999=>"001010011",
  33000=>"000011001",
  33001=>"110111111",
  33002=>"010000000",
  33003=>"000100111",
  33004=>"000100110",
  33005=>"000000011",
  33006=>"110100100",
  33007=>"011010000",
  33008=>"101010000",
  33009=>"110110111",
  33010=>"000000011",
  33011=>"100100111",
  33012=>"010000011",
  33013=>"111001101",
  33014=>"000011011",
  33015=>"011000110",
  33016=>"100100111",
  33017=>"010000000",
  33018=>"110110111",
  33019=>"101111001",
  33020=>"011011000",
  33021=>"011110110",
  33022=>"011011000",
  33023=>"011011011",
  33024=>"010000000",
  33025=>"011011010",
  33026=>"000000111",
  33027=>"001000010",
  33028=>"100001001",
  33029=>"000100111",
  33030=>"001111011",
  33031=>"000011010",
  33032=>"010000111",
  33033=>"111011101",
  33034=>"011001111",
  33035=>"001000111",
  33036=>"000000111",
  33037=>"000001010",
  33038=>"101011010",
  33039=>"110111000",
  33040=>"111011010",
  33041=>"000000000",
  33042=>"101000000",
  33043=>"010000000",
  33044=>"011111001",
  33045=>"000000100",
  33046=>"000000100",
  33047=>"100011110",
  33048=>"010001111",
  33049=>"101111010",
  33050=>"000101011",
  33051=>"100000110",
  33052=>"111111001",
  33053=>"000111111",
  33054=>"000000010",
  33055=>"000100100",
  33056=>"111000000",
  33057=>"010010011",
  33058=>"111100100",
  33059=>"111110010",
  33060=>"000110000",
  33061=>"010110000",
  33062=>"011000010",
  33063=>"000011011",
  33064=>"000000000",
  33065=>"000111011",
  33066=>"111011010",
  33067=>"001100000",
  33068=>"011001011",
  33069=>"111000010",
  33070=>"000001010",
  33071=>"100111110",
  33072=>"000000000",
  33073=>"000000001",
  33074=>"000101100",
  33075=>"010000000",
  33076=>"000000101",
  33077=>"101000111",
  33078=>"110010010",
  33079=>"111010000",
  33080=>"011010000",
  33081=>"001001000",
  33082=>"000100001",
  33083=>"000000000",
  33084=>"000000000",
  33085=>"111101110",
  33086=>"001100100",
  33087=>"011011101",
  33088=>"100101111",
  33089=>"111111101",
  33090=>"000000101",
  33091=>"000000010",
  33092=>"101101001",
  33093=>"000000100",
  33094=>"000000001",
  33095=>"010111000",
  33096=>"100001001",
  33097=>"110111100",
  33098=>"110000001",
  33099=>"000010001",
  33100=>"000000000",
  33101=>"110111111",
  33102=>"011100110",
  33103=>"010110100",
  33104=>"010000101",
  33105=>"111000011",
  33106=>"011011101",
  33107=>"000001100",
  33108=>"000010010",
  33109=>"100110100",
  33110=>"100111110",
  33111=>"011000111",
  33112=>"000001101",
  33113=>"000001001",
  33114=>"000111001",
  33115=>"011011100",
  33116=>"011010110",
  33117=>"000001000",
  33118=>"111111111",
  33119=>"000100111",
  33120=>"111101111",
  33121=>"000101011",
  33122=>"101000111",
  33123=>"000100100",
  33124=>"100010000",
  33125=>"100001111",
  33126=>"110100110",
  33127=>"111000100",
  33128=>"101001101",
  33129=>"010000111",
  33130=>"101011111",
  33131=>"110001101",
  33132=>"000000000",
  33133=>"001010010",
  33134=>"000000011",
  33135=>"000001000",
  33136=>"001100000",
  33137=>"000001010",
  33138=>"011011011",
  33139=>"000000111",
  33140=>"111101001",
  33141=>"001000101",
  33142=>"101001010",
  33143=>"111100100",
  33144=>"001000011",
  33145=>"111111011",
  33146=>"111111010",
  33147=>"000101111",
  33148=>"100110110",
  33149=>"000100001",
  33150=>"100101101",
  33151=>"000100101",
  33152=>"010011000",
  33153=>"000000000",
  33154=>"010000001",
  33155=>"101111110",
  33156=>"000000111",
  33157=>"001101010",
  33158=>"010011000",
  33159=>"001011011",
  33160=>"000100010",
  33161=>"000000010",
  33162=>"111011111",
  33163=>"000000111",
  33164=>"101000000",
  33165=>"011111111",
  33166=>"000000000",
  33167=>"001000100",
  33168=>"001001101",
  33169=>"111111000",
  33170=>"011011000",
  33171=>"000000111",
  33172=>"100011110",
  33173=>"000000010",
  33174=>"111011010",
  33175=>"000111000",
  33176=>"110010100",
  33177=>"011111111",
  33178=>"111100111",
  33179=>"011001001",
  33180=>"111101101",
  33181=>"101101111",
  33182=>"010011111",
  33183=>"000111111",
  33184=>"101011101",
  33185=>"111000000",
  33186=>"000010000",
  33187=>"010000101",
  33188=>"000111111",
  33189=>"110110000",
  33190=>"111110001",
  33191=>"011101010",
  33192=>"000000010",
  33193=>"111000000",
  33194=>"101101111",
  33195=>"000000000",
  33196=>"101111010",
  33197=>"100000101",
  33198=>"110110000",
  33199=>"111111111",
  33200=>"000101010",
  33201=>"001101111",
  33202=>"101101111",
  33203=>"100100010",
  33204=>"010110001",
  33205=>"100100111",
  33206=>"001011000",
  33207=>"111011101",
  33208=>"100100001",
  33209=>"000110111",
  33210=>"110000000",
  33211=>"011011000",
  33212=>"010111001",
  33213=>"001111111",
  33214=>"100100101",
  33215=>"000000010",
  33216=>"000000100",
  33217=>"101001110",
  33218=>"101111010",
  33219=>"000000011",
  33220=>"010011000",
  33221=>"110110010",
  33222=>"100011011",
  33223=>"011111100",
  33224=>"000111011",
  33225=>"010111000",
  33226=>"111111000",
  33227=>"000110100",
  33228=>"101000001",
  33229=>"100011011",
  33230=>"101111010",
  33231=>"111000000",
  33232=>"111101111",
  33233=>"011111110",
  33234=>"101010010",
  33235=>"000000111",
  33236=>"001000011",
  33237=>"100001000",
  33238=>"010101011",
  33239=>"000000100",
  33240=>"000000010",
  33241=>"111101000",
  33242=>"011111110",
  33243=>"001000001",
  33244=>"000000010",
  33245=>"111001101",
  33246=>"001000001",
  33247=>"000001010",
  33248=>"101000101",
  33249=>"000000011",
  33250=>"001100100",
  33251=>"111111011",
  33252=>"100000100",
  33253=>"101101000",
  33254=>"110000000",
  33255=>"111011000",
  33256=>"011101010",
  33257=>"111111110",
  33258=>"110011011",
  33259=>"100000101",
  33260=>"000100000",
  33261=>"010001010",
  33262=>"010000010",
  33263=>"010100000",
  33264=>"000010000",
  33265=>"001011111",
  33266=>"111000110",
  33267=>"001101101",
  33268=>"110001001",
  33269=>"111111111",
  33270=>"000000011",
  33271=>"011101011",
  33272=>"010010000",
  33273=>"001001100",
  33274=>"000111110",
  33275=>"000111111",
  33276=>"000000000",
  33277=>"010011000",
  33278=>"000001011",
  33279=>"101000100",
  33280=>"000000000",
  33281=>"010010010",
  33282=>"100001001",
  33283=>"010011110",
  33284=>"100111011",
  33285=>"111110100",
  33286=>"100111101",
  33287=>"000100111",
  33288=>"000000100",
  33289=>"000001000",
  33290=>"000000010",
  33291=>"111110100",
  33292=>"101110100",
  33293=>"101110101",
  33294=>"111111111",
  33295=>"111111111",
  33296=>"001101011",
  33297=>"000011010",
  33298=>"000010000",
  33299=>"111011110",
  33300=>"110111111",
  33301=>"000000011",
  33302=>"000000110",
  33303=>"111110010",
  33304=>"101001001",
  33305=>"101101100",
  33306=>"100000110",
  33307=>"000011011",
  33308=>"110111011",
  33309=>"100010000",
  33310=>"110110010",
  33311=>"000000000",
  33312=>"000001011",
  33313=>"110110101",
  33314=>"100100001",
  33315=>"000000000",
  33316=>"111110000",
  33317=>"011110000",
  33318=>"000001010",
  33319=>"011110110",
  33320=>"000000100",
  33321=>"000010110",
  33322=>"000100110",
  33323=>"100100000",
  33324=>"011111100",
  33325=>"011000000",
  33326=>"111100000",
  33327=>"100100001",
  33328=>"110100100",
  33329=>"000111111",
  33330=>"100100101",
  33331=>"100100000",
  33332=>"000001011",
  33333=>"001001011",
  33334=>"011110100",
  33335=>"111111110",
  33336=>"110100100",
  33337=>"100011010",
  33338=>"100001011",
  33339=>"010100000",
  33340=>"001001000",
  33341=>"001111111",
  33342=>"000000001",
  33343=>"010100000",
  33344=>"011111001",
  33345=>"100100100",
  33346=>"110111111",
  33347=>"000000000",
  33348=>"111001000",
  33349=>"000000000",
  33350=>"001100110",
  33351=>"111101100",
  33352=>"101101100",
  33353=>"010111111",
  33354=>"100000000",
  33355=>"100000001",
  33356=>"100101000",
  33357=>"001011011",
  33358=>"011010000",
  33359=>"000011001",
  33360=>"100111000",
  33361=>"110010011",
  33362=>"011100001",
  33363=>"000000000",
  33364=>"111111001",
  33365=>"001101000",
  33366=>"000100100",
  33367=>"000011011",
  33368=>"111111111",
  33369=>"001111111",
  33370=>"001011000",
  33371=>"000100101",
  33372=>"000001111",
  33373=>"001001011",
  33374=>"111000011",
  33375=>"111100111",
  33376=>"111110100",
  33377=>"011011011",
  33378=>"100000011",
  33379=>"110011011",
  33380=>"000000000",
  33381=>"010110100",
  33382=>"011101100",
  33383=>"111101110",
  33384=>"111111100",
  33385=>"011111110",
  33386=>"011110110",
  33387=>"111011111",
  33388=>"000100000",
  33389=>"000001011",
  33390=>"000000001",
  33391=>"011011011",
  33392=>"011011010",
  33393=>"011110010",
  33394=>"000000000",
  33395=>"000100000",
  33396=>"111111111",
  33397=>"000010000",
  33398=>"000001011",
  33399=>"001011010",
  33400=>"100000000",
  33401=>"111111100",
  33402=>"110100100",
  33403=>"010000000",
  33404=>"000000000",
  33405=>"111111100",
  33406=>"111110000",
  33407=>"101001011",
  33408=>"110100110",
  33409=>"100110100",
  33410=>"000110110",
  33411=>"001100001",
  33412=>"111100000",
  33413=>"001100000",
  33414=>"110110010",
  33415=>"000011011",
  33416=>"001111101",
  33417=>"100000001",
  33418=>"001100100",
  33419=>"101100001",
  33420=>"101011000",
  33421=>"100100001",
  33422=>"101001111",
  33423=>"001001001",
  33424=>"000010000",
  33425=>"001011011",
  33426=>"000000000",
  33427=>"011001011",
  33428=>"011011000",
  33429=>"100001011",
  33430=>"001011000",
  33431=>"100000111",
  33432=>"000110100",
  33433=>"100000011",
  33434=>"111001001",
  33435=>"000000011",
  33436=>"001011011",
  33437=>"110111111",
  33438=>"000010001",
  33439=>"000001001",
  33440=>"000010101",
  33441=>"110000011",
  33442=>"001000101",
  33443=>"111001000",
  33444=>"111110100",
  33445=>"111101010",
  33446=>"001000010",
  33447=>"011110100",
  33448=>"000000000",
  33449=>"001000001",
  33450=>"111000001",
  33451=>"000000001",
  33452=>"001001000",
  33453=>"100010000",
  33454=>"111111111",
  33455=>"001010011",
  33456=>"000000110",
  33457=>"000000000",
  33458=>"110000000",
  33459=>"000000000",
  33460=>"000111100",
  33461=>"011101000",
  33462=>"001101101",
  33463=>"001100101",
  33464=>"000100100",
  33465=>"000000110",
  33466=>"111101011",
  33467=>"010111010",
  33468=>"000000100",
  33469=>"111110100",
  33470=>"000000100",
  33471=>"000000001",
  33472=>"000001010",
  33473=>"000001011",
  33474=>"010110111",
  33475=>"011111100",
  33476=>"001000000",
  33477=>"010000001",
  33478=>"111111111",
  33479=>"100110110",
  33480=>"000000101",
  33481=>"101001001",
  33482=>"111010001",
  33483=>"001011000",
  33484=>"001011011",
  33485=>"111011111",
  33486=>"000000001",
  33487=>"011110001",
  33488=>"000110100",
  33489=>"011010000",
  33490=>"001001001",
  33491=>"111110100",
  33492=>"100000001",
  33493=>"001011110",
  33494=>"110000010",
  33495=>"101111110",
  33496=>"101110100",
  33497=>"001000100",
  33498=>"111000000",
  33499=>"110001011",
  33500=>"111110000",
  33501=>"101001010",
  33502=>"001010000",
  33503=>"011110000",
  33504=>"000001001",
  33505=>"000001001",
  33506=>"111000100",
  33507=>"000001001",
  33508=>"000000000",
  33509=>"000001000",
  33510=>"001111100",
  33511=>"000000000",
  33512=>"000110110",
  33513=>"000000000",
  33514=>"010111111",
  33515=>"000000110",
  33516=>"000011110",
  33517=>"111001001",
  33518=>"000000000",
  33519=>"000000100",
  33520=>"000100100",
  33521=>"000111111",
  33522=>"110000110",
  33523=>"010000000",
  33524=>"111111111",
  33525=>"100100000",
  33526=>"100001101",
  33527=>"011110101",
  33528=>"110010010",
  33529=>"111111111",
  33530=>"100101011",
  33531=>"000010100",
  33532=>"111111110",
  33533=>"000000110",
  33534=>"011111111",
  33535=>"110110110",
  33536=>"100110110",
  33537=>"001101101",
  33538=>"111010000",
  33539=>"000000000",
  33540=>"001001000",
  33541=>"101111111",
  33542=>"111010000",
  33543=>"111000011",
  33544=>"001001001",
  33545=>"101000000",
  33546=>"110100110",
  33547=>"111111001",
  33548=>"111111100",
  33549=>"111001000",
  33550=>"010000000",
  33551=>"110010011",
  33552=>"100101011",
  33553=>"000000000",
  33554=>"000000000",
  33555=>"111101101",
  33556=>"111110000",
  33557=>"111111000",
  33558=>"000000001",
  33559=>"110110010",
  33560=>"111111111",
  33561=>"000101111",
  33562=>"111111111",
  33563=>"111111000",
  33564=>"001100000",
  33565=>"011000001",
  33566=>"001000010",
  33567=>"000000000",
  33568=>"111111111",
  33569=>"111010111",
  33570=>"000000000",
  33571=>"111111101",
  33572=>"001000000",
  33573=>"111111111",
  33574=>"111010000",
  33575=>"000100011",
  33576=>"000011000",
  33577=>"111101111",
  33578=>"000000000",
  33579=>"111111111",
  33580=>"111111001",
  33581=>"111111111",
  33582=>"000100111",
  33583=>"001000001",
  33584=>"100000111",
  33585=>"000000000",
  33586=>"010010111",
  33587=>"010111111",
  33588=>"011001000",
  33589=>"111101101",
  33590=>"100000000",
  33591=>"010110110",
  33592=>"000000100",
  33593=>"111111000",
  33594=>"000000000",
  33595=>"001000110",
  33596=>"111011011",
  33597=>"111001001",
  33598=>"000000001",
  33599=>"001001010",
  33600=>"111101111",
  33601=>"101101110",
  33602=>"000000111",
  33603=>"100000101",
  33604=>"111101110",
  33605=>"000000000",
  33606=>"011011011",
  33607=>"000101111",
  33608=>"101111111",
  33609=>"110100111",
  33610=>"000000000",
  33611=>"111101001",
  33612=>"100100010",
  33613=>"000000000",
  33614=>"000000000",
  33615=>"111101111",
  33616=>"000000000",
  33617=>"111010111",
  33618=>"011111111",
  33619=>"000000000",
  33620=>"000101001",
  33621=>"000011000",
  33622=>"001001000",
  33623=>"010000000",
  33624=>"001011001",
  33625=>"100000000",
  33626=>"011001000",
  33627=>"000000101",
  33628=>"000000000",
  33629=>"000000000",
  33630=>"111111110",
  33631=>"001000000",
  33632=>"101101111",
  33633=>"111111111",
  33634=>"000000110",
  33635=>"000000000",
  33636=>"000000000",
  33637=>"101000001",
  33638=>"111111000",
  33639=>"011011000",
  33640=>"000000000",
  33641=>"111010111",
  33642=>"000010001",
  33643=>"111111111",
  33644=>"111111110",
  33645=>"111111111",
  33646=>"111110111",
  33647=>"000011100",
  33648=>"000000000",
  33649=>"111010111",
  33650=>"001000000",
  33651=>"111111111",
  33652=>"000000111",
  33653=>"000000000",
  33654=>"110000000",
  33655=>"100000111",
  33656=>"111111010",
  33657=>"101011000",
  33658=>"111111011",
  33659=>"001000000",
  33660=>"011000000",
  33661=>"000000000",
  33662=>"111111111",
  33663=>"001000000",
  33664=>"000000011",
  33665=>"111000000",
  33666=>"111000000",
  33667=>"010000000",
  33668=>"000001010",
  33669=>"110101101",
  33670=>"100100111",
  33671=>"100100001",
  33672=>"000100001",
  33673=>"101101101",
  33674=>"000000000",
  33675=>"000000100",
  33676=>"111111110",
  33677=>"101011110",
  33678=>"000000100",
  33679=>"000000000",
  33680=>"000000000",
  33681=>"010010111",
  33682=>"010000111",
  33683=>"110111011",
  33684=>"010101100",
  33685=>"000000000",
  33686=>"111111111",
  33687=>"000000001",
  33688=>"101101101",
  33689=>"111111101",
  33690=>"010111100",
  33691=>"111001111",
  33692=>"010111100",
  33693=>"111111101",
  33694=>"001000001",
  33695=>"100000000",
  33696=>"100000000",
  33697=>"000011000",
  33698=>"101000001",
  33699=>"111111010",
  33700=>"110101101",
  33701=>"001001001",
  33702=>"000000001",
  33703=>"111111110",
  33704=>"110000001",
  33705=>"110111100",
  33706=>"111111000",
  33707=>"000010110",
  33708=>"011001000",
  33709=>"000000000",
  33710=>"101110010",
  33711=>"110100111",
  33712=>"000001010",
  33713=>"111101011",
  33714=>"000000000",
  33715=>"000000000",
  33716=>"000100000",
  33717=>"111111011",
  33718=>"000010000",
  33719=>"110110001",
  33720=>"100011110",
  33721=>"010101101",
  33722=>"000111111",
  33723=>"011111001",
  33724=>"111111111",
  33725=>"111000000",
  33726=>"001000100",
  33727=>"111110111",
  33728=>"101110001",
  33729=>"101101101",
  33730=>"000001000",
  33731=>"000000100",
  33732=>"010010000",
  33733=>"001011111",
  33734=>"111101000",
  33735=>"110110110",
  33736=>"000100000",
  33737=>"000000000",
  33738=>"000101000",
  33739=>"111101111",
  33740=>"011101110",
  33741=>"110100000",
  33742=>"001000000",
  33743=>"000000000",
  33744=>"000000000",
  33745=>"001001001",
  33746=>"101110111",
  33747=>"000000011",
  33748=>"000001111",
  33749=>"111001100",
  33750=>"111111110",
  33751=>"000000111",
  33752=>"111111001",
  33753=>"111111111",
  33754=>"001001001",
  33755=>"000000010",
  33756=>"000001001",
  33757=>"100000000",
  33758=>"110101001",
  33759=>"111001111",
  33760=>"101011111",
  33761=>"010001111",
  33762=>"000000000",
  33763=>"101011011",
  33764=>"000000001",
  33765=>"111111000",
  33766=>"000100000",
  33767=>"101111101",
  33768=>"000000001",
  33769=>"111110111",
  33770=>"001001000",
  33771=>"111101110",
  33772=>"010000000",
  33773=>"000000111",
  33774=>"000000000",
  33775=>"000000110",
  33776=>"111111000",
  33777=>"100110111",
  33778=>"000101101",
  33779=>"001001000",
  33780=>"001001001",
  33781=>"100001011",
  33782=>"000000101",
  33783=>"000000101",
  33784=>"111000110",
  33785=>"000000111",
  33786=>"111111111",
  33787=>"111110111",
  33788=>"001001111",
  33789=>"111111000",
  33790=>"001000001",
  33791=>"010000001",
  33792=>"100100110",
  33793=>"111111000",
  33794=>"000010110",
  33795=>"111001000",
  33796=>"011010000",
  33797=>"001111111",
  33798=>"111101000",
  33799=>"010010000",
  33800=>"101111011",
  33801=>"001000001",
  33802=>"110111111",
  33803=>"111001000",
  33804=>"000110111",
  33805=>"110101001",
  33806=>"001011000",
  33807=>"000101110",
  33808=>"111111000",
  33809=>"111000000",
  33810=>"110110111",
  33811=>"111001000",
  33812=>"000110111",
  33813=>"000111111",
  33814=>"010100000",
  33815=>"111000100",
  33816=>"010101111",
  33817=>"110011111",
  33818=>"111000000",
  33819=>"111001000",
  33820=>"000011000",
  33821=>"000001110",
  33822=>"000001011",
  33823=>"001001111",
  33824=>"110000101",
  33825=>"001000000",
  33826=>"001000000",
  33827=>"111111000",
  33828=>"100100110",
  33829=>"111100000",
  33830=>"000010111",
  33831=>"000000000",
  33832=>"000111111",
  33833=>"111001000",
  33834=>"000000000",
  33835=>"111000101",
  33836=>"011100111",
  33837=>"110110010",
  33838=>"010111111",
  33839=>"011111111",
  33840=>"101000000",
  33841=>"111000010",
  33842=>"000110000",
  33843=>"000000000",
  33844=>"111000000",
  33845=>"111111111",
  33846=>"110100000",
  33847=>"101001001",
  33848=>"110110110",
  33849=>"111101111",
  33850=>"000000000",
  33851=>"110000000",
  33852=>"001100000",
  33853=>"001000001",
  33854=>"001100000",
  33855=>"011011000",
  33856=>"000111111",
  33857=>"101111000",
  33858=>"111001000",
  33859=>"100110111",
  33860=>"000000000",
  33861=>"000111100",
  33862=>"111111000",
  33863=>"001111111",
  33864=>"101100000",
  33865=>"101101001",
  33866=>"000110110",
  33867=>"011000000",
  33868=>"111000000",
  33869=>"011011110",
  33870=>"111011011",
  33871=>"000001111",
  33872=>"001001001",
  33873=>"111110101",
  33874=>"111001000",
  33875=>"000010010",
  33876=>"011111000",
  33877=>"000100000",
  33878=>"011001001",
  33879=>"010111110",
  33880=>"000000001",
  33881=>"100000000",
  33882=>"000000000",
  33883=>"111001001",
  33884=>"000000000",
  33885=>"000110011",
  33886=>"000111111",
  33887=>"011111111",
  33888=>"111001000",
  33889=>"000010110",
  33890=>"111000000",
  33891=>"001011101",
  33892=>"000000010",
  33893=>"001001111",
  33894=>"111101111",
  33895=>"000000010",
  33896=>"000000000",
  33897=>"000000000",
  33898=>"011111001",
  33899=>"001011010",
  33900=>"111101000",
  33901=>"111111111",
  33902=>"000000111",
  33903=>"110111000",
  33904=>"011110100",
  33905=>"000000000",
  33906=>"111001001",
  33907=>"000110000",
  33908=>"110000000",
  33909=>"110111000",
  33910=>"000000000",
  33911=>"111111100",
  33912=>"000111010",
  33913=>"111001000",
  33914=>"000000000",
  33915=>"010110110",
  33916=>"011001000",
  33917=>"000011110",
  33918=>"000010110",
  33919=>"000010111",
  33920=>"111101000",
  33921=>"111001001",
  33922=>"101000000",
  33923=>"000000100",
  33924=>"000000000",
  33925=>"001000001",
  33926=>"111011000",
  33927=>"101000001",
  33928=>"010011001",
  33929=>"111001000",
  33930=>"000111111",
  33931=>"111111000",
  33932=>"111000000",
  33933=>"001100000",
  33934=>"000011100",
  33935=>"111011101",
  33936=>"010011011",
  33937=>"000001000",
  33938=>"111000000",
  33939=>"110111000",
  33940=>"000000010",
  33941=>"101001000",
  33942=>"110100110",
  33943=>"000000000",
  33944=>"111001010",
  33945=>"000011000",
  33946=>"001001011",
  33947=>"000111110",
  33948=>"111101000",
  33949=>"110011101",
  33950=>"101011101",
  33951=>"111001010",
  33952=>"111000111",
  33953=>"010011000",
  33954=>"000111111",
  33955=>"111001001",
  33956=>"111100000",
  33957=>"110100010",
  33958=>"000000111",
  33959=>"111101000",
  33960=>"111110000",
  33961=>"110000000",
  33962=>"000011111",
  33963=>"110110000",
  33964=>"110010110",
  33965=>"000100111",
  33966=>"000011011",
  33967=>"000111111",
  33968=>"000000000",
  33969=>"111001000",
  33970=>"000110000",
  33971=>"001001011",
  33972=>"110001001",
  33973=>"000100000",
  33974=>"110000000",
  33975=>"001110011",
  33976=>"000001001",
  33977=>"000000100",
  33978=>"101101011",
  33979=>"000000010",
  33980=>"010111111",
  33981=>"111111000",
  33982=>"110100000",
  33983=>"101000100",
  33984=>"000110111",
  33985=>"010001001",
  33986=>"100000000",
  33987=>"111111111",
  33988=>"011111110",
  33989=>"000100101",
  33990=>"000001000",
  33991=>"000000101",
  33992=>"011111000",
  33993=>"111000101",
  33994=>"001000000",
  33995=>"111010000",
  33996=>"011010000",
  33997=>"100100001",
  33998=>"101001001",
  33999=>"011000000",
  34000=>"111100101",
  34001=>"111010010",
  34002=>"100000000",
  34003=>"000000000",
  34004=>"001111000",
  34005=>"110000011",
  34006=>"001111111",
  34007=>"110111010",
  34008=>"000111111",
  34009=>"000000000",
  34010=>"111101111",
  34011=>"111000000",
  34012=>"000000001",
  34013=>"111101111",
  34014=>"000000001",
  34015=>"110101001",
  34016=>"000111111",
  34017=>"001111111",
  34018=>"000000010",
  34019=>"010110010",
  34020=>"000010110",
  34021=>"111000000",
  34022=>"111011011",
  34023=>"001001111",
  34024=>"100001000",
  34025=>"110110010",
  34026=>"110111110",
  34027=>"000000000",
  34028=>"000111111",
  34029=>"011111111",
  34030=>"000010000",
  34031=>"111000000",
  34032=>"000000000",
  34033=>"001011000",
  34034=>"000001000",
  34035=>"000100100",
  34036=>"001011000",
  34037=>"000001111",
  34038=>"100101011",
  34039=>"000000110",
  34040=>"101111000",
  34041=>"111110000",
  34042=>"110110101",
  34043=>"001001110",
  34044=>"000111011",
  34045=>"000001000",
  34046=>"111101011",
  34047=>"010111011",
  34048=>"000100110",
  34049=>"011101100",
  34050=>"000011100",
  34051=>"011111101",
  34052=>"110001011",
  34053=>"111101101",
  34054=>"011100101",
  34055=>"000010000",
  34056=>"101100000",
  34057=>"000111101",
  34058=>"001000000",
  34059=>"101000100",
  34060=>"111111111",
  34061=>"100101110",
  34062=>"110100100",
  34063=>"000000000",
  34064=>"101100100",
  34065=>"101100000",
  34066=>"111111011",
  34067=>"111101101",
  34068=>"000011000",
  34069=>"000100000",
  34070=>"000000100",
  34071=>"111111111",
  34072=>"000000101",
  34073=>"100001101",
  34074=>"000000000",
  34075=>"000111110",
  34076=>"010011110",
  34077=>"001010011",
  34078=>"000111101",
  34079=>"111111111",
  34080=>"000000000",
  34081=>"101100000",
  34082=>"011111000",
  34083=>"101000000",
  34084=>"001111010",
  34085=>"100000110",
  34086=>"000100000",
  34087=>"000000000",
  34088=>"100111111",
  34089=>"000111011",
  34090=>"100010010",
  34091=>"110111111",
  34092=>"100100100",
  34093=>"000000000",
  34094=>"010010010",
  34095=>"001111100",
  34096=>"000111111",
  34097=>"100000110",
  34098=>"111100101",
  34099=>"000000100",
  34100=>"100000111",
  34101=>"000000000",
  34102=>"100100001",
  34103=>"000100100",
  34104=>"011000111",
  34105=>"010000000",
  34106=>"001111010",
  34107=>"111111111",
  34108=>"010111010",
  34109=>"111101111",
  34110=>"100000111",
  34111=>"001001001",
  34112=>"111110111",
  34113=>"110100111",
  34114=>"111101000",
  34115=>"000000100",
  34116=>"100000100",
  34117=>"100111111",
  34118=>"111111111",
  34119=>"111011011",
  34120=>"010110101",
  34121=>"000010000",
  34122=>"001111100",
  34123=>"000111111",
  34124=>"110100100",
  34125=>"010011001",
  34126=>"011110100",
  34127=>"001100100",
  34128=>"000000000",
  34129=>"101111111",
  34130=>"011111111",
  34131=>"010111111",
  34132=>"101000000",
  34133=>"000101000",
  34134=>"000110100",
  34135=>"000011111",
  34136=>"000001111",
  34137=>"111110110",
  34138=>"010000001",
  34139=>"110011000",
  34140=>"100100101",
  34141=>"010010000",
  34142=>"000011110",
  34143=>"000000000",
  34144=>"101101111",
  34145=>"111111111",
  34146=>"100110000",
  34147=>"011000010",
  34148=>"111111111",
  34149=>"001001001",
  34150=>"000000000",
  34151=>"000101111",
  34152=>"000000100",
  34153=>"100000010",
  34154=>"111011010",
  34155=>"110000000",
  34156=>"001111010",
  34157=>"111011111",
  34158=>"000000000",
  34159=>"100000100",
  34160=>"001000001",
  34161=>"110111100",
  34162=>"001000000",
  34163=>"111111011",
  34164=>"111111010",
  34165=>"010000010",
  34166=>"100000000",
  34167=>"000111000",
  34168=>"111000110",
  34169=>"111110010",
  34170=>"111000100",
  34171=>"011000000",
  34172=>"011001000",
  34173=>"010011010",
  34174=>"000011111",
  34175=>"111100110",
  34176=>"000100100",
  34177=>"011011011",
  34178=>"100000000",
  34179=>"100000000",
  34180=>"111000000",
  34181=>"101010010",
  34182=>"000100100",
  34183=>"001000100",
  34184=>"110110110",
  34185=>"000100000",
  34186=>"000000000",
  34187=>"111111011",
  34188=>"111111111",
  34189=>"000000101",
  34190=>"011000000",
  34191=>"000111000",
  34192=>"110011111",
  34193=>"101000010",
  34194=>"111000000",
  34195=>"111111011",
  34196=>"001100011",
  34197=>"101110100",
  34198=>"101101000",
  34199=>"110110010",
  34200=>"111101011",
  34201=>"111000001",
  34202=>"000011000",
  34203=>"111111111",
  34204=>"110100001",
  34205=>"111100111",
  34206=>"101100111",
  34207=>"111111111",
  34208=>"001100111",
  34209=>"000000000",
  34210=>"000000000",
  34211=>"000100101",
  34212=>"000000010",
  34213=>"000000000",
  34214=>"110110110",
  34215=>"101000000",
  34216=>"101001000",
  34217=>"010010011",
  34218=>"100000000",
  34219=>"111011111",
  34220=>"010001000",
  34221=>"000000000",
  34222=>"101000000",
  34223=>"101001010",
  34224=>"111011111",
  34225=>"000010010",
  34226=>"111001100",
  34227=>"011001000",
  34228=>"101001001",
  34229=>"001000101",
  34230=>"100010000",
  34231=>"010010000",
  34232=>"110100101",
  34233=>"111101101",
  34234=>"111011010",
  34235=>"011001000",
  34236=>"000000011",
  34237=>"010011011",
  34238=>"110100110",
  34239=>"000000110",
  34240=>"000000000",
  34241=>"000000100",
  34242=>"110000000",
  34243=>"001011001",
  34244=>"000000010",
  34245=>"000011100",
  34246=>"011111000",
  34247=>"110011000",
  34248=>"010110101",
  34249=>"111111111",
  34250=>"111000100",
  34251=>"000000000",
  34252=>"111101110",
  34253=>"111110101",
  34254=>"111100010",
  34255=>"111111111",
  34256=>"111010000",
  34257=>"011011011",
  34258=>"100110111",
  34259=>"000101001",
  34260=>"101000000",
  34261=>"000010011",
  34262=>"111111011",
  34263=>"111111101",
  34264=>"001101100",
  34265=>"100000000",
  34266=>"010001001",
  34267=>"111111111",
  34268=>"000001000",
  34269=>"111110101",
  34270=>"111111111",
  34271=>"101111111",
  34272=>"000000100",
  34273=>"000010000",
  34274=>"100000011",
  34275=>"001001000",
  34276=>"000010000",
  34277=>"000000000",
  34278=>"111111111",
  34279=>"000010010",
  34280=>"111111110",
  34281=>"000000101",
  34282=>"000001001",
  34283=>"111010111",
  34284=>"000000000",
  34285=>"110000110",
  34286=>"111111111",
  34287=>"110000000",
  34288=>"110000111",
  34289=>"000011111",
  34290=>"111111111",
  34291=>"110011011",
  34292=>"001011111",
  34293=>"000000000",
  34294=>"111011001",
  34295=>"111001111",
  34296=>"100000000",
  34297=>"001000000",
  34298=>"000100111",
  34299=>"110000000",
  34300=>"011111001",
  34301=>"111000011",
  34302=>"100100101",
  34303=>"111111011",
  34304=>"000101110",
  34305=>"111111111",
  34306=>"011000101",
  34307=>"100101100",
  34308=>"001001010",
  34309=>"000001001",
  34310=>"110011000",
  34311=>"000000011",
  34312=>"000000001",
  34313=>"011000000",
  34314=>"000000001",
  34315=>"000010000",
  34316=>"000000000",
  34317=>"000010111",
  34318=>"111010000",
  34319=>"001001000",
  34320=>"111001000",
  34321=>"111010000",
  34322=>"011101111",
  34323=>"111111000",
  34324=>"111111111",
  34325=>"100110000",
  34326=>"100111111",
  34327=>"010110000",
  34328=>"101001101",
  34329=>"111010111",
  34330=>"000000011",
  34331=>"011110111",
  34332=>"111111101",
  34333=>"000100101",
  34334=>"000111111",
  34335=>"000000111",
  34336=>"111000000",
  34337=>"111011111",
  34338=>"010011111",
  34339=>"000000111",
  34340=>"101101000",
  34341=>"001001111",
  34342=>"010110101",
  34343=>"111101001",
  34344=>"110000000",
  34345=>"110000000",
  34346=>"100101111",
  34347=>"010111010",
  34348=>"011101111",
  34349=>"110110011",
  34350=>"000101111",
  34351=>"100000010",
  34352=>"110000000",
  34353=>"001001000",
  34354=>"111010100",
  34355=>"000100000",
  34356=>"000000111",
  34357=>"000001110",
  34358=>"001000100",
  34359=>"111000000",
  34360=>"011000000",
  34361=>"000001101",
  34362=>"000101111",
  34363=>"000010001",
  34364=>"001001001",
  34365=>"010111110",
  34366=>"000001101",
  34367=>"101111110",
  34368=>"111001000",
  34369=>"000000111",
  34370=>"001101000",
  34371=>"010100000",
  34372=>"111000001",
  34373=>"000000000",
  34374=>"000000111",
  34375=>"000000110",
  34376=>"001001111",
  34377=>"101101011",
  34378=>"000001111",
  34379=>"000000000",
  34380=>"010000000",
  34381=>"010011001",
  34382=>"100110000",
  34383=>"010010101",
  34384=>"101110110",
  34385=>"000010111",
  34386=>"010011011",
  34387=>"100100000",
  34388=>"111111101",
  34389=>"101111100",
  34390=>"001110101",
  34391=>"000010011",
  34392=>"010111111",
  34393=>"001101111",
  34394=>"000111111",
  34395=>"110000000",
  34396=>"111000101",
  34397=>"000001111",
  34398=>"111010111",
  34399=>"000000100",
  34400=>"110010000",
  34401=>"010000010",
  34402=>"010000001",
  34403=>"001101111",
  34404=>"101101101",
  34405=>"101000100",
  34406=>"111001000",
  34407=>"101110110",
  34408=>"000000101",
  34409=>"000001111",
  34410=>"111000010",
  34411=>"010000110",
  34412=>"001111100",
  34413=>"110010111",
  34414=>"111001111",
  34415=>"001001100",
  34416=>"100000000",
  34417=>"000000000",
  34418=>"110000000",
  34419=>"000011000",
  34420=>"000000000",
  34421=>"000000111",
  34422=>"000001111",
  34423=>"010011000",
  34424=>"010101101",
  34425=>"100100111",
  34426=>"111000000",
  34427=>"100100010",
  34428=>"111011001",
  34429=>"000001000",
  34430=>"010000000",
  34431=>"000000001",
  34432=>"111000000",
  34433=>"011111111",
  34434=>"011010011",
  34435=>"111101110",
  34436=>"010111001",
  34437=>"111100111",
  34438=>"100100111",
  34439=>"100001001",
  34440=>"101101000",
  34441=>"111010110",
  34442=>"000110001",
  34443=>"000001010",
  34444=>"110110111",
  34445=>"110000000",
  34446=>"011000000",
  34447=>"101000000",
  34448=>"100001001",
  34449=>"110011000",
  34450=>"000000000",
  34451=>"000001001",
  34452=>"110110000",
  34453=>"111000001",
  34454=>"001111111",
  34455=>"001000100",
  34456=>"111010001",
  34457=>"000111101",
  34458=>"000010000",
  34459=>"010000111",
  34460=>"000011111",
  34461=>"111010010",
  34462=>"101000000",
  34463=>"000001111",
  34464=>"100100011",
  34465=>"000000011",
  34466=>"101001111",
  34467=>"011011111",
  34468=>"111111110",
  34469=>"011010000",
  34470=>"011011010",
  34471=>"000001000",
  34472=>"111110000",
  34473=>"110110010",
  34474=>"111101000",
  34475=>"010001001",
  34476=>"000111011",
  34477=>"000001101",
  34478=>"011011001",
  34479=>"111000000",
  34480=>"011111111",
  34481=>"110100111",
  34482=>"000101111",
  34483=>"110110111",
  34484=>"110011000",
  34485=>"000000101",
  34486=>"011000100",
  34487=>"100001001",
  34488=>"100100100",
  34489=>"001000000",
  34490=>"111111010",
  34491=>"000001110",
  34492=>"000110111",
  34493=>"111000001",
  34494=>"001011110",
  34495=>"010000101",
  34496=>"111111000",
  34497=>"111000000",
  34498=>"110111111",
  34499=>"000001001",
  34500=>"000000000",
  34501=>"100100110",
  34502=>"111111101",
  34503=>"000010010",
  34504=>"010000000",
  34505=>"111101101",
  34506=>"101101111",
  34507=>"101000110",
  34508=>"101000000",
  34509=>"111100100",
  34510=>"000000000",
  34511=>"000000000",
  34512=>"010111000",
  34513=>"100101111",
  34514=>"101000110",
  34515=>"101001000",
  34516=>"111001101",
  34517=>"101101101",
  34518=>"000010111",
  34519=>"111011010",
  34520=>"111111000",
  34521=>"011111000",
  34522=>"101101111",
  34523=>"111000000",
  34524=>"111110110",
  34525=>"010010111",
  34526=>"101010000",
  34527=>"000000101",
  34528=>"000000000",
  34529=>"000000101",
  34530=>"110111111",
  34531=>"111001101",
  34532=>"000000000",
  34533=>"010110110",
  34534=>"011000000",
  34535=>"100101101",
  34536=>"000000011",
  34537=>"000011101",
  34538=>"000000100",
  34539=>"101111010",
  34540=>"000000000",
  34541=>"000000101",
  34542=>"000000100",
  34543=>"000000110",
  34544=>"000000010",
  34545=>"001001010",
  34546=>"010001010",
  34547=>"000001110",
  34548=>"001101111",
  34549=>"001111110",
  34550=>"000000000",
  34551=>"001001101",
  34552=>"011000000",
  34553=>"001000010",
  34554=>"000110110",
  34555=>"000000010",
  34556=>"100001111",
  34557=>"010110000",
  34558=>"111001100",
  34559=>"101101110",
  34560=>"010010000",
  34561=>"101101111",
  34562=>"101001011",
  34563=>"000111011",
  34564=>"110111000",
  34565=>"000100000",
  34566=>"111110010",
  34567=>"001010000",
  34568=>"110110000",
  34569=>"000000111",
  34570=>"000000110",
  34571=>"111101000",
  34572=>"001101111",
  34573=>"110110111",
  34574=>"111001011",
  34575=>"101111001",
  34576=>"000010111",
  34577=>"000111111",
  34578=>"000001111",
  34579=>"101011000",
  34580=>"101101111",
  34581=>"101001100",
  34582=>"110111011",
  34583=>"000000000",
  34584=>"101000111",
  34585=>"000000000",
  34586=>"111010101",
  34587=>"010100100",
  34588=>"000010111",
  34589=>"111001001",
  34590=>"100010011",
  34591=>"010011000",
  34592=>"101000000",
  34593=>"110101111",
  34594=>"000001000",
  34595=>"010100000",
  34596=>"100000000",
  34597=>"111011001",
  34598=>"101100110",
  34599=>"000000011",
  34600=>"000001001",
  34601=>"011101000",
  34602=>"000000100",
  34603=>"000101111",
  34604=>"000000000",
  34605=>"000000111",
  34606=>"010001000",
  34607=>"110111111",
  34608=>"010111100",
  34609=>"110100100",
  34610=>"000000000",
  34611=>"011110100",
  34612=>"101001111",
  34613=>"010110111",
  34614=>"011001001",
  34615=>"101111111",
  34616=>"000011111",
  34617=>"000111000",
  34618=>"010010000",
  34619=>"000010000",
  34620=>"100001001",
  34621=>"000111101",
  34622=>"010000011",
  34623=>"100110010",
  34624=>"111001101",
  34625=>"000010001",
  34626=>"111110111",
  34627=>"100111100",
  34628=>"110010000",
  34629=>"111100100",
  34630=>"110111000",
  34631=>"101100000",
  34632=>"001110111",
  34633=>"000010110",
  34634=>"101000101",
  34635=>"001010101",
  34636=>"000000000",
  34637=>"011011000",
  34638=>"111111000",
  34639=>"111110001",
  34640=>"111001000",
  34641=>"110000110",
  34642=>"111011000",
  34643=>"111011110",
  34644=>"100000111",
  34645=>"100110111",
  34646=>"010100000",
  34647=>"101101111",
  34648=>"110000001",
  34649=>"001111110",
  34650=>"011111110",
  34651=>"011111000",
  34652=>"000010010",
  34653=>"010011001",
  34654=>"101000111",
  34655=>"011111111",
  34656=>"100000010",
  34657=>"000000101",
  34658=>"000001111",
  34659=>"100111011",
  34660=>"011011100",
  34661=>"011101000",
  34662=>"000000110",
  34663=>"011111001",
  34664=>"101111000",
  34665=>"000010111",
  34666=>"101110111",
  34667=>"000001000",
  34668=>"010000000",
  34669=>"010000000",
  34670=>"000010110",
  34671=>"000100000",
  34672=>"110000100",
  34673=>"011001000",
  34674=>"110100110",
  34675=>"101011111",
  34676=>"100001111",
  34677=>"000000100",
  34678=>"101100000",
  34679=>"111000000",
  34680=>"000110111",
  34681=>"000010010",
  34682=>"111111111",
  34683=>"000000000",
  34684=>"100010001",
  34685=>"010110101",
  34686=>"111111011",
  34687=>"011000000",
  34688=>"111000000",
  34689=>"111100111",
  34690=>"010000010",
  34691=>"010110000",
  34692=>"100000111",
  34693=>"010000000",
  34694=>"010010010",
  34695=>"100110001",
  34696=>"011011001",
  34697=>"010001001",
  34698=>"010000101",
  34699=>"101001110",
  34700=>"111000110",
  34701=>"001011010",
  34702=>"000000011",
  34703=>"101000000",
  34704=>"100011111",
  34705=>"000111111",
  34706=>"000010111",
  34707=>"001000000",
  34708=>"101000010",
  34709=>"101101111",
  34710=>"001010101",
  34711=>"010100000",
  34712=>"111111111",
  34713=>"110110110",
  34714=>"111010110",
  34715=>"000000101",
  34716=>"000000000",
  34717=>"100101101",
  34718=>"000000000",
  34719=>"000001111",
  34720=>"100010011",
  34721=>"000111010",
  34722=>"011000000",
  34723=>"110111111",
  34724=>"101000000",
  34725=>"010110000",
  34726=>"011100111",
  34727=>"111000100",
  34728=>"000101111",
  34729=>"000000000",
  34730=>"111101011",
  34731=>"111101110",
  34732=>"111101110",
  34733=>"110101011",
  34734=>"011011000",
  34735=>"101011111",
  34736=>"101000111",
  34737=>"000110110",
  34738=>"000010110",
  34739=>"111110110",
  34740=>"101110110",
  34741=>"101010000",
  34742=>"111100000",
  34743=>"010000100",
  34744=>"010010000",
  34745=>"011010110",
  34746=>"010010010",
  34747=>"001001000",
  34748=>"011000100",
  34749=>"111000110",
  34750=>"100011011",
  34751=>"001000011",
  34752=>"010011011",
  34753=>"000000110",
  34754=>"111010000",
  34755=>"011101100",
  34756=>"000000000",
  34757=>"110000001",
  34758=>"000111111",
  34759=>"111000111",
  34760=>"010011100",
  34761=>"101101100",
  34762=>"001101000",
  34763=>"000010011",
  34764=>"110010011",
  34765=>"001110000",
  34766=>"111100000",
  34767=>"000110111",
  34768=>"111000101",
  34769=>"010110011",
  34770=>"101001100",
  34771=>"010011000",
  34772=>"111001010",
  34773=>"011011000",
  34774=>"010000001",
  34775=>"000000000",
  34776=>"000000000",
  34777=>"110111110",
  34778=>"111010110",
  34779=>"101101110",
  34780=>"011111101",
  34781=>"011011000",
  34782=>"101001001",
  34783=>"110101111",
  34784=>"001101111",
  34785=>"000101111",
  34786=>"010001001",
  34787=>"011100100",
  34788=>"011001001",
  34789=>"001101000",
  34790=>"000000000",
  34791=>"100110000",
  34792=>"111111001",
  34793=>"111000111",
  34794=>"000011011",
  34795=>"100100100",
  34796=>"001000111",
  34797=>"111111001",
  34798=>"111100111",
  34799=>"000000000",
  34800=>"111000000",
  34801=>"011000100",
  34802=>"000010111",
  34803=>"010011001",
  34804=>"001001000",
  34805=>"101101101",
  34806=>"111000010",
  34807=>"011111101",
  34808=>"000011000",
  34809=>"101000000",
  34810=>"011011111",
  34811=>"101000001",
  34812=>"010010100",
  34813=>"100101100",
  34814=>"111111000",
  34815=>"111111111",
  34816=>"110110110",
  34817=>"111111111",
  34818=>"101000010",
  34819=>"001101111",
  34820=>"001000000",
  34821=>"001101111",
  34822=>"010000100",
  34823=>"000000110",
  34824=>"001001000",
  34825=>"110000100",
  34826=>"011111011",
  34827=>"011100010",
  34828=>"101101100",
  34829=>"111000000",
  34830=>"111001000",
  34831=>"000000000",
  34832=>"100000101",
  34833=>"111111111",
  34834=>"111001001",
  34835=>"010111111",
  34836=>"001000000",
  34837=>"010000000",
  34838=>"111111111",
  34839=>"111011111",
  34840=>"011110010",
  34841=>"000000000",
  34842=>"000000100",
  34843=>"000000101",
  34844=>"100001111",
  34845=>"010111011",
  34846=>"010111011",
  34847=>"111111000",
  34848=>"000001000",
  34849=>"111111111",
  34850=>"111001111",
  34851=>"111011111",
  34852=>"001001001",
  34853=>"100010001",
  34854=>"010111010",
  34855=>"010100111",
  34856=>"010111111",
  34857=>"000000000",
  34858=>"111111000",
  34859=>"111111001",
  34860=>"110111111",
  34861=>"000010000",
  34862=>"100101111",
  34863=>"100100111",
  34864=>"111100111",
  34865=>"000000000",
  34866=>"111111111",
  34867=>"000111000",
  34868=>"111111111",
  34869=>"111101000",
  34870=>"011111010",
  34871=>"010111100",
  34872=>"000000111",
  34873=>"101101001",
  34874=>"110100000",
  34875=>"000000001",
  34876=>"000000000",
  34877=>"111111111",
  34878=>"111100101",
  34879=>"101101101",
  34880=>"000000000",
  34881=>"010010011",
  34882=>"000000000",
  34883=>"000111011",
  34884=>"111101001",
  34885=>"100000101",
  34886=>"000000100",
  34887=>"000111111",
  34888=>"100000000",
  34889=>"111111111",
  34890=>"100100101",
  34891=>"100000100",
  34892=>"000000000",
  34893=>"100100100",
  34894=>"000000000",
  34895=>"011010101",
  34896=>"110111110",
  34897=>"111111111",
  34898=>"011100000",
  34899=>"100101001",
  34900=>"010111011",
  34901=>"011111111",
  34902=>"100100111",
  34903=>"111111111",
  34904=>"010010111",
  34905=>"000000000",
  34906=>"000001001",
  34907=>"000000000",
  34908=>"101000010",
  34909=>"011011011",
  34910=>"000001000",
  34911=>"011111110",
  34912=>"101000100",
  34913=>"111111011",
  34914=>"000000000",
  34915=>"000110000",
  34916=>"101001000",
  34917=>"101101000",
  34918=>"111101100",
  34919=>"010000000",
  34920=>"000101000",
  34921=>"000101111",
  34922=>"111101101",
  34923=>"000000000",
  34924=>"111000011",
  34925=>"110111000",
  34926=>"000000100",
  34927=>"100001110",
  34928=>"101000000",
  34929=>"000000000",
  34930=>"111111010",
  34931=>"010010000",
  34932=>"111101000",
  34933=>"100000111",
  34934=>"000111000",
  34935=>"010000000",
  34936=>"000000000",
  34937=>"101001101",
  34938=>"111101000",
  34939=>"000000000",
  34940=>"111111101",
  34941=>"000001111",
  34942=>"000010000",
  34943=>"101000110",
  34944=>"000000101",
  34945=>"101100001",
  34946=>"000100101",
  34947=>"000001101",
  34948=>"101001101",
  34949=>"000000000",
  34950=>"000000010",
  34951=>"100001000",
  34952=>"111100100",
  34953=>"110000010",
  34954=>"001010000",
  34955=>"000000101",
  34956=>"111011000",
  34957=>"000100101",
  34958=>"000000000",
  34959=>"101000000",
  34960=>"000101001",
  34961=>"010010110",
  34962=>"000000000",
  34963=>"110010100",
  34964=>"101011000",
  34965=>"001000100",
  34966=>"011111110",
  34967=>"111100000",
  34968=>"000110101",
  34969=>"010011011",
  34970=>"101000000",
  34971=>"100101100",
  34972=>"101101101",
  34973=>"000000000",
  34974=>"000000111",
  34975=>"101101101",
  34976=>"000001001",
  34977=>"110111011",
  34978=>"011010011",
  34979=>"001000111",
  34980=>"000110001",
  34981=>"000100000",
  34982=>"000000000",
  34983=>"111111000",
  34984=>"110010110",
  34985=>"011111111",
  34986=>"100000101",
  34987=>"100000101",
  34988=>"101111111",
  34989=>"001000100",
  34990=>"011011111",
  34991=>"001010000",
  34992=>"000000110",
  34993=>"011111011",
  34994=>"111101101",
  34995=>"111000000",
  34996=>"011011001",
  34997=>"011000001",
  34998=>"101000101",
  34999=>"001001001",
  35000=>"000000000",
  35001=>"101011000",
  35002=>"000000111",
  35003=>"111111111",
  35004=>"100110111",
  35005=>"111001001",
  35006=>"110100101",
  35007=>"111011111",
  35008=>"000111010",
  35009=>"010000011",
  35010=>"101111100",
  35011=>"000000001",
  35012=>"000000101",
  35013=>"010110111",
  35014=>"000000101",
  35015=>"110011010",
  35016=>"011111101",
  35017=>"001111011",
  35018=>"111111000",
  35019=>"111000000",
  35020=>"000000000",
  35021=>"111111001",
  35022=>"100000101",
  35023=>"000101001",
  35024=>"101111000",
  35025=>"011111101",
  35026=>"110000000",
  35027=>"000000100",
  35028=>"101100100",
  35029=>"111111111",
  35030=>"010010000",
  35031=>"101001101",
  35032=>"000010000",
  35033=>"111101000",
  35034=>"001001101",
  35035=>"000100100",
  35036=>"011111111",
  35037=>"011011011",
  35038=>"000000000",
  35039=>"000001000",
  35040=>"111100100",
  35041=>"100100101",
  35042=>"000010111",
  35043=>"011011000",
  35044=>"000000010",
  35045=>"111111111",
  35046=>"001000000",
  35047=>"101011010",
  35048=>"111101001",
  35049=>"000111111",
  35050=>"110111111",
  35051=>"000000000",
  35052=>"000000000",
  35053=>"000000101",
  35054=>"100000001",
  35055=>"000000101",
  35056=>"001001101",
  35057=>"111011111",
  35058=>"100000000",
  35059=>"010111100",
  35060=>"001011000",
  35061=>"010111111",
  35062=>"000100000",
  35063=>"001101011",
  35064=>"101100000",
  35065=>"111111001",
  35066=>"110011011",
  35067=>"000111101",
  35068=>"111000000",
  35069=>"000101000",
  35070=>"100000000",
  35071=>"000000000",
  35072=>"110111001",
  35073=>"000000001",
  35074=>"101110111",
  35075=>"000000011",
  35076=>"000000100",
  35077=>"000110110",
  35078=>"000111110",
  35079=>"111101010",
  35080=>"000100001",
  35081=>"110110000",
  35082=>"011111110",
  35083=>"000110111",
  35084=>"001001001",
  35085=>"111111000",
  35086=>"000111111",
  35087=>"110000111",
  35088=>"110000110",
  35089=>"000010111",
  35090=>"000001000",
  35091=>"111000010",
  35092=>"000000100",
  35093=>"111001001",
  35094=>"101001000",
  35095=>"110000111",
  35096=>"111000001",
  35097=>"111111111",
  35098=>"000001100",
  35099=>"110110000",
  35100=>"111111001",
  35101=>"111000001",
  35102=>"111110110",
  35103=>"001001001",
  35104=>"000110110",
  35105=>"100000101",
  35106=>"110100000",
  35107=>"000111111",
  35108=>"100101101",
  35109=>"100110000",
  35110=>"001000001",
  35111=>"000100110",
  35112=>"000100110",
  35113=>"111000001",
  35114=>"000001000",
  35115=>"001100000",
  35116=>"000011111",
  35117=>"111011100",
  35118=>"111111100",
  35119=>"000000001",
  35120=>"111111000",
  35121=>"000011011",
  35122=>"111000001",
  35123=>"111111111",
  35124=>"000110000",
  35125=>"001001001",
  35126=>"001001011",
  35127=>"001001001",
  35128=>"011001110",
  35129=>"001101000",
  35130=>"001001000",
  35131=>"011001001",
  35132=>"001001000",
  35133=>"000001000",
  35134=>"000110010",
  35135=>"001111011",
  35136=>"110000000",
  35137=>"111110000",
  35138=>"000100111",
  35139=>"010011000",
  35140=>"111001000",
  35141=>"111110110",
  35142=>"111111011",
  35143=>"110010001",
  35144=>"111001000",
  35145=>"110111000",
  35146=>"000110011",
  35147=>"111010001",
  35148=>"000111110",
  35149=>"011011011",
  35150=>"100011101",
  35151=>"111111111",
  35152=>"000000010",
  35153=>"110010010",
  35154=>"111110000",
  35155=>"011111100",
  35156=>"001000001",
  35157=>"011000001",
  35158=>"111111101",
  35159=>"110110110",
  35160=>"110000001",
  35161=>"000001011",
  35162=>"000001001",
  35163=>"011001111",
  35164=>"000000000",
  35165=>"110110000",
  35166=>"111001001",
  35167=>"000110110",
  35168=>"000000100",
  35169=>"000111111",
  35170=>"100110110",
  35171=>"000000001",
  35172=>"000100100",
  35173=>"010001001",
  35174=>"000110000",
  35175=>"110110000",
  35176=>"110110000",
  35177=>"111000011",
  35178=>"001000110",
  35179=>"110100111",
  35180=>"111011001",
  35181=>"000111110",
  35182=>"110111000",
  35183=>"110110101",
  35184=>"000111001",
  35185=>"111011011",
  35186=>"011000000",
  35187=>"001000000",
  35188=>"111111000",
  35189=>"100000000",
  35190=>"000101110",
  35191=>"101000001",
  35192=>"011011001",
  35193=>"111000000",
  35194=>"111101101",
  35195=>"110011001",
  35196=>"110100100",
  35197=>"010110011",
  35198=>"000000000",
  35199=>"000110010",
  35200=>"000100010",
  35201=>"110000000",
  35202=>"110001000",
  35203=>"110110110",
  35204=>"011100000",
  35205=>"111110111",
  35206=>"111011000",
  35207=>"000000011",
  35208=>"010111011",
  35209=>"111111000",
  35210=>"001110101",
  35211=>"010000101",
  35212=>"000001011",
  35213=>"000000010",
  35214=>"111001011",
  35215=>"101000000",
  35216=>"110001011",
  35217=>"110100000",
  35218=>"110110010",
  35219=>"101000100",
  35220=>"010110111",
  35221=>"110100110",
  35222=>"000100110",
  35223=>"110100100",
  35224=>"110110111",
  35225=>"111111110",
  35226=>"111010010",
  35227=>"000000001",
  35228=>"110011110",
  35229=>"000111101",
  35230=>"100100111",
  35231=>"000110110",
  35232=>"100101111",
  35233=>"001001001",
  35234=>"010001111",
  35235=>"101000001",
  35236=>"111111000",
  35237=>"000011011",
  35238=>"001010111",
  35239=>"101001001",
  35240=>"111001000",
  35241=>"111001110",
  35242=>"011001010",
  35243=>"110110000",
  35244=>"100000111",
  35245=>"111101100",
  35246=>"001010011",
  35247=>"001011111",
  35248=>"100001111",
  35249=>"010011000",
  35250=>"000110010",
  35251=>"000000110",
  35252=>"100110110",
  35253=>"100000010",
  35254=>"011100001",
  35255=>"101011111",
  35256=>"010110000",
  35257=>"010100100",
  35258=>"110111000",
  35259=>"000110110",
  35260=>"000110100",
  35261=>"110011110",
  35262=>"110110001",
  35263=>"110001000",
  35264=>"000111111",
  35265=>"011011000",
  35266=>"100000111",
  35267=>"000111000",
  35268=>"110010001",
  35269=>"100101011",
  35270=>"110111011",
  35271=>"000010000",
  35272=>"110000110",
  35273=>"110001001",
  35274=>"000001001",
  35275=>"111111001",
  35276=>"000010000",
  35277=>"001011010",
  35278=>"010110011",
  35279=>"000001011",
  35280=>"000110110",
  35281=>"011111011",
  35282=>"000101111",
  35283=>"110111000",
  35284=>"100001001",
  35285=>"001011001",
  35286=>"000010000",
  35287=>"111010000",
  35288=>"011001111",
  35289=>"001001001",
  35290=>"110110011",
  35291=>"110110110",
  35292=>"001001001",
  35293=>"100000011",
  35294=>"111001111",
  35295=>"110110011",
  35296=>"000000000",
  35297=>"000000000",
  35298=>"010001111",
  35299=>"111100100",
  35300=>"001000000",
  35301=>"000001000",
  35302=>"011110100",
  35303=>"111011001",
  35304=>"100000110",
  35305=>"001111110",
  35306=>"100111110",
  35307=>"111111010",
  35308=>"110001001",
  35309=>"001001001",
  35310=>"000000000",
  35311=>"000000010",
  35312=>"111001001",
  35313=>"010001100",
  35314=>"000000110",
  35315=>"111111011",
  35316=>"100100111",
  35317=>"011011011",
  35318=>"000001110",
  35319=>"111101101",
  35320=>"111000000",
  35321=>"000000111",
  35322=>"111101111",
  35323=>"000010111",
  35324=>"010010000",
  35325=>"111001000",
  35326=>"000111101",
  35327=>"111001001",
  35328=>"111011000",
  35329=>"010001000",
  35330=>"110000111",
  35331=>"101001000",
  35332=>"011100001",
  35333=>"101101100",
  35334=>"111101011",
  35335=>"000000100",
  35336=>"100000000",
  35337=>"000000000",
  35338=>"001000111",
  35339=>"000000000",
  35340=>"000001111",
  35341=>"110101111",
  35342=>"111101101",
  35343=>"000010001",
  35344=>"100100000",
  35345=>"100000001",
  35346=>"100110111",
  35347=>"010000000",
  35348=>"001110000",
  35349=>"111101101",
  35350=>"011111011",
  35351=>"111000110",
  35352=>"101100010",
  35353=>"111111111",
  35354=>"000001001",
  35355=>"010111111",
  35356=>"111111000",
  35357=>"111001000",
  35358=>"110000000",
  35359=>"000111100",
  35360=>"111111000",
  35361=>"000000010",
  35362=>"001101111",
  35363=>"000101100",
  35364=>"000000000",
  35365=>"111110000",
  35366=>"111011000",
  35367=>"000011111",
  35368=>"010010000",
  35369=>"001101100",
  35370=>"101000111",
  35371=>"011101111",
  35372=>"110011110",
  35373=>"001010010",
  35374=>"011011010",
  35375=>"001101011",
  35376=>"000010011",
  35377=>"000000001",
  35378=>"000101011",
  35379=>"010000101",
  35380=>"111000000",
  35381=>"111111111",
  35382=>"110000010",
  35383=>"000111000",
  35384=>"111100101",
  35385=>"000000111",
  35386=>"111000101",
  35387=>"111010110",
  35388=>"110110110",
  35389=>"111111111",
  35390=>"000100000",
  35391=>"110111110",
  35392=>"011000111",
  35393=>"111111000",
  35394=>"000000000",
  35395=>"111101011",
  35396=>"111000110",
  35397=>"101101001",
  35398=>"000011101",
  35399=>"100000001",
  35400=>"110001001",
  35401=>"101111010",
  35402=>"101101110",
  35403=>"011101000",
  35404=>"011111000",
  35405=>"100000100",
  35406=>"010000000",
  35407=>"110010010",
  35408=>"010001000",
  35409=>"110111111",
  35410=>"100000101",
  35411=>"011101001",
  35412=>"011111011",
  35413=>"010111001",
  35414=>"000100000",
  35415=>"111001001",
  35416=>"001001000",
  35417=>"001000000",
  35418=>"100100000",
  35419=>"001100000",
  35420=>"000000101",
  35421=>"010001111",
  35422=>"010010011",
  35423=>"111110001",
  35424=>"001000000",
  35425=>"001111010",
  35426=>"101001111",
  35427=>"011100000",
  35428=>"100000001",
  35429=>"011111011",
  35430=>"010010000",
  35431=>"000111001",
  35432=>"101111011",
  35433=>"111000000",
  35434=>"000100000",
  35435=>"010010011",
  35436=>"000000111",
  35437=>"101000101",
  35438=>"101101011",
  35439=>"110110010",
  35440=>"100000000",
  35441=>"010011001",
  35442=>"011000110",
  35443=>"101101101",
  35444=>"000000000",
  35445=>"000000111",
  35446=>"111001101",
  35447=>"000101101",
  35448=>"010111000",
  35449=>"000111010",
  35450=>"111110011",
  35451=>"101000111",
  35452=>"100110111",
  35453=>"111100000",
  35454=>"111111111",
  35455=>"111101100",
  35456=>"000000000",
  35457=>"000100000",
  35458=>"011010001",
  35459=>"100011111",
  35460=>"101001001",
  35461=>"000111110",
  35462=>"111111000",
  35463=>"000011110",
  35464=>"001001001",
  35465=>"111111000",
  35466=>"101000111",
  35467=>"000100111",
  35468=>"001011000",
  35469=>"101111110",
  35470=>"010010001",
  35471=>"101001100",
  35472=>"111111110",
  35473=>"011101000",
  35474=>"000110000",
  35475=>"001011010",
  35476=>"000111111",
  35477=>"000000000",
  35478=>"010010010",
  35479=>"110000101",
  35480=>"000000000",
  35481=>"110111010",
  35482=>"000010010",
  35483=>"000000100",
  35484=>"000100000",
  35485=>"101001000",
  35486=>"000000000",
  35487=>"011000111",
  35488=>"000100000",
  35489=>"010111001",
  35490=>"111100000",
  35491=>"010000000",
  35492=>"100100101",
  35493=>"000100000",
  35494=>"100001000",
  35495=>"000011000",
  35496=>"000000010",
  35497=>"001000000",
  35498=>"000101111",
  35499=>"000000001",
  35500=>"010110111",
  35501=>"000000001",
  35502=>"111000000",
  35503=>"101001101",
  35504=>"000101001",
  35505=>"110000100",
  35506=>"000000100",
  35507=>"111001001",
  35508=>"011111011",
  35509=>"101111000",
  35510=>"001001100",
  35511=>"010010000",
  35512=>"001011000",
  35513=>"000110111",
  35514=>"110111000",
  35515=>"010010011",
  35516=>"111011000",
  35517=>"111011111",
  35518=>"111110110",
  35519=>"101111011",
  35520=>"111011011",
  35521=>"000001000",
  35522=>"111111000",
  35523=>"110001000",
  35524=>"111111000",
  35525=>"000000010",
  35526=>"000000101",
  35527=>"000101111",
  35528=>"111000000",
  35529=>"111111111",
  35530=>"111101000",
  35531=>"001100101",
  35532=>"011011000",
  35533=>"001011111",
  35534=>"000001010",
  35535=>"010110101",
  35536=>"111010111",
  35537=>"110000101",
  35538=>"000010010",
  35539=>"010010010",
  35540=>"000110111",
  35541=>"111011000",
  35542=>"101000111",
  35543=>"111010000",
  35544=>"010000000",
  35545=>"101000101",
  35546=>"000001011",
  35547=>"101000100",
  35548=>"010111100",
  35549=>"101000001",
  35550=>"000101000",
  35551=>"110010000",
  35552=>"010111100",
  35553=>"100100001",
  35554=>"110100110",
  35555=>"111001001",
  35556=>"000010000",
  35557=>"111011000",
  35558=>"101100000",
  35559=>"000000101",
  35560=>"001001000",
  35561=>"111111010",
  35562=>"100000000",
  35563=>"111000011",
  35564=>"111000000",
  35565=>"000000000",
  35566=>"000001000",
  35567=>"100001001",
  35568=>"000001111",
  35569=>"100001100",
  35570=>"000000010",
  35571=>"110100100",
  35572=>"110101011",
  35573=>"101001100",
  35574=>"000000000",
  35575=>"000101010",
  35576=>"000111111",
  35577=>"001101110",
  35578=>"111100100",
  35579=>"101111110",
  35580=>"000001110",
  35581=>"001111000",
  35582=>"100000010",
  35583=>"111000000",
  35584=>"101000000",
  35585=>"000000001",
  35586=>"000000100",
  35587=>"010000000",
  35588=>"000000010",
  35589=>"010000000",
  35590=>"010010010",
  35591=>"010011111",
  35592=>"111000000",
  35593=>"111101100",
  35594=>"000001001",
  35595=>"011001101",
  35596=>"101000000",
  35597=>"000111000",
  35598=>"000011010",
  35599=>"000100000",
  35600=>"000100000",
  35601=>"111111111",
  35602=>"111010101",
  35603=>"000111111",
  35604=>"000001100",
  35605=>"111111111",
  35606=>"000000001",
  35607=>"010111111",
  35608=>"111111000",
  35609=>"101000001",
  35610=>"111000000",
  35611=>"000000000",
  35612=>"111000111",
  35613=>"111111011",
  35614=>"110111001",
  35615=>"111111101",
  35616=>"000000111",
  35617=>"000101111",
  35618=>"110111111",
  35619=>"001100000",
  35620=>"111101100",
  35621=>"100111000",
  35622=>"111000000",
  35623=>"000001000",
  35624=>"011111111",
  35625=>"101100000",
  35626=>"010000010",
  35627=>"111110000",
  35628=>"110110110",
  35629=>"100101001",
  35630=>"111111111",
  35631=>"000101101",
  35632=>"000000000",
  35633=>"000100000",
  35634=>"000101111",
  35635=>"010111111",
  35636=>"101000000",
  35637=>"011100111",
  35638=>"001011000",
  35639=>"000000000",
  35640=>"100000101",
  35641=>"010111111",
  35642=>"000110111",
  35643=>"000000000",
  35644=>"011111110",
  35645=>"111000101",
  35646=>"001100000",
  35647=>"111001001",
  35648=>"111111111",
  35649=>"010000000",
  35650=>"000100000",
  35651=>"111101101",
  35652=>"101011111",
  35653=>"101111000",
  35654=>"111111000",
  35655=>"000000111",
  35656=>"000000001",
  35657=>"100000001",
  35658=>"000000100",
  35659=>"111100100",
  35660=>"110111111",
  35661=>"011001111",
  35662=>"000000101",
  35663=>"111100000",
  35664=>"000000101",
  35665=>"111111111",
  35666=>"111011111",
  35667=>"110100100",
  35668=>"001000001",
  35669=>"100111001",
  35670=>"000100000",
  35671=>"100111111",
  35672=>"000001001",
  35673=>"000111001",
  35674=>"001011011",
  35675=>"000011111",
  35676=>"000000000",
  35677=>"010011110",
  35678=>"100000000",
  35679=>"100001101",
  35680=>"111000000",
  35681=>"001101100",
  35682=>"101000000",
  35683=>"000010111",
  35684=>"111101001",
  35685=>"000001111",
  35686=>"100001101",
  35687=>"111110111",
  35688=>"111111111",
  35689=>"000000111",
  35690=>"000110111",
  35691=>"000000011",
  35692=>"000111111",
  35693=>"010010010",
  35694=>"000000100",
  35695=>"000000110",
  35696=>"001001000",
  35697=>"000000000",
  35698=>"000111001",
  35699=>"000111010",
  35700=>"100111011",
  35701=>"111000011",
  35702=>"110111110",
  35703=>"111111111",
  35704=>"001001100",
  35705=>"000000000",
  35706=>"000000001",
  35707=>"000101111",
  35708=>"001001000",
  35709=>"110011001",
  35710=>"111001100",
  35711=>"101000000",
  35712=>"000000101",
  35713=>"011010000",
  35714=>"000110111",
  35715=>"000110010",
  35716=>"011111111",
  35717=>"000111111",
  35718=>"101110000",
  35719=>"101101001",
  35720=>"100010010",
  35721=>"000100000",
  35722=>"000000000",
  35723=>"000000111",
  35724=>"000000111",
  35725=>"111101100",
  35726=>"110011000",
  35727=>"111000001",
  35728=>"010100110",
  35729=>"010001000",
  35730=>"000000000",
  35731=>"000000000",
  35732=>"111011001",
  35733=>"101101101",
  35734=>"101111000",
  35735=>"111111000",
  35736=>"111000001",
  35737=>"001111111",
  35738=>"000111101",
  35739=>"101000000",
  35740=>"010111000",
  35741=>"110111111",
  35742=>"010111110",
  35743=>"010010010",
  35744=>"011101101",
  35745=>"111111111",
  35746=>"000000011",
  35747=>"000000011",
  35748=>"100111111",
  35749=>"000111110",
  35750=>"110100010",
  35751=>"000100111",
  35752=>"110100000",
  35753=>"111001100",
  35754=>"000000111",
  35755=>"000000000",
  35756=>"111110110",
  35757=>"101000000",
  35758=>"000000001",
  35759=>"001000000",
  35760=>"000000101",
  35761=>"000110110",
  35762=>"000011010",
  35763=>"000000101",
  35764=>"110000000",
  35765=>"100110101",
  35766=>"010000111",
  35767=>"110111111",
  35768=>"111111001",
  35769=>"111110111",
  35770=>"110010101",
  35771=>"010101100",
  35772=>"010000011",
  35773=>"010010111",
  35774=>"110111110",
  35775=>"000000001",
  35776=>"000000111",
  35777=>"111000100",
  35778=>"011111000",
  35779=>"111001000",
  35780=>"000000010",
  35781=>"011101001",
  35782=>"110111111",
  35783=>"111111010",
  35784=>"010010010",
  35785=>"000000000",
  35786=>"110111101",
  35787=>"000000000",
  35788=>"110111000",
  35789=>"100000100",
  35790=>"001011000",
  35791=>"100011100",
  35792=>"111010111",
  35793=>"011001000",
  35794=>"000000000",
  35795=>"000100000",
  35796=>"101000111",
  35797=>"000011011",
  35798=>"110111010",
  35799=>"110110111",
  35800=>"000000001",
  35801=>"000000101",
  35802=>"100011011",
  35803=>"000110010",
  35804=>"001110000",
  35805=>"101100100",
  35806=>"111010111",
  35807=>"111101111",
  35808=>"111000000",
  35809=>"111101000",
  35810=>"010011000",
  35811=>"001011010",
  35812=>"100000000",
  35813=>"000000101",
  35814=>"111000111",
  35815=>"000000100",
  35816=>"101100101",
  35817=>"000000000",
  35818=>"001000000",
  35819=>"000111111",
  35820=>"100100001",
  35821=>"011000111",
  35822=>"111101111",
  35823=>"111000101",
  35824=>"011000100",
  35825=>"011110000",
  35826=>"011000000",
  35827=>"011011001",
  35828=>"000101101",
  35829=>"000000001",
  35830=>"110000100",
  35831=>"100110000",
  35832=>"111111111",
  35833=>"001111111",
  35834=>"111100100",
  35835=>"111001000",
  35836=>"010010100",
  35837=>"000000000",
  35838=>"010110111",
  35839=>"010111000",
  35840=>"011111110",
  35841=>"010000000",
  35842=>"001000101",
  35843=>"000000000",
  35844=>"001111011",
  35845=>"000000000",
  35846=>"011111010",
  35847=>"000000000",
  35848=>"000000100",
  35849=>"010000000",
  35850=>"000011000",
  35851=>"111001101",
  35852=>"000000000",
  35853=>"000000101",
  35854=>"000001000",
  35855=>"000000101",
  35856=>"100100100",
  35857=>"111010010",
  35858=>"110110111",
  35859=>"111000000",
  35860=>"111111111",
  35861=>"111111000",
  35862=>"011101111",
  35863=>"011000011",
  35864=>"000000011",
  35865=>"111101101",
  35866=>"000000000",
  35867=>"010011000",
  35868=>"000100100",
  35869=>"111000000",
  35870=>"110111111",
  35871=>"000000000",
  35872=>"000011111",
  35873=>"101001000",
  35874=>"000011111",
  35875=>"011111010",
  35876=>"011000000",
  35877=>"011100000",
  35878=>"111001000",
  35879=>"101111111",
  35880=>"111100000",
  35881=>"001111111",
  35882=>"010110000",
  35883=>"000010110",
  35884=>"000011010",
  35885=>"100000000",
  35886=>"111000111",
  35887=>"000000000",
  35888=>"000000010",
  35889=>"011111001",
  35890=>"000000000",
  35891=>"100000001",
  35892=>"010011010",
  35893=>"000000000",
  35894=>"001011011",
  35895=>"000001000",
  35896=>"000000000",
  35897=>"000000001",
  35898=>"000000000",
  35899=>"000000000",
  35900=>"000000000",
  35901=>"101100111",
  35902=>"100000100",
  35903=>"010011000",
  35904=>"111111111",
  35905=>"011011011",
  35906=>"010111110",
  35907=>"110110100",
  35908=>"011011000",
  35909=>"000000111",
  35910=>"000011011",
  35911=>"111111000",
  35912=>"000000000",
  35913=>"100110000",
  35914=>"111111001",
  35915=>"111001000",
  35916=>"111110111",
  35917=>"110111111",
  35918=>"011111111",
  35919=>"111101111",
  35920=>"010001000",
  35921=>"111011101",
  35922=>"000000000",
  35923=>"001100000",
  35924=>"010011000",
  35925=>"110111111",
  35926=>"000000000",
  35927=>"111100001",
  35928=>"000010000",
  35929=>"000010000",
  35930=>"000100000",
  35931=>"110000000",
  35932=>"110000000",
  35933=>"000000000",
  35934=>"111111111",
  35935=>"000011011",
  35936=>"000010000",
  35937=>"000000000",
  35938=>"000010111",
  35939=>"000001000",
  35940=>"100101100",
  35941=>"100000100",
  35942=>"000000110",
  35943=>"000000000",
  35944=>"001111000",
  35945=>"000100111",
  35946=>"111001000",
  35947=>"111111101",
  35948=>"000000000",
  35949=>"000100000",
  35950=>"000000000",
  35951=>"000000010",
  35952=>"000011011",
  35953=>"000000010",
  35954=>"000110110",
  35955=>"101110110",
  35956=>"101111111",
  35957=>"101000000",
  35958=>"011111011",
  35959=>"100101111",
  35960=>"000000000",
  35961=>"010111111",
  35962=>"100000000",
  35963=>"000100000",
  35964=>"000100111",
  35965=>"100100000",
  35966=>"111111110",
  35967=>"100000100",
  35968=>"001111101",
  35969=>"100000000",
  35970=>"010001010",
  35971=>"101111111",
  35972=>"110000000",
  35973=>"000000110",
  35974=>"110000010",
  35975=>"010100000",
  35976=>"010111100",
  35977=>"100000000",
  35978=>"100000111",
  35979=>"111111101",
  35980=>"000000000",
  35981=>"010000000",
  35982=>"110111011",
  35983=>"000000000",
  35984=>"001001000",
  35985=>"110111010",
  35986=>"000001111",
  35987=>"111101000",
  35988=>"111001000",
  35989=>"000000111",
  35990=>"111001111",
  35991=>"001011111",
  35992=>"000001000",
  35993=>"111111111",
  35994=>"101100000",
  35995=>"000000000",
  35996=>"001010111",
  35997=>"010000011",
  35998=>"000011010",
  35999=>"100000010",
  36000=>"001111001",
  36001=>"110011111",
  36002=>"000101000",
  36003=>"000111101",
  36004=>"000111110",
  36005=>"000000000",
  36006=>"110111111",
  36007=>"110111000",
  36008=>"110110111",
  36009=>"000000001",
  36010=>"000000000",
  36011=>"011011010",
  36012=>"101100111",
  36013=>"111111111",
  36014=>"000011011",
  36015=>"111101111",
  36016=>"110100101",
  36017=>"000001000",
  36018=>"000000001",
  36019=>"000000110",
  36020=>"100100000",
  36021=>"000011011",
  36022=>"100010111",
  36023=>"101001011",
  36024=>"010000000",
  36025=>"010100000",
  36026=>"110001000",
  36027=>"010010000",
  36028=>"111101001",
  36029=>"111111111",
  36030=>"000110101",
  36031=>"000000000",
  36032=>"000000000",
  36033=>"000010000",
  36034=>"001000000",
  36035=>"011011000",
  36036=>"111001111",
  36037=>"111000000",
  36038=>"000001111",
  36039=>"001000001",
  36040=>"001000111",
  36041=>"000111011",
  36042=>"111111111",
  36043=>"000000000",
  36044=>"111000000",
  36045=>"010011111",
  36046=>"000011010",
  36047=>"000011111",
  36048=>"100101111",
  36049=>"110111111",
  36050=>"111000001",
  36051=>"000000011",
  36052=>"101111100",
  36053=>"100111000",
  36054=>"000000001",
  36055=>"000000000",
  36056=>"000000000",
  36057=>"111000000",
  36058=>"110111110",
  36059=>"010100100",
  36060=>"100111110",
  36061=>"011000100",
  36062=>"010000111",
  36063=>"000000001",
  36064=>"010111000",
  36065=>"100000000",
  36066=>"111111111",
  36067=>"011101000",
  36068=>"101001000",
  36069=>"000111000",
  36070=>"000011111",
  36071=>"100110110",
  36072=>"111100000",
  36073=>"000010110",
  36074=>"100110010",
  36075=>"001111011",
  36076=>"000000000",
  36077=>"000011111",
  36078=>"000010010",
  36079=>"100000000",
  36080=>"100000000",
  36081=>"011111000",
  36082=>"101100100",
  36083=>"100001000",
  36084=>"001111011",
  36085=>"000001000",
  36086=>"000000000",
  36087=>"111101101",
  36088=>"000111000",
  36089=>"110000000",
  36090=>"111111111",
  36091=>"000000000",
  36092=>"010010000",
  36093=>"000001000",
  36094=>"011010000",
  36095=>"000001011",
  36096=>"000000110",
  36097=>"000110110",
  36098=>"001011101",
  36099=>"100111110",
  36100=>"111110100",
  36101=>"111011001",
  36102=>"101000000",
  36103=>"110000001",
  36104=>"100101111",
  36105=>"011011000",
  36106=>"010011111",
  36107=>"010011110",
  36108=>"100100100",
  36109=>"001011000",
  36110=>"011000000",
  36111=>"100000101",
  36112=>"011000000",
  36113=>"001011001",
  36114=>"101101010",
  36115=>"010010011",
  36116=>"000100011",
  36117=>"100110110",
  36118=>"000100100",
  36119=>"011011011",
  36120=>"001010010",
  36121=>"010000011",
  36122=>"100110111",
  36123=>"001011111",
  36124=>"011011011",
  36125=>"011011000",
  36126=>"101001111",
  36127=>"100000100",
  36128=>"000011001",
  36129=>"111110111",
  36130=>"000000011",
  36131=>"101011001",
  36132=>"110110110",
  36133=>"111100111",
  36134=>"010011000",
  36135=>"111111100",
  36136=>"011100110",
  36137=>"100000001",
  36138=>"100100000",
  36139=>"011000011",
  36140=>"000100110",
  36141=>"110110110",
  36142=>"100000100",
  36143=>"001100100",
  36144=>"111000100",
  36145=>"000010000",
  36146=>"101100111",
  36147=>"011000011",
  36148=>"001011111",
  36149=>"111110010",
  36150=>"011001000",
  36151=>"100000100",
  36152=>"100110111",
  36153=>"110000100",
  36154=>"001001000",
  36155=>"001001111",
  36156=>"000000100",
  36157=>"001001000",
  36158=>"000000100",
  36159=>"100111011",
  36160=>"011010110",
  36161=>"111010011",
  36162=>"111011001",
  36163=>"001011111",
  36164=>"110100110",
  36165=>"111011000",
  36166=>"101110010",
  36167=>"011101000",
  36168=>"100100111",
  36169=>"110101100",
  36170=>"000010000",
  36171=>"110100110",
  36172=>"001011001",
  36173=>"010100110",
  36174=>"000100100",
  36175=>"111100110",
  36176=>"001011000",
  36177=>"101101111",
  36178=>"101100110",
  36179=>"010010110",
  36180=>"101000001",
  36181=>"111100100",
  36182=>"000000000",
  36183=>"001011000",
  36184=>"100100100",
  36185=>"100100001",
  36186=>"100101101",
  36187=>"110110110",
  36188=>"100101100",
  36189=>"000010000",
  36190=>"110100111",
  36191=>"111001000",
  36192=>"100110011",
  36193=>"010100100",
  36194=>"000001101",
  36195=>"110110110",
  36196=>"011101111",
  36197=>"110100111",
  36198=>"100110100",
  36199=>"011001000",
  36200=>"100000101",
  36201=>"111101100",
  36202=>"110011011",
  36203=>"110010110",
  36204=>"110110110",
  36205=>"011011011",
  36206=>"100100100",
  36207=>"100100111",
  36208=>"110100000",
  36209=>"100110110",
  36210=>"001011111",
  36211=>"000000000",
  36212=>"111111011",
  36213=>"000001001",
  36214=>"110110001",
  36215=>"100011011",
  36216=>"010011010",
  36217=>"110000011",
  36218=>"010100110",
  36219=>"000100001",
  36220=>"110110100",
  36221=>"101001000",
  36222=>"001001000",
  36223=>"011011000",
  36224=>"110010001",
  36225=>"010010011",
  36226=>"011011110",
  36227=>"100101101",
  36228=>"000000011",
  36229=>"110010110",
  36230=>"000000000",
  36231=>"010000000",
  36232=>"101000100",
  36233=>"101100010",
  36234=>"000000000",
  36235=>"110011011",
  36236=>"110010000",
  36237=>"011001011",
  36238=>"110100111",
  36239=>"000100101",
  36240=>"000100000",
  36241=>"000000111",
  36242=>"011011001",
  36243=>"110010010",
  36244=>"010100110",
  36245=>"001001001",
  36246=>"000100100",
  36247=>"010010000",
  36248=>"111111110",
  36249=>"100000011",
  36250=>"011011001",
  36251=>"011011100",
  36252=>"110100100",
  36253=>"011111111",
  36254=>"111011110",
  36255=>"000001000",
  36256=>"110100010",
  36257=>"011000011",
  36258=>"000100000",
  36259=>"010110010",
  36260=>"011111100",
  36261=>"100000011",
  36262=>"101111111",
  36263=>"000000000",
  36264=>"001011011",
  36265=>"000100111",
  36266=>"011011111",
  36267=>"001011011",
  36268=>"101100011",
  36269=>"000000101",
  36270=>"110110100",
  36271=>"100100000",
  36272=>"110110000",
  36273=>"100110000",
  36274=>"111011111",
  36275=>"001111111",
  36276=>"111111101",
  36277=>"110011111",
  36278=>"111100000",
  36279=>"100100011",
  36280=>"100101110",
  36281=>"110110111",
  36282=>"100110000",
  36283=>"110011011",
  36284=>"110111011",
  36285=>"111011010",
  36286=>"010011001",
  36287=>"000000000",
  36288=>"100100110",
  36289=>"011011010",
  36290=>"111011011",
  36291=>"001100100",
  36292=>"100100100",
  36293=>"100000100",
  36294=>"111010110",
  36295=>"111000101",
  36296=>"000111001",
  36297=>"111110010",
  36298=>"111010000",
  36299=>"100110111",
  36300=>"110011001",
  36301=>"001001101",
  36302=>"011011011",
  36303=>"000011011",
  36304=>"001001000",
  36305=>"000000100",
  36306=>"111100110",
  36307=>"111110110",
  36308=>"100110111",
  36309=>"011101100",
  36310=>"100100100",
  36311=>"100011111",
  36312=>"100100110",
  36313=>"000100010",
  36314=>"011111111",
  36315=>"011011001",
  36316=>"100000110",
  36317=>"000110111",
  36318=>"110110010",
  36319=>"100000100",
  36320=>"100100110",
  36321=>"000000111",
  36322=>"000001001",
  36323=>"100110111",
  36324=>"000000011",
  36325=>"111100000",
  36326=>"110000100",
  36327=>"000000110",
  36328=>"111011111",
  36329=>"011011010",
  36330=>"111111001",
  36331=>"100101000",
  36332=>"100100011",
  36333=>"011111111",
  36334=>"011011011",
  36335=>"000010011",
  36336=>"011010000",
  36337=>"000100110",
  36338=>"100111101",
  36339=>"100100100",
  36340=>"111110001",
  36341=>"001011001",
  36342=>"000000010",
  36343=>"010000110",
  36344=>"110010111",
  36345=>"100000011",
  36346=>"110100111",
  36347=>"110110000",
  36348=>"011110110",
  36349=>"110110110",
  36350=>"000000010",
  36351=>"000100111",
  36352=>"010011111",
  36353=>"101001011",
  36354=>"101101001",
  36355=>"111110010",
  36356=>"110111011",
  36357=>"110000000",
  36358=>"111000111",
  36359=>"000000000",
  36360=>"000111001",
  36361=>"001001111",
  36362=>"101101111",
  36363=>"100101011",
  36364=>"000111110",
  36365=>"010110110",
  36366=>"100000100",
  36367=>"111000001",
  36368=>"101101000",
  36369=>"001001111",
  36370=>"100100000",
  36371=>"001011010",
  36372=>"111101100",
  36373=>"000000110",
  36374=>"100111111",
  36375=>"111000010",
  36376=>"100000000",
  36377=>"000001111",
  36378=>"100001000",
  36379=>"101001101",
  36380=>"111000000",
  36381=>"011101100",
  36382=>"111110001",
  36383=>"101111000",
  36384=>"000000100",
  36385=>"110011111",
  36386=>"000011100",
  36387=>"000010100",
  36388=>"010111111",
  36389=>"110000111",
  36390=>"000000000",
  36391=>"100001110",
  36392=>"000010010",
  36393=>"100111110",
  36394=>"000000100",
  36395=>"000010010",
  36396=>"000011111",
  36397=>"000000111",
  36398=>"010011111",
  36399=>"110010010",
  36400=>"101101101",
  36401=>"100111110",
  36402=>"010010111",
  36403=>"101000001",
  36404=>"101101111",
  36405=>"110110111",
  36406=>"100000011",
  36407=>"101001001",
  36408=>"110000000",
  36409=>"101000000",
  36410=>"010101011",
  36411=>"010001111",
  36412=>"000000100",
  36413=>"010111010",
  36414=>"011001100",
  36415=>"111011100",
  36416=>"000110110",
  36417=>"100010110",
  36418=>"110111111",
  36419=>"100000010",
  36420=>"000110000",
  36421=>"001000000",
  36422=>"010101101",
  36423=>"111101001",
  36424=>"010001011",
  36425=>"111101111",
  36426=>"101000001",
  36427=>"101101101",
  36428=>"111000000",
  36429=>"110110110",
  36430=>"001011011",
  36431=>"110111111",
  36432=>"001000000",
  36433=>"010010000",
  36434=>"001000111",
  36435=>"010000001",
  36436=>"111101111",
  36437=>"110111110",
  36438=>"010011101",
  36439=>"111001111",
  36440=>"111000101",
  36441=>"000001011",
  36442=>"000100100",
  36443=>"100010000",
  36444=>"010000000",
  36445=>"100001010",
  36446=>"111001111",
  36447=>"001000101",
  36448=>"010010010",
  36449=>"000000111",
  36450=>"011000111",
  36451=>"000000111",
  36452=>"101001111",
  36453=>"101100111",
  36454=>"111110100",
  36455=>"111010111",
  36456=>"011000101",
  36457=>"111000000",
  36458=>"010111111",
  36459=>"110111000",
  36460=>"100111110",
  36461=>"001000010",
  36462=>"000101011",
  36463=>"011000111",
  36464=>"001000111",
  36465=>"000000100",
  36466=>"000000100",
  36467=>"000010000",
  36468=>"111010011",
  36469=>"100101111",
  36470=>"111000010",
  36471=>"111000000",
  36472=>"110111111",
  36473=>"010011111",
  36474=>"001001100",
  36475=>"101001010",
  36476=>"000100000",
  36477=>"011101110",
  36478=>"111110110",
  36479=>"001101101",
  36480=>"110110000",
  36481=>"001111000",
  36482=>"011000000",
  36483=>"000010110",
  36484=>"101001101",
  36485=>"100111000",
  36486=>"111001010",
  36487=>"000000011",
  36488=>"101100111",
  36489=>"001000011",
  36490=>"111001001",
  36491=>"110010000",
  36492=>"000000000",
  36493=>"000000111",
  36494=>"001001000",
  36495=>"110000000",
  36496=>"011111110",
  36497=>"011111011",
  36498=>"000000010",
  36499=>"001100101",
  36500=>"000101000",
  36501=>"000000000",
  36502=>"001001101",
  36503=>"000010011",
  36504=>"000111101",
  36505=>"100010011",
  36506=>"001101001",
  36507=>"010001111",
  36508=>"111100110",
  36509=>"011101111",
  36510=>"010010000",
  36511=>"000100110",
  36512=>"000111110",
  36513=>"101000000",
  36514=>"000110100",
  36515=>"010101100",
  36516=>"110010111",
  36517=>"000110100",
  36518=>"000110000",
  36519=>"010111000",
  36520=>"001000111",
  36521=>"000001111",
  36522=>"111101000",
  36523=>"111000000",
  36524=>"000000100",
  36525=>"111000000",
  36526=>"111100100",
  36527=>"000100010",
  36528=>"110010011",
  36529=>"001000110",
  36530=>"101101101",
  36531=>"000000000",
  36532=>"100011001",
  36533=>"111011101",
  36534=>"000011011",
  36535=>"110110101",
  36536=>"011010101",
  36537=>"000101101",
  36538=>"010000101",
  36539=>"111111000",
  36540=>"110000000",
  36541=>"000100111",
  36542=>"001001000",
  36543=>"000000000",
  36544=>"101000000",
  36545=>"111001101",
  36546=>"001000110",
  36547=>"011010110",
  36548=>"000110000",
  36549=>"001010011",
  36550=>"010100000",
  36551=>"000010111",
  36552=>"000010100",
  36553=>"000110010",
  36554=>"110111111",
  36555=>"000000111",
  36556=>"111100100",
  36557=>"001001000",
  36558=>"011000001",
  36559=>"000010111",
  36560=>"000000010",
  36561=>"000110110",
  36562=>"001101111",
  36563=>"000111111",
  36564=>"111100000",
  36565=>"100001101",
  36566=>"111001010",
  36567=>"000011000",
  36568=>"000000000",
  36569=>"000110010",
  36570=>"000110110",
  36571=>"111000000",
  36572=>"001111111",
  36573=>"100000011",
  36574=>"010000101",
  36575=>"001000000",
  36576=>"100111111",
  36577=>"101000001",
  36578=>"111101001",
  36579=>"001100000",
  36580=>"100101001",
  36581=>"100001011",
  36582=>"000010011",
  36583=>"001001010",
  36584=>"010010111",
  36585=>"100001101",
  36586=>"101111110",
  36587=>"100110000",
  36588=>"000110110",
  36589=>"000110110",
  36590=>"000000000",
  36591=>"000101000",
  36592=>"001011111",
  36593=>"100011111",
  36594=>"000001101",
  36595=>"010100101",
  36596=>"110110100",
  36597=>"111100111",
  36598=>"000000111",
  36599=>"001001111",
  36600=>"000000000",
  36601=>"101110110",
  36602=>"100100000",
  36603=>"101111111",
  36604=>"111110001",
  36605=>"000101011",
  36606=>"111111101",
  36607=>"000000000",
  36608=>"110111000",
  36609=>"100000110",
  36610=>"001000101",
  36611=>"111101101",
  36612=>"111011001",
  36613=>"000001111",
  36614=>"010111110",
  36615=>"110000010",
  36616=>"111000101",
  36617=>"010110000",
  36618=>"111111011",
  36619=>"111111111",
  36620=>"101001001",
  36621=>"111011111",
  36622=>"011111111",
  36623=>"000001110",
  36624=>"111111001",
  36625=>"000111010",
  36626=>"100101101",
  36627=>"000000011",
  36628=>"000011011",
  36629=>"011111000",
  36630=>"000000000",
  36631=>"111101000",
  36632=>"010111001",
  36633=>"101001111",
  36634=>"011010111",
  36635=>"010111110",
  36636=>"000011101",
  36637=>"010000010",
  36638=>"111101101",
  36639=>"001000000",
  36640=>"001000001",
  36641=>"001000100",
  36642=>"111000010",
  36643=>"000100101",
  36644=>"001001101",
  36645=>"100011111",
  36646=>"110110110",
  36647=>"001111111",
  36648=>"011110011",
  36649=>"010000011",
  36650=>"111111011",
  36651=>"010001100",
  36652=>"011001000",
  36653=>"001000001",
  36654=>"000000000",
  36655=>"111001111",
  36656=>"000000010",
  36657=>"111011001",
  36658=>"000001000",
  36659=>"001001001",
  36660=>"111110111",
  36661=>"111110011",
  36662=>"010000000",
  36663=>"010000110",
  36664=>"111001111",
  36665=>"000000000",
  36666=>"001001000",
  36667=>"000000001",
  36668=>"110110110",
  36669=>"111111111",
  36670=>"000010010",
  36671=>"111111011",
  36672=>"011010000",
  36673=>"111111000",
  36674=>"101101111",
  36675=>"111110111",
  36676=>"001000111",
  36677=>"010101000",
  36678=>"000010001",
  36679=>"111000100",
  36680=>"001001011",
  36681=>"110110000",
  36682=>"000001111",
  36683=>"101001001",
  36684=>"000000000",
  36685=>"100101110",
  36686=>"011001110",
  36687=>"001101001",
  36688=>"110110110",
  36689=>"000010100",
  36690=>"110111111",
  36691=>"111001001",
  36692=>"000010010",
  36693=>"100101100",
  36694=>"111101110",
  36695=>"110111001",
  36696=>"100101110",
  36697=>"110100101",
  36698=>"110100000",
  36699=>"101101111",
  36700=>"000000110",
  36701=>"001000000",
  36702=>"001001000",
  36703=>"011111111",
  36704=>"000011111",
  36705=>"110110110",
  36706=>"010000000",
  36707=>"100000000",
  36708=>"111101100",
  36709=>"001011001",
  36710=>"010110111",
  36711=>"010000001",
  36712=>"010111111",
  36713=>"010111111",
  36714=>"001000000",
  36715=>"101110111",
  36716=>"010011111",
  36717=>"110111010",
  36718=>"111000000",
  36719=>"000000101",
  36720=>"010110100",
  36721=>"111111110",
  36722=>"000110000",
  36723=>"101111111",
  36724=>"111111010",
  36725=>"000100011",
  36726=>"111110110",
  36727=>"110110110",
  36728=>"101000000",
  36729=>"111101000",
  36730=>"000000011",
  36731=>"111101001",
  36732=>"010100110",
  36733=>"011001000",
  36734=>"111110111",
  36735=>"110110110",
  36736=>"001111110",
  36737=>"111010000",
  36738=>"111110111",
  36739=>"111011100",
  36740=>"110111111",
  36741=>"000000001",
  36742=>"001111111",
  36743=>"100111101",
  36744=>"011001011",
  36745=>"110110110",
  36746=>"010111010",
  36747=>"001000000",
  36748=>"001000000",
  36749=>"110000000",
  36750=>"111111111",
  36751=>"001000001",
  36752=>"001100100",
  36753=>"000101000",
  36754=>"101101111",
  36755=>"100000000",
  36756=>"101111111",
  36757=>"110110101",
  36758=>"111001000",
  36759=>"110001001",
  36760=>"010110010",
  36761=>"101100111",
  36762=>"001000000",
  36763=>"000000100",
  36764=>"000000000",
  36765=>"101100101",
  36766=>"111001111",
  36767=>"110110000",
  36768=>"100000000",
  36769=>"000010000",
  36770=>"010000011",
  36771=>"111100000",
  36772=>"011011101",
  36773=>"000011110",
  36774=>"011111010",
  36775=>"000010110",
  36776=>"000101111",
  36777=>"110101111",
  36778=>"101000000",
  36779=>"110000000",
  36780=>"001000101",
  36781=>"111010000",
  36782=>"001001011",
  36783=>"000000000",
  36784=>"000000000",
  36785=>"001011011",
  36786=>"000010000",
  36787=>"111101000",
  36788=>"010111001",
  36789=>"100000000",
  36790=>"100100100",
  36791=>"101111111",
  36792=>"111110011",
  36793=>"101111111",
  36794=>"111111110",
  36795=>"111000011",
  36796=>"000110111",
  36797=>"011111111",
  36798=>"101001111",
  36799=>"000000000",
  36800=>"001000000",
  36801=>"111000000",
  36802=>"111111010",
  36803=>"111101100",
  36804=>"010111110",
  36805=>"001001011",
  36806=>"000000111",
  36807=>"100000000",
  36808=>"101100000",
  36809=>"101110110",
  36810=>"100000111",
  36811=>"101000000",
  36812=>"110010010",
  36813=>"110010110",
  36814=>"000010000",
  36815=>"000111111",
  36816=>"001010000",
  36817=>"010111110",
  36818=>"110100111",
  36819=>"100100110",
  36820=>"101000001",
  36821=>"000000000",
  36822=>"110110000",
  36823=>"110100000",
  36824=>"000000000",
  36825=>"000110111",
  36826=>"011001010",
  36827=>"101111001",
  36828=>"000000010",
  36829=>"001011001",
  36830=>"001000001",
  36831=>"111100000",
  36832=>"010010010",
  36833=>"010111111",
  36834=>"111110000",
  36835=>"101111111",
  36836=>"011000000",
  36837=>"000000000",
  36838=>"110000111",
  36839=>"010000000",
  36840=>"111110111",
  36841=>"000000111",
  36842=>"110110110",
  36843=>"110110010",
  36844=>"110111110",
  36845=>"111101001",
  36846=>"001001000",
  36847=>"110110110",
  36848=>"000110110",
  36849=>"111001001",
  36850=>"111111101",
  36851=>"111111010",
  36852=>"010100100",
  36853=>"000001000",
  36854=>"110111111",
  36855=>"110111100",
  36856=>"000000000",
  36857=>"111111010",
  36858=>"000111110",
  36859=>"000111111",
  36860=>"000111111",
  36861=>"010010100",
  36862=>"001100110",
  36863=>"000000000",
  36864=>"010110110",
  36865=>"010011111",
  36866=>"000000000",
  36867=>"000000010",
  36868=>"010110111",
  36869=>"000000011",
  36870=>"111111111",
  36871=>"111111010",
  36872=>"000000000",
  36873=>"001001101",
  36874=>"000000001",
  36875=>"001100100",
  36876=>"000000000",
  36877=>"000000001",
  36878=>"010110100",
  36879=>"111111111",
  36880=>"000000000",
  36881=>"001111101",
  36882=>"111111110",
  36883=>"111100111",
  36884=>"100000011",
  36885=>"001001111",
  36886=>"111100100",
  36887=>"010111000",
  36888=>"111001111",
  36889=>"111110000",
  36890=>"011000000",
  36891=>"111101000",
  36892=>"111111001",
  36893=>"000111101",
  36894=>"101100011",
  36895=>"001111100",
  36896=>"000000000",
  36897=>"011000000",
  36898=>"111001101",
  36899=>"000000000",
  36900=>"010111011",
  36901=>"111111101",
  36902=>"110111010",
  36903=>"111000000",
  36904=>"000010000",
  36905=>"100111000",
  36906=>"110111000",
  36907=>"100000000",
  36908=>"011111011",
  36909=>"010101101",
  36910=>"000111110",
  36911=>"110000000",
  36912=>"111111101",
  36913=>"101100001",
  36914=>"101000000",
  36915=>"001011110",
  36916=>"001100111",
  36917=>"011111111",
  36918=>"111010000",
  36919=>"100000110",
  36920=>"000000111",
  36921=>"111111111",
  36922=>"111101000",
  36923=>"111011001",
  36924=>"111110001",
  36925=>"111111111",
  36926=>"111101101",
  36927=>"000001000",
  36928=>"101101100",
  36929=>"100111110",
  36930=>"001101010",
  36931=>"000000111",
  36932=>"111110101",
  36933=>"101101101",
  36934=>"111000100",
  36935=>"000011111",
  36936=>"000010000",
  36937=>"111000010",
  36938=>"111111111",
  36939=>"110100000",
  36940=>"000000000",
  36941=>"111111111",
  36942=>"111001011",
  36943=>"110001101",
  36944=>"000110111",
  36945=>"111111111",
  36946=>"111010111",
  36947=>"011111110",
  36948=>"111111111",
  36949=>"001001000",
  36950=>"101111110",
  36951=>"101101101",
  36952=>"001000000",
  36953=>"111111110",
  36954=>"100001001",
  36955=>"000110100",
  36956=>"111111000",
  36957=>"101101100",
  36958=>"111101111",
  36959=>"001000111",
  36960=>"000000000",
  36961=>"000000000",
  36962=>"111001111",
  36963=>"111111110",
  36964=>"111111111",
  36965=>"000100100",
  36966=>"110111111",
  36967=>"100111101",
  36968=>"101101111",
  36969=>"010000000",
  36970=>"001111000",
  36971=>"110110111",
  36972=>"000000000",
  36973=>"000100000",
  36974=>"000111111",
  36975=>"101011000",
  36976=>"010111111",
  36977=>"111111010",
  36978=>"111101100",
  36979=>"001000000",
  36980=>"111110111",
  36981=>"100100100",
  36982=>"000000110",
  36983=>"010000101",
  36984=>"000010010",
  36985=>"111111000",
  36986=>"011111111",
  36987=>"000000000",
  36988=>"111011111",
  36989=>"101101011",
  36990=>"001000111",
  36991=>"101001111",
  36992=>"110111111",
  36993=>"000000000",
  36994=>"010010100",
  36995=>"001000111",
  36996=>"111111111",
  36997=>"000111111",
  36998=>"100110111",
  36999=>"000010000",
  37000=>"100110111",
  37001=>"001011011",
  37002=>"100101100",
  37003=>"000101110",
  37004=>"000000101",
  37005=>"101100110",
  37006=>"100000001",
  37007=>"001000000",
  37008=>"110011001",
  37009=>"000100101",
  37010=>"111111001",
  37011=>"000000111",
  37012=>"111111101",
  37013=>"000101111",
  37014=>"110111010",
  37015=>"111110110",
  37016=>"111110000",
  37017=>"000010101",
  37018=>"000010000",
  37019=>"000000001",
  37020=>"110100100",
  37021=>"000100000",
  37022=>"010111010",
  37023=>"001111111",
  37024=>"000000000",
  37025=>"111011111",
  37026=>"000000001",
  37027=>"110000000",
  37028=>"011111110",
  37029=>"011111101",
  37030=>"101001001",
  37031=>"000010000",
  37032=>"000111111",
  37033=>"001000000",
  37034=>"011001111",
  37035=>"011101011",
  37036=>"000000101",
  37037=>"101101111",
  37038=>"111011011",
  37039=>"000000100",
  37040=>"000000111",
  37041=>"000000000",
  37042=>"000101000",
  37043=>"001000000",
  37044=>"111000001",
  37045=>"011101111",
  37046=>"000110100",
  37047=>"111110111",
  37048=>"010110100",
  37049=>"101101101",
  37050=>"110110100",
  37051=>"111101101",
  37052=>"111110110",
  37053=>"000000000",
  37054=>"000000000",
  37055=>"000001111",
  37056=>"000000110",
  37057=>"111111101",
  37058=>"010011000",
  37059=>"001001001",
  37060=>"111111000",
  37061=>"111111111",
  37062=>"010111000",
  37063=>"110111110",
  37064=>"111111001",
  37065=>"100100000",
  37066=>"111010111",
  37067=>"000001001",
  37068=>"110110111",
  37069=>"111111111",
  37070=>"111101111",
  37071=>"001000001",
  37072=>"000111111",
  37073=>"001001001",
  37074=>"111100111",
  37075=>"111111011",
  37076=>"010111111",
  37077=>"011001101",
  37078=>"000000000",
  37079=>"110111011",
  37080=>"110110010",
  37081=>"010011010",
  37082=>"000000001",
  37083=>"000000000",
  37084=>"111101001",
  37085=>"000000000",
  37086=>"111011000",
  37087=>"111011111",
  37088=>"000001111",
  37089=>"000001111",
  37090=>"001000100",
  37091=>"000000000",
  37092=>"000100000",
  37093=>"010100011",
  37094=>"101000000",
  37095=>"011011110",
  37096=>"000000000",
  37097=>"001001110",
  37098=>"000000100",
  37099=>"101001111",
  37100=>"000000000",
  37101=>"011110001",
  37102=>"000111110",
  37103=>"110101111",
  37104=>"001100101",
  37105=>"000010111",
  37106=>"111111000",
  37107=>"111111001",
  37108=>"111111001",
  37109=>"000000001",
  37110=>"010011111",
  37111=>"101000111",
  37112=>"110111000",
  37113=>"001101100",
  37114=>"011111111",
  37115=>"001111111",
  37116=>"111111010",
  37117=>"001000000",
  37118=>"000111000",
  37119=>"111111110",
  37120=>"010000101",
  37121=>"010000000",
  37122=>"101100100",
  37123=>"100000000",
  37124=>"011001011",
  37125=>"001001110",
  37126=>"111000111",
  37127=>"000111111",
  37128=>"000011011",
  37129=>"000010011",
  37130=>"000000001",
  37131=>"100000000",
  37132=>"000000100",
  37133=>"010000000",
  37134=>"000111111",
  37135=>"100100111",
  37136=>"100011000",
  37137=>"000000000",
  37138=>"000100011",
  37139=>"100100000",
  37140=>"001011010",
  37141=>"100000100",
  37142=>"111111101",
  37143=>"011000011",
  37144=>"000000000",
  37145=>"111100011",
  37146=>"000100111",
  37147=>"111011010",
  37148=>"100100000",
  37149=>"000000111",
  37150=>"000011000",
  37151=>"000010011",
  37152=>"000101111",
  37153=>"111011011",
  37154=>"010110100",
  37155=>"000000000",
  37156=>"011011001",
  37157=>"001110110",
  37158=>"100100100",
  37159=>"011100111",
  37160=>"100100111",
  37161=>"010111111",
  37162=>"111011010",
  37163=>"110100010",
  37164=>"001011000",
  37165=>"000001000",
  37166=>"000000100",
  37167=>"010110011",
  37168=>"000111111",
  37169=>"000100011",
  37170=>"000101111",
  37171=>"000101100",
  37172=>"001000110",
  37173=>"100000100",
  37174=>"111110110",
  37175=>"011011000",
  37176=>"000000000",
  37177=>"000000000",
  37178=>"111100110",
  37179=>"100101000",
  37180=>"010001110",
  37181=>"111111111",
  37182=>"000000100",
  37183=>"011011011",
  37184=>"100100111",
  37185=>"101111001",
  37186=>"111011011",
  37187=>"011111011",
  37188=>"000010000",
  37189=>"100100100",
  37190=>"011111011",
  37191=>"111011011",
  37192=>"100011110",
  37193=>"011011000",
  37194=>"000000000",
  37195=>"111001100",
  37196=>"000111111",
  37197=>"100111111",
  37198=>"000110110",
  37199=>"000010100",
  37200=>"100110000",
  37201=>"111011001",
  37202=>"011110101",
  37203=>"000100001",
  37204=>"100100110",
  37205=>"100000111",
  37206=>"110100110",
  37207=>"000000011",
  37208=>"000000111",
  37209=>"100110000",
  37210=>"100110110",
  37211=>"010010000",
  37212=>"111011000",
  37213=>"100001001",
  37214=>"011111011",
  37215=>"111011110",
  37216=>"111000010",
  37217=>"101000010",
  37218=>"100000000",
  37219=>"011000000",
  37220=>"000001000",
  37221=>"000100111",
  37222=>"101000101",
  37223=>"111111101",
  37224=>"010011111",
  37225=>"011000010",
  37226=>"011000100",
  37227=>"111101111",
  37228=>"100100111",
  37229=>"111100000",
  37230=>"010100110",
  37231=>"001000010",
  37232=>"000000000",
  37233=>"110000000",
  37234=>"011011000",
  37235=>"011101100",
  37236=>"111010000",
  37237=>"111100000",
  37238=>"011011011",
  37239=>"111111011",
  37240=>"010000011",
  37241=>"011011000",
  37242=>"000100101",
  37243=>"100101010",
  37244=>"000010011",
  37245=>"001000010",
  37246=>"100111111",
  37247=>"000000000",
  37248=>"000011010",
  37249=>"111110011",
  37250=>"111111010",
  37251=>"000111000",
  37252=>"001111000",
  37253=>"000100100",
  37254=>"010001001",
  37255=>"001001000",
  37256=>"000111101",
  37257=>"101100001",
  37258=>"000100100",
  37259=>"111000111",
  37260=>"010010000",
  37261=>"000000101",
  37262=>"111111011",
  37263=>"010101100",
  37264=>"000110110",
  37265=>"000000100",
  37266=>"100100111",
  37267=>"011000000",
  37268=>"001001000",
  37269=>"111111100",
  37270=>"000000010",
  37271=>"000000011",
  37272=>"000011111",
  37273=>"000101111",
  37274=>"110100100",
  37275=>"111110111",
  37276=>"111111111",
  37277=>"000011111",
  37278=>"000100010",
  37279=>"110100100",
  37280=>"000100001",
  37281=>"100110000",
  37282=>"111011111",
  37283=>"000000011",
  37284=>"111100001",
  37285=>"000000000",
  37286=>"100111111",
  37287=>"100000000",
  37288=>"111100000",
  37289=>"000011011",
  37290=>"111100100",
  37291=>"000000000",
  37292=>"111001100",
  37293=>"001011111",
  37294=>"011110000",
  37295=>"000011111",
  37296=>"100000111",
  37297=>"001110000",
  37298=>"111101010",
  37299=>"000000011",
  37300=>"000111000",
  37301=>"011011100",
  37302=>"000111111",
  37303=>"000100011",
  37304=>"000001011",
  37305=>"001011001",
  37306=>"011111000",
  37307=>"010011010",
  37308=>"000000000",
  37309=>"000111011",
  37310=>"111111000",
  37311=>"111111000",
  37312=>"000000100",
  37313=>"010000000",
  37314=>"000011111",
  37315=>"100100110",
  37316=>"011000010",
  37317=>"111111000",
  37318=>"000011011",
  37319=>"111101000",
  37320=>"111111000",
  37321=>"100110000",
  37322=>"000011000",
  37323=>"011011011",
  37324=>"111111000",
  37325=>"100010011",
  37326=>"000000110",
  37327=>"111111100",
  37328=>"000000000",
  37329=>"000000000",
  37330=>"110100000",
  37331=>"111111000",
  37332=>"000000000",
  37333=>"100111111",
  37334=>"111000010",
  37335=>"010000000",
  37336=>"100100111",
  37337=>"000011011",
  37338=>"110100000",
  37339=>"100100100",
  37340=>"111111101",
  37341=>"000011001",
  37342=>"100111111",
  37343=>"010000000",
  37344=>"111011011",
  37345=>"101100100",
  37346=>"111000000",
  37347=>"100001000",
  37348=>"010101111",
  37349=>"011011011",
  37350=>"000010100",
  37351=>"001111011",
  37352=>"000100000",
  37353=>"011000001",
  37354=>"100000000",
  37355=>"000000001",
  37356=>"001000000",
  37357=>"110100000",
  37358=>"111100101",
  37359=>"011000000",
  37360=>"000100100",
  37361=>"001001110",
  37362=>"111011100",
  37363=>"000000010",
  37364=>"111101000",
  37365=>"000000000",
  37366=>"000000111",
  37367=>"111100111",
  37368=>"101000110",
  37369=>"000111111",
  37370=>"011000000",
  37371=>"101111010",
  37372=>"100000000",
  37373=>"000011011",
  37374=>"000110110",
  37375=>"001011010",
  37376=>"000000100",
  37377=>"101101111",
  37378=>"101000101",
  37379=>"000000000",
  37380=>"101000000",
  37381=>"100000001",
  37382=>"111000110",
  37383=>"111111111",
  37384=>"111101000",
  37385=>"101101100",
  37386=>"010100111",
  37387=>"100000001",
  37388=>"101000110",
  37389=>"000001000",
  37390=>"011000110",
  37391=>"000011111",
  37392=>"011000000",
  37393=>"000101000",
  37394=>"111101011",
  37395=>"101100000",
  37396=>"111111111",
  37397=>"000010000",
  37398=>"100000010",
  37399=>"101111101",
  37400=>"000101001",
  37401=>"111101101",
  37402=>"111001000",
  37403=>"000100111",
  37404=>"100101000",
  37405=>"010011111",
  37406=>"000101000",
  37407=>"000010000",
  37408=>"110111101",
  37409=>"000000111",
  37410=>"010110111",
  37411=>"111000000",
  37412=>"100110110",
  37413=>"100001111",
  37414=>"000010000",
  37415=>"111010100",
  37416=>"000010000",
  37417=>"011111011",
  37418=>"101100010",
  37419=>"110010000",
  37420=>"001111000",
  37421=>"111100000",
  37422=>"100101111",
  37423=>"111001000",
  37424=>"000101000",
  37425=>"000000000",
  37426=>"110110010",
  37427=>"000101000",
  37428=>"101010111",
  37429=>"000010010",
  37430=>"101110110",
  37431=>"000000010",
  37432=>"010111001",
  37433=>"000001011",
  37434=>"110010010",
  37435=>"101110100",
  37436=>"110001001",
  37437=>"101010100",
  37438=>"100000100",
  37439=>"011111011",
  37440=>"111101111",
  37441=>"000111001",
  37442=>"011101101",
  37443=>"100000101",
  37444=>"111101111",
  37445=>"000101000",
  37446=>"000111111",
  37447=>"111111011",
  37448=>"010110000",
  37449=>"111101111",
  37450=>"100100110",
  37451=>"000010000",
  37452=>"010000001",
  37453=>"000000011",
  37454=>"100000100",
  37455=>"010110100",
  37456=>"001101111",
  37457=>"111111110",
  37458=>"011101101",
  37459=>"110011000",
  37460=>"101100101",
  37461=>"111110111",
  37462=>"001011001",
  37463=>"101000111",
  37464=>"111000101",
  37465=>"100001000",
  37466=>"011001000",
  37467=>"001001100",
  37468=>"000000101",
  37469=>"011001000",
  37470=>"111010000",
  37471=>"001000100",
  37472=>"111001000",
  37473=>"000000000",
  37474=>"101000001",
  37475=>"110100000",
  37476=>"110000011",
  37477=>"110100100",
  37478=>"010101111",
  37479=>"010111000",
  37480=>"101111000",
  37481=>"100101000",
  37482=>"110000010",
  37483=>"010100111",
  37484=>"010111111",
  37485=>"010011001",
  37486=>"100100101",
  37487=>"000111111",
  37488=>"001000111",
  37489=>"100100100",
  37490=>"101111001",
  37491=>"011000100",
  37492=>"110010010",
  37493=>"111101000",
  37494=>"101101010",
  37495=>"010000000",
  37496=>"110000000",
  37497=>"000110010",
  37498=>"000111101",
  37499=>"000011000",
  37500=>"011001010",
  37501=>"011110000",
  37502=>"010110000",
  37503=>"101001111",
  37504=>"000000000",
  37505=>"001000111",
  37506=>"000000101",
  37507=>"010010110",
  37508=>"101000000",
  37509=>"110111000",
  37510=>"000100110",
  37511=>"000000100",
  37512=>"101001111",
  37513=>"000101001",
  37514=>"011011011",
  37515=>"101001000",
  37516=>"000000101",
  37517=>"101001101",
  37518=>"000000000",
  37519=>"101000000",
  37520=>"001011010",
  37521=>"100000100",
  37522=>"101000100",
  37523=>"000001110",
  37524=>"011101000",
  37525=>"100100000",
  37526=>"111101111",
  37527=>"100111011",
  37528=>"010010001",
  37529=>"101000000",
  37530=>"010111111",
  37531=>"111111000",
  37532=>"111100101",
  37533=>"000000101",
  37534=>"100111000",
  37535=>"101101111",
  37536=>"110111110",
  37537=>"101111011",
  37538=>"110011000",
  37539=>"100010111",
  37540=>"010110000",
  37541=>"000100101",
  37542=>"001110000",
  37543=>"000101000",
  37544=>"000100100",
  37545=>"101101111",
  37546=>"111101100",
  37547=>"101000101",
  37548=>"000111111",
  37549=>"110000011",
  37550=>"011011111",
  37551=>"111010100",
  37552=>"000000000",
  37553=>"000001010",
  37554=>"111100110",
  37555=>"000000010",
  37556=>"010011001",
  37557=>"011111110",
  37558=>"011011000",
  37559=>"000001001",
  37560=>"100000110",
  37561=>"100001000",
  37562=>"000000101",
  37563=>"011111101",
  37564=>"010000000",
  37565=>"111001100",
  37566=>"110001000",
  37567=>"000000000",
  37568=>"010110010",
  37569=>"000000010",
  37570=>"101011010",
  37571=>"110100010",
  37572=>"000000000",
  37573=>"100110000",
  37574=>"000110101",
  37575=>"001000010",
  37576=>"110101000",
  37577=>"000100100",
  37578=>"111100100",
  37579=>"100000100",
  37580=>"001000000",
  37581=>"111110010",
  37582=>"111000111",
  37583=>"000001000",
  37584=>"011110111",
  37585=>"010111110",
  37586=>"100100000",
  37587=>"100100101",
  37588=>"000000111",
  37589=>"110100111",
  37590=>"111001101",
  37591=>"001001111",
  37592=>"010010000",
  37593=>"001001111",
  37594=>"000010010",
  37595=>"110000000",
  37596=>"001011010",
  37597=>"111011100",
  37598=>"010111111",
  37599=>"001100111",
  37600=>"111000111",
  37601=>"100000000",
  37602=>"100010000",
  37603=>"001000011",
  37604=>"000000000",
  37605=>"111001000",
  37606=>"000101000",
  37607=>"110110010",
  37608=>"111101111",
  37609=>"010000000",
  37610=>"011010011",
  37611=>"111000000",
  37612=>"101001000",
  37613=>"000000010",
  37614=>"111101110",
  37615=>"000000111",
  37616=>"000000000",
  37617=>"110011000",
  37618=>"111110111",
  37619=>"100110000",
  37620=>"000110001",
  37621=>"111011101",
  37622=>"000000111",
  37623=>"010011011",
  37624=>"000010111",
  37625=>"110010000",
  37626=>"000010010",
  37627=>"010011010",
  37628=>"000010011",
  37629=>"101100101",
  37630=>"000001110",
  37631=>"000111111",
  37632=>"011000000",
  37633=>"110110110",
  37634=>"000000000",
  37635=>"100100100",
  37636=>"110010011",
  37637=>"001100111",
  37638=>"110110000",
  37639=>"110101101",
  37640=>"011111111",
  37641=>"000000100",
  37642=>"111111111",
  37643=>"011010111",
  37644=>"110101111",
  37645=>"000000000",
  37646=>"001101011",
  37647=>"010010000",
  37648=>"000110111",
  37649=>"011011110",
  37650=>"100010000",
  37651=>"110110100",
  37652=>"111111010",
  37653=>"001101110",
  37654=>"011100111",
  37655=>"111110110",
  37656=>"000000100",
  37657=>"011000000",
  37658=>"011011100",
  37659=>"000010000",
  37660=>"010001001",
  37661=>"111011101",
  37662=>"001100000",
  37663=>"000111011",
  37664=>"111011110",
  37665=>"011011011",
  37666=>"111111000",
  37667=>"101111100",
  37668=>"110101111",
  37669=>"010100111",
  37670=>"000001001",
  37671=>"110110110",
  37672=>"100011011",
  37673=>"010010101",
  37674=>"000100000",
  37675=>"001001000",
  37676=>"000101011",
  37677=>"011100101",
  37678=>"011000110",
  37679=>"111111001",
  37680=>"010000001",
  37681=>"111011001",
  37682=>"111101001",
  37683=>"111010000",
  37684=>"111111110",
  37685=>"110100000",
  37686=>"000000001",
  37687=>"111101000",
  37688=>"110000011",
  37689=>"110100111",
  37690=>"000100111",
  37691=>"011100100",
  37692=>"011000000",
  37693=>"000011011",
  37694=>"000000000",
  37695=>"001001011",
  37696=>"110111011",
  37697=>"000000110",
  37698=>"011111111",
  37699=>"011110110",
  37700=>"000010010",
  37701=>"010000000",
  37702=>"000000000",
  37703=>"011011111",
  37704=>"001101110",
  37705=>"100100110",
  37706=>"100100011",
  37707=>"100010010",
  37708=>"011000000",
  37709=>"011001101",
  37710=>"110110100",
  37711=>"110011111",
  37712=>"100001001",
  37713=>"001010101",
  37714=>"010000100",
  37715=>"001000110",
  37716=>"010010000",
  37717=>"100111110",
  37718=>"000001011",
  37719=>"001000100",
  37720=>"001111110",
  37721=>"100101101",
  37722=>"000000000",
  37723=>"111001011",
  37724=>"011110100",
  37725=>"001001011",
  37726=>"000110110",
  37727=>"101101011",
  37728=>"000011011",
  37729=>"100000100",
  37730=>"100100100",
  37731=>"000000011",
  37732=>"100100001",
  37733=>"000110110",
  37734=>"111110111",
  37735=>"010001001",
  37736=>"110000110",
  37737=>"111100110",
  37738=>"011010111",
  37739=>"110110011",
  37740=>"011111011",
  37741=>"010011001",
  37742=>"101111100",
  37743=>"111011011",
  37744=>"110110010",
  37745=>"111101111",
  37746=>"111110110",
  37747=>"000001000",
  37748=>"111000010",
  37749=>"010100100",
  37750=>"010000000",
  37751=>"111001100",
  37752=>"000000100",
  37753=>"001010000",
  37754=>"110000000",
  37755=>"000000000",
  37756=>"001001111",
  37757=>"110100001",
  37758=>"110100010",
  37759=>"000001000",
  37760=>"111000010",
  37761=>"000000000",
  37762=>"011011100",
  37763=>"011111011",
  37764=>"011010000",
  37765=>"001010010",
  37766=>"000000000",
  37767=>"000000000",
  37768=>"100101000",
  37769=>"010000010",
  37770=>"100000111",
  37771=>"001000111",
  37772=>"000001011",
  37773=>"111111011",
  37774=>"011111111",
  37775=>"000000000",
  37776=>"110100100",
  37777=>"101011011",
  37778=>"000000110",
  37779=>"101110111",
  37780=>"100001000",
  37781=>"001000110",
  37782=>"010010010",
  37783=>"011111011",
  37784=>"011111001",
  37785=>"100110001",
  37786=>"000010000",
  37787=>"000000101",
  37788=>"000011011",
  37789=>"001011011",
  37790=>"011110110",
  37791=>"001001011",
  37792=>"111100100",
  37793=>"010111000",
  37794=>"111110101",
  37795=>"110000111",
  37796=>"011110110",
  37797=>"010110110",
  37798=>"110000001",
  37799=>"001010010",
  37800=>"011000000",
  37801=>"000110111",
  37802=>"011001000",
  37803=>"010100000",
  37804=>"111111000",
  37805=>"111111111",
  37806=>"111111111",
  37807=>"000100100",
  37808=>"000000000",
  37809=>"000000000",
  37810=>"110111100",
  37811=>"000100111",
  37812=>"101100001",
  37813=>"111100111",
  37814=>"101001000",
  37815=>"001001000",
  37816=>"001010000",
  37817=>"001000000",
  37818=>"001000000",
  37819=>"011111011",
  37820=>"100100000",
  37821=>"001111011",
  37822=>"001001001",
  37823=>"100000000",
  37824=>"110010000",
  37825=>"010000000",
  37826=>"111000101",
  37827=>"011101001",
  37828=>"001100111",
  37829=>"110000111",
  37830=>"111111111",
  37831=>"010001101",
  37832=>"000001100",
  37833=>"010010010",
  37834=>"111001110",
  37835=>"000000010",
  37836=>"001000000",
  37837=>"111111100",
  37838=>"100111000",
  37839=>"110110011",
  37840=>"010010000",
  37841=>"011101001",
  37842=>"000001011",
  37843=>"011111110",
  37844=>"111011001",
  37845=>"111111111",
  37846=>"100000100",
  37847=>"010000000",
  37848=>"010100100",
  37849=>"000000110",
  37850=>"110110110",
  37851=>"100000000",
  37852=>"111001010",
  37853=>"000001000",
  37854=>"011010010",
  37855=>"011010001",
  37856=>"000111001",
  37857=>"111100000",
  37858=>"010110100",
  37859=>"001000000",
  37860=>"000000000",
  37861=>"011001000",
  37862=>"111001100",
  37863=>"000000000",
  37864=>"000001010",
  37865=>"011011110",
  37866=>"000000000",
  37867=>"001011111",
  37868=>"100101011",
  37869=>"111111100",
  37870=>"001011010",
  37871=>"001000100",
  37872=>"010010000",
  37873=>"001111100",
  37874=>"001000000",
  37875=>"001101011",
  37876=>"111111111",
  37877=>"100101101",
  37878=>"000000000",
  37879=>"100110001",
  37880=>"000110000",
  37881=>"110100100",
  37882=>"111111011",
  37883=>"110110110",
  37884=>"110111101",
  37885=>"011011000",
  37886=>"101111101",
  37887=>"000010000",
  37888=>"100100110",
  37889=>"111111000",
  37890=>"000000100",
  37891=>"111010000",
  37892=>"000000000",
  37893=>"111111111",
  37894=>"101000000",
  37895=>"111111100",
  37896=>"010011011",
  37897=>"000000001",
  37898=>"100001100",
  37899=>"000000000",
  37900=>"111111001",
  37901=>"000111111",
  37902=>"110100000",
  37903=>"000000000",
  37904=>"101110111",
  37905=>"111100100",
  37906=>"101000000",
  37907=>"000000000",
  37908=>"101000000",
  37909=>"101101101",
  37910=>"011000000",
  37911=>"111111111",
  37912=>"111010011",
  37913=>"000110000",
  37914=>"000000000",
  37915=>"100111010",
  37916=>"001000100",
  37917=>"000101000",
  37918=>"000100110",
  37919=>"000000001",
  37920=>"011101100",
  37921=>"000010011",
  37922=>"111101100",
  37923=>"011000000",
  37924=>"000100000",
  37925=>"000000000",
  37926=>"111000101",
  37927=>"111001101",
  37928=>"101100101",
  37929=>"101101111",
  37930=>"101000000",
  37931=>"010111111",
  37932=>"000101101",
  37933=>"111110011",
  37934=>"011101111",
  37935=>"101000100",
  37936=>"100100111",
  37937=>"101110111",
  37938=>"000000100",
  37939=>"011101111",
  37940=>"101000000",
  37941=>"000110100",
  37942=>"100100001",
  37943=>"000000000",
  37944=>"010111111",
  37945=>"101101101",
  37946=>"101000111",
  37947=>"011000111",
  37948=>"001000011",
  37949=>"100111111",
  37950=>"000000010",
  37951=>"101010001",
  37952=>"111111011",
  37953=>"011000000",
  37954=>"111001101",
  37955=>"000001110",
  37956=>"000111111",
  37957=>"101100000",
  37958=>"100111011",
  37959=>"111111111",
  37960=>"000111111",
  37961=>"000000111",
  37962=>"111111000",
  37963=>"001000000",
  37964=>"000001101",
  37965=>"101111000",
  37966=>"010111111",
  37967=>"000001111",
  37968=>"000100101",
  37969=>"110111111",
  37970=>"100001101",
  37971=>"101000000",
  37972=>"110000000",
  37973=>"010101110",
  37974=>"000000000",
  37975=>"000000000",
  37976=>"100111111",
  37977=>"000000000",
  37978=>"000110011",
  37979=>"111111010",
  37980=>"001011011",
  37981=>"100110010",
  37982=>"011111111",
  37983=>"000000000",
  37984=>"000001000",
  37985=>"111111000",
  37986=>"000110101",
  37987=>"001111110",
  37988=>"000000000",
  37989=>"100000000",
  37990=>"001100000",
  37991=>"000101111",
  37992=>"111010001",
  37993=>"000000000",
  37994=>"001000000",
  37995=>"000010111",
  37996=>"000000000",
  37997=>"000111100",
  37998=>"000000000",
  37999=>"111111111",
  38000=>"100111111",
  38001=>"000000000",
  38002=>"001001000",
  38003=>"100000000",
  38004=>"000101111",
  38005=>"111110110",
  38006=>"000000000",
  38007=>"000000000",
  38008=>"001010011",
  38009=>"111111010",
  38010=>"001110110",
  38011=>"101000111",
  38012=>"011001000",
  38013=>"001011011",
  38014=>"100111111",
  38015=>"000001010",
  38016=>"000010000",
  38017=>"000000000",
  38018=>"000001011",
  38019=>"101000010",
  38020=>"000000000",
  38021=>"101010101",
  38022=>"001000010",
  38023=>"100000000",
  38024=>"000111000",
  38025=>"000100101",
  38026=>"100000000",
  38027=>"101010111",
  38028=>"000011111",
  38029=>"111111111",
  38030=>"011000010",
  38031=>"001000000",
  38032=>"111010111",
  38033=>"000101000",
  38034=>"000000000",
  38035=>"111011000",
  38036=>"010000000",
  38037=>"000001000",
  38038=>"010111011",
  38039=>"000000101",
  38040=>"001000100",
  38041=>"111011011",
  38042=>"001111111",
  38043=>"111000000",
  38044=>"100000000",
  38045=>"111111111",
  38046=>"111000011",
  38047=>"000000000",
  38048=>"000001111",
  38049=>"010111111",
  38050=>"000011111",
  38051=>"100001111",
  38052=>"000011010",
  38053=>"001100100",
  38054=>"111101001",
  38055=>"000000000",
  38056=>"111010000",
  38057=>"111000101",
  38058=>"000111011",
  38059=>"000010001",
  38060=>"110111000",
  38061=>"111100111",
  38062=>"000011111",
  38063=>"101111001",
  38064=>"000000000",
  38065=>"100110110",
  38066=>"111000000",
  38067=>"011011011",
  38068=>"111111111",
  38069=>"100000001",
  38070=>"000101001",
  38071=>"000111011",
  38072=>"100100000",
  38073=>"000000000",
  38074=>"000001111",
  38075=>"000000010",
  38076=>"000000000",
  38077=>"110111111",
  38078=>"001111010",
  38079=>"110000100",
  38080=>"000000000",
  38081=>"000101010",
  38082=>"111111100",
  38083=>"000001001",
  38084=>"001000110",
  38085=>"010010110",
  38086=>"111111111",
  38087=>"001111001",
  38088=>"000110011",
  38089=>"100000000",
  38090=>"000000010",
  38091=>"111000000",
  38092=>"000000000",
  38093=>"010100100",
  38094=>"011111011",
  38095=>"111111111",
  38096=>"000111001",
  38097=>"000110110",
  38098=>"010111001",
  38099=>"101100101",
  38100=>"001000000",
  38101=>"001011011",
  38102=>"000000101",
  38103=>"000010101",
  38104=>"001000100",
  38105=>"110111000",
  38106=>"000000011",
  38107=>"000010110",
  38108=>"010011010",
  38109=>"110110111",
  38110=>"101000000",
  38111=>"000100101",
  38112=>"101000000",
  38113=>"000011111",
  38114=>"111011111",
  38115=>"011011001",
  38116=>"000000001",
  38117=>"000000010",
  38118=>"011001101",
  38119=>"000111010",
  38120=>"111111011",
  38121=>"110111111",
  38122=>"101100000",
  38123=>"000000011",
  38124=>"000011010",
  38125=>"100100000",
  38126=>"000111000",
  38127=>"010000000",
  38128=>"111100111",
  38129=>"010000011",
  38130=>"000000110",
  38131=>"111011001",
  38132=>"000001011",
  38133=>"000010111",
  38134=>"111010110",
  38135=>"111010011",
  38136=>"000000000",
  38137=>"000011101",
  38138=>"100000000",
  38139=>"010010000",
  38140=>"111111101",
  38141=>"011010010",
  38142=>"100000000",
  38143=>"111001000",
  38144=>"110011000",
  38145=>"111111111",
  38146=>"010111111",
  38147=>"111101100",
  38148=>"010010111",
  38149=>"110111111",
  38150=>"000000101",
  38151=>"101000000",
  38152=>"111000101",
  38153=>"101100001",
  38154=>"000000000",
  38155=>"101101111",
  38156=>"111111011",
  38157=>"101101101",
  38158=>"010000011",
  38159=>"010100000",
  38160=>"001000100",
  38161=>"111101101",
  38162=>"010011010",
  38163=>"111000100",
  38164=>"010111010",
  38165=>"001010000",
  38166=>"100011011",
  38167=>"000000000",
  38168=>"010111000",
  38169=>"000001010",
  38170=>"111101111",
  38171=>"111010000",
  38172=>"111111010",
  38173=>"101110111",
  38174=>"011111101",
  38175=>"111000101",
  38176=>"111111111",
  38177=>"001111010",
  38178=>"111101110",
  38179=>"111111111",
  38180=>"001000100",
  38181=>"100000110",
  38182=>"100101001",
  38183=>"111000111",
  38184=>"000100100",
  38185=>"101101001",
  38186=>"000000101",
  38187=>"111111111",
  38188=>"100000100",
  38189=>"000011111",
  38190=>"000000010",
  38191=>"100001000",
  38192=>"001101111",
  38193=>"110010110",
  38194=>"111101111",
  38195=>"111111000",
  38196=>"111111000",
  38197=>"110001000",
  38198=>"111110100",
  38199=>"111010000",
  38200=>"101101001",
  38201=>"011011000",
  38202=>"111111111",
  38203=>"000000101",
  38204=>"111111111",
  38205=>"000000000",
  38206=>"011111010",
  38207=>"000000100",
  38208=>"000000000",
  38209=>"111101111",
  38210=>"001001101",
  38211=>"011011001",
  38212=>"111101101",
  38213=>"000010010",
  38214=>"111111111",
  38215=>"111111111",
  38216=>"010000010",
  38217=>"101100101",
  38218=>"111111111",
  38219=>"110110100",
  38220=>"110111101",
  38221=>"110000011",
  38222=>"001000000",
  38223=>"000011011",
  38224=>"111101111",
  38225=>"000010000",
  38226=>"101000000",
  38227=>"110100111",
  38228=>"111111111",
  38229=>"010000000",
  38230=>"111100100",
  38231=>"111101111",
  38232=>"101101100",
  38233=>"111000110",
  38234=>"111011111",
  38235=>"001000111",
  38236=>"111000000",
  38237=>"111111110",
  38238=>"100111000",
  38239=>"000110100",
  38240=>"101101101",
  38241=>"101101100",
  38242=>"011111010",
  38243=>"011010010",
  38244=>"011000011",
  38245=>"000000011",
  38246=>"101000000",
  38247=>"110000001",
  38248=>"010010000",
  38249=>"111000000",
  38250=>"000000000",
  38251=>"100101000",
  38252=>"111011111",
  38253=>"111110010",
  38254=>"000011011",
  38255=>"101111111",
  38256=>"011001001",
  38257=>"101001000",
  38258=>"001011000",
  38259=>"110111111",
  38260=>"110100101",
  38261=>"011111011",
  38262=>"100100100",
  38263=>"001100111",
  38264=>"111101100",
  38265=>"001000000",
  38266=>"000000000",
  38267=>"011011011",
  38268=>"011011001",
  38269=>"011011111",
  38270=>"011111000",
  38271=>"010111110",
  38272=>"110111101",
  38273=>"000001011",
  38274=>"101000101",
  38275=>"101000001",
  38276=>"010001000",
  38277=>"000001000",
  38278=>"001001111",
  38279=>"000010100",
  38280=>"010000110",
  38281=>"000001101",
  38282=>"110000100",
  38283=>"111111111",
  38284=>"101111111",
  38285=>"000000010",
  38286=>"111011011",
  38287=>"110111111",
  38288=>"010000110",
  38289=>"111001001",
  38290=>"010111101",
  38291=>"001101000",
  38292=>"111100001",
  38293=>"011001001",
  38294=>"001010000",
  38295=>"111100100",
  38296=>"000001000",
  38297=>"111101000",
  38298=>"011011010",
  38299=>"010111111",
  38300=>"101101111",
  38301=>"100100000",
  38302=>"000101101",
  38303=>"011011011",
  38304=>"110110110",
  38305=>"111111101",
  38306=>"001000111",
  38307=>"111111010",
  38308=>"011001001",
  38309=>"001100111",
  38310=>"100101101",
  38311=>"111000101",
  38312=>"000000001",
  38313=>"111101101",
  38314=>"000011000",
  38315=>"111111010",
  38316=>"100111111",
  38317=>"111001111",
  38318=>"011011010",
  38319=>"100000101",
  38320=>"111011010",
  38321=>"110001001",
  38322=>"111111111",
  38323=>"111111011",
  38324=>"101000100",
  38325=>"111111111",
  38326=>"100000111",
  38327=>"100111110",
  38328=>"101111111",
  38329=>"110000010",
  38330=>"111000000",
  38331=>"001100000",
  38332=>"101100111",
  38333=>"000111111",
  38334=>"111001111",
  38335=>"111101101",
  38336=>"111111000",
  38337=>"111000111",
  38338=>"010101101",
  38339=>"011101011",
  38340=>"100101111",
  38341=>"000110011",
  38342=>"111100000",
  38343=>"000010000",
  38344=>"101100010",
  38345=>"000010011",
  38346=>"000111011",
  38347=>"111110000",
  38348=>"111000000",
  38349=>"111111100",
  38350=>"111101101",
  38351=>"011000000",
  38352=>"010111010",
  38353=>"011001011",
  38354=>"000111101",
  38355=>"010010000",
  38356=>"010011010",
  38357=>"111111111",
  38358=>"111111100",
  38359=>"111101000",
  38360=>"000000000",
  38361=>"011001001",
  38362=>"011011011",
  38363=>"010111111",
  38364=>"001000111",
  38365=>"100100100",
  38366=>"101101111",
  38367=>"001001001",
  38368=>"010011011",
  38369=>"010111010",
  38370=>"000000010",
  38371=>"110001111",
  38372=>"111101111",
  38373=>"000111101",
  38374=>"111111110",
  38375=>"111101001",
  38376=>"101101000",
  38377=>"111111111",
  38378=>"000010001",
  38379=>"101101111",
  38380=>"111111111",
  38381=>"111111111",
  38382=>"110110111",
  38383=>"000010110",
  38384=>"010010011",
  38385=>"000110110",
  38386=>"100101100",
  38387=>"011001011",
  38388=>"110000101",
  38389=>"000110000",
  38390=>"101111101",
  38391=>"101101000",
  38392=>"001111011",
  38393=>"101101001",
  38394=>"000111000",
  38395=>"001101000",
  38396=>"000000000",
  38397=>"000000111",
  38398=>"011001110",
  38399=>"010010111",
  38400=>"000000000",
  38401=>"011000111",
  38402=>"000000101",
  38403=>"010000000",
  38404=>"100110111",
  38405=>"100100110",
  38406=>"011000100",
  38407=>"000000010",
  38408=>"000111110",
  38409=>"000101101",
  38410=>"001001001",
  38411=>"111111100",
  38412=>"111111101",
  38413=>"011101011",
  38414=>"100111001",
  38415=>"111011000",
  38416=>"010000011",
  38417=>"010111100",
  38418=>"010100100",
  38419=>"111100010",
  38420=>"110111110",
  38421=>"111100100",
  38422=>"011100101",
  38423=>"000010100",
  38424=>"000000011",
  38425=>"111111001",
  38426=>"011111011",
  38427=>"100100001",
  38428=>"000000001",
  38429=>"000100111",
  38430=>"110000000",
  38431=>"101111000",
  38432=>"101101111",
  38433=>"111111000",
  38434=>"010011001",
  38435=>"000111111",
  38436=>"100110100",
  38437=>"010010000",
  38438=>"010011110",
  38439=>"000001111",
  38440=>"111011000",
  38441=>"111000000",
  38442=>"100100000",
  38443=>"000010000",
  38444=>"110101011",
  38445=>"100000010",
  38446=>"010010011",
  38447=>"110111101",
  38448=>"100111111",
  38449=>"100110111",
  38450=>"000110011",
  38451=>"000000000",
  38452=>"000000100",
  38453=>"000000001",
  38454=>"000000000",
  38455=>"000000100",
  38456=>"010010111",
  38457=>"000000000",
  38458=>"000000110",
  38459=>"000101111",
  38460=>"001000111",
  38461=>"100111101",
  38462=>"000101111",
  38463=>"111000110",
  38464=>"111111111",
  38465=>"000000111",
  38466=>"000000110",
  38467=>"011001010",
  38468=>"011111111",
  38469=>"000000000",
  38470=>"001001011",
  38471=>"110011101",
  38472=>"000111111",
  38473=>"000111111",
  38474=>"000011111",
  38475=>"000000011",
  38476=>"000100111",
  38477=>"111111011",
  38478=>"101001001",
  38479=>"011011111",
  38480=>"001000000",
  38481=>"111100000",
  38482=>"111011010",
  38483=>"111100001",
  38484=>"111010000",
  38485=>"111100001",
  38486=>"001001111",
  38487=>"000000101",
  38488=>"111110101",
  38489=>"000011000",
  38490=>"111111000",
  38491=>"111011001",
  38492=>"010111111",
  38493=>"000001001",
  38494=>"111011000",
  38495=>"000000001",
  38496=>"000000000",
  38497=>"111100000",
  38498=>"000000100",
  38499=>"001011011",
  38500=>"000100000",
  38501=>"000110100",
  38502=>"000111100",
  38503=>"011001111",
  38504=>"011111100",
  38505=>"100000000",
  38506=>"111100111",
  38507=>"000101011",
  38508=>"011111111",
  38509=>"000010010",
  38510=>"101101011",
  38511=>"000000000",
  38512=>"001011111",
  38513=>"000000111",
  38514=>"000100000",
  38515=>"100000000",
  38516=>"010110000",
  38517=>"000000000",
  38518=>"000001010",
  38519=>"010010000",
  38520=>"100000101",
  38521=>"111111111",
  38522=>"101111011",
  38523=>"100110100",
  38524=>"000100000",
  38525=>"000100100",
  38526=>"001111111",
  38527=>"000000100",
  38528=>"011011000",
  38529=>"000100000",
  38530=>"000111011",
  38531=>"100101011",
  38532=>"111000000",
  38533=>"100100000",
  38534=>"010001011",
  38535=>"000011000",
  38536=>"101001111",
  38537=>"100000000",
  38538=>"010111101",
  38539=>"000001111",
  38540=>"011000000",
  38541=>"101011000",
  38542=>"111011011",
  38543=>"000000000",
  38544=>"001101011",
  38545=>"100111101",
  38546=>"101111110",
  38547=>"001010111",
  38548=>"010110001",
  38549=>"000000111",
  38550=>"111000001",
  38551=>"001001000",
  38552=>"100111011",
  38553=>"000000000",
  38554=>"011011000",
  38555=>"000000010",
  38556=>"100000100",
  38557=>"101111111",
  38558=>"011100101",
  38559=>"111010110",
  38560=>"111100100",
  38561=>"000000011",
  38562=>"001111111",
  38563=>"111111000",
  38564=>"110101111",
  38565=>"110111010",
  38566=>"101000010",
  38567=>"000000000",
  38568=>"110000010",
  38569=>"000010010",
  38570=>"001111101",
  38571=>"000011111",
  38572=>"011011000",
  38573=>"001101111",
  38574=>"000001011",
  38575=>"111011001",
  38576=>"111111100",
  38577=>"100010000",
  38578=>"000100000",
  38579=>"000100000",
  38580=>"001011000",
  38581=>"101110000",
  38582=>"011111000",
  38583=>"000000000",
  38584=>"000001111",
  38585=>"101110100",
  38586=>"010001000",
  38587=>"011011111",
  38588=>"000001010",
  38589=>"101101111",
  38590=>"001001001",
  38591=>"111110101",
  38592=>"000000001",
  38593=>"000000000",
  38594=>"000101101",
  38595=>"111110000",
  38596=>"011000111",
  38597=>"110001001",
  38598=>"111100101",
  38599=>"000100111",
  38600=>"000001101",
  38601=>"111011010",
  38602=>"111010000",
  38603=>"000000111",
  38604=>"000000111",
  38605=>"000000000",
  38606=>"000000001",
  38607=>"101101001",
  38608=>"100101111",
  38609=>"101101111",
  38610=>"101111011",
  38611=>"000010111",
  38612=>"101111010",
  38613=>"000100000",
  38614=>"000000101",
  38615=>"011011001",
  38616=>"011011000",
  38617=>"001000010",
  38618=>"101101000",
  38619=>"111001000",
  38620=>"100000111",
  38621=>"111111000",
  38622=>"111111000",
  38623=>"111000000",
  38624=>"010111010",
  38625=>"000000101",
  38626=>"110000000",
  38627=>"111110110",
  38628=>"000000001",
  38629=>"100000000",
  38630=>"111111000",
  38631=>"010000101",
  38632=>"000000001",
  38633=>"000100010",
  38634=>"000000010",
  38635=>"100000101",
  38636=>"010010110",
  38637=>"000000100",
  38638=>"000000000",
  38639=>"000100111",
  38640=>"100111111",
  38641=>"011000110",
  38642=>"111000000",
  38643=>"000111111",
  38644=>"101100110",
  38645=>"100001101",
  38646=>"000000011",
  38647=>"111001000",
  38648=>"000010010",
  38649=>"000011100",
  38650=>"111010000",
  38651=>"101100100",
  38652=>"000001111",
  38653=>"101010010",
  38654=>"111111110",
  38655=>"100000110",
  38656=>"101101100",
  38657=>"000000011",
  38658=>"100100110",
  38659=>"010010001",
  38660=>"101101101",
  38661=>"010010111",
  38662=>"011011001",
  38663=>"000001000",
  38664=>"011000000",
  38665=>"100100100",
  38666=>"100010000",
  38667=>"000000110",
  38668=>"011010011",
  38669=>"111111110",
  38670=>"000110101",
  38671=>"110111111",
  38672=>"000000100",
  38673=>"111110100",
  38674=>"110110100",
  38675=>"111001001",
  38676=>"000100000",
  38677=>"001101111",
  38678=>"110100000",
  38679=>"001001011",
  38680=>"110100100",
  38681=>"011100110",
  38682=>"010110100",
  38683=>"100100000",
  38684=>"000000110",
  38685=>"111010111",
  38686=>"001111111",
  38687=>"000000011",
  38688=>"100100000",
  38689=>"000000100",
  38690=>"111110000",
  38691=>"000000001",
  38692=>"010110100",
  38693=>"001110110",
  38694=>"101001011",
  38695=>"111111111",
  38696=>"010011011",
  38697=>"000001100",
  38698=>"000001001",
  38699=>"000100100",
  38700=>"000010111",
  38701=>"000000001",
  38702=>"001111110",
  38703=>"001010111",
  38704=>"111111110",
  38705=>"001111101",
  38706=>"101000111",
  38707=>"110110110",
  38708=>"000000001",
  38709=>"111011111",
  38710=>"110110100",
  38711=>"001011011",
  38712=>"111110100",
  38713=>"011000010",
  38714=>"010110011",
  38715=>"110100000",
  38716=>"010010111",
  38717=>"011011011",
  38718=>"000100000",
  38719=>"101001001",
  38720=>"110100100",
  38721=>"001101001",
  38722=>"100011111",
  38723=>"100111101",
  38724=>"000000001",
  38725=>"011000001",
  38726=>"100001000",
  38727=>"100100001",
  38728=>"000001111",
  38729=>"010000000",
  38730=>"000000111",
  38731=>"001001000",
  38732=>"001001101",
  38733=>"010110101",
  38734=>"011011010",
  38735=>"111110000",
  38736=>"110101000",
  38737=>"111110100",
  38738=>"000000110",
  38739=>"101100000",
  38740=>"100101001",
  38741=>"000011010",
  38742=>"000010000",
  38743=>"100000100",
  38744=>"110110110",
  38745=>"000010101",
  38746=>"100010001",
  38747=>"001111100",
  38748=>"100100100",
  38749=>"000100101",
  38750=>"001011001",
  38751=>"000011110",
  38752=>"110110000",
  38753=>"100011011",
  38754=>"110100100",
  38755=>"100000100",
  38756=>"001011011",
  38757=>"010010001",
  38758=>"001000000",
  38759=>"001011010",
  38760=>"000011011",
  38761=>"111110110",
  38762=>"111010110",
  38763=>"011000100",
  38764=>"000101000",
  38765=>"110100001",
  38766=>"001100110",
  38767=>"011000110",
  38768=>"000001001",
  38769=>"011111011",
  38770=>"100100000",
  38771=>"000100001",
  38772=>"111000100",
  38773=>"110100100",
  38774=>"000101111",
  38775=>"001001011",
  38776=>"110100110",
  38777=>"001100100",
  38778=>"110000110",
  38779=>"111011011",
  38780=>"010001011",
  38781=>"011010110",
  38782=>"011011011",
  38783=>"101100000",
  38784=>"001011101",
  38785=>"011110110",
  38786=>"100100001",
  38787=>"001000100",
  38788=>"100100101",
  38789=>"111111111",
  38790=>"100100000",
  38791=>"100010000",
  38792=>"011011101",
  38793=>"100111010",
  38794=>"010110000",
  38795=>"111001000",
  38796=>"100101001",
  38797=>"111100001",
  38798=>"001010001",
  38799=>"100000000",
  38800=>"111011110",
  38801=>"011000001",
  38802=>"001001000",
  38803=>"001111011",
  38804=>"001111001",
  38805=>"100100100",
  38806=>"000000000",
  38807=>"000000111",
  38808=>"011010010",
  38809=>"000110111",
  38810=>"110110010",
  38811=>"110100000",
  38812=>"000001011",
  38813=>"110111101",
  38814=>"000110111",
  38815=>"011011000",
  38816=>"000010010",
  38817=>"110100110",
  38818=>"011011010",
  38819=>"111111110",
  38820=>"100110010",
  38821=>"111101111",
  38822=>"011011110",
  38823=>"001001001",
  38824=>"101100000",
  38825=>"110110100",
  38826=>"110110100",
  38827=>"100100100",
  38828=>"100100000",
  38829=>"001011011",
  38830=>"110010110",
  38831=>"110000110",
  38832=>"001011010",
  38833=>"110100000",
  38834=>"000010111",
  38835=>"010100111",
  38836=>"101111100",
  38837=>"000000010",
  38838=>"001111110",
  38839=>"001111100",
  38840=>"000001001",
  38841=>"001001000",
  38842=>"111011100",
  38843=>"110110000",
  38844=>"000110111",
  38845=>"110110010",
  38846=>"001010000",
  38847=>"110000100",
  38848=>"110110110",
  38849=>"111100000",
  38850=>"110001011",
  38851=>"000101110",
  38852=>"000001000",
  38853=>"100100000",
  38854=>"011111111",
  38855=>"110101111",
  38856=>"011010011",
  38857=>"000101011",
  38858=>"111101100",
  38859=>"100000000",
  38860=>"001001001",
  38861=>"100000101",
  38862=>"000100100",
  38863=>"111110100",
  38864=>"100111101",
  38865=>"011110110",
  38866=>"010001110",
  38867=>"111111111",
  38868=>"100111000",
  38869=>"100000100",
  38870=>"100110110",
  38871=>"111010110",
  38872=>"001011011",
  38873=>"111011000",
  38874=>"011101000",
  38875=>"110100100",
  38876=>"100111101",
  38877=>"110100100",
  38878=>"111110101",
  38879=>"111011110",
  38880=>"110000010",
  38881=>"110110100",
  38882=>"111011011",
  38883=>"101111011",
  38884=>"110100000",
  38885=>"001011111",
  38886=>"011001011",
  38887=>"000001011",
  38888=>"111111110",
  38889=>"100101100",
  38890=>"000000100",
  38891=>"111100100",
  38892=>"001001011",
  38893=>"000011111",
  38894=>"001000000",
  38895=>"001000100",
  38896=>"001011101",
  38897=>"010110110",
  38898=>"001001110",
  38899=>"011111110",
  38900=>"001011010",
  38901=>"110100000",
  38902=>"101100100",
  38903=>"000000000",
  38904=>"111100111",
  38905=>"000111111",
  38906=>"011110110",
  38907=>"001011111",
  38908=>"100011010",
  38909=>"000111100",
  38910=>"111111011",
  38911=>"100000000",
  38912=>"001100111",
  38913=>"000000000",
  38914=>"000000000",
  38915=>"101101000",
  38916=>"001011111",
  38917=>"110000000",
  38918=>"100010111",
  38919=>"100000000",
  38920=>"010011001",
  38921=>"111000000",
  38922=>"100000111",
  38923=>"000000101",
  38924=>"000000111",
  38925=>"000000000",
  38926=>"010101000",
  38927=>"100111111",
  38928=>"111000000",
  38929=>"000000000",
  38930=>"000101000",
  38931=>"100000000",
  38932=>"110000000",
  38933=>"111000000",
  38934=>"011111111",
  38935=>"000110110",
  38936=>"101000000",
  38937=>"111011111",
  38938=>"111111000",
  38939=>"000000000",
  38940=>"010111111",
  38941=>"000001001",
  38942=>"000000101",
  38943=>"000000001",
  38944=>"000011001",
  38945=>"010000110",
  38946=>"111111111",
  38947=>"000010010",
  38948=>"111010000",
  38949=>"000111111",
  38950=>"111001001",
  38951=>"000000110",
  38952=>"111101001",
  38953=>"111111000",
  38954=>"111110110",
  38955=>"000101000",
  38956=>"111111101",
  38957=>"110110111",
  38958=>"010000101",
  38959=>"000000000",
  38960=>"111111111",
  38961=>"111111110",
  38962=>"000010100",
  38963=>"000000101",
  38964=>"000100000",
  38965=>"100010101",
  38966=>"011100111",
  38967=>"000000111",
  38968=>"000111101",
  38969=>"000000101",
  38970=>"000100110",
  38971=>"100111000",
  38972=>"011010011",
  38973=>"001000010",
  38974=>"000000000",
  38975=>"111011011",
  38976=>"100000101",
  38977=>"000011111",
  38978=>"111000000",
  38979=>"111111001",
  38980=>"010000000",
  38981=>"001000101",
  38982=>"000000111",
  38983=>"011000001",
  38984=>"000100111",
  38985=>"000000101",
  38986=>"000000000",
  38987=>"111010000",
  38988=>"000001111",
  38989=>"111111110",
  38990=>"101110000",
  38991=>"000101100",
  38992=>"111000000",
  38993=>"011000110",
  38994=>"010001001",
  38995=>"001100000",
  38996=>"001000010",
  38997=>"001000111",
  38998=>"001000111",
  38999=>"001101110",
  39000=>"111111001",
  39001=>"000010100",
  39002=>"111110000",
  39003=>"110110001",
  39004=>"000001010",
  39005=>"001111000",
  39006=>"111011010",
  39007=>"111100110",
  39008=>"111111000",
  39009=>"101000000",
  39010=>"111000101",
  39011=>"001001101",
  39012=>"110111001",
  39013=>"000011011",
  39014=>"111100110",
  39015=>"110101111",
  39016=>"010111111",
  39017=>"000011111",
  39018=>"000001000",
  39019=>"010000111",
  39020=>"011111001",
  39021=>"111111000",
  39022=>"000000000",
  39023=>"000101111",
  39024=>"110100000",
  39025=>"000010010",
  39026=>"100100110",
  39027=>"111101000",
  39028=>"000000001",
  39029=>"010000000",
  39030=>"111111001",
  39031=>"111001000",
  39032=>"010100010",
  39033=>"110000101",
  39034=>"111010111",
  39035=>"101101001",
  39036=>"001001000",
  39037=>"100101001",
  39038=>"101111010",
  39039=>"111111011",
  39040=>"000111000",
  39041=>"000000010",
  39042=>"000000011",
  39043=>"001000110",
  39044=>"101000011",
  39045=>"001111011",
  39046=>"100111111",
  39047=>"111000010",
  39048=>"011001000",
  39049=>"110000000",
  39050=>"111010000",
  39051=>"001000000",
  39052=>"111001000",
  39053=>"101110111",
  39054=>"000000110",
  39055=>"001000000",
  39056=>"110100100",
  39057=>"110111001",
  39058=>"001111111",
  39059=>"001000101",
  39060=>"000000010",
  39061=>"111001000",
  39062=>"110110010",
  39063=>"011111000",
  39064=>"001111111",
  39065=>"000100011",
  39066=>"000000111",
  39067=>"111000000",
  39068=>"100000101",
  39069=>"011001001",
  39070=>"101111111",
  39071=>"000001111",
  39072=>"111100110",
  39073=>"010000011",
  39074=>"110000000",
  39075=>"111000000",
  39076=>"010000001",
  39077=>"011111100",
  39078=>"111010101",
  39079=>"010011000",
  39080=>"110000001",
  39081=>"100111111",
  39082=>"011110100",
  39083=>"101000000",
  39084=>"101111010",
  39085=>"111000000",
  39086=>"000110001",
  39087=>"111001000",
  39088=>"001111101",
  39089=>"101110110",
  39090=>"010010010",
  39091=>"000001001",
  39092=>"111111011",
  39093=>"111111000",
  39094=>"100000011",
  39095=>"010110010",
  39096=>"010010011",
  39097=>"000000110",
  39098=>"110000000",
  39099=>"010111111",
  39100=>"100110000",
  39101=>"111101001",
  39102=>"001000000",
  39103=>"000000010",
  39104=>"000001111",
  39105=>"001101111",
  39106=>"110111001",
  39107=>"011000111",
  39108=>"000010110",
  39109=>"000001111",
  39110=>"100111100",
  39111=>"000000101",
  39112=>"011011111",
  39113=>"000001000",
  39114=>"001000011",
  39115=>"111000000",
  39116=>"110000011",
  39117=>"000000000",
  39118=>"011101001",
  39119=>"001000111",
  39120=>"000000000",
  39121=>"110110001",
  39122=>"110000111",
  39123=>"110111110",
  39124=>"101000110",
  39125=>"101001011",
  39126=>"000000101",
  39127=>"111010000",
  39128=>"000111111",
  39129=>"111000101",
  39130=>"111001001",
  39131=>"000000000",
  39132=>"000110110",
  39133=>"111111101",
  39134=>"111111111",
  39135=>"000111100",
  39136=>"000000111",
  39137=>"101000111",
  39138=>"000111111",
  39139=>"111011110",
  39140=>"001001111",
  39141=>"111000011",
  39142=>"111111101",
  39143=>"010110111",
  39144=>"111100001",
  39145=>"000000010",
  39146=>"001000100",
  39147=>"000001000",
  39148=>"111000000",
  39149=>"000011011",
  39150=>"011000000",
  39151=>"010101111",
  39152=>"000000001",
  39153=>"110000001",
  39154=>"010000001",
  39155=>"100000010",
  39156=>"000001110",
  39157=>"111111000",
  39158=>"000000010",
  39159=>"100000000",
  39160=>"000000111",
  39161=>"111111110",
  39162=>"001000110",
  39163=>"000001101",
  39164=>"000010111",
  39165=>"101001011",
  39166=>"110111011",
  39167=>"000000010",
  39168=>"111000101",
  39169=>"101111000",
  39170=>"000000111",
  39171=>"101101001",
  39172=>"011000100",
  39173=>"111100100",
  39174=>"000101111",
  39175=>"111011110",
  39176=>"000000000",
  39177=>"011110000",
  39178=>"011010000",
  39179=>"101010000",
  39180=>"001001111",
  39181=>"100000111",
  39182=>"001001000",
  39183=>"101000001",
  39184=>"000010110",
  39185=>"000000000",
  39186=>"000000010",
  39187=>"000010000",
  39188=>"110010100",
  39189=>"100101111",
  39190=>"100100000",
  39191=>"101111000",
  39192=>"000010011",
  39193=>"100010010",
  39194=>"111011001",
  39195=>"010011100",
  39196=>"111111000",
  39197=>"110110010",
  39198=>"010001000",
  39199=>"000001101",
  39200=>"111001101",
  39201=>"101010101",
  39202=>"110000101",
  39203=>"100111110",
  39204=>"000100100",
  39205=>"000100100",
  39206=>"010000010",
  39207=>"011111000",
  39208=>"111010110",
  39209=>"110110001",
  39210=>"101111110",
  39211=>"010110010",
  39212=>"011011100",
  39213=>"111010010",
  39214=>"101111000",
  39215=>"100110111",
  39216=>"111010000",
  39217=>"000001100",
  39218=>"000010000",
  39219=>"010010000",
  39220=>"101000101",
  39221=>"110000100",
  39222=>"001001000",
  39223=>"100010000",
  39224=>"010100000",
  39225=>"000000000",
  39226=>"000101000",
  39227=>"101111111",
  39228=>"011101101",
  39229=>"101100111",
  39230=>"010000001",
  39231=>"100100100",
  39232=>"111111011",
  39233=>"111000111",
  39234=>"100111111",
  39235=>"111110101",
  39236=>"101101011",
  39237=>"000000111",
  39238=>"001000000",
  39239=>"000111000",
  39240=>"110110001",
  39241=>"010100100",
  39242=>"110100111",
  39243=>"100101101",
  39244=>"011000000",
  39245=>"000101110",
  39246=>"000110001",
  39247=>"111111010",
  39248=>"000001111",
  39249=>"100101111",
  39250=>"111010110",
  39251=>"111100000",
  39252=>"111111100",
  39253=>"000000111",
  39254=>"000001001",
  39255=>"011111111",
  39256=>"000010111",
  39257=>"010111100",
  39258=>"000100100",
  39259=>"000110001",
  39260=>"001011111",
  39261=>"000001000",
  39262=>"100101100",
  39263=>"101001000",
  39264=>"000000000",
  39265=>"010001001",
  39266=>"000000111",
  39267=>"111111001",
  39268=>"110001000",
  39269=>"000001000",
  39270=>"001000000",
  39271=>"101100100",
  39272=>"011000000",
  39273=>"111101011",
  39274=>"010010010",
  39275=>"011101111",
  39276=>"111011011",
  39277=>"101000100",
  39278=>"111111111",
  39279=>"110010010",
  39280=>"001100000",
  39281=>"000010011",
  39282=>"000110100",
  39283=>"000000101",
  39284=>"101111011",
  39285=>"000001000",
  39286=>"110011000",
  39287=>"010100101",
  39288=>"100100000",
  39289=>"111101101",
  39290=>"011011101",
  39291=>"000001011",
  39292=>"110110001",
  39293=>"111100000",
  39294=>"111110101",
  39295=>"111000111",
  39296=>"011000000",
  39297=>"000001001",
  39298=>"000001001",
  39299=>"101101101",
  39300=>"000010111",
  39301=>"101100110",
  39302=>"101001001",
  39303=>"100011110",
  39304=>"000101000",
  39305=>"000000000",
  39306=>"100100100",
  39307=>"001111111",
  39308=>"111000100",
  39309=>"000001011",
  39310=>"111111101",
  39311=>"000001000",
  39312=>"111110000",
  39313=>"101000111",
  39314=>"100000001",
  39315=>"111000110",
  39316=>"111011000",
  39317=>"000010010",
  39318=>"011111110",
  39319=>"001001000",
  39320=>"010010000",
  39321=>"111110101",
  39322=>"010000110",
  39323=>"111001010",
  39324=>"100100010",
  39325=>"001000000",
  39326=>"111010010",
  39327=>"111011000",
  39328=>"100000101",
  39329=>"110010101",
  39330=>"010111101",
  39331=>"101000000",
  39332=>"011111110",
  39333=>"000000111",
  39334=>"000100111",
  39335=>"000111010",
  39336=>"001010010",
  39337=>"100111000",
  39338=>"111000111",
  39339=>"000001000",
  39340=>"011111111",
  39341=>"000100101",
  39342=>"011100101",
  39343=>"010110111",
  39344=>"101000111",
  39345=>"001011001",
  39346=>"101101000",
  39347=>"100100001",
  39348=>"110000111",
  39349=>"001101000",
  39350=>"000100100",
  39351=>"010111001",
  39352=>"000001101",
  39353=>"111110001",
  39354=>"001000010",
  39355=>"010010000",
  39356=>"000100111",
  39357=>"110000000",
  39358=>"001000101",
  39359=>"010010111",
  39360=>"000101100",
  39361=>"000000001",
  39362=>"100100000",
  39363=>"100000100",
  39364=>"000100101",
  39365=>"111110111",
  39366=>"111011101",
  39367=>"100101100",
  39368=>"000000011",
  39369=>"111101101",
  39370=>"111101011",
  39371=>"001000000",
  39372=>"000000000",
  39373=>"011001100",
  39374=>"010111111",
  39375=>"111110111",
  39376=>"000101111",
  39377=>"101110101",
  39378=>"100010010",
  39379=>"100100101",
  39380=>"011011111",
  39381=>"000110001",
  39382=>"011011101",
  39383=>"001011010",
  39384=>"101001011",
  39385=>"010011000",
  39386=>"011111100",
  39387=>"111000111",
  39388=>"011001100",
  39389=>"111101111",
  39390=>"000010000",
  39391=>"001110110",
  39392=>"001101111",
  39393=>"010000101",
  39394=>"111001111",
  39395=>"100100000",
  39396=>"010000000",
  39397=>"111101000",
  39398=>"000011000",
  39399=>"110110111",
  39400=>"100000011",
  39401=>"001011111",
  39402=>"110000111",
  39403=>"010110100",
  39404=>"000000110",
  39405=>"000100111",
  39406=>"000000000",
  39407=>"011000000",
  39408=>"000000000",
  39409=>"111111111",
  39410=>"111011101",
  39411=>"011001000",
  39412=>"101001100",
  39413=>"001111110",
  39414=>"000001011",
  39415=>"111011000",
  39416=>"010010000",
  39417=>"011001000",
  39418=>"101001111",
  39419=>"110111001",
  39420=>"000000000",
  39421=>"111110000",
  39422=>"010001001",
  39423=>"011001001",
  39424=>"111011100",
  39425=>"000100111",
  39426=>"101000000",
  39427=>"000000000",
  39428=>"000101011",
  39429=>"110000101",
  39430=>"111101111",
  39431=>"011010111",
  39432=>"111101011",
  39433=>"000000000",
  39434=>"000000001",
  39435=>"111111000",
  39436=>"000000000",
  39437=>"111100000",
  39438=>"110100111",
  39439=>"010000111",
  39440=>"011000111",
  39441=>"010000111",
  39442=>"000111111",
  39443=>"010000000",
  39444=>"110010110",
  39445=>"101000000",
  39446=>"000000010",
  39447=>"000100010",
  39448=>"111000001",
  39449=>"110111101",
  39450=>"110101111",
  39451=>"000011011",
  39452=>"111111101",
  39453=>"000101111",
  39454=>"101100000",
  39455=>"000000111",
  39456=>"001111100",
  39457=>"110010111",
  39458=>"000000100",
  39459=>"000000110",
  39460=>"000000100",
  39461=>"011001100",
  39462=>"011001101",
  39463=>"011111000",
  39464=>"111000111",
  39465=>"111000000",
  39466=>"010110010",
  39467=>"010111111",
  39468=>"011000101",
  39469=>"001101101",
  39470=>"001000000",
  39471=>"010000011",
  39472=>"111101011",
  39473=>"100100110",
  39474=>"110010010",
  39475=>"000111110",
  39476=>"000000000",
  39477=>"111111001",
  39478=>"100100011",
  39479=>"000010010",
  39480=>"111110010",
  39481=>"000010000",
  39482=>"010010100",
  39483=>"001100111",
  39484=>"110011011",
  39485=>"111111110",
  39486=>"110100100",
  39487=>"111001001",
  39488=>"111101000",
  39489=>"001000000",
  39490=>"000000010",
  39491=>"101100111",
  39492=>"010111010",
  39493=>"000010010",
  39494=>"010100101",
  39495=>"111000111",
  39496=>"100000011",
  39497=>"111000001",
  39498=>"000001000",
  39499=>"111000000",
  39500=>"100110100",
  39501=>"100111011",
  39502=>"000011011",
  39503=>"100111000",
  39504=>"000000000",
  39505=>"111011100",
  39506=>"111111000",
  39507=>"011011001",
  39508=>"101000010",
  39509=>"100100100",
  39510=>"000000011",
  39511=>"111000101",
  39512=>"111101001",
  39513=>"000001001",
  39514=>"100110111",
  39515=>"011110010",
  39516=>"000111000",
  39517=>"010000001",
  39518=>"011010011",
  39519=>"001000101",
  39520=>"111110111",
  39521=>"000000001",
  39522=>"111000000",
  39523=>"000010000",
  39524=>"000101010",
  39525=>"011111100",
  39526=>"100000000",
  39527=>"010011101",
  39528=>"101010110",
  39529=>"010000000",
  39530=>"110100000",
  39531=>"000001110",
  39532=>"000000100",
  39533=>"000111010",
  39534=>"000000001",
  39535=>"101001101",
  39536=>"010000001",
  39537=>"000000000",
  39538=>"001001111",
  39539=>"010000000",
  39540=>"111000011",
  39541=>"001000101",
  39542=>"000111010",
  39543=>"111000001",
  39544=>"001000001",
  39545=>"000111111",
  39546=>"000100010",
  39547=>"000000000",
  39548=>"100011011",
  39549=>"110100100",
  39550=>"000000000",
  39551=>"101101111",
  39552=>"010011000",
  39553=>"111000000",
  39554=>"111101000",
  39555=>"000000000",
  39556=>"010000000",
  39557=>"110110000",
  39558=>"100101001",
  39559=>"001100110",
  39560=>"000000100",
  39561=>"100111011",
  39562=>"011111010",
  39563=>"000000100",
  39564=>"111101101",
  39565=>"010111100",
  39566=>"000010110",
  39567=>"000000101",
  39568=>"000100011",
  39569=>"111100101",
  39570=>"110110000",
  39571=>"110111111",
  39572=>"000010101",
  39573=>"000000000",
  39574=>"000000111",
  39575=>"100100110",
  39576=>"000010011",
  39577=>"001001001",
  39578=>"000111000",
  39579=>"000000000",
  39580=>"000100101",
  39581=>"111011001",
  39582=>"111111101",
  39583=>"000000000",
  39584=>"000000111",
  39585=>"001000000",
  39586=>"000100011",
  39587=>"001000000",
  39588=>"100111111",
  39589=>"110110110",
  39590=>"001101111",
  39591=>"000110111",
  39592=>"111010000",
  39593=>"000010110",
  39594=>"101000101",
  39595=>"110000010",
  39596=>"001111111",
  39597=>"111001000",
  39598=>"000001011",
  39599=>"001111000",
  39600=>"111000001",
  39601=>"100101111",
  39602=>"111011000",
  39603=>"000000000",
  39604=>"000111111",
  39605=>"100101111",
  39606=>"000011111",
  39607=>"010111111",
  39608=>"011110100",
  39609=>"000111011",
  39610=>"010000100",
  39611=>"100010010",
  39612=>"111000111",
  39613=>"111111111",
  39614=>"011101111",
  39615=>"000000000",
  39616=>"000000000",
  39617=>"111101000",
  39618=>"100101111",
  39619=>"001001111",
  39620=>"000011011",
  39621=>"100101111",
  39622=>"000000011",
  39623=>"011000000",
  39624=>"000000101",
  39625=>"000000110",
  39626=>"010111111",
  39627=>"000101111",
  39628=>"000000100",
  39629=>"000110110",
  39630=>"000000000",
  39631=>"010111111",
  39632=>"111111000",
  39633=>"110000110",
  39634=>"010111101",
  39635=>"101111111",
  39636=>"110011010",
  39637=>"001101101",
  39638=>"001000110",
  39639=>"111100111",
  39640=>"010111010",
  39641=>"000011010",
  39642=>"011001010",
  39643=>"001000100",
  39644=>"001000011",
  39645=>"111111100",
  39646=>"000010000",
  39647=>"101100011",
  39648=>"000000011",
  39649=>"111000000",
  39650=>"111101100",
  39651=>"111001011",
  39652=>"110000000",
  39653=>"010001101",
  39654=>"000101000",
  39655=>"000101110",
  39656=>"111110000",
  39657=>"111111100",
  39658=>"000000100",
  39659=>"000000111",
  39660=>"000011111",
  39661=>"111111000",
  39662=>"100000000",
  39663=>"000000111",
  39664=>"111111010",
  39665=>"001001101",
  39666=>"000111101",
  39667=>"110110111",
  39668=>"110100100",
  39669=>"000001000",
  39670=>"000110000",
  39671=>"000000001",
  39672=>"010010010",
  39673=>"101000000",
  39674=>"111111000",
  39675=>"000111111",
  39676=>"110010010",
  39677=>"011111111",
  39678=>"011110111",
  39679=>"001110101",
  39680=>"000001101",
  39681=>"111100100",
  39682=>"111000000",
  39683=>"001000000",
  39684=>"001010001",
  39685=>"111011010",
  39686=>"010000000",
  39687=>"100100110",
  39688=>"100010111",
  39689=>"000000100",
  39690=>"100100110",
  39691=>"000001100",
  39692=>"100111111",
  39693=>"111000000",
  39694=>"100011000",
  39695=>"010000000",
  39696=>"001010111",
  39697=>"111011001",
  39698=>"010001000",
  39699=>"011111101",
  39700=>"001000011",
  39701=>"100001111",
  39702=>"001011011",
  39703=>"101111010",
  39704=>"111101101",
  39705=>"100001100",
  39706=>"110111111",
  39707=>"111000100",
  39708=>"010111100",
  39709=>"000000000",
  39710=>"011101011",
  39711=>"000000010",
  39712=>"110000000",
  39713=>"111100101",
  39714=>"000000000",
  39715=>"000011011",
  39716=>"000100100",
  39717=>"100100001",
  39718=>"000000110",
  39719=>"000010111",
  39720=>"111001111",
  39721=>"111111101",
  39722=>"000000001",
  39723=>"000111001",
  39724=>"100110110",
  39725=>"000000111",
  39726=>"000100101",
  39727=>"010000000",
  39728=>"000000010",
  39729=>"111001001",
  39730=>"000101110",
  39731=>"111000000",
  39732=>"000101000",
  39733=>"110000001",
  39734=>"000110101",
  39735=>"111001000",
  39736=>"100000000",
  39737=>"111101001",
  39738=>"010111010",
  39739=>"010010111",
  39740=>"101111111",
  39741=>"111011010",
  39742=>"100000100",
  39743=>"110010010",
  39744=>"111100010",
  39745=>"100111010",
  39746=>"100100000",
  39747=>"010110011",
  39748=>"011110111",
  39749=>"111001000",
  39750=>"000010011",
  39751=>"010011000",
  39752=>"100011011",
  39753=>"010010101",
  39754=>"111101101",
  39755=>"111101101",
  39756=>"111101000",
  39757=>"001000000",
  39758=>"100100000",
  39759=>"001001011",
  39760=>"101101101",
  39761=>"011000001",
  39762=>"011010111",
  39763=>"000011001",
  39764=>"000000000",
  39765=>"011110110",
  39766=>"000011011",
  39767=>"000010111",
  39768=>"100100100",
  39769=>"000011001",
  39770=>"110110110",
  39771=>"000011011",
  39772=>"100000101",
  39773=>"110001001",
  39774=>"111100101",
  39775=>"000011111",
  39776=>"000010000",
  39777=>"000001111",
  39778=>"000100100",
  39779=>"101001101",
  39780=>"111101001",
  39781=>"011011010",
  39782=>"000010111",
  39783=>"111000000",
  39784=>"111110001",
  39785=>"111100010",
  39786=>"101100010",
  39787=>"111111111",
  39788=>"010001000",
  39789=>"000000000",
  39790=>"111100000",
  39791=>"101101111",
  39792=>"100001100",
  39793=>"111100110",
  39794=>"000001101",
  39795=>"000010011",
  39796=>"001111010",
  39797=>"111000100",
  39798=>"111100100",
  39799=>"110100100",
  39800=>"000000000",
  39801=>"010111111",
  39802=>"010000100",
  39803=>"100001001",
  39804=>"010111010",
  39805=>"110110100",
  39806=>"101000000",
  39807=>"010010010",
  39808=>"010010010",
  39809=>"010110010",
  39810=>"000000000",
  39811=>"000111111",
  39812=>"000000000",
  39813=>"000111110",
  39814=>"001011011",
  39815=>"000001001",
  39816=>"111110110",
  39817=>"101100100",
  39818=>"101001111",
  39819=>"010011010",
  39820=>"111000000",
  39821=>"000000000",
  39822=>"111000000",
  39823=>"100000000",
  39824=>"101100101",
  39825=>"010001000",
  39826=>"111000000",
  39827=>"100000000",
  39828=>"000011010",
  39829=>"110111111",
  39830=>"111101101",
  39831=>"001101000",
  39832=>"000000000",
  39833=>"101100000",
  39834=>"000000010",
  39835=>"000000000",
  39836=>"000110101",
  39837=>"111100000",
  39838=>"111111000",
  39839=>"000010011",
  39840=>"011111011",
  39841=>"111011110",
  39842=>"000111101",
  39843=>"011110000",
  39844=>"001100101",
  39845=>"100110110",
  39846=>"000110110",
  39847=>"111000000",
  39848=>"000111000",
  39849=>"100101111",
  39850=>"111110100",
  39851=>"111000000",
  39852=>"011010010",
  39853=>"111100000",
  39854=>"110110111",
  39855=>"000000100",
  39856=>"111101000",
  39857=>"011000100",
  39858=>"101101101",
  39859=>"000110110",
  39860=>"011011011",
  39861=>"000000100",
  39862=>"000000100",
  39863=>"100000000",
  39864=>"100000111",
  39865=>"100110010",
  39866=>"101110100",
  39867=>"111111001",
  39868=>"000010111",
  39869=>"110000000",
  39870=>"001000000",
  39871=>"000101011",
  39872=>"000000000",
  39873=>"101101000",
  39874=>"111000000",
  39875=>"001110010",
  39876=>"000000011",
  39877=>"100100000",
  39878=>"000110011",
  39879=>"000000010",
  39880=>"000111111",
  39881=>"100010010",
  39882=>"101101001",
  39883=>"111101101",
  39884=>"111100000",
  39885=>"111110110",
  39886=>"001101000",
  39887=>"001000100",
  39888=>"111000000",
  39889=>"110111011",
  39890=>"100100000",
  39891=>"000101001",
  39892=>"010010000",
  39893=>"111001101",
  39894=>"000111111",
  39895=>"110011000",
  39896=>"000011010",
  39897=>"101000011",
  39898=>"111111010",
  39899=>"110010101",
  39900=>"000011111",
  39901=>"000001111",
  39902=>"000000000",
  39903=>"111010010",
  39904=>"101000000",
  39905=>"111100101",
  39906=>"100000000",
  39907=>"000101110",
  39908=>"101100000",
  39909=>"000111000",
  39910=>"000000011",
  39911=>"000010011",
  39912=>"000100110",
  39913=>"000011111",
  39914=>"000001001",
  39915=>"101101000",
  39916=>"111000000",
  39917=>"000100001",
  39918=>"000000001",
  39919=>"100000000",
  39920=>"010011111",
  39921=>"001011001",
  39922=>"000010000",
  39923=>"000110010",
  39924=>"101100000",
  39925=>"101101100",
  39926=>"000000000",
  39927=>"001111001",
  39928=>"000010111",
  39929=>"000111100",
  39930=>"010000001",
  39931=>"000100001",
  39932=>"101100010",
  39933=>"000000000",
  39934=>"000001011",
  39935=>"111000000",
  39936=>"011011101",
  39937=>"111110010",
  39938=>"101000000",
  39939=>"110100000",
  39940=>"000001001",
  39941=>"111111000",
  39942=>"010001011",
  39943=>"110111101",
  39944=>"000110000",
  39945=>"111111111",
  39946=>"000110111",
  39947=>"010111010",
  39948=>"111000101",
  39949=>"000000000",
  39950=>"101011001",
  39951=>"000101000",
  39952=>"000010110",
  39953=>"111000011",
  39954=>"000000000",
  39955=>"011001111",
  39956=>"101011111",
  39957=>"101000000",
  39958=>"000010001",
  39959=>"111000010",
  39960=>"000000000",
  39961=>"100000000",
  39962=>"000010111",
  39963=>"000110111",
  39964=>"111001110",
  39965=>"010010001",
  39966=>"111111000",
  39967=>"000000000",
  39968=>"100111111",
  39969=>"010010010",
  39970=>"001000000",
  39971=>"000111111",
  39972=>"001111011",
  39973=>"101100100",
  39974=>"001101101",
  39975=>"111101111",
  39976=>"111111111",
  39977=>"000010110",
  39978=>"001101001",
  39979=>"010000000",
  39980=>"010000100",
  39981=>"000001000",
  39982=>"111101111",
  39983=>"110110000",
  39984=>"111010010",
  39985=>"011111011",
  39986=>"010000000",
  39987=>"100001101",
  39988=>"110111111",
  39989=>"101110111",
  39990=>"110110011",
  39991=>"000010000",
  39992=>"010000000",
  39993=>"111111111",
  39994=>"101000000",
  39995=>"111100101",
  39996=>"100110100",
  39997=>"111001000",
  39998=>"000000111",
  39999=>"000011011",
  40000=>"111111111",
  40001=>"101111000",
  40002=>"111101110",
  40003=>"001111011",
  40004=>"000101001",
  40005=>"000001000",
  40006=>"000011110",
  40007=>"000000000",
  40008=>"000000000",
  40009=>"000000000",
  40010=>"111101001",
  40011=>"111111111",
  40012=>"110000000",
  40013=>"000011001",
  40014=>"001100110",
  40015=>"001000000",
  40016=>"000000101",
  40017=>"111000000",
  40018=>"000000101",
  40019=>"011001100",
  40020=>"011111000",
  40021=>"011100111",
  40022=>"000100100",
  40023=>"000000000",
  40024=>"100101000",
  40025=>"110100100",
  40026=>"000100100",
  40027=>"101100101",
  40028=>"110111000",
  40029=>"001001001",
  40030=>"110111111",
  40031=>"100110111",
  40032=>"000100000",
  40033=>"000111111",
  40034=>"111101000",
  40035=>"000111101",
  40036=>"101110101",
  40037=>"001001011",
  40038=>"000000000",
  40039=>"000010000",
  40040=>"010111111",
  40041=>"000000010",
  40042=>"010110000",
  40043=>"100000000",
  40044=>"111000111",
  40045=>"111111111",
  40046=>"000000000",
  40047=>"101000000",
  40048=>"000110100",
  40049=>"110100111",
  40050=>"011011110",
  40051=>"000101111",
  40052=>"011111111",
  40053=>"111000000",
  40054=>"000011111",
  40055=>"111001000",
  40056=>"100010010",
  40057=>"111011000",
  40058=>"011001011",
  40059=>"100000000",
  40060=>"001110110",
  40061=>"110100000",
  40062=>"111100001",
  40063=>"000010111",
  40064=>"101001000",
  40065=>"111100000",
  40066=>"011001001",
  40067=>"110010000",
  40068=>"010111101",
  40069=>"000000000",
  40070=>"111001000",
  40071=>"000001001",
  40072=>"000001001",
  40073=>"111001000",
  40074=>"000111111",
  40075=>"000000000",
  40076=>"000110010",
  40077=>"100010111",
  40078=>"101101100",
  40079=>"101001000",
  40080=>"001100101",
  40081=>"001100101",
  40082=>"111111011",
  40083=>"000001010",
  40084=>"000011111",
  40085=>"111010010",
  40086=>"100111010",
  40087=>"010011001",
  40088=>"111111110",
  40089=>"000000001",
  40090=>"111001000",
  40091=>"100000110",
  40092=>"001001110",
  40093=>"101111101",
  40094=>"101000010",
  40095=>"000000000",
  40096=>"011000000",
  40097=>"011010010",
  40098=>"111000000",
  40099=>"000000000",
  40100=>"001101111",
  40101=>"111001100",
  40102=>"010000101",
  40103=>"000010110",
  40104=>"111111000",
  40105=>"000000000",
  40106=>"011011101",
  40107=>"000100000",
  40108=>"000010100",
  40109=>"000111001",
  40110=>"110110101",
  40111=>"111101001",
  40112=>"000111000",
  40113=>"000000000",
  40114=>"001111000",
  40115=>"000100100",
  40116=>"001100001",
  40117=>"111000101",
  40118=>"000001000",
  40119=>"000010110",
  40120=>"000001011",
  40121=>"000100110",
  40122=>"000000000",
  40123=>"110000010",
  40124=>"010111000",
  40125=>"111110110",
  40126=>"100100111",
  40127=>"000000000",
  40128=>"000000000",
  40129=>"111000000",
  40130=>"111000000",
  40131=>"001011101",
  40132=>"001001000",
  40133=>"100001000",
  40134=>"000000011",
  40135=>"010111000",
  40136=>"000110011",
  40137=>"000000001",
  40138=>"000000000",
  40139=>"111010000",
  40140=>"000000010",
  40141=>"000011011",
  40142=>"000010010",
  40143=>"100101011",
  40144=>"000010010",
  40145=>"000110100",
  40146=>"000000010",
  40147=>"100011010",
  40148=>"101000000",
  40149=>"000110000",
  40150=>"000110110",
  40151=>"111100000",
  40152=>"111000000",
  40153=>"000000101",
  40154=>"100000000",
  40155=>"011000000",
  40156=>"100001110",
  40157=>"000000000",
  40158=>"111000000",
  40159=>"000010110",
  40160=>"000000000",
  40161=>"101000000",
  40162=>"000100100",
  40163=>"001111111",
  40164=>"000000110",
  40165=>"000111111",
  40166=>"111001111",
  40167=>"111101111",
  40168=>"010000000",
  40169=>"000010001",
  40170=>"011111111",
  40171=>"000101110",
  40172=>"100000111",
  40173=>"000110000",
  40174=>"010000000",
  40175=>"010001101",
  40176=>"111111111",
  40177=>"101111100",
  40178=>"111000000",
  40179=>"000001001",
  40180=>"000100011",
  40181=>"000001101",
  40182=>"000010000",
  40183=>"010000000",
  40184=>"111000000",
  40185=>"001011111",
  40186=>"110010000",
  40187=>"100111011",
  40188=>"001001101",
  40189=>"010011111",
  40190=>"110110100",
  40191=>"111001000",
  40192=>"110001001",
  40193=>"101111111",
  40194=>"101000111",
  40195=>"110000000",
  40196=>"100010011",
  40197=>"000000010",
  40198=>"000011111",
  40199=>"110011001",
  40200=>"000001001",
  40201=>"000000000",
  40202=>"010010110",
  40203=>"000110010",
  40204=>"000000010",
  40205=>"010000000",
  40206=>"001011110",
  40207=>"011001000",
  40208=>"111111111",
  40209=>"111000111",
  40210=>"111101000",
  40211=>"111011000",
  40212=>"000110111",
  40213=>"111001001",
  40214=>"011000001",
  40215=>"111111100",
  40216=>"001001101",
  40217=>"001010111",
  40218=>"000100101",
  40219=>"000011111",
  40220=>"000100010",
  40221=>"000111111",
  40222=>"100000110",
  40223=>"011101101",
  40224=>"001000111",
  40225=>"000110111",
  40226=>"111111101",
  40227=>"111111000",
  40228=>"000011011",
  40229=>"101000001",
  40230=>"111010110",
  40231=>"000000000",
  40232=>"111111111",
  40233=>"111111101",
  40234=>"001000000",
  40235=>"010010010",
  40236=>"000100011",
  40237=>"011111111",
  40238=>"100000000",
  40239=>"001110101",
  40240=>"110000111",
  40241=>"110001001",
  40242=>"000010001",
  40243=>"101100110",
  40244=>"000000000",
  40245=>"110111101",
  40246=>"110100001",
  40247=>"111111101",
  40248=>"010010110",
  40249=>"101001101",
  40250=>"100111111",
  40251=>"111001101",
  40252=>"010100011",
  40253=>"010000111",
  40254=>"000000111",
  40255=>"111001100",
  40256=>"101101101",
  40257=>"100000000",
  40258=>"000000000",
  40259=>"001100011",
  40260=>"000000000",
  40261=>"111011101",
  40262=>"000010110",
  40263=>"011000101",
  40264=>"111100001",
  40265=>"000111111",
  40266=>"111101101",
  40267=>"000000000",
  40268=>"111101100",
  40269=>"000110110",
  40270=>"101010000",
  40271=>"010110111",
  40272=>"000000111",
  40273=>"010010110",
  40274=>"000000111",
  40275=>"000001001",
  40276=>"100000010",
  40277=>"001110111",
  40278=>"001100100",
  40279=>"111111111",
  40280=>"111001111",
  40281=>"001111010",
  40282=>"111100000",
  40283=>"000000100",
  40284=>"010000000",
  40285=>"001100101",
  40286=>"000101000",
  40287=>"000000100",
  40288=>"101001000",
  40289=>"000010010",
  40290=>"000000000",
  40291=>"111001001",
  40292=>"010100111",
  40293=>"000000001",
  40294=>"000110111",
  40295=>"111001001",
  40296=>"010000000",
  40297=>"000111111",
  40298=>"111111101",
  40299=>"011000000",
  40300=>"000000000",
  40301=>"110111111",
  40302=>"111010010",
  40303=>"000111111",
  40304=>"100100110",
  40305=>"000101010",
  40306=>"011000000",
  40307=>"111000000",
  40308=>"111111101",
  40309=>"000000001",
  40310=>"000110111",
  40311=>"101111001",
  40312=>"010011101",
  40313=>"010111001",
  40314=>"000000001",
  40315=>"010010111",
  40316=>"101100100",
  40317=>"011001010",
  40318=>"000000111",
  40319=>"000000111",
  40320=>"110000000",
  40321=>"111110110",
  40322=>"011110000",
  40323=>"001000110",
  40324=>"010011000",
  40325=>"111101101",
  40326=>"111000000",
  40327=>"001000000",
  40328=>"011001011",
  40329=>"100001110",
  40330=>"011010111",
  40331=>"111010011",
  40332=>"010111111",
  40333=>"001010111",
  40334=>"111111001",
  40335=>"000001000",
  40336=>"110100100",
  40337=>"110001101",
  40338=>"011101010",
  40339=>"000000000",
  40340=>"000000010",
  40341=>"101000111",
  40342=>"010001000",
  40343=>"011111100",
  40344=>"101011001",
  40345=>"000010010",
  40346=>"110000000",
  40347=>"000000000",
  40348=>"000000111",
  40349=>"001001010",
  40350=>"110000000",
  40351=>"111000000",
  40352=>"111111100",
  40353=>"100100000",
  40354=>"001010011",
  40355=>"101011000",
  40356=>"000000000",
  40357=>"110100000",
  40358=>"111111001",
  40359=>"001000111",
  40360=>"000000000",
  40361=>"111111101",
  40362=>"001000000",
  40363=>"000000010",
  40364=>"011111010",
  40365=>"000010111",
  40366=>"000001000",
  40367=>"111000010",
  40368=>"111001000",
  40369=>"001101001",
  40370=>"000000010",
  40371=>"000101110",
  40372=>"010010010",
  40373=>"010000000",
  40374=>"111111100",
  40375=>"000000000",
  40376=>"011001010",
  40377=>"101100001",
  40378=>"000000111",
  40379=>"011000101",
  40380=>"010000011",
  40381=>"011111111",
  40382=>"111100000",
  40383=>"000010011",
  40384=>"000000000",
  40385=>"100000000",
  40386=>"001011000",
  40387=>"100011011",
  40388=>"000000000",
  40389=>"000111010",
  40390=>"000000000",
  40391=>"111000000",
  40392=>"001110111",
  40393=>"111101000",
  40394=>"101011101",
  40395=>"111101001",
  40396=>"011100100",
  40397=>"001001000",
  40398=>"010101101",
  40399=>"111000000",
  40400=>"111011000",
  40401=>"111001001",
  40402=>"001000101",
  40403=>"011111101",
  40404=>"000000000",
  40405=>"111111111",
  40406=>"100010000",
  40407=>"111111101",
  40408=>"111110100",
  40409=>"000101101",
  40410=>"100101000",
  40411=>"000100000",
  40412=>"000001001",
  40413=>"111000000",
  40414=>"011000000",
  40415=>"011000000",
  40416=>"000000111",
  40417=>"100110111",
  40418=>"111011011",
  40419=>"110110111",
  40420=>"001101100",
  40421=>"000011011",
  40422=>"000000000",
  40423=>"111111000",
  40424=>"000000110",
  40425=>"010000100",
  40426=>"000010111",
  40427=>"101000000",
  40428=>"000010111",
  40429=>"111010000",
  40430=>"000000010",
  40431=>"111110100",
  40432=>"111101100",
  40433=>"000110111",
  40434=>"111011101",
  40435=>"100100100",
  40436=>"101110101",
  40437=>"001101111",
  40438=>"000101000",
  40439=>"000000000",
  40440=>"000000110",
  40441=>"111010000",
  40442=>"000110000",
  40443=>"101001011",
  40444=>"111101100",
  40445=>"000111010",
  40446=>"001110110",
  40447=>"000111111",
  40448=>"000100100",
  40449=>"010000010",
  40450=>"010100100",
  40451=>"100110010",
  40452=>"011111000",
  40453=>"000100111",
  40454=>"101000010",
  40455=>"111000101",
  40456=>"010000000",
  40457=>"000000000",
  40458=>"100110001",
  40459=>"000100000",
  40460=>"000000000",
  40461=>"001010111",
  40462=>"111100001",
  40463=>"111101000",
  40464=>"101101000",
  40465=>"000000000",
  40466=>"101101101",
  40467=>"110110001",
  40468=>"111000010",
  40469=>"011111111",
  40470=>"101100101",
  40471=>"101101101",
  40472=>"000001000",
  40473=>"001000000",
  40474=>"111010000",
  40475=>"100000000",
  40476=>"001101111",
  40477=>"000011111",
  40478=>"000000000",
  40479=>"111000111",
  40480=>"000100101",
  40481=>"111011000",
  40482=>"100100111",
  40483=>"000000100",
  40484=>"111101100",
  40485=>"000001110",
  40486=>"000000111",
  40487=>"110101111",
  40488=>"111111111",
  40489=>"100101101",
  40490=>"001101101",
  40491=>"000001000",
  40492=>"000101100",
  40493=>"100110110",
  40494=>"010010011",
  40495=>"000001000",
  40496=>"011111010",
  40497=>"111100000",
  40498=>"100000110",
  40499=>"111111101",
  40500=>"000100100",
  40501=>"111101001",
  40502=>"000000101",
  40503=>"010010011",
  40504=>"111010001",
  40505=>"110110110",
  40506=>"100101101",
  40507=>"001011101",
  40508=>"110111111",
  40509=>"111111110",
  40510=>"000000000",
  40511=>"011011000",
  40512=>"000000001",
  40513=>"010000100",
  40514=>"111111011",
  40515=>"110100000",
  40516=>"010010111",
  40517=>"000000000",
  40518=>"010110100",
  40519=>"000100010",
  40520=>"011011000",
  40521=>"010001001",
  40522=>"001000010",
  40523=>"101111000",
  40524=>"111110001",
  40525=>"111001001",
  40526=>"110111000",
  40527=>"011010001",
  40528=>"000000111",
  40529=>"011000010",
  40530=>"010111111",
  40531=>"100100100",
  40532=>"010000000",
  40533=>"100011010",
  40534=>"101101100",
  40535=>"001000110",
  40536=>"000000110",
  40537=>"001001000",
  40538=>"100000000",
  40539=>"110100011",
  40540=>"000110010",
  40541=>"011111101",
  40542=>"010010010",
  40543=>"011010100",
  40544=>"000000000",
  40545=>"001000010",
  40546=>"000101000",
  40547=>"001001000",
  40548=>"110111110",
  40549=>"111001011",
  40550=>"010001100",
  40551=>"010000100",
  40552=>"111011111",
  40553=>"101000101",
  40554=>"011011000",
  40555=>"110001101",
  40556=>"101000011",
  40557=>"101111111",
  40558=>"000100000",
  40559=>"010100000",
  40560=>"111001001",
  40561=>"111100000",
  40562=>"000000110",
  40563=>"001101111",
  40564=>"001011111",
  40565=>"000101111",
  40566=>"000001000",
  40567=>"000010100",
  40568=>"000000001",
  40569=>"001101101",
  40570=>"011111101",
  40571=>"111111000",
  40572=>"000100100",
  40573=>"000001101",
  40574=>"000100001",
  40575=>"010010000",
  40576=>"000000000",
  40577=>"111000000",
  40578=>"000001111",
  40579=>"111111111",
  40580=>"111111011",
  40581=>"101000111",
  40582=>"100100101",
  40583=>"000100000",
  40584=>"010000000",
  40585=>"110111111",
  40586=>"111111000",
  40587=>"001000000",
  40588=>"010000010",
  40589=>"100100000",
  40590=>"110001001",
  40591=>"001101101",
  40592=>"101101101",
  40593=>"101001001",
  40594=>"111101001",
  40595=>"001000000",
  40596=>"111111111",
  40597=>"000000000",
  40598=>"010111111",
  40599=>"011011100",
  40600=>"011101000",
  40601=>"010101111",
  40602=>"000011110",
  40603=>"000011000",
  40604=>"111010010",
  40605=>"001000101",
  40606=>"111101010",
  40607=>"111101000",
  40608=>"011111111",
  40609=>"011001111",
  40610=>"111101101",
  40611=>"111000000",
  40612=>"100110110",
  40613=>"000000001",
  40614=>"000001000",
  40615=>"011011001",
  40616=>"110111011",
  40617=>"010000010",
  40618=>"101101101",
  40619=>"000000000",
  40620=>"111110111",
  40621=>"010000100",
  40622=>"100001111",
  40623=>"110111010",
  40624=>"111110000",
  40625=>"010000011",
  40626=>"101111111",
  40627=>"110001000",
  40628=>"111101001",
  40629=>"000111100",
  40630=>"000000100",
  40631=>"000001001",
  40632=>"111111011",
  40633=>"011011110",
  40634=>"000101001",
  40635=>"001110010",
  40636=>"000101101",
  40637=>"101100000",
  40638=>"011110000",
  40639=>"100000010",
  40640=>"111000000",
  40641=>"001101000",
  40642=>"110111111",
  40643=>"111100001",
  40644=>"000000000",
  40645=>"001011110",
  40646=>"111011000",
  40647=>"100000001",
  40648=>"011011010",
  40649=>"010010011",
  40650=>"001000101",
  40651=>"000000001",
  40652=>"010110111",
  40653=>"110000001",
  40654=>"000000000",
  40655=>"000101001",
  40656=>"010010111",
  40657=>"100110011",
  40658=>"100010000",
  40659=>"011111011",
  40660=>"000001000",
  40661=>"101001110",
  40662=>"001000111",
  40663=>"100111010",
  40664=>"001000000",
  40665=>"110010011",
  40666=>"110100101",
  40667=>"101000000",
  40668=>"101101000",
  40669=>"010100010",
  40670=>"000101100",
  40671=>"010110010",
  40672=>"010010000",
  40673=>"000111000",
  40674=>"111101000",
  40675=>"110011011",
  40676=>"100101001",
  40677=>"111001111",
  40678=>"110110101",
  40679=>"011000110",
  40680=>"111111101",
  40681=>"110000000",
  40682=>"001010111",
  40683=>"000001100",
  40684=>"000000000",
  40685=>"111001000",
  40686=>"110100000",
  40687=>"111111100",
  40688=>"000000101",
  40689=>"000100001",
  40690=>"000010010",
  40691=>"001001000",
  40692=>"100001001",
  40693=>"101011010",
  40694=>"000000000",
  40695=>"010000000",
  40696=>"001000000",
  40697=>"111001111",
  40698=>"111100100",
  40699=>"100000110",
  40700=>"000011001",
  40701=>"011100000",
  40702=>"110110000",
  40703=>"000101111",
  40704=>"111101111",
  40705=>"100000000",
  40706=>"000110010",
  40707=>"000000000",
  40708=>"001101000",
  40709=>"000100111",
  40710=>"001010000",
  40711=>"111000001",
  40712=>"000000000",
  40713=>"011111000",
  40714=>"000111111",
  40715=>"001001001",
  40716=>"111001000",
  40717=>"100000000",
  40718=>"001011110",
  40719=>"010000111",
  40720=>"000011101",
  40721=>"000000110",
  40722=>"000000000",
  40723=>"110000111",
  40724=>"110101101",
  40725=>"111001111",
  40726=>"111100000",
  40727=>"000011000",
  40728=>"000010101",
  40729=>"001000001",
  40730=>"100000101",
  40731=>"111111010",
  40732=>"100000110",
  40733=>"010011010",
  40734=>"000100010",
  40735=>"000000000",
  40736=>"111111111",
  40737=>"000000001",
  40738=>"011000001",
  40739=>"100000001",
  40740=>"011110110",
  40741=>"100100111",
  40742=>"001001000",
  40743=>"001111111",
  40744=>"111011101",
  40745=>"111101000",
  40746=>"000000000",
  40747=>"001000100",
  40748=>"000000000",
  40749=>"111000110",
  40750=>"011011000",
  40751=>"001110000",
  40752=>"000000001",
  40753=>"011111011",
  40754=>"000101101",
  40755=>"000111000",
  40756=>"000111111",
  40757=>"110111111",
  40758=>"111111111",
  40759=>"000000000",
  40760=>"010000101",
  40761=>"000000000",
  40762=>"000010111",
  40763=>"100010001",
  40764=>"111100000",
  40765=>"000011011",
  40766=>"110010010",
  40767=>"000000000",
  40768=>"111111110",
  40769=>"000000011",
  40770=>"000100000",
  40771=>"000001111",
  40772=>"000000001",
  40773=>"101101101",
  40774=>"110000110",
  40775=>"110111110",
  40776=>"000000000",
  40777=>"011010000",
  40778=>"000000000",
  40779=>"000000111",
  40780=>"100110111",
  40781=>"100110011",
  40782=>"100111111",
  40783=>"000111111",
  40784=>"000000000",
  40785=>"001010011",
  40786=>"000000110",
  40787=>"011011111",
  40788=>"111111111",
  40789=>"000000000",
  40790=>"100100111",
  40791=>"111111000",
  40792=>"000000000",
  40793=>"010001001",
  40794=>"000000000",
  40795=>"011000100",
  40796=>"001000000",
  40797=>"010010000",
  40798=>"001111011",
  40799=>"110111111",
  40800=>"110000100",
  40801=>"010000000",
  40802=>"111011000",
  40803=>"001000000",
  40804=>"000000000",
  40805=>"000011111",
  40806=>"011111111",
  40807=>"010010010",
  40808=>"000000000",
  40809=>"111100111",
  40810=>"111000000",
  40811=>"100000000",
  40812=>"111111011",
  40813=>"001011111",
  40814=>"111000000",
  40815=>"111000101",
  40816=>"111110011",
  40817=>"000000111",
  40818=>"111111111",
  40819=>"111111111",
  40820=>"101101111",
  40821=>"100100111",
  40822=>"111101000",
  40823=>"111111111",
  40824=>"010111110",
  40825=>"000000001",
  40826=>"000001111",
  40827=>"101111000",
  40828=>"111111110",
  40829=>"101111110",
  40830=>"111000000",
  40831=>"000111000",
  40832=>"111000111",
  40833=>"000000000",
  40834=>"000000000",
  40835=>"000000000",
  40836=>"111111100",
  40837=>"100011111",
  40838=>"011000010",
  40839=>"110100000",
  40840=>"000101000",
  40841=>"000100000",
  40842=>"111111111",
  40843=>"101000111",
  40844=>"000000111",
  40845=>"000000000",
  40846=>"111111100",
  40847=>"100000101",
  40848=>"111001010",
  40849=>"001000000",
  40850=>"000000000",
  40851=>"000000111",
  40852=>"000100100",
  40853=>"111000000",
  40854=>"000000000",
  40855=>"111110010",
  40856=>"111111101",
  40857=>"000111001",
  40858=>"000011001",
  40859=>"111111000",
  40860=>"101000111",
  40861=>"001000000",
  40862=>"000101101",
  40863=>"000010001",
  40864=>"101100000",
  40865=>"111111101",
  40866=>"001000000",
  40867=>"000000000",
  40868=>"000000010",
  40869=>"110000001",
  40870=>"001000001",
  40871=>"000000000",
  40872=>"000000000",
  40873=>"000101100",
  40874=>"000000000",
  40875=>"110100111",
  40876=>"101101111",
  40877=>"100110000",
  40878=>"011111110",
  40879=>"111111111",
  40880=>"000000000",
  40881=>"000000010",
  40882=>"111011000",
  40883=>"111110100",
  40884=>"011110100",
  40885=>"000010111",
  40886=>"010010000",
  40887=>"101101010",
  40888=>"011001000",
  40889=>"111001011",
  40890=>"111110101",
  40891=>"000000000",
  40892=>"100000011",
  40893=>"000111011",
  40894=>"000000000",
  40895=>"000000100",
  40896=>"010001111",
  40897=>"000000111",
  40898=>"101001000",
  40899=>"100111000",
  40900=>"000111111",
  40901=>"100001000",
  40902=>"011111000",
  40903=>"011010000",
  40904=>"000101101",
  40905=>"111111111",
  40906=>"110101111",
  40907=>"000000100",
  40908=>"111111111",
  40909=>"110111000",
  40910=>"000000000",
  40911=>"111110000",
  40912=>"111111000",
  40913=>"111011000",
  40914=>"100101111",
  40915=>"011011010",
  40916=>"000000001",
  40917=>"111011011",
  40918=>"111111010",
  40919=>"000111011",
  40920=>"000000000",
  40921=>"000111101",
  40922=>"001001000",
  40923=>"010111111",
  40924=>"110100000",
  40925=>"011111111",
  40926=>"111111111",
  40927=>"001000001",
  40928=>"000011010",
  40929=>"111111111",
  40930=>"111111111",
  40931=>"111110111",
  40932=>"010010010",
  40933=>"110100000",
  40934=>"001111110",
  40935=>"100100001",
  40936=>"111101111",
  40937=>"111000000",
  40938=>"111111111",
  40939=>"111111111",
  40940=>"000000000",
  40941=>"101111111",
  40942=>"111000000",
  40943=>"110101111",
  40944=>"001111011",
  40945=>"001000000",
  40946=>"000000100",
  40947=>"001000011",
  40948=>"111101001",
  40949=>"000111111",
  40950=>"011011111",
  40951=>"000000000",
  40952=>"000000000",
  40953=>"111001000",
  40954=>"011110101",
  40955=>"111100010",
  40956=>"000001000",
  40957=>"011100101",
  40958=>"001111110",
  40959=>"111111110",
  40960=>"011001001",
  40961=>"000000111",
  40962=>"110011111",
  40963=>"000001001",
  40964=>"100000000",
  40965=>"000000000",
  40966=>"000001010",
  40967=>"010000011",
  40968=>"100000000",
  40969=>"101101101",
  40970=>"010101001",
  40971=>"000000110",
  40972=>"010010000",
  40973=>"110101100",
  40974=>"000011011",
  40975=>"111111000",
  40976=>"100011111",
  40977=>"001001000",
  40978=>"010011110",
  40979=>"000101111",
  40980=>"000001110",
  40981=>"011000000",
  40982=>"111101101",
  40983=>"111000000",
  40984=>"111011000",
  40985=>"110101010",
  40986=>"111000001",
  40987=>"111000100",
  40988=>"000001010",
  40989=>"000000000",
  40990=>"111000000",
  40991=>"001101000",
  40992=>"110111110",
  40993=>"111111000",
  40994=>"000010000",
  40995=>"000000000",
  40996=>"110011001",
  40997=>"001011111",
  40998=>"010001101",
  40999=>"111110001",
  41000=>"110101010",
  41001=>"010110001",
  41002=>"101110010",
  41003=>"000000011",
  41004=>"001011111",
  41005=>"000000110",
  41006=>"101001001",
  41007=>"001001010",
  41008=>"000000011",
  41009=>"111111100",
  41010=>"000000110",
  41011=>"101000000",
  41012=>"001111111",
  41013=>"101111111",
  41014=>"111000000",
  41015=>"111111001",
  41016=>"101000010",
  41017=>"001001111",
  41018=>"000001000",
  41019=>"110000110",
  41020=>"011111001",
  41021=>"001101001",
  41022=>"111111101",
  41023=>"001011011",
  41024=>"011011111",
  41025=>"000111111",
  41026=>"100110111",
  41027=>"000101111",
  41028=>"010010001",
  41029=>"111111000",
  41030=>"001010111",
  41031=>"111011110",
  41032=>"000000010",
  41033=>"000011110",
  41034=>"011011000",
  41035=>"011001000",
  41036=>"001111111",
  41037=>"011101110",
  41038=>"011111100",
  41039=>"101111111",
  41040=>"101000000",
  41041=>"001000000",
  41042=>"001111111",
  41043=>"011000100",
  41044=>"000001011",
  41045=>"111001100",
  41046=>"000011011",
  41047=>"001000111",
  41048=>"100000001",
  41049=>"110110110",
  41050=>"000110100",
  41051=>"111111111",
  41052=>"111100000",
  41053=>"001001001",
  41054=>"110111011",
  41055=>"001000100",
  41056=>"111111111",
  41057=>"110000100",
  41058=>"110111110",
  41059=>"011111111",
  41060=>"100101100",
  41061=>"000100100",
  41062=>"000111110",
  41063=>"111101001",
  41064=>"000101000",
  41065=>"110000000",
  41066=>"011000111",
  41067=>"000000001",
  41068=>"010001000",
  41069=>"000000011",
  41070=>"000000100",
  41071=>"001001000",
  41072=>"100111101",
  41073=>"111101000",
  41074=>"110100110",
  41075=>"000001111",
  41076=>"100111110",
  41077=>"000000000",
  41078=>"011111111",
  41079=>"111111010",
  41080=>"100000110",
  41081=>"111111111",
  41082=>"010111111",
  41083=>"000000000",
  41084=>"011001010",
  41085=>"100000000",
  41086=>"000000010",
  41087=>"000000000",
  41088=>"111110010",
  41089=>"100010010",
  41090=>"100111000",
  41091=>"001111010",
  41092=>"000000010",
  41093=>"001111001",
  41094=>"000100111",
  41095=>"110100111",
  41096=>"011111100",
  41097=>"000001001",
  41098=>"110010110",
  41099=>"010011001",
  41100=>"111101100",
  41101=>"000010111",
  41102=>"000010010",
  41103=>"010001010",
  41104=>"111101111",
  41105=>"000000111",
  41106=>"100001000",
  41107=>"010001000",
  41108=>"111000000",
  41109=>"101000101",
  41110=>"110111100",
  41111=>"001011001",
  41112=>"111101110",
  41113=>"000110111",
  41114=>"001000001",
  41115=>"000110000",
  41116=>"101000100",
  41117=>"001000000",
  41118=>"100000000",
  41119=>"000001000",
  41120=>"100111000",
  41121=>"101010000",
  41122=>"101111111",
  41123=>"110010110",
  41124=>"111001100",
  41125=>"011111111",
  41126=>"100110110",
  41127=>"011111111",
  41128=>"111000000",
  41129=>"000101111",
  41130=>"001110110",
  41131=>"000000101",
  41132=>"100101011",
  41133=>"101000101",
  41134=>"010001011",
  41135=>"110110111",
  41136=>"000000000",
  41137=>"011011111",
  41138=>"111101101",
  41139=>"000001100",
  41140=>"110100111",
  41141=>"111111111",
  41142=>"000111100",
  41143=>"000010110",
  41144=>"100101101",
  41145=>"111001000",
  41146=>"111111000",
  41147=>"110101111",
  41148=>"000110010",
  41149=>"000010111",
  41150=>"100100000",
  41151=>"100000000",
  41152=>"000000000",
  41153=>"110000110",
  41154=>"000101111",
  41155=>"110100100",
  41156=>"010111010",
  41157=>"111111100",
  41158=>"101000011",
  41159=>"010010000",
  41160=>"000111110",
  41161=>"001101000",
  41162=>"111111101",
  41163=>"111111000",
  41164=>"011101111",
  41165=>"100100111",
  41166=>"111010111",
  41167=>"111011110",
  41168=>"000001101",
  41169=>"010111011",
  41170=>"011111000",
  41171=>"000100000",
  41172=>"010111011",
  41173=>"100000100",
  41174=>"000000110",
  41175=>"111000001",
  41176=>"000000111",
  41177=>"111000000",
  41178=>"111111100",
  41179=>"000000000",
  41180=>"111001011",
  41181=>"001001000",
  41182=>"000101001",
  41183=>"111011001",
  41184=>"110011101",
  41185=>"000000000",
  41186=>"000000001",
  41187=>"000010110",
  41188=>"010100111",
  41189=>"000000000",
  41190=>"001011101",
  41191=>"111001011",
  41192=>"111111000",
  41193=>"010010011",
  41194=>"000100000",
  41195=>"101111110",
  41196=>"001000110",
  41197=>"000000000",
  41198=>"000000000",
  41199=>"000110000",
  41200=>"000000100",
  41201=>"110000000",
  41202=>"111101000",
  41203=>"001000001",
  41204=>"111100100",
  41205=>"001000001",
  41206=>"000010111",
  41207=>"010111101",
  41208=>"110010101",
  41209=>"000000101",
  41210=>"100000000",
  41211=>"111011000",
  41212=>"111010000",
  41213=>"000000011",
  41214=>"100000011",
  41215=>"110110111",
  41216=>"001000010",
  41217=>"111111111",
  41218=>"001011001",
  41219=>"100110110",
  41220=>"001011111",
  41221=>"001011010",
  41222=>"110111100",
  41223=>"000011010",
  41224=>"001001001",
  41225=>"011011001",
  41226=>"000101001",
  41227=>"011011010",
  41228=>"011001001",
  41229=>"110111010",
  41230=>"111000000",
  41231=>"000011000",
  41232=>"000000010",
  41233=>"110011111",
  41234=>"100001110",
  41235=>"010000100",
  41236=>"100010100",
  41237=>"100110000",
  41238=>"010011011",
  41239=>"000001011",
  41240=>"000000000",
  41241=>"000000100",
  41242=>"110010110",
  41243=>"011001011",
  41244=>"000000100",
  41245=>"100100000",
  41246=>"010010011",
  41247=>"000000110",
  41248=>"011011001",
  41249=>"000011011",
  41250=>"001111111",
  41251=>"000001011",
  41252=>"011011010",
  41253=>"000010110",
  41254=>"011110000",
  41255=>"010010011",
  41256=>"001111011",
  41257=>"000100110",
  41258=>"011010011",
  41259=>"100001011",
  41260=>"101100000",
  41261=>"100110111",
  41262=>"110011111",
  41263=>"000100010",
  41264=>"000001000",
  41265=>"000111001",
  41266=>"011010100",
  41267=>"000100100",
  41268=>"000001000",
  41269=>"100100000",
  41270=>"101100000",
  41271=>"110001011",
  41272=>"000010011",
  41273=>"011000110",
  41274=>"100100110",
  41275=>"001000001",
  41276=>"001001011",
  41277=>"000110111",
  41278=>"011011011",
  41279=>"110010001",
  41280=>"011001001",
  41281=>"000011110",
  41282=>"111101110",
  41283=>"011011011",
  41284=>"001100110",
  41285=>"000000010",
  41286=>"011000000",
  41287=>"101101000",
  41288=>"111110101",
  41289=>"110000011",
  41290=>"010010011",
  41291=>"100110000",
  41292=>"111011001",
  41293=>"000011011",
  41294=>"011000000",
  41295=>"011011110",
  41296=>"011010000",
  41297=>"100111111",
  41298=>"111111100",
  41299=>"100111011",
  41300=>"011010110",
  41301=>"000001001",
  41302=>"001011101",
  41303=>"010001011",
  41304=>"001111101",
  41305=>"100110100",
  41306=>"100111111",
  41307=>"111111001",
  41308=>"001001000",
  41309=>"001101101",
  41310=>"111110010",
  41311=>"011011011",
  41312=>"010011011",
  41313=>"010000000",
  41314=>"011001001",
  41315=>"100100010",
  41316=>"011001011",
  41317=>"111100101",
  41318=>"011100000",
  41319=>"100100100",
  41320=>"000101000",
  41321=>"001110100",
  41322=>"110010111",
  41323=>"011110011",
  41324=>"000010000",
  41325=>"100100100",
  41326=>"010001011",
  41327=>"110011010",
  41328=>"011110011",
  41329=>"000001011",
  41330=>"000010010",
  41331=>"000100000",
  41332=>"101111111",
  41333=>"010010010",
  41334=>"011110110",
  41335=>"110000000",
  41336=>"000010011",
  41337=>"100100101",
  41338=>"110011110",
  41339=>"100101001",
  41340=>"111011011",
  41341=>"101000000",
  41342=>"011100001",
  41343=>"111001000",
  41344=>"010011011",
  41345=>"000000001",
  41346=>"100001011",
  41347=>"100100000",
  41348=>"101101100",
  41349=>"110000000",
  41350=>"000000111",
  41351=>"111010000",
  41352=>"001111010",
  41353=>"000100000",
  41354=>"101100101",
  41355=>"101001000",
  41356=>"000000000",
  41357=>"011011011",
  41358=>"110001111",
  41359=>"001001000",
  41360=>"101111110",
  41361=>"011011001",
  41362=>"111011010",
  41363=>"011011011",
  41364=>"101001001",
  41365=>"011001011",
  41366=>"100110100",
  41367=>"001001001",
  41368=>"010010010",
  41369=>"001100100",
  41370=>"011001001",
  41371=>"111111011",
  41372=>"111000111",
  41373=>"011011011",
  41374=>"101011000",
  41375=>"011010010",
  41376=>"111011010",
  41377=>"100100110",
  41378=>"111000000",
  41379=>"000100100",
  41380=>"100110100",
  41381=>"010000000",
  41382=>"001000111",
  41383=>"001011100",
  41384=>"100100111",
  41385=>"011011111",
  41386=>"001011011",
  41387=>"011001001",
  41388=>"000000111",
  41389=>"000001000",
  41390=>"011000010",
  41391=>"100111110",
  41392=>"011001001",
  41393=>"000010110",
  41394=>"100011111",
  41395=>"000001001",
  41396=>"100101101",
  41397=>"100100101",
  41398=>"100010111",
  41399=>"011011011",
  41400=>"010000000",
  41401=>"000000001",
  41402=>"101100110",
  41403=>"111011000",
  41404=>"100110100",
  41405=>"001001111",
  41406=>"000000001",
  41407=>"000100110",
  41408=>"101001011",
  41409=>"100110001",
  41410=>"111011000",
  41411=>"000110001",
  41412=>"000100111",
  41413=>"110011110",
  41414=>"101001001",
  41415=>"100000001",
  41416=>"100010010",
  41417=>"001000010",
  41418=>"110110111",
  41419=>"000000100",
  41420=>"011011000",
  41421=>"011010001",
  41422=>"100100100",
  41423=>"010011001",
  41424=>"111110100",
  41425=>"111110111",
  41426=>"000111110",
  41427=>"111100001",
  41428=>"011011011",
  41429=>"000000000",
  41430=>"011001011",
  41431=>"111110001",
  41432=>"000010110",
  41433=>"110110100",
  41434=>"001001001",
  41435=>"100100100",
  41436=>"111111011",
  41437=>"010100111",
  41438=>"001110110",
  41439=>"110010000",
  41440=>"111111110",
  41441=>"111100111",
  41442=>"101100000",
  41443=>"011011011",
  41444=>"010010000",
  41445=>"000110110",
  41446=>"111001001",
  41447=>"011111011",
  41448=>"011111000",
  41449=>"000000000",
  41450=>"110110000",
  41451=>"001000011",
  41452=>"010011011",
  41453=>"100110110",
  41454=>"000001100",
  41455=>"000001011",
  41456=>"000000000",
  41457=>"000001111",
  41458=>"011001001",
  41459=>"000000000",
  41460=>"001011011",
  41461=>"000100100",
  41462=>"000000000",
  41463=>"010100001",
  41464=>"011011011",
  41465=>"100000000",
  41466=>"111111111",
  41467=>"111100100",
  41468=>"001001001",
  41469=>"000000000",
  41470=>"111000000",
  41471=>"111010011",
  41472=>"001001011",
  41473=>"111111111",
  41474=>"111101111",
  41475=>"101101000",
  41476=>"111111111",
  41477=>"111001110",
  41478=>"011111001",
  41479=>"001010111",
  41480=>"010111111",
  41481=>"001000011",
  41482=>"001100100",
  41483=>"000111001",
  41484=>"011010000",
  41485=>"010111010",
  41486=>"100110110",
  41487=>"110000010",
  41488=>"000001011",
  41489=>"010100111",
  41490=>"111101101",
  41491=>"001001000",
  41492=>"111111111",
  41493=>"101000101",
  41494=>"101100111",
  41495=>"110100100",
  41496=>"101101110",
  41497=>"001111000",
  41498=>"000011010",
  41499=>"000111101",
  41500=>"000000110",
  41501=>"111000000",
  41502=>"100101101",
  41503=>"000111010",
  41504=>"001101111",
  41505=>"111111010",
  41506=>"000100001",
  41507=>"111111010",
  41508=>"101011110",
  41509=>"100100110",
  41510=>"100100011",
  41511=>"000000100",
  41512=>"100111110",
  41513=>"011011111",
  41514=>"001001000",
  41515=>"000000000",
  41516=>"010011001",
  41517=>"110111001",
  41518=>"111101010",
  41519=>"101101110",
  41520=>"100001111",
  41521=>"000111111",
  41522=>"001000010",
  41523=>"100000001",
  41524=>"101000000",
  41525=>"000111111",
  41526=>"000000100",
  41527=>"000000000",
  41528=>"101101111",
  41529=>"000000010",
  41530=>"011010111",
  41531=>"000000101",
  41532=>"010111110",
  41533=>"010111000",
  41534=>"000000000",
  41535=>"110101111",
  41536=>"000100000",
  41537=>"000000110",
  41538=>"101101111",
  41539=>"001000010",
  41540=>"110000110",
  41541=>"001000000",
  41542=>"110010000",
  41543=>"000101000",
  41544=>"111111000",
  41545=>"101111111",
  41546=>"100000101",
  41547=>"101001110",
  41548=>"000000110",
  41549=>"000111111",
  41550=>"001111111",
  41551=>"000011111",
  41552=>"000000111",
  41553=>"110000100",
  41554=>"001101000",
  41555=>"011000000",
  41556=>"101101100",
  41557=>"011011011",
  41558=>"111111111",
  41559=>"000000000",
  41560=>"010110100",
  41561=>"000010100",
  41562=>"100100111",
  41563=>"001010111",
  41564=>"001001111",
  41565=>"000010010",
  41566=>"110011101",
  41567=>"100010111",
  41568=>"000010010",
  41569=>"000111111",
  41570=>"100000111",
  41571=>"001011110",
  41572=>"000111111",
  41573=>"011100000",
  41574=>"110111000",
  41575=>"110000011",
  41576=>"011110000",
  41577=>"110000100",
  41578=>"010000000",
  41579=>"111110000",
  41580=>"110110000",
  41581=>"100100100",
  41582=>"011000110",
  41583=>"000000000",
  41584=>"000111111",
  41585=>"100101100",
  41586=>"000001001",
  41587=>"001000001",
  41588=>"000000000",
  41589=>"111000000",
  41590=>"000000000",
  41591=>"000000101",
  41592=>"101001000",
  41593=>"110111100",
  41594=>"011000001",
  41595=>"001000000",
  41596=>"000011011",
  41597=>"111100010",
  41598=>"111001110",
  41599=>"101000011",
  41600=>"110000000",
  41601=>"111101000",
  41602=>"010010011",
  41603=>"111111000",
  41604=>"001111000",
  41605=>"111000000",
  41606=>"010001011",
  41607=>"000110110",
  41608=>"000110110",
  41609=>"100001101",
  41610=>"111100100",
  41611=>"010010000",
  41612=>"110011001",
  41613=>"000010010",
  41614=>"111110101",
  41615=>"001001001",
  41616=>"110110110",
  41617=>"111111010",
  41618=>"101100110",
  41619=>"100101001",
  41620=>"001101011",
  41621=>"101000101",
  41622=>"000000001",
  41623=>"010111011",
  41624=>"000111101",
  41625=>"101000100",
  41626=>"000111110",
  41627=>"000000010",
  41628=>"010010010",
  41629=>"101101110",
  41630=>"110000100",
  41631=>"111101000",
  41632=>"011101100",
  41633=>"100000001",
  41634=>"111010000",
  41635=>"101101000",
  41636=>"000111100",
  41637=>"110000000",
  41638=>"110000111",
  41639=>"000010010",
  41640=>"010010101",
  41641=>"000001001",
  41642=>"011011111",
  41643=>"101000010",
  41644=>"111110000",
  41645=>"000000110",
  41646=>"000100110",
  41647=>"000010000",
  41648=>"010101101",
  41649=>"011011100",
  41650=>"000111111",
  41651=>"000001011",
  41652=>"011011010",
  41653=>"111100110",
  41654=>"011011000",
  41655=>"111101010",
  41656=>"110111011",
  41657=>"000110011",
  41658=>"111000111",
  41659=>"000111010",
  41660=>"000110000",
  41661=>"010111111",
  41662=>"011001010",
  41663=>"000101111",
  41664=>"000001000",
  41665=>"000100000",
  41666=>"011000010",
  41667=>"100101011",
  41668=>"000000000",
  41669=>"000000000",
  41670=>"111011111",
  41671=>"001000010",
  41672=>"000000111",
  41673=>"001000000",
  41674=>"111000000",
  41675=>"010110111",
  41676=>"000101111",
  41677=>"000110110",
  41678=>"001000000",
  41679=>"010111000",
  41680=>"111111011",
  41681=>"110010110",
  41682=>"000000000",
  41683=>"011000000",
  41684=>"001110110",
  41685=>"111110000",
  41686=>"101100111",
  41687=>"010000000",
  41688=>"111000001",
  41689=>"011010010",
  41690=>"110100001",
  41691=>"101000111",
  41692=>"101001110",
  41693=>"010000000",
  41694=>"111001000",
  41695=>"001100110",
  41696=>"001111111",
  41697=>"101101000",
  41698=>"100001101",
  41699=>"011011011",
  41700=>"101101101",
  41701=>"110110000",
  41702=>"011010000",
  41703=>"000000110",
  41704=>"111000001",
  41705=>"000000101",
  41706=>"100000000",
  41707=>"000000011",
  41708=>"010010001",
  41709=>"001000101",
  41710=>"110001000",
  41711=>"111000000",
  41712=>"000000100",
  41713=>"000000011",
  41714=>"010101001",
  41715=>"110110110",
  41716=>"110110110",
  41717=>"101000101",
  41718=>"000000000",
  41719=>"000001111",
  41720=>"101000101",
  41721=>"010000000",
  41722=>"111111111",
  41723=>"000000000",
  41724=>"010010111",
  41725=>"100010001",
  41726=>"011010110",
  41727=>"000101000",
  41728=>"000000110",
  41729=>"000100010",
  41730=>"000101110",
  41731=>"000000000",
  41732=>"011001111",
  41733=>"101101001",
  41734=>"110110110",
  41735=>"111110000",
  41736=>"000000111",
  41737=>"111000000",
  41738=>"000000110",
  41739=>"000000000",
  41740=>"000000111",
  41741=>"101111001",
  41742=>"000000110",
  41743=>"001000111",
  41744=>"111111000",
  41745=>"111111000",
  41746=>"000111011",
  41747=>"100111110",
  41748=>"000110110",
  41749=>"110111111",
  41750=>"011110111",
  41751=>"110111000",
  41752=>"110000000",
  41753=>"010111000",
  41754=>"111111111",
  41755=>"110010100",
  41756=>"111101111",
  41757=>"000110110",
  41758=>"111111110",
  41759=>"000001101",
  41760=>"000101110",
  41761=>"000100000",
  41762=>"011000000",
  41763=>"000100110",
  41764=>"000010100",
  41765=>"101011110",
  41766=>"000000111",
  41767=>"000111110",
  41768=>"011110000",
  41769=>"011000110",
  41770=>"101101101",
  41771=>"110010000",
  41772=>"000001111",
  41773=>"101110111",
  41774=>"101111110",
  41775=>"010110001",
  41776=>"001001100",
  41777=>"000101111",
  41778=>"111000010",
  41779=>"111000000",
  41780=>"000010111",
  41781=>"010000000",
  41782=>"000100100",
  41783=>"000000000",
  41784=>"111111011",
  41785=>"000001111",
  41786=>"111001000",
  41787=>"111111011",
  41788=>"000111111",
  41789=>"111001000",
  41790=>"001001111",
  41791=>"001110101",
  41792=>"111010110",
  41793=>"101001000",
  41794=>"101000000",
  41795=>"100111011",
  41796=>"000101110",
  41797=>"000001111",
  41798=>"111000101",
  41799=>"001001000",
  41800=>"000110110",
  41801=>"111111000",
  41802=>"001000111",
  41803=>"001101100",
  41804=>"110111111",
  41805=>"011001011",
  41806=>"100010110",
  41807=>"000000110",
  41808=>"001111111",
  41809=>"111111000",
  41810=>"000001110",
  41811=>"000011011",
  41812=>"000000000",
  41813=>"111111111",
  41814=>"000010111",
  41815=>"111110000",
  41816=>"100111110",
  41817=>"110111111",
  41818=>"000100101",
  41819=>"100110111",
  41820=>"001111110",
  41821=>"001101101",
  41822=>"111111111",
  41823=>"011111101",
  41824=>"000110111",
  41825=>"000000000",
  41826=>"000000011",
  41827=>"011011111",
  41828=>"000001001",
  41829=>"111111000",
  41830=>"000110000",
  41831=>"001000000",
  41832=>"111111000",
  41833=>"111111000",
  41834=>"000000011",
  41835=>"001001110",
  41836=>"000111110",
  41837=>"111000000",
  41838=>"000100100",
  41839=>"000000000",
  41840=>"000011011",
  41841=>"111000000",
  41842=>"100010011",
  41843=>"001001111",
  41844=>"100100111",
  41845=>"000001111",
  41846=>"111000000",
  41847=>"000000111",
  41848=>"111101111",
  41849=>"010001111",
  41850=>"000000110",
  41851=>"000100111",
  41852=>"001011011",
  41853=>"000000100",
  41854=>"101111111",
  41855=>"000001111",
  41856=>"001010110",
  41857=>"000010000",
  41858=>"011110111",
  41859=>"111000000",
  41860=>"000000000",
  41861=>"100001000",
  41862=>"100011110",
  41863=>"000000000",
  41864=>"000010000",
  41865=>"000000000",
  41866=>"000000001",
  41867=>"001000100",
  41868=>"110111000",
  41869=>"111111000",
  41870=>"111100101",
  41871=>"000001010",
  41872=>"000000011",
  41873=>"000000110",
  41874=>"111111001",
  41875=>"111010000",
  41876=>"000000000",
  41877=>"111111000",
  41878=>"111111111",
  41879=>"000101101",
  41880=>"000110111",
  41881=>"011111000",
  41882=>"000000010",
  41883=>"111000100",
  41884=>"000001001",
  41885=>"010111001",
  41886=>"001110111",
  41887=>"000000100",
  41888=>"001111110",
  41889=>"111110110",
  41890=>"000001000",
  41891=>"110101000",
  41892=>"111111110",
  41893=>"001011111",
  41894=>"101001111",
  41895=>"001111111",
  41896=>"111111110",
  41897=>"110111111",
  41898=>"111000011",
  41899=>"000000011",
  41900=>"111100001",
  41901=>"000000010",
  41902=>"000101100",
  41903=>"001101111",
  41904=>"000111111",
  41905=>"011001000",
  41906=>"010001111",
  41907=>"010001010",
  41908=>"000111100",
  41909=>"111111111",
  41910=>"000000101",
  41911=>"000001010",
  41912=>"000111111",
  41913=>"001001010",
  41914=>"000001111",
  41915=>"000001111",
  41916=>"111001111",
  41917=>"111110001",
  41918=>"110011011",
  41919=>"111110110",
  41920=>"000111000",
  41921=>"000000100",
  41922=>"111111111",
  41923=>"000001111",
  41924=>"000001111",
  41925=>"000010111",
  41926=>"000110001",
  41927=>"101101110",
  41928=>"010000001",
  41929=>"010101111",
  41930=>"111111100",
  41931=>"000000110",
  41932=>"000111011",
  41933=>"001111100",
  41934=>"110110111",
  41935=>"111110111",
  41936=>"111010011",
  41937=>"000011111",
  41938=>"011000010",
  41939=>"101111101",
  41940=>"000111111",
  41941=>"000001010",
  41942=>"000011111",
  41943=>"111101100",
  41944=>"000100111",
  41945=>"000000111",
  41946=>"001101101",
  41947=>"111000000",
  41948=>"110111111",
  41949=>"000001000",
  41950=>"000101111",
  41951=>"111101111",
  41952=>"111000001",
  41953=>"000000000",
  41954=>"111101011",
  41955=>"001011111",
  41956=>"001001110",
  41957=>"110111011",
  41958=>"111001111",
  41959=>"011111111",
  41960=>"111111111",
  41961=>"000000100",
  41962=>"000000001",
  41963=>"001000000",
  41964=>"000111111",
  41965=>"011101000",
  41966=>"111000000",
  41967=>"000000110",
  41968=>"000000101",
  41969=>"001111111",
  41970=>"000001110",
  41971=>"110111110",
  41972=>"000001011",
  41973=>"001000100",
  41974=>"100000111",
  41975=>"111000010",
  41976=>"111111000",
  41977=>"111111111",
  41978=>"111000010",
  41979=>"000110111",
  41980=>"000010111",
  41981=>"000111000",
  41982=>"000000011",
  41983=>"000000110",
  41984=>"011000101",
  41985=>"000000100",
  41986=>"111101100",
  41987=>"000000010",
  41988=>"001001111",
  41989=>"110101111",
  41990=>"110111101",
  41991=>"000011010",
  41992=>"000110111",
  41993=>"110000000",
  41994=>"001011100",
  41995=>"111001000",
  41996=>"001010011",
  41997=>"000010011",
  41998=>"000000010",
  41999=>"111111011",
  42000=>"000110010",
  42001=>"000000101",
  42002=>"000000000",
  42003=>"111111101",
  42004=>"111110101",
  42005=>"111101001",
  42006=>"100111111",
  42007=>"010010111",
  42008=>"100000111",
  42009=>"000100110",
  42010=>"000000000",
  42011=>"000001010",
  42012=>"100100111",
  42013=>"101000101",
  42014=>"010100101",
  42015=>"000100101",
  42016=>"000000100",
  42017=>"010110010",
  42018=>"000000000",
  42019=>"000111010",
  42020=>"000100110",
  42021=>"111011011",
  42022=>"000011000",
  42023=>"000010000",
  42024=>"111111000",
  42025=>"010010111",
  42026=>"011001000",
  42027=>"101101011",
  42028=>"000011011",
  42029=>"010010101",
  42030=>"010111111",
  42031=>"000110010",
  42032=>"101100110",
  42033=>"001111110",
  42034=>"000000010",
  42035=>"000100100",
  42036=>"000001000",
  42037=>"110110000",
  42038=>"100101001",
  42039=>"001000000",
  42040=>"010111111",
  42041=>"000001000",
  42042=>"011000100",
  42043=>"101101000",
  42044=>"000001101",
  42045=>"000111110",
  42046=>"101101111",
  42047=>"011110100",
  42048=>"101001001",
  42049=>"010000111",
  42050=>"111101001",
  42051=>"001001100",
  42052=>"110110110",
  42053=>"001000000",
  42054=>"000101111",
  42055=>"000010110",
  42056=>"000011110",
  42057=>"111110010",
  42058=>"111111011",
  42059=>"011000100",
  42060=>"000000000",
  42061=>"001101111",
  42062=>"110111111",
  42063=>"111111111",
  42064=>"000000000",
  42065=>"110011110",
  42066=>"010010000",
  42067=>"010011001",
  42068=>"000101101",
  42069=>"000001011",
  42070=>"001111100",
  42071=>"101000100",
  42072=>"110100000",
  42073=>"000011111",
  42074=>"100101110",
  42075=>"000000011",
  42076=>"111101101",
  42077=>"100001011",
  42078=>"111111111",
  42079=>"100001001",
  42080=>"000110011",
  42081=>"001101101",
  42082=>"010101111",
  42083=>"000110100",
  42084=>"000110111",
  42085=>"011011001",
  42086=>"000110100",
  42087=>"111000000",
  42088=>"011100100",
  42089=>"010000110",
  42090=>"010000000",
  42091=>"010110000",
  42092=>"000011010",
  42093=>"100110100",
  42094=>"000001100",
  42095=>"000101000",
  42096=>"101111111",
  42097=>"010010001",
  42098=>"001100100",
  42099=>"000000000",
  42100=>"111111111",
  42101=>"001000000",
  42102=>"000110111",
  42103=>"011000110",
  42104=>"111001111",
  42105=>"000010100",
  42106=>"000000101",
  42107=>"111000000",
  42108=>"001011011",
  42109=>"010100000",
  42110=>"000101011",
  42111=>"001000100",
  42112=>"010010000",
  42113=>"111100000",
  42114=>"010010010",
  42115=>"000010000",
  42116=>"111111000",
  42117=>"000001110",
  42118=>"111100000",
  42119=>"100110110",
  42120=>"111111010",
  42121=>"011000000",
  42122=>"011010111",
  42123=>"010010000",
  42124=>"111000100",
  42125=>"101001000",
  42126=>"111000100",
  42127=>"011001000",
  42128=>"100110110",
  42129=>"001101101",
  42130=>"000000010",
  42131=>"111111111",
  42132=>"101010110",
  42133=>"010000000",
  42134=>"111111100",
  42135=>"000111010",
  42136=>"100010010",
  42137=>"101000110",
  42138=>"011101100",
  42139=>"101101010",
  42140=>"000000000",
  42141=>"100000100",
  42142=>"111010110",
  42143=>"111101000",
  42144=>"101101111",
  42145=>"101100100",
  42146=>"000110000",
  42147=>"010000000",
  42148=>"010100011",
  42149=>"010110000",
  42150=>"000000001",
  42151=>"000010010",
  42152=>"010010110",
  42153=>"011010110",
  42154=>"111111111",
  42155=>"101101000",
  42156=>"000010001",
  42157=>"000000110",
  42158=>"100101011",
  42159=>"010010010",
  42160=>"000100000",
  42161=>"101011011",
  42162=>"001011000",
  42163=>"000001110",
  42164=>"000010011",
  42165=>"010000101",
  42166=>"011011000",
  42167=>"011001000",
  42168=>"000110110",
  42169=>"011000011",
  42170=>"011111111",
  42171=>"001000000",
  42172=>"011111010",
  42173=>"111110011",
  42174=>"000011001",
  42175=>"000000001",
  42176=>"000000000",
  42177=>"101101100",
  42178=>"111010010",
  42179=>"001011001",
  42180=>"000000000",
  42181=>"100100100",
  42182=>"000010010",
  42183=>"000001000",
  42184=>"111100010",
  42185=>"101111111",
  42186=>"111110000",
  42187=>"110101101",
  42188=>"000000100",
  42189=>"100110010",
  42190=>"101000000",
  42191=>"000000101",
  42192=>"111000000",
  42193=>"100110111",
  42194=>"011011000",
  42195=>"100111000",
  42196=>"000001000",
  42197=>"000000100",
  42198=>"111010010",
  42199=>"010111000",
  42200=>"000000111",
  42201=>"000001011",
  42202=>"101110100",
  42203=>"111000000",
  42204=>"001001110",
  42205=>"111100101",
  42206=>"110010010",
  42207=>"110000010",
  42208=>"111000000",
  42209=>"111000100",
  42210=>"111000010",
  42211=>"000111111",
  42212=>"101101111",
  42213=>"100011000",
  42214=>"111111010",
  42215=>"011111101",
  42216=>"101101000",
  42217=>"000000101",
  42218=>"100101001",
  42219=>"111001001",
  42220=>"001000000",
  42221=>"111011000",
  42222=>"001000000",
  42223=>"000000111",
  42224=>"110110000",
  42225=>"011001001",
  42226=>"000101111",
  42227=>"010110110",
  42228=>"000110111",
  42229=>"111101101",
  42230=>"010000100",
  42231=>"111110111",
  42232=>"010000000",
  42233=>"110010010",
  42234=>"011011000",
  42235=>"101101011",
  42236=>"101111011",
  42237=>"110111100",
  42238=>"100111111",
  42239=>"010100000",
  42240=>"100100100",
  42241=>"010010101",
  42242=>"010111111",
  42243=>"111111111",
  42244=>"011011011",
  42245=>"111111010",
  42246=>"000010000",
  42247=>"100000111",
  42248=>"111111011",
  42249=>"101100111",
  42250=>"001001000",
  42251=>"000100000",
  42252=>"010111011",
  42253=>"000000000",
  42254=>"111100101",
  42255=>"000000001",
  42256=>"011111111",
  42257=>"001000000",
  42258=>"101011010",
  42259=>"111000100",
  42260=>"000010010",
  42261=>"111111111",
  42262=>"000100010",
  42263=>"101000100",
  42264=>"010000111",
  42265=>"010101000",
  42266=>"010000000",
  42267=>"101000100",
  42268=>"101111011",
  42269=>"100001101",
  42270=>"001101000",
  42271=>"110100101",
  42272=>"010111110",
  42273=>"010010010",
  42274=>"111100101",
  42275=>"001000000",
  42276=>"000011011",
  42277=>"011001000",
  42278=>"000011010",
  42279=>"110100100",
  42280=>"010111111",
  42281=>"101001101",
  42282=>"101100100",
  42283=>"000000000",
  42284=>"111011111",
  42285=>"101000001",
  42286=>"000000000",
  42287=>"000000000",
  42288=>"000111111",
  42289=>"011110000",
  42290=>"100000100",
  42291=>"000011001",
  42292=>"000000000",
  42293=>"000000011",
  42294=>"100000001",
  42295=>"000101100",
  42296=>"110110100",
  42297=>"100101111",
  42298=>"111111011",
  42299=>"000100110",
  42300=>"001011011",
  42301=>"000111111",
  42302=>"000000010",
  42303=>"000000100",
  42304=>"111000110",
  42305=>"100000000",
  42306=>"100111000",
  42307=>"011110000",
  42308=>"110111111",
  42309=>"000000111",
  42310=>"111001111",
  42311=>"111101111",
  42312=>"101011010",
  42313=>"011010010",
  42314=>"111100101",
  42315=>"001000000",
  42316=>"111011101",
  42317=>"000100000",
  42318=>"100111111",
  42319=>"000111101",
  42320=>"100000111",
  42321=>"110111111",
  42322=>"110111010",
  42323=>"010111101",
  42324=>"111000000",
  42325=>"111011010",
  42326=>"000001001",
  42327=>"111101001",
  42328=>"000001011",
  42329=>"000110100",
  42330=>"011011011",
  42331=>"000111000",
  42332=>"000111010",
  42333=>"010110000",
  42334=>"111111010",
  42335=>"011110110",
  42336=>"000100100",
  42337=>"000101001",
  42338=>"001000000",
  42339=>"111111111",
  42340=>"000011010",
  42341=>"111111100",
  42342=>"010000010",
  42343=>"100101100",
  42344=>"011001000",
  42345=>"000000000",
  42346=>"011000000",
  42347=>"111111111",
  42348=>"000000010",
  42349=>"000011100",
  42350=>"000000000",
  42351=>"111011010",
  42352=>"100110110",
  42353=>"001000000",
  42354=>"000000100",
  42355=>"100100000",
  42356=>"101111000",
  42357=>"101000011",
  42358=>"110011000",
  42359=>"110100000",
  42360=>"111001000",
  42361=>"011011001",
  42362=>"000000000",
  42363=>"111111000",
  42364=>"110001111",
  42365=>"101001100",
  42366=>"111101110",
  42367=>"010010011",
  42368=>"000000000",
  42369=>"110011010",
  42370=>"011001111",
  42371=>"100000110",
  42372=>"011001011",
  42373=>"101001000",
  42374=>"101100010",
  42375=>"000100100",
  42376=>"001011011",
  42377=>"100001001",
  42378=>"100000111",
  42379=>"111111111",
  42380=>"010011000",
  42381=>"100110111",
  42382=>"010000010",
  42383=>"001001011",
  42384=>"000000000",
  42385=>"010111100",
  42386=>"000000000",
  42387=>"111101001",
  42388=>"000001101",
  42389=>"000111111",
  42390=>"111111111",
  42391=>"000101100",
  42392=>"000000000",
  42393=>"010101000",
  42394=>"011111111",
  42395=>"000000111",
  42396=>"010101101",
  42397=>"111000000",
  42398=>"101000000",
  42399=>"111000000",
  42400=>"111110010",
  42401=>"110010000",
  42402=>"111101010",
  42403=>"111111111",
  42404=>"111010000",
  42405=>"011001000",
  42406=>"101111111",
  42407=>"000011010",
  42408=>"100000000",
  42409=>"000011111",
  42410=>"000010010",
  42411=>"100100110",
  42412=>"000000110",
  42413=>"000111101",
  42414=>"011111000",
  42415=>"010010000",
  42416=>"001000000",
  42417=>"010111000",
  42418=>"100000000",
  42419=>"100010011",
  42420=>"110101001",
  42421=>"110000011",
  42422=>"010000010",
  42423=>"010011100",
  42424=>"110111100",
  42425=>"011001001",
  42426=>"000100111",
  42427=>"001010111",
  42428=>"110110001",
  42429=>"010111111",
  42430=>"100100000",
  42431=>"100000101",
  42432=>"010010000",
  42433=>"000000000",
  42434=>"010010001",
  42435=>"001001000",
  42436=>"000100101",
  42437=>"110001110",
  42438=>"000100111",
  42439=>"111011000",
  42440=>"110010011",
  42441=>"100000000",
  42442=>"101110100",
  42443=>"101000100",
  42444=>"000100100",
  42445=>"010110110",
  42446=>"000000001",
  42447=>"111111001",
  42448=>"010000100",
  42449=>"100110000",
  42450=>"011111111",
  42451=>"111101111",
  42452=>"000000000",
  42453=>"011001000",
  42454=>"001000000",
  42455=>"000011111",
  42456=>"101100000",
  42457=>"000000001",
  42458=>"011010011",
  42459=>"111000000",
  42460=>"001001111",
  42461=>"100101101",
  42462=>"100000101",
  42463=>"000000000",
  42464=>"110010000",
  42465=>"000010011",
  42466=>"101100000",
  42467=>"011001000",
  42468=>"011000000",
  42469=>"010011111",
  42470=>"000100010",
  42471=>"100011100",
  42472=>"000000000",
  42473=>"000000101",
  42474=>"100000000",
  42475=>"111111111",
  42476=>"000111000",
  42477=>"000101110",
  42478=>"000110010",
  42479=>"001000000",
  42480=>"000100111",
  42481=>"110110110",
  42482=>"111101011",
  42483=>"001001011",
  42484=>"000011011",
  42485=>"111011100",
  42486=>"001000000",
  42487=>"100000000",
  42488=>"000100000",
  42489=>"111111111",
  42490=>"000000000",
  42491=>"011000000",
  42492=>"000000000",
  42493=>"000010000",
  42494=>"110100110",
  42495=>"000000000",
  42496=>"000110101",
  42497=>"111111001",
  42498=>"000010011",
  42499=>"000000000",
  42500=>"011000100",
  42501=>"100000001",
  42502=>"000000000",
  42503=>"011000000",
  42504=>"101101100",
  42505=>"000000000",
  42506=>"010111111",
  42507=>"111001100",
  42508=>"010111011",
  42509=>"010111001",
  42510=>"111100100",
  42511=>"110111011",
  42512=>"100000100",
  42513=>"010111111",
  42514=>"000011011",
  42515=>"111000000",
  42516=>"001111010",
  42517=>"000000000",
  42518=>"111100000",
  42519=>"011111100",
  42520=>"000000111",
  42521=>"010011111",
  42522=>"000000000",
  42523=>"000111111",
  42524=>"000111011",
  42525=>"000000000",
  42526=>"111111000",
  42527=>"011111000",
  42528=>"100000000",
  42529=>"111111111",
  42530=>"111000000",
  42531=>"111000000",
  42532=>"111111100",
  42533=>"000011010",
  42534=>"010111111",
  42535=>"000101001",
  42536=>"011111111",
  42537=>"011111111",
  42538=>"000000111",
  42539=>"000000000",
  42540=>"010111111",
  42541=>"000111000",
  42542=>"101000011",
  42543=>"111101101",
  42544=>"100000000",
  42545=>"010110000",
  42546=>"000000110",
  42547=>"011000001",
  42548=>"000010010",
  42549=>"111111111",
  42550=>"000011000",
  42551=>"000000000",
  42552=>"011000000",
  42553=>"111001000",
  42554=>"000000001",
  42555=>"110000000",
  42556=>"000001001",
  42557=>"001111111",
  42558=>"111000000",
  42559=>"000000000",
  42560=>"010111010",
  42561=>"010000110",
  42562=>"000000000",
  42563=>"111000000",
  42564=>"010111111",
  42565=>"000000000",
  42566=>"111111011",
  42567=>"000000111",
  42568=>"011011110",
  42569=>"000000000",
  42570=>"000000010",
  42571=>"101100100",
  42572=>"000000100",
  42573=>"000011001",
  42574=>"110011000",
  42575=>"011111111",
  42576=>"010111010",
  42577=>"001111111",
  42578=>"000100000",
  42579=>"111001000",
  42580=>"000000000",
  42581=>"001101000",
  42582=>"111111001",
  42583=>"111000000",
  42584=>"001110000",
  42585=>"010111111",
  42586=>"010010010",
  42587=>"010101100",
  42588=>"000000000",
  42589=>"110000000",
  42590=>"111111010",
  42591=>"111101000",
  42592=>"100000100",
  42593=>"100000000",
  42594=>"101011010",
  42595=>"001111001",
  42596=>"010111001",
  42597=>"011111111",
  42598=>"000000000",
  42599=>"000000001",
  42600=>"000000000",
  42601=>"000000000",
  42602=>"011100100",
  42603=>"101011010",
  42604=>"000001111",
  42605=>"000000000",
  42606=>"101100101",
  42607=>"010010000",
  42608=>"111110110",
  42609=>"000000111",
  42610=>"001111000",
  42611=>"111001111",
  42612=>"001100100",
  42613=>"000101000",
  42614=>"111101000",
  42615=>"000010000",
  42616=>"101001101",
  42617=>"110111000",
  42618=>"010010111",
  42619=>"010011001",
  42620=>"011001001",
  42621=>"100000000",
  42622=>"100000000",
  42623=>"100000000",
  42624=>"110000000",
  42625=>"000010010",
  42626=>"000000000",
  42627=>"111110111",
  42628=>"010100000",
  42629=>"000000100",
  42630=>"000000010",
  42631=>"011110100",
  42632=>"100111111",
  42633=>"001001000",
  42634=>"000000000",
  42635=>"101101001",
  42636=>"100000000",
  42637=>"100001101",
  42638=>"000000101",
  42639=>"110000000",
  42640=>"010011110",
  42641=>"010010000",
  42642=>"011101111",
  42643=>"101110110",
  42644=>"011110000",
  42645=>"000010000",
  42646=>"000111010",
  42647=>"000000000",
  42648=>"000101111",
  42649=>"010010001",
  42650=>"000111111",
  42651=>"000000000",
  42652=>"100000101",
  42653=>"000000000",
  42654=>"000000111",
  42655=>"101000100",
  42656=>"111010110",
  42657=>"111111110",
  42658=>"111011000",
  42659=>"111111111",
  42660=>"001100000",
  42661=>"110111000",
  42662=>"110110111",
  42663=>"011101100",
  42664=>"111011010",
  42665=>"101000100",
  42666=>"111111111",
  42667=>"111111111",
  42668=>"111111111",
  42669=>"100100101",
  42670=>"100111010",
  42671=>"101111011",
  42672=>"100000000",
  42673=>"100111110",
  42674=>"010100000",
  42675=>"011000000",
  42676=>"010111000",
  42677=>"010011111",
  42678=>"110000000",
  42679=>"000010011",
  42680=>"000110110",
  42681=>"110001001",
  42682=>"000000111",
  42683=>"011111111",
  42684=>"000000111",
  42685=>"000111001",
  42686=>"110100100",
  42687=>"000011110",
  42688=>"011111011",
  42689=>"000000101",
  42690=>"111111101",
  42691=>"111100111",
  42692=>"010001111",
  42693=>"101110111",
  42694=>"110111000",
  42695=>"000000000",
  42696=>"111111111",
  42697=>"000110000",
  42698=>"110111111",
  42699=>"000111011",
  42700=>"111100100",
  42701=>"100110100",
  42702=>"111111111",
  42703=>"000000000",
  42704=>"101000001",
  42705=>"000110100",
  42706=>"101001001",
  42707=>"000111001",
  42708=>"101101001",
  42709=>"001011111",
  42710=>"000000000",
  42711=>"100001000",
  42712=>"011000000",
  42713=>"010110010",
  42714=>"111011101",
  42715=>"000110110",
  42716=>"110011000",
  42717=>"011001100",
  42718=>"000000000",
  42719=>"111111111",
  42720=>"010111011",
  42721=>"010111111",
  42722=>"000000000",
  42723=>"111111111",
  42724=>"111000101",
  42725=>"101100000",
  42726=>"101000000",
  42727=>"011101000",
  42728=>"011111111",
  42729=>"111111110",
  42730=>"000011011",
  42731=>"111111111",
  42732=>"000011111",
  42733=>"111000000",
  42734=>"100111010",
  42735=>"100000000",
  42736=>"100111111",
  42737=>"101001001",
  42738=>"111101000",
  42739=>"110111010",
  42740=>"101001101",
  42741=>"011111111",
  42742=>"001000100",
  42743=>"000000100",
  42744=>"111100000",
  42745=>"011000000",
  42746=>"000011111",
  42747=>"111111000",
  42748=>"000111000",
  42749=>"111000000",
  42750=>"011111001",
  42751=>"000000000",
  42752=>"011100100",
  42753=>"111010000",
  42754=>"111100101",
  42755=>"001000111",
  42756=>"010000000",
  42757=>"000001111",
  42758=>"001111111",
  42759=>"010111111",
  42760=>"000001111",
  42761=>"000101111",
  42762=>"111010000",
  42763=>"001101100",
  42764=>"000000111",
  42765=>"111111111",
  42766=>"000111110",
  42767=>"101111110",
  42768=>"111111000",
  42769=>"011110000",
  42770=>"010000110",
  42771=>"001000001",
  42772=>"111110110",
  42773=>"000000111",
  42774=>"101011111",
  42775=>"011010000",
  42776=>"000000111",
  42777=>"001111111",
  42778=>"100111111",
  42779=>"111110000",
  42780=>"110111111",
  42781=>"100000000",
  42782=>"101000000",
  42783=>"100111111",
  42784=>"111001001",
  42785=>"111111111",
  42786=>"000110111",
  42787=>"000111111",
  42788=>"000000100",
  42789=>"011000010",
  42790=>"011000010",
  42791=>"000011001",
  42792=>"110000110",
  42793=>"111111000",
  42794=>"000110110",
  42795=>"000011111",
  42796=>"111111010",
  42797=>"111000000",
  42798=>"111000000",
  42799=>"000011111",
  42800=>"000000000",
  42801=>"100100000",
  42802=>"111111111",
  42803=>"001100000",
  42804=>"111111000",
  42805=>"000000000",
  42806=>"011000010",
  42807=>"000001111",
  42808=>"101010111",
  42809=>"000000001",
  42810=>"000010000",
  42811=>"000111110",
  42812=>"000001110",
  42813=>"111000110",
  42814=>"000000001",
  42815=>"000001100",
  42816=>"100000000",
  42817=>"001101111",
  42818=>"000111111",
  42819=>"000101111",
  42820=>"000000000",
  42821=>"101000000",
  42822=>"110010000",
  42823=>"111110011",
  42824=>"110001111",
  42825=>"101111010",
  42826=>"100001111",
  42827=>"001001011",
  42828=>"001000101",
  42829=>"100000000",
  42830=>"011001101",
  42831=>"000100000",
  42832=>"000000000",
  42833=>"111101111",
  42834=>"101111111",
  42835=>"001000000",
  42836=>"011010000",
  42837=>"010110011",
  42838=>"110011011",
  42839=>"000000000",
  42840=>"001111111",
  42841=>"000000011",
  42842=>"111111000",
  42843=>"000000111",
  42844=>"110000000",
  42845=>"001111111",
  42846=>"111000000",
  42847=>"001000110",
  42848=>"000111111",
  42849=>"010111111",
  42850=>"000101111",
  42851=>"111001000",
  42852=>"100001101",
  42853=>"011011111",
  42854=>"111111100",
  42855=>"000100000",
  42856=>"000000111",
  42857=>"101000100",
  42858=>"011111111",
  42859=>"010010111",
  42860=>"110010110",
  42861=>"111111000",
  42862=>"000001111",
  42863=>"111111111",
  42864=>"111111011",
  42865=>"000011000",
  42866=>"000000000",
  42867=>"000000000",
  42868=>"000000000",
  42869=>"000101001",
  42870=>"111111111",
  42871=>"000111111",
  42872=>"111000000",
  42873=>"101010111",
  42874=>"011110111",
  42875=>"000000111",
  42876=>"100001000",
  42877=>"100000000",
  42878=>"110000011",
  42879=>"000000111",
  42880=>"000000000",
  42881=>"000000111",
  42882=>"100111111",
  42883=>"111111110",
  42884=>"000000010",
  42885=>"000000101",
  42886=>"110100000",
  42887=>"000000000",
  42888=>"011010111",
  42889=>"111000000",
  42890=>"011011000",
  42891=>"000000101",
  42892=>"111001111",
  42893=>"001101111",
  42894=>"100110111",
  42895=>"000001111",
  42896=>"111111011",
  42897=>"111011111",
  42898=>"011000000",
  42899=>"111100000",
  42900=>"111000000",
  42901=>"000111111",
  42902=>"001100010",
  42903=>"101100111",
  42904=>"000000100",
  42905=>"000001000",
  42906=>"010110111",
  42907=>"000001000",
  42908=>"100100111",
  42909=>"100101111",
  42910=>"010010011",
  42911=>"000111111",
  42912=>"000001011",
  42913=>"010000000",
  42914=>"110101111",
  42915=>"000110101",
  42916=>"111101110",
  42917=>"110000010",
  42918=>"101000110",
  42919=>"000000000",
  42920=>"111111011",
  42921=>"101100010",
  42922=>"000101111",
  42923=>"001011000",
  42924=>"111110111",
  42925=>"000001111",
  42926=>"100001011",
  42927=>"000000111",
  42928=>"001100000",
  42929=>"100100111",
  42930=>"101101000",
  42931=>"000110111",
  42932=>"111100000",
  42933=>"011000000",
  42934=>"100011001",
  42935=>"011100000",
  42936=>"000110111",
  42937=>"111011000",
  42938=>"000000000",
  42939=>"111110111",
  42940=>"000100111",
  42941=>"000111111",
  42942=>"000000110",
  42943=>"000000000",
  42944=>"010010000",
  42945=>"000001000",
  42946=>"001001000",
  42947=>"001011011",
  42948=>"000000000",
  42949=>"011000100",
  42950=>"010000000",
  42951=>"001111010",
  42952=>"000111111",
  42953=>"001001011",
  42954=>"001111100",
  42955=>"000011000",
  42956=>"011000000",
  42957=>"100100010",
  42958=>"000000000",
  42959=>"000001111",
  42960=>"000000000",
  42961=>"011011111",
  42962=>"000000111",
  42963=>"111100010",
  42964=>"000110111",
  42965=>"110011000",
  42966=>"111000000",
  42967=>"100000000",
  42968=>"111000000",
  42969=>"001111111",
  42970=>"000000100",
  42971=>"000001111",
  42972=>"111010110",
  42973=>"100100111",
  42974=>"101111010",
  42975=>"111111000",
  42976=>"111100101",
  42977=>"100110111",
  42978=>"000000001",
  42979=>"010011011",
  42980=>"011000000",
  42981=>"000000111",
  42982=>"001000111",
  42983=>"110000111",
  42984=>"000000010",
  42985=>"111101001",
  42986=>"111010000",
  42987=>"101111111",
  42988=>"000010101",
  42989=>"001000000",
  42990=>"011000000",
  42991=>"000100100",
  42992=>"001111101",
  42993=>"011101000",
  42994=>"001101011",
  42995=>"111101100",
  42996=>"001000011",
  42997=>"111000000",
  42998=>"000000111",
  42999=>"111101000",
  43000=>"011000111",
  43001=>"110000110",
  43002=>"100111111",
  43003=>"111000010",
  43004=>"000100010",
  43005=>"000001011",
  43006=>"001001111",
  43007=>"000011010",
  43008=>"111010010",
  43009=>"111001000",
  43010=>"101101111",
  43011=>"111010000",
  43012=>"110111110",
  43013=>"001111110",
  43014=>"000111100",
  43015=>"001011110",
  43016=>"010011001",
  43017=>"000101110",
  43018=>"101001001",
  43019=>"000000100",
  43020=>"011000000",
  43021=>"100101001",
  43022=>"011110100",
  43023=>"001000000",
  43024=>"000110001",
  43025=>"001000000",
  43026=>"101010010",
  43027=>"011111001",
  43028=>"101101101",
  43029=>"000000101",
  43030=>"111010111",
  43031=>"000000000",
  43032=>"000111101",
  43033=>"110111101",
  43034=>"011111101",
  43035=>"010101100",
  43036=>"000000100",
  43037=>"111100101",
  43038=>"001011100",
  43039=>"111000000",
  43040=>"010111111",
  43041=>"100000001",
  43042=>"111101101",
  43043=>"000011000",
  43044=>"010011010",
  43045=>"011011111",
  43046=>"100101111",
  43047=>"111111111",
  43048=>"100101111",
  43049=>"000000010",
  43050=>"111100000",
  43051=>"100000000",
  43052=>"011000010",
  43053=>"000000000",
  43054=>"111000000",
  43055=>"010010000",
  43056=>"000010100",
  43057=>"010111011",
  43058=>"001010111",
  43059=>"111111101",
  43060=>"001000000",
  43061=>"000001100",
  43062=>"001011000",
  43063=>"110010000",
  43064=>"101011001",
  43065=>"111111000",
  43066=>"100100011",
  43067=>"000000111",
  43068=>"111010011",
  43069=>"001010111",
  43070=>"100101101",
  43071=>"010011101",
  43072=>"101010111",
  43073=>"101111111",
  43074=>"011111111",
  43075=>"100010011",
  43076=>"010111011",
  43077=>"000000111",
  43078=>"111111011",
  43079=>"011011011",
  43080=>"100010011",
  43081=>"111001101",
  43082=>"011100000",
  43083=>"011000110",
  43084=>"010101111",
  43085=>"010110111",
  43086=>"000110111",
  43087=>"101101000",
  43088=>"010010001",
  43089=>"111111111",
  43090=>"011000000",
  43091=>"011011001",
  43092=>"010100110",
  43093=>"111110001",
  43094=>"101010001",
  43095=>"001101101",
  43096=>"111111011",
  43097=>"011010110",
  43098=>"111100000",
  43099=>"110000000",
  43100=>"011000101",
  43101=>"101100110",
  43102=>"111101111",
  43103=>"001010100",
  43104=>"010010110",
  43105=>"011011000",
  43106=>"100100110",
  43107=>"111011000",
  43108=>"111000000",
  43109=>"110010110",
  43110=>"111001001",
  43111=>"100100100",
  43112=>"010010111",
  43113=>"000111111",
  43114=>"000111111",
  43115=>"000000000",
  43116=>"000011001",
  43117=>"000000000",
  43118=>"110111111",
  43119=>"000011011",
  43120=>"011011111",
  43121=>"000111111",
  43122=>"110110011",
  43123=>"011111111",
  43124=>"000111000",
  43125=>"000000000",
  43126=>"010111001",
  43127=>"001101101",
  43128=>"001101111",
  43129=>"101011100",
  43130=>"111101100",
  43131=>"001011011",
  43132=>"100010001",
  43133=>"101110110",
  43134=>"000010111",
  43135=>"111010111",
  43136=>"000111110",
  43137=>"001010000",
  43138=>"000101100",
  43139=>"111011000",
  43140=>"000010010",
  43141=>"000000000",
  43142=>"110110111",
  43143=>"111011110",
  43144=>"110110110",
  43145=>"011010111",
  43146=>"100111000",
  43147=>"011000010",
  43148=>"110101111",
  43149=>"100110111",
  43150=>"111010111",
  43151=>"000110010",
  43152=>"111110011",
  43153=>"100111111",
  43154=>"110100011",
  43155=>"111111101",
  43156=>"010111000",
  43157=>"000101101",
  43158=>"101110000",
  43159=>"001001010",
  43160=>"111111010",
  43161=>"011000000",
  43162=>"111110111",
  43163=>"000110000",
  43164=>"010111101",
  43165=>"000010011",
  43166=>"110100001",
  43167=>"001000000",
  43168=>"000010101",
  43169=>"011110100",
  43170=>"000000000",
  43171=>"101111111",
  43172=>"010110111",
  43173=>"010110001",
  43174=>"110010101",
  43175=>"111101101",
  43176=>"111111001",
  43177=>"000001111",
  43178=>"100100000",
  43179=>"000010001",
  43180=>"111101011",
  43181=>"000100111",
  43182=>"000010000",
  43183=>"111000001",
  43184=>"110000000",
  43185=>"001000011",
  43186=>"101111111",
  43187=>"110111001",
  43188=>"111010110",
  43189=>"000000011",
  43190=>"111001000",
  43191=>"001111100",
  43192=>"000010110",
  43193=>"110011001",
  43194=>"010111111",
  43195=>"111101000",
  43196=>"101000000",
  43197=>"001111111",
  43198=>"110110110",
  43199=>"101001101",
  43200=>"111100000",
  43201=>"111000000",
  43202=>"011010000",
  43203=>"010010010",
  43204=>"000000000",
  43205=>"011000000",
  43206=>"101011000",
  43207=>"111000000",
  43208=>"101111101",
  43209=>"111110101",
  43210=>"010000000",
  43211=>"011010111",
  43212=>"000000000",
  43213=>"101010100",
  43214=>"110000000",
  43215=>"010111000",
  43216=>"010110000",
  43217=>"110110110",
  43218=>"111111101",
  43219=>"001000000",
  43220=>"111000101",
  43221=>"100010000",
  43222=>"111101000",
  43223=>"010010000",
  43224=>"101000000",
  43225=>"111000101",
  43226=>"110100001",
  43227=>"111101101",
  43228=>"000010101",
  43229=>"000000000",
  43230=>"111011111",
  43231=>"001101000",
  43232=>"000111000",
  43233=>"000000000",
  43234=>"101100000",
  43235=>"011011011",
  43236=>"000101101",
  43237=>"010010010",
  43238=>"000011111",
  43239=>"000010000",
  43240=>"100111111",
  43241=>"010000101",
  43242=>"101101100",
  43243=>"111101000",
  43244=>"000101101",
  43245=>"000111100",
  43246=>"000101111",
  43247=>"000010000",
  43248=>"000000000",
  43249=>"111000001",
  43250=>"001000101",
  43251=>"011011000",
  43252=>"001001010",
  43253=>"111000001",
  43254=>"000000100",
  43255=>"111111111",
  43256=>"101100101",
  43257=>"111111101",
  43258=>"010110101",
  43259=>"111111000",
  43260=>"010010000",
  43261=>"111000110",
  43262=>"011011101",
  43263=>"010000000",
  43264=>"001101000",
  43265=>"000010010",
  43266=>"001000111",
  43267=>"000000101",
  43268=>"001011000",
  43269=>"110111111",
  43270=>"001111000",
  43271=>"000001111",
  43272=>"000000000",
  43273=>"000000000",
  43274=>"110100100",
  43275=>"110111000",
  43276=>"000000000",
  43277=>"110110100",
  43278=>"011111111",
  43279=>"111111111",
  43280=>"000000000",
  43281=>"000100000",
  43282=>"000000010",
  43283=>"011010000",
  43284=>"101010000",
  43285=>"111001111",
  43286=>"110100111",
  43287=>"010111101",
  43288=>"000000000",
  43289=>"111110110",
  43290=>"000010011",
  43291=>"000000111",
  43292=>"000000101",
  43293=>"000000010",
  43294=>"011010011",
  43295=>"000010010",
  43296=>"110000111",
  43297=>"000010000",
  43298=>"111001111",
  43299=>"000000000",
  43300=>"001000001",
  43301=>"100110100",
  43302=>"000100000",
  43303=>"111101001",
  43304=>"101010111",
  43305=>"100100000",
  43306=>"000100000",
  43307=>"010000000",
  43308=>"000010100",
  43309=>"011010000",
  43310=>"111010010",
  43311=>"111111011",
  43312=>"110110000",
  43313=>"100001011",
  43314=>"011010000",
  43315=>"000101101",
  43316=>"111111000",
  43317=>"110000110",
  43318=>"111111011",
  43319=>"010111111",
  43320=>"000011011",
  43321=>"000000101",
  43322=>"000000111",
  43323=>"111101100",
  43324=>"100110110",
  43325=>"111111010",
  43326=>"000000000",
  43327=>"011011100",
  43328=>"000111101",
  43329=>"010111000",
  43330=>"100101001",
  43331=>"111111000",
  43332=>"010000000",
  43333=>"000100000",
  43334=>"000111100",
  43335=>"101111111",
  43336=>"010011011",
  43337=>"000010000",
  43338=>"010000000",
  43339=>"000001010",
  43340=>"010010000",
  43341=>"011011010",
  43342=>"000100000",
  43343=>"000001000",
  43344=>"000111111",
  43345=>"111110000",
  43346=>"011010100",
  43347=>"000110000",
  43348=>"100000010",
  43349=>"110000001",
  43350=>"010011110",
  43351=>"010000111",
  43352=>"000110111",
  43353=>"000001111",
  43354=>"111111011",
  43355=>"100100111",
  43356=>"010000000",
  43357=>"010000011",
  43358=>"111001000",
  43359=>"101100101",
  43360=>"000110111",
  43361=>"000111111",
  43362=>"111100111",
  43363=>"001101110",
  43364=>"000010000",
  43365=>"111100110",
  43366=>"100110011",
  43367=>"111011011",
  43368=>"101000011",
  43369=>"101101111",
  43370=>"110101101",
  43371=>"000111111",
  43372=>"010000101",
  43373=>"101101101",
  43374=>"111101001",
  43375=>"000111111",
  43376=>"001111110",
  43377=>"000000111",
  43378=>"010101110",
  43379=>"011000000",
  43380=>"010100000",
  43381=>"100101101",
  43382=>"000101100",
  43383=>"010110111",
  43384=>"000100100",
  43385=>"011101111",
  43386=>"011111111",
  43387=>"001001001",
  43388=>"100100010",
  43389=>"000010000",
  43390=>"001101111",
  43391=>"000000110",
  43392=>"000001101",
  43393=>"011100000",
  43394=>"010010010",
  43395=>"000000001",
  43396=>"000010000",
  43397=>"001001111",
  43398=>"001011000",
  43399=>"100100110",
  43400=>"100100011",
  43401=>"111101100",
  43402=>"101101000",
  43403=>"000010111",
  43404=>"000110111",
  43405=>"101101111",
  43406=>"010101111",
  43407=>"000001001",
  43408=>"011001011",
  43409=>"001111111",
  43410=>"100000000",
  43411=>"000111111",
  43412=>"100101111",
  43413=>"000000111",
  43414=>"010011110",
  43415=>"000010000",
  43416=>"111101001",
  43417=>"011011000",
  43418=>"100010010",
  43419=>"111101101",
  43420=>"111101100",
  43421=>"111011110",
  43422=>"101000010",
  43423=>"000000000",
  43424=>"010000100",
  43425=>"101000000",
  43426=>"101101111",
  43427=>"000110000",
  43428=>"010111111",
  43429=>"011100110",
  43430=>"000000110",
  43431=>"000110100",
  43432=>"010010000",
  43433=>"100100001",
  43434=>"101000000",
  43435=>"110101000",
  43436=>"000000011",
  43437=>"000100100",
  43438=>"110100100",
  43439=>"101111000",
  43440=>"000000010",
  43441=>"110101011",
  43442=>"011110000",
  43443=>"100110110",
  43444=>"100111011",
  43445=>"110011010",
  43446=>"000001001",
  43447=>"011000010",
  43448=>"001001011",
  43449=>"001001011",
  43450=>"000011011",
  43451=>"011110000",
  43452=>"000000000",
  43453=>"111111111",
  43454=>"000100101",
  43455=>"000011010",
  43456=>"010010000",
  43457=>"000001101",
  43458=>"101010000",
  43459=>"011010111",
  43460=>"010111000",
  43461=>"111111110",
  43462=>"000111111",
  43463=>"111100111",
  43464=>"100100000",
  43465=>"000001011",
  43466=>"111100101",
  43467=>"000100110",
  43468=>"001100000",
  43469=>"101001011",
  43470=>"100000010",
  43471=>"111000101",
  43472=>"100111000",
  43473=>"000110110",
  43474=>"101010111",
  43475=>"010000111",
  43476=>"000010111",
  43477=>"000000000",
  43478=>"010000101",
  43479=>"101000011",
  43480=>"110111000",
  43481=>"000111111",
  43482=>"001000001",
  43483=>"101101101",
  43484=>"001000110",
  43485=>"001000000",
  43486=>"000111111",
  43487=>"000010000",
  43488=>"100101000",
  43489=>"111101000",
  43490=>"111001001",
  43491=>"011001001",
  43492=>"000000000",
  43493=>"000010101",
  43494=>"111101101",
  43495=>"111010100",
  43496=>"100101101",
  43497=>"111000000",
  43498=>"111001001",
  43499=>"000000110",
  43500=>"000000000",
  43501=>"101010000",
  43502=>"111000000",
  43503=>"111000011",
  43504=>"100000011",
  43505=>"111011010",
  43506=>"010000000",
  43507=>"001110110",
  43508=>"110110000",
  43509=>"111001101",
  43510=>"000010010",
  43511=>"100100010",
  43512=>"111110110",
  43513=>"000000101",
  43514=>"111110110",
  43515=>"101100001",
  43516=>"111000100",
  43517=>"010101000",
  43518=>"100100111",
  43519=>"111001100",
  43520=>"011011001",
  43521=>"000001100",
  43522=>"100000101",
  43523=>"010100100",
  43524=>"010001011",
  43525=>"111110000",
  43526=>"101000111",
  43527=>"000010011",
  43528=>"000011111",
  43529=>"000000111",
  43530=>"101001001",
  43531=>"001000011",
  43532=>"000000000",
  43533=>"100111101",
  43534=>"100001011",
  43535=>"110001111",
  43536=>"100110101",
  43537=>"100100010",
  43538=>"111110111",
  43539=>"111100100",
  43540=>"110101111",
  43541=>"000100000",
  43542=>"110100101",
  43543=>"101101111",
  43544=>"000000000",
  43545=>"011000000",
  43546=>"000011000",
  43547=>"011011111",
  43548=>"000100111",
  43549=>"010011000",
  43550=>"111101101",
  43551=>"100100000",
  43552=>"000000100",
  43553=>"111100010",
  43554=>"111101001",
  43555=>"000011000",
  43556=>"011011001",
  43557=>"110111011",
  43558=>"000010010",
  43559=>"000001110",
  43560=>"101000101",
  43561=>"000111111",
  43562=>"100000000",
  43563=>"100000100",
  43564=>"111000101",
  43565=>"000101111",
  43566=>"011000101",
  43567=>"010100100",
  43568=>"001000110",
  43569=>"101100011",
  43570=>"000010111",
  43571=>"000100001",
  43572=>"000000111",
  43573=>"000000000",
  43574=>"100100111",
  43575=>"000000000",
  43576=>"011000011",
  43577=>"101100111",
  43578=>"100000110",
  43579=>"000100000",
  43580=>"010010000",
  43581=>"111111000",
  43582=>"100100011",
  43583=>"011111110",
  43584=>"011111111",
  43585=>"110111111",
  43586=>"111111011",
  43587=>"010010000",
  43588=>"011111101",
  43589=>"111101101",
  43590=>"001011111",
  43591=>"010000110",
  43592=>"101001111",
  43593=>"000000000",
  43594=>"001000101",
  43595=>"111000011",
  43596=>"111111111",
  43597=>"101001001",
  43598=>"100000000",
  43599=>"101111111",
  43600=>"100000100",
  43601=>"110111111",
  43602=>"101111111",
  43603=>"001101101",
  43604=>"000011011",
  43605=>"011111111",
  43606=>"111010110",
  43607=>"000111111",
  43608=>"100000011",
  43609=>"011110100",
  43610=>"100100000",
  43611=>"110110000",
  43612=>"000101100",
  43613=>"001000001",
  43614=>"010111111",
  43615=>"100010001",
  43616=>"000111010",
  43617=>"011111000",
  43618=>"101111010",
  43619=>"001000111",
  43620=>"000000001",
  43621=>"100001010",
  43622=>"000000111",
  43623=>"100000000",
  43624=>"111101000",
  43625=>"111010111",
  43626=>"111011101",
  43627=>"010001101",
  43628=>"010010101",
  43629=>"000100100",
  43630=>"100000000",
  43631=>"111000001",
  43632=>"100111011",
  43633=>"000001011",
  43634=>"000001011",
  43635=>"111111001",
  43636=>"111111111",
  43637=>"000000101",
  43638=>"010000011",
  43639=>"101101111",
  43640=>"011001011",
  43641=>"111111000",
  43642=>"111101101",
  43643=>"111101100",
  43644=>"100000011",
  43645=>"110100100",
  43646=>"000101010",
  43647=>"111110110",
  43648=>"111101100",
  43649=>"111000010",
  43650=>"011011110",
  43651=>"111011101",
  43652=>"000101101",
  43653=>"111001011",
  43654=>"011011111",
  43655=>"000000100",
  43656=>"100100100",
  43657=>"011111100",
  43658=>"100100111",
  43659=>"010000000",
  43660=>"000000000",
  43661=>"001111100",
  43662=>"011010010",
  43663=>"001000000",
  43664=>"010000000",
  43665=>"010010000",
  43666=>"000000000",
  43667=>"101101111",
  43668=>"000000111",
  43669=>"000001111",
  43670=>"010111111",
  43671=>"000011011",
  43672=>"110111000",
  43673=>"100000111",
  43674=>"000000010",
  43675=>"000011010",
  43676=>"000100010",
  43677=>"011000000",
  43678=>"010000110",
  43679=>"000000110",
  43680=>"001110100",
  43681=>"010000010",
  43682=>"100111111",
  43683=>"111111111",
  43684=>"111111000",
  43685=>"011011001",
  43686=>"110110011",
  43687=>"111111011",
  43688=>"010000101",
  43689=>"000010111",
  43690=>"100111111",
  43691=>"010000000",
  43692=>"111111011",
  43693=>"101000110",
  43694=>"100000010",
  43695=>"111100101",
  43696=>"000100000",
  43697=>"000100000",
  43698=>"000000000",
  43699=>"111001000",
  43700=>"110110100",
  43701=>"111100000",
  43702=>"100110100",
  43703=>"000000000",
  43704=>"110110110",
  43705=>"000001001",
  43706=>"110000100",
  43707=>"111000000",
  43708=>"111000011",
  43709=>"110011010",
  43710=>"111111001",
  43711=>"101100110",
  43712=>"100000000",
  43713=>"101000101",
  43714=>"000000101",
  43715=>"001110100",
  43716=>"101001001",
  43717=>"100000111",
  43718=>"010110100",
  43719=>"100000101",
  43720=>"100000010",
  43721=>"000100000",
  43722=>"111101000",
  43723=>"111101000",
  43724=>"111100000",
  43725=>"001000111",
  43726=>"101101111",
  43727=>"010111000",
  43728=>"000000011",
  43729=>"110110111",
  43730=>"000000000",
  43731=>"111111111",
  43732=>"000001101",
  43733=>"100110000",
  43734=>"100110111",
  43735=>"000111111",
  43736=>"100100111",
  43737=>"111000000",
  43738=>"101101001",
  43739=>"000000000",
  43740=>"111011111",
  43741=>"000011111",
  43742=>"111111111",
  43743=>"100101110",
  43744=>"000000000",
  43745=>"000000100",
  43746=>"100100111",
  43747=>"001111100",
  43748=>"101000000",
  43749=>"010010011",
  43750=>"010110111",
  43751=>"010001000",
  43752=>"000111101",
  43753=>"100111111",
  43754=>"111100100",
  43755=>"110100100",
  43756=>"000011010",
  43757=>"101011010",
  43758=>"000000000",
  43759=>"000010000",
  43760=>"111111100",
  43761=>"000000011",
  43762=>"010001101",
  43763=>"010001011",
  43764=>"111110111",
  43765=>"100101111",
  43766=>"000000000",
  43767=>"110000001",
  43768=>"000000111",
  43769=>"100001000",
  43770=>"100100101",
  43771=>"000000111",
  43772=>"111010000",
  43773=>"000000000",
  43774=>"110110100",
  43775=>"100000011",
  43776=>"111000100",
  43777=>"010011010",
  43778=>"000000101",
  43779=>"110010000",
  43780=>"111001100",
  43781=>"100100111",
  43782=>"111000011",
  43783=>"111011111",
  43784=>"011101111",
  43785=>"101100100",
  43786=>"000010010",
  43787=>"100101000",
  43788=>"000000100",
  43789=>"000000010",
  43790=>"101001000",
  43791=>"101001111",
  43792=>"111001001",
  43793=>"101000000",
  43794=>"101101111",
  43795=>"000000001",
  43796=>"000000010",
  43797=>"000000100",
  43798=>"000010011",
  43799=>"001111000",
  43800=>"000000000",
  43801=>"000000100",
  43802=>"100100000",
  43803=>"111000000",
  43804=>"100110101",
  43805=>"111111111",
  43806=>"001000001",
  43807=>"011010010",
  43808=>"000000110",
  43809=>"110101111",
  43810=>"000010110",
  43811=>"000000111",
  43812=>"001001111",
  43813=>"110000001",
  43814=>"000010000",
  43815=>"111111111",
  43816=>"100100010",
  43817=>"100000000",
  43818=>"101101001",
  43819=>"100000111",
  43820=>"000011101",
  43821=>"010010000",
  43822=>"010010010",
  43823=>"010000000",
  43824=>"111101101",
  43825=>"011000110",
  43826=>"101000111",
  43827=>"100000101",
  43828=>"010010010",
  43829=>"000111111",
  43830=>"000011010",
  43831=>"011010000",
  43832=>"100001111",
  43833=>"011011000",
  43834=>"101101101",
  43835=>"101100111",
  43836=>"111111011",
  43837=>"111111011",
  43838=>"001000000",
  43839=>"010100110",
  43840=>"000000111",
  43841=>"000000100",
  43842=>"111000000",
  43843=>"111001100",
  43844=>"111111000",
  43845=>"111100101",
  43846=>"000100100",
  43847=>"111001000",
  43848=>"111111111",
  43849=>"111111011",
  43850=>"010010000",
  43851=>"111011101",
  43852=>"101000101",
  43853=>"000100110",
  43854=>"110110000",
  43855=>"000100111",
  43856=>"010010010",
  43857=>"111111010",
  43858=>"111111010",
  43859=>"101101100",
  43860=>"000011111",
  43861=>"100110110",
  43862=>"100111111",
  43863=>"000100010",
  43864=>"101110110",
  43865=>"001100100",
  43866=>"000001001",
  43867=>"111100111",
  43868=>"110100000",
  43869=>"111011011",
  43870=>"111101011",
  43871=>"110100001",
  43872=>"000000000",
  43873=>"001000000",
  43874=>"100001101",
  43875=>"000100000",
  43876=>"110000001",
  43877=>"111011111",
  43878=>"011010011",
  43879=>"111100010",
  43880=>"001111111",
  43881=>"101000110",
  43882=>"101101111",
  43883=>"111101101",
  43884=>"101111111",
  43885=>"101100000",
  43886=>"010000000",
  43887=>"010100101",
  43888=>"000000000",
  43889=>"111100101",
  43890=>"000010110",
  43891=>"010111011",
  43892=>"010010000",
  43893=>"001000101",
  43894=>"010000001",
  43895=>"000000100",
  43896=>"001000000",
  43897=>"011000000",
  43898=>"011011100",
  43899=>"010000011",
  43900=>"110111110",
  43901=>"111100110",
  43902=>"001101111",
  43903=>"001101000",
  43904=>"101000111",
  43905=>"110011011",
  43906=>"100000111",
  43907=>"011000011",
  43908=>"000000000",
  43909=>"101111111",
  43910=>"000100110",
  43911=>"000010001",
  43912=>"010110000",
  43913=>"010111111",
  43914=>"001000000",
  43915=>"111000100",
  43916=>"011100010",
  43917=>"000000111",
  43918=>"100100101",
  43919=>"000000000",
  43920=>"110100110",
  43921=>"001100000",
  43922=>"001101111",
  43923=>"010111111",
  43924=>"001010000",
  43925=>"000000100",
  43926=>"000110001",
  43927=>"000100100",
  43928=>"000101111",
  43929=>"100111111",
  43930=>"100000101",
  43931=>"100101101",
  43932=>"011101101",
  43933=>"100100101",
  43934=>"000001111",
  43935=>"110111111",
  43936=>"011011011",
  43937=>"101011111",
  43938=>"010011101",
  43939=>"101100110",
  43940=>"111011000",
  43941=>"100000111",
  43942=>"111111000",
  43943=>"000101100",
  43944=>"010111101",
  43945=>"000111100",
  43946=>"101101100",
  43947=>"000101100",
  43948=>"000010010",
  43949=>"001100101",
  43950=>"010000011",
  43951=>"110011000",
  43952=>"011000000",
  43953=>"011011011",
  43954=>"111100000",
  43955=>"110001100",
  43956=>"111011110",
  43957=>"100100111",
  43958=>"000000011",
  43959=>"100100101",
  43960=>"111111111",
  43961=>"001011001",
  43962=>"110000011",
  43963=>"010101101",
  43964=>"000000111",
  43965=>"101101001",
  43966=>"100001011",
  43967=>"000010111",
  43968=>"001100000",
  43969=>"000100111",
  43970=>"110010000",
  43971=>"000000000",
  43972=>"010100110",
  43973=>"010001000",
  43974=>"000101011",
  43975=>"000000000",
  43976=>"010111111",
  43977=>"000011010",
  43978=>"000010100",
  43979=>"000100111",
  43980=>"011100100",
  43981=>"111011010",
  43982=>"000000000",
  43983=>"010101111",
  43984=>"001101011",
  43985=>"010000011",
  43986=>"110100000",
  43987=>"000000011",
  43988=>"101001000",
  43989=>"110110000",
  43990=>"111111100",
  43991=>"000010110",
  43992=>"000110101",
  43993=>"011111000",
  43994=>"100100110",
  43995=>"101100101",
  43996=>"000000000",
  43997=>"111010111",
  43998=>"000000010",
  43999=>"111101011",
  44000=>"000101111",
  44001=>"010001000",
  44002=>"111110000",
  44003=>"110001001",
  44004=>"101100100",
  44005=>"111111110",
  44006=>"110111111",
  44007=>"000100100",
  44008=>"111001000",
  44009=>"001000001",
  44010=>"010011000",
  44011=>"100100000",
  44012=>"010010100",
  44013=>"000111110",
  44014=>"001000000",
  44015=>"111101101",
  44016=>"100101111",
  44017=>"011101000",
  44018=>"010010000",
  44019=>"110100111",
  44020=>"010000001",
  44021=>"000010011",
  44022=>"101100101",
  44023=>"100000110",
  44024=>"101101111",
  44025=>"100111111",
  44026=>"111000000",
  44027=>"000100000",
  44028=>"000101111",
  44029=>"111100000",
  44030=>"110000000",
  44031=>"100010000",
  44032=>"010000100",
  44033=>"100101000",
  44034=>"001001001",
  44035=>"000001111",
  44036=>"110111001",
  44037=>"000010010",
  44038=>"000111111",
  44039=>"101111111",
  44040=>"010000000",
  44041=>"111111000",
  44042=>"000000010",
  44043=>"111110101",
  44044=>"000110110",
  44045=>"010011010",
  44046=>"111111111",
  44047=>"110000000",
  44048=>"111101011",
  44049=>"001111111",
  44050=>"001000010",
  44051=>"000101111",
  44052=>"000000001",
  44053=>"000111111",
  44054=>"111100000",
  44055=>"110111111",
  44056=>"000000001",
  44057=>"111111111",
  44058=>"111101110",
  44059=>"111111011",
  44060=>"111111111",
  44061=>"111111000",
  44062=>"000000000",
  44063=>"000000101",
  44064=>"010100000",
  44065=>"010000001",
  44066=>"111010111",
  44067=>"111000000",
  44068=>"100101000",
  44069=>"100000001",
  44070=>"111100000",
  44071=>"110000000",
  44072=>"111110011",
  44073=>"111111000",
  44074=>"111111111",
  44075=>"110111110",
  44076=>"000111000",
  44077=>"000000000",
  44078=>"111111000",
  44079=>"110111000",
  44080=>"101011000",
  44081=>"000000000",
  44082=>"000000100",
  44083=>"000111111",
  44084=>"111111000",
  44085=>"111110101",
  44086=>"001001011",
  44087=>"000111011",
  44088=>"000000101",
  44089=>"000000111",
  44090=>"000000111",
  44091=>"111111111",
  44092=>"110000001",
  44093=>"001111111",
  44094=>"000111111",
  44095=>"011000000",
  44096=>"111111111",
  44097=>"000000000",
  44098=>"000010000",
  44099=>"111011000",
  44100=>"001000000",
  44101=>"000000000",
  44102=>"111110110",
  44103=>"000111111",
  44104=>"000000000",
  44105=>"011000000",
  44106=>"000010000",
  44107=>"111111111",
  44108=>"001111111",
  44109=>"000100000",
  44110=>"000000000",
  44111=>"110011011",
  44112=>"111110110",
  44113=>"000011111",
  44114=>"000000011",
  44115=>"000100110",
  44116=>"000010000",
  44117=>"100001001",
  44118=>"101110000",
  44119=>"000111111",
  44120=>"000000101",
  44121=>"001000101",
  44122=>"101101000",
  44123=>"000111111",
  44124=>"000011000",
  44125=>"000001011",
  44126=>"010000000",
  44127=>"011111100",
  44128=>"111110111",
  44129=>"001000000",
  44130=>"000111111",
  44131=>"110011001",
  44132=>"100100001",
  44133=>"100011001",
  44134=>"000000001",
  44135=>"010101001",
  44136=>"111011111",
  44137=>"000110111",
  44138=>"000000010",
  44139=>"000100101",
  44140=>"111101001",
  44141=>"000110111",
  44142=>"111111110",
  44143=>"110111110",
  44144=>"110111110",
  44145=>"001111111",
  44146=>"100110110",
  44147=>"000000010",
  44148=>"000000101",
  44149=>"000000101",
  44150=>"111111111",
  44151=>"000000001",
  44152=>"000111111",
  44153=>"000000000",
  44154=>"000000000",
  44155=>"101000111",
  44156=>"011111111",
  44157=>"000001011",
  44158=>"000000000",
  44159=>"111001000",
  44160=>"110000001",
  44161=>"111111010",
  44162=>"111000000",
  44163=>"101000000",
  44164=>"101001000",
  44165=>"000000000",
  44166=>"011000000",
  44167=>"101111101",
  44168=>"001100110",
  44169=>"111111111",
  44170=>"111010010",
  44171=>"000101001",
  44172=>"111101000",
  44173=>"110110100",
  44174=>"000111101",
  44175=>"111111100",
  44176=>"000000111",
  44177=>"100000100",
  44178=>"000001001",
  44179=>"111111101",
  44180=>"001101111",
  44181=>"111111001",
  44182=>"010010010",
  44183=>"100000000",
  44184=>"111111111",
  44185=>"000001001",
  44186=>"111111111",
  44187=>"111111110",
  44188=>"100110000",
  44189=>"111111111",
  44190=>"000010101",
  44191=>"111111111",
  44192=>"000000000",
  44193=>"111111010",
  44194=>"111111111",
  44195=>"111010101",
  44196=>"000010011",
  44197=>"101111111",
  44198=>"000001000",
  44199=>"111111101",
  44200=>"110010000",
  44201=>"010000000",
  44202=>"011011011",
  44203=>"101101111",
  44204=>"010000011",
  44205=>"000000001",
  44206=>"001001001",
  44207=>"000010010",
  44208=>"000000010",
  44209=>"110110100",
  44210=>"000000011",
  44211=>"111111111",
  44212=>"000000011",
  44213=>"000000000",
  44214=>"100100110",
  44215=>"010101000",
  44216=>"000000100",
  44217=>"100111110",
  44218=>"111001001",
  44219=>"111111101",
  44220=>"111100101",
  44221=>"000000000",
  44222=>"110110010",
  44223=>"111111000",
  44224=>"000010010",
  44225=>"101111111",
  44226=>"010000000",
  44227=>"001011001",
  44228=>"110111110",
  44229=>"010010001",
  44230=>"000000011",
  44231=>"000110010",
  44232=>"111111111",
  44233=>"000000010",
  44234=>"011011010",
  44235=>"000000101",
  44236=>"110101110",
  44237=>"111111101",
  44238=>"111111111",
  44239=>"111111111",
  44240=>"000000000",
  44241=>"000010000",
  44242=>"111111111",
  44243=>"110110101",
  44244=>"111101111",
  44245=>"111111111",
  44246=>"000000000",
  44247=>"101001110",
  44248=>"001111001",
  44249=>"011000000",
  44250=>"000001011",
  44251=>"111111111",
  44252=>"111011000",
  44253=>"000000000",
  44254=>"110111100",
  44255=>"000000001",
  44256=>"111111000",
  44257=>"111110000",
  44258=>"000000000",
  44259=>"111111111",
  44260=>"000111101",
  44261=>"110111101",
  44262=>"100000111",
  44263=>"001000000",
  44264=>"000000000",
  44265=>"110111000",
  44266=>"000001011",
  44267=>"011001000",
  44268=>"111110000",
  44269=>"111001000",
  44270=>"010011001",
  44271=>"111111011",
  44272=>"111111111",
  44273=>"010001100",
  44274=>"011110000",
  44275=>"000000000",
  44276=>"000100011",
  44277=>"111111001",
  44278=>"101101111",
  44279=>"101111100",
  44280=>"111101101",
  44281=>"000000000",
  44282=>"111111111",
  44283=>"110010001",
  44284=>"111111111",
  44285=>"111111111",
  44286=>"101011111",
  44287=>"111111111",
  44288=>"000010000",
  44289=>"011010100",
  44290=>"100000000",
  44291=>"110000000",
  44292=>"011111001",
  44293=>"110000001",
  44294=>"000000111",
  44295=>"011111111",
  44296=>"000100111",
  44297=>"111010111",
  44298=>"110110101",
  44299=>"001111010",
  44300=>"000111100",
  44301=>"100000011",
  44302=>"000100100",
  44303=>"000000000",
  44304=>"001010110",
  44305=>"010000011",
  44306=>"000100101",
  44307=>"000000111",
  44308=>"100000100",
  44309=>"111101111",
  44310=>"111011010",
  44311=>"111000010",
  44312=>"011000111",
  44313=>"101011000",
  44314=>"000011111",
  44315=>"000000100",
  44316=>"111010000",
  44317=>"101100111",
  44318=>"100101000",
  44319=>"000010010",
  44320=>"000000110",
  44321=>"000100010",
  44322=>"111001000",
  44323=>"000000010",
  44324=>"010110110",
  44325=>"111110000",
  44326=>"000110011",
  44327=>"111101101",
  44328=>"010011111",
  44329=>"000011010",
  44330=>"001000011",
  44331=>"111111010",
  44332=>"101111101",
  44333=>"111101111",
  44334=>"110000111",
  44335=>"111100000",
  44336=>"111000110",
  44337=>"111001100",
  44338=>"110111000",
  44339=>"101011111",
  44340=>"011000111",
  44341=>"000111111",
  44342=>"010000011",
  44343=>"100101001",
  44344=>"100011111",
  44345=>"000000010",
  44346=>"001000000",
  44347=>"111111111",
  44348=>"100110110",
  44349=>"010010010",
  44350=>"000000100",
  44351=>"111111111",
  44352=>"000000010",
  44353=>"101111100",
  44354=>"110000000",
  44355=>"011011100",
  44356=>"101101111",
  44357=>"001001000",
  44358=>"101000011",
  44359=>"110000000",
  44360=>"110101111",
  44361=>"010111111",
  44362=>"000100000",
  44363=>"000010110",
  44364=>"111111111",
  44365=>"000011000",
  44366=>"100110100",
  44367=>"000000000",
  44368=>"010011000",
  44369=>"000000001",
  44370=>"111011000",
  44371=>"001010111",
  44372=>"000000010",
  44373=>"101110100",
  44374=>"010001001",
  44375=>"100000010",
  44376=>"000001001",
  44377=>"001111011",
  44378=>"000011010",
  44379=>"110000000",
  44380=>"111111000",
  44381=>"100100100",
  44382=>"111101111",
  44383=>"100101111",
  44384=>"111101101",
  44385=>"001000000",
  44386=>"001101000",
  44387=>"000111111",
  44388=>"000011001",
  44389=>"110110000",
  44390=>"111111111",
  44391=>"001001000",
  44392=>"101111010",
  44393=>"010101011",
  44394=>"000010111",
  44395=>"111000100",
  44396=>"111110101",
  44397=>"101111111",
  44398=>"101100001",
  44399=>"111010101",
  44400=>"010011101",
  44401=>"100011111",
  44402=>"011000010",
  44403=>"100100100",
  44404=>"100111111",
  44405=>"101000000",
  44406=>"111010010",
  44407=>"101101101",
  44408=>"011000101",
  44409=>"111010000",
  44410=>"111000000",
  44411=>"000010000",
  44412=>"101110010",
  44413=>"000000011",
  44414=>"111011111",
  44415=>"100101011",
  44416=>"010000000",
  44417=>"000011000",
  44418=>"111000111",
  44419=>"111001111",
  44420=>"111111111",
  44421=>"000000101",
  44422=>"011011000",
  44423=>"000011011",
  44424=>"110110110",
  44425=>"001011000",
  44426=>"000000000",
  44427=>"001000111",
  44428=>"111100100",
  44429=>"001000001",
  44430=>"000101111",
  44431=>"100000000",
  44432=>"011011101",
  44433=>"000010111",
  44434=>"000000011",
  44435=>"000010111",
  44436=>"000100111",
  44437=>"010111111",
  44438=>"111111110",
  44439=>"100000000",
  44440=>"101001110",
  44441=>"000001011",
  44442=>"100010000",
  44443=>"001000101",
  44444=>"100000111",
  44445=>"000000000",
  44446=>"111000110",
  44447=>"000111111",
  44448=>"011011001",
  44449=>"111111011",
  44450=>"000000111",
  44451=>"110000111",
  44452=>"111010010",
  44453=>"000000000",
  44454=>"000001111",
  44455=>"000101000",
  44456=>"110000011",
  44457=>"011000000",
  44458=>"011010000",
  44459=>"010100100",
  44460=>"000010000",
  44461=>"011111000",
  44462=>"000100101",
  44463=>"101101101",
  44464=>"111011101",
  44465=>"000110110",
  44466=>"001001111",
  44467=>"011001000",
  44468=>"110110111",
  44469=>"110100011",
  44470=>"001001100",
  44471=>"101111000",
  44472=>"001011001",
  44473=>"000110011",
  44474=>"010010000",
  44475=>"001111111",
  44476=>"100101101",
  44477=>"011011111",
  44478=>"101011100",
  44479=>"011111000",
  44480=>"111111100",
  44481=>"011011000",
  44482=>"010010101",
  44483=>"001100000",
  44484=>"111101111",
  44485=>"110110001",
  44486=>"010010111",
  44487=>"000100111",
  44488=>"100111111",
  44489=>"000100111",
  44490=>"100111011",
  44491=>"000100111",
  44492=>"111100100",
  44493=>"000000010",
  44494=>"010111010",
  44495=>"111101111",
  44496=>"001010000",
  44497=>"001010000",
  44498=>"000000111",
  44499=>"000110000",
  44500=>"111000101",
  44501=>"010011011",
  44502=>"000011010",
  44503=>"111010111",
  44504=>"100101111",
  44505=>"110100000",
  44506=>"001000000",
  44507=>"111000001",
  44508=>"100111011",
  44509=>"101100000",
  44510=>"111101111",
  44511=>"010000111",
  44512=>"111000100",
  44513=>"000111001",
  44514=>"101000101",
  44515=>"010001100",
  44516=>"000000000",
  44517=>"111101000",
  44518=>"010111001",
  44519=>"011011101",
  44520=>"111100100",
  44521=>"111111111",
  44522=>"011011000",
  44523=>"111000101",
  44524=>"011001011",
  44525=>"111010000",
  44526=>"000000000",
  44527=>"001010000",
  44528=>"100100111",
  44529=>"011111100",
  44530=>"000010011",
  44531=>"111111111",
  44532=>"000101011",
  44533=>"001111101",
  44534=>"000000000",
  44535=>"111101001",
  44536=>"010111001",
  44537=>"110001110",
  44538=>"010010110",
  44539=>"011010111",
  44540=>"110111011",
  44541=>"111101111",
  44542=>"100111001",
  44543=>"000010000",
  44544=>"001000000",
  44545=>"000001111",
  44546=>"000110000",
  44547=>"111000101",
  44548=>"110111110",
  44549=>"111110000",
  44550=>"110000000",
  44551=>"001000011",
  44552=>"011011000",
  44553=>"000000000",
  44554=>"011011101",
  44555=>"111110100",
  44556=>"000001111",
  44557=>"011010000",
  44558=>"000011011",
  44559=>"110000000",
  44560=>"101000110",
  44561=>"111111000",
  44562=>"011101101",
  44563=>"000011011",
  44564=>"001000011",
  44565=>"000111111",
  44566=>"110000000",
  44567=>"110010010",
  44568=>"000000000",
  44569=>"000000110",
  44570=>"011010000",
  44571=>"010000100",
  44572=>"101100111",
  44573=>"011100100",
  44574=>"000000000",
  44575=>"000000101",
  44576=>"000000000",
  44577=>"000000010",
  44578=>"010101001",
  44579=>"111011010",
  44580=>"100100100",
  44581=>"101111110",
  44582=>"011011111",
  44583=>"111111010",
  44584=>"110110111",
  44585=>"101000111",
  44586=>"111111000",
  44587=>"111111111",
  44588=>"111011001",
  44589=>"000010010",
  44590=>"111110000",
  44591=>"110010000",
  44592=>"010000010",
  44593=>"101100100",
  44594=>"011000000",
  44595=>"111000010",
  44596=>"000010000",
  44597=>"101111011",
  44598=>"001011011",
  44599=>"000000000",
  44600=>"011000000",
  44601=>"001101000",
  44602=>"000000100",
  44603=>"010010000",
  44604=>"111011011",
  44605=>"111101010",
  44606=>"000111011",
  44607=>"011001111",
  44608=>"010101000",
  44609=>"000101111",
  44610=>"111001111",
  44611=>"011011111",
  44612=>"101000000",
  44613=>"001000000",
  44614=>"000000000",
  44615=>"000000101",
  44616=>"101100110",
  44617=>"101001000",
  44618=>"001000000",
  44619=>"101011010",
  44620=>"111010111",
  44621=>"101111011",
  44622=>"001001111",
  44623=>"000011111",
  44624=>"000111111",
  44625=>"001000000",
  44626=>"001101111",
  44627=>"011100000",
  44628=>"000101111",
  44629=>"111000000",
  44630=>"001001001",
  44631=>"111111111",
  44632=>"100110110",
  44633=>"000100101",
  44634=>"000110110",
  44635=>"011100011",
  44636=>"111111101",
  44637=>"110001001",
  44638=>"010111000",
  44639=>"010110010",
  44640=>"000110010",
  44641=>"111111000",
  44642=>"000010111",
  44643=>"000001001",
  44644=>"101101000",
  44645=>"111000101",
  44646=>"111111010",
  44647=>"000100101",
  44648=>"010000000",
  44649=>"010000001",
  44650=>"000000000",
  44651=>"001111101",
  44652=>"111110000",
  44653=>"111000000",
  44654=>"000000111",
  44655=>"000010010",
  44656=>"110111110",
  44657=>"011010000",
  44658=>"110110100",
  44659=>"110011001",
  44660=>"000000111",
  44661=>"111100010",
  44662=>"110100110",
  44663=>"001111111",
  44664=>"000010111",
  44665=>"000000000",
  44666=>"010000110",
  44667=>"111000000",
  44668=>"001000101",
  44669=>"111000000",
  44670=>"000001000",
  44671=>"000100111",
  44672=>"000000010",
  44673=>"110000000",
  44674=>"111111000",
  44675=>"101111101",
  44676=>"000000001",
  44677=>"111110010",
  44678=>"100110111",
  44679=>"100100011",
  44680=>"001101101",
  44681=>"000110111",
  44682=>"000111111",
  44683=>"010111000",
  44684=>"110111111",
  44685=>"000111110",
  44686=>"111101000",
  44687=>"000010000",
  44688=>"111101100",
  44689=>"100100101",
  44690=>"010100100",
  44691=>"001000100",
  44692=>"000110011",
  44693=>"111110000",
  44694=>"001000000",
  44695=>"011001000",
  44696=>"111101111",
  44697=>"101111111",
  44698=>"000001001",
  44699=>"000000000",
  44700=>"000000000",
  44701=>"111111111",
  44702=>"001000000",
  44703=>"000111111",
  44704=>"101100001",
  44705=>"010000000",
  44706=>"101101000",
  44707=>"111111100",
  44708=>"101000111",
  44709=>"011011100",
  44710=>"001101011",
  44711=>"111110111",
  44712=>"111111100",
  44713=>"101001111",
  44714=>"000000000",
  44715=>"110110110",
  44716=>"110101111",
  44717=>"000111111",
  44718=>"001001001",
  44719=>"000111111",
  44720=>"111100010",
  44721=>"000001111",
  44722=>"000000000",
  44723=>"000110100",
  44724=>"111100101",
  44725=>"000111110",
  44726=>"000101011",
  44727=>"110001111",
  44728=>"111110000",
  44729=>"000011110",
  44730=>"111111000",
  44731=>"110001111",
  44732=>"111111110",
  44733=>"000111111",
  44734=>"110111011",
  44735=>"011000000",
  44736=>"000000111",
  44737=>"110110000",
  44738=>"010000100",
  44739=>"000110100",
  44740=>"111000011",
  44741=>"100100001",
  44742=>"011000110",
  44743=>"000010110",
  44744=>"001111010",
  44745=>"100111111",
  44746=>"100101010",
  44747=>"111111010",
  44748=>"011001000",
  44749=>"100000111",
  44750=>"000000001",
  44751=>"010000111",
  44752=>"111101111",
  44753=>"100011111",
  44754=>"000011111",
  44755=>"010100010",
  44756=>"000010111",
  44757=>"100000000",
  44758=>"101100101",
  44759=>"010100000",
  44760=>"101100111",
  44761=>"011111101",
  44762=>"101110111",
  44763=>"110111010",
  44764=>"011000001",
  44765=>"000111111",
  44766=>"000101100",
  44767=>"010000010",
  44768=>"000010111",
  44769=>"000111111",
  44770=>"111111111",
  44771=>"000111111",
  44772=>"000010111",
  44773=>"101001011",
  44774=>"111011111",
  44775=>"100000111",
  44776=>"110011100",
  44777=>"000010010",
  44778=>"110100100",
  44779=>"110001100",
  44780=>"000110000",
  44781=>"011011111",
  44782=>"010000000",
  44783=>"000000010",
  44784=>"000000000",
  44785=>"001001110",
  44786=>"101000001",
  44787=>"111011000",
  44788=>"110000000",
  44789=>"000101001",
  44790=>"000010011",
  44791=>"000100000",
  44792=>"111000000",
  44793=>"111000000",
  44794=>"101101111",
  44795=>"000111111",
  44796=>"001011111",
  44797=>"110100100",
  44798=>"111111100",
  44799=>"000100111",
  44800=>"011011101",
  44801=>"110011001",
  44802=>"001000000",
  44803=>"110000011",
  44804=>"010100100",
  44805=>"000000110",
  44806=>"110110011",
  44807=>"110111111",
  44808=>"000001001",
  44809=>"000111101",
  44810=>"000100110",
  44811=>"111111100",
  44812=>"001111111",
  44813=>"000000111",
  44814=>"000000010",
  44815=>"111111001",
  44816=>"100111000",
  44817=>"111000000",
  44818=>"000101000",
  44819=>"111001000",
  44820=>"111111011",
  44821=>"111001111",
  44822=>"011111110",
  44823=>"111111111",
  44824=>"001001001",
  44825=>"001110111",
  44826=>"101001101",
  44827=>"000110000",
  44828=>"101000001",
  44829=>"111111000",
  44830=>"110111111",
  44831=>"001111010",
  44832=>"100110000",
  44833=>"000000000",
  44834=>"000000100",
  44835=>"111101111",
  44836=>"110001001",
  44837=>"010011110",
  44838=>"111001001",
  44839=>"001110110",
  44840=>"111110101",
  44841=>"001111111",
  44842=>"001101111",
  44843=>"100000000",
  44844=>"111000100",
  44845=>"111000110",
  44846=>"110000101",
  44847=>"000100100",
  44848=>"111000000",
  44849=>"110100100",
  44850=>"000000001",
  44851=>"011110110",
  44852=>"101110000",
  44853=>"110111110",
  44854=>"000011011",
  44855=>"110111001",
  44856=>"111111111",
  44857=>"000001001",
  44858=>"000000101",
  44859=>"110000000",
  44860=>"000100110",
  44861=>"111111111",
  44862=>"111000001",
  44863=>"010011111",
  44864=>"001000100",
  44865=>"101100000",
  44866=>"000000101",
  44867=>"001110011",
  44868=>"000001000",
  44869=>"010110001",
  44870=>"101011000",
  44871=>"000001000",
  44872=>"111000000",
  44873=>"000000110",
  44874=>"110001111",
  44875=>"000000110",
  44876=>"111001001",
  44877=>"101001000",
  44878=>"001001011",
  44879=>"111001001",
  44880=>"000010110",
  44881=>"111110111",
  44882=>"010101001",
  44883=>"011000100",
  44884=>"010000000",
  44885=>"101111111",
  44886=>"100011001",
  44887=>"001010110",
  44888=>"101001110",
  44889=>"000101111",
  44890=>"000101101",
  44891=>"101001001",
  44892=>"100000000",
  44893=>"000000000",
  44894=>"000110110",
  44895=>"000000100",
  44896=>"001000000",
  44897=>"100010011",
  44898=>"001000000",
  44899=>"100111111",
  44900=>"000000000",
  44901=>"000001010",
  44902=>"000111111",
  44903=>"000111001",
  44904=>"000100111",
  44905=>"111000001",
  44906=>"000000111",
  44907=>"111110110",
  44908=>"111010011",
  44909=>"011000000",
  44910=>"011000111",
  44911=>"111001111",
  44912=>"110100100",
  44913=>"000001101",
  44914=>"001111100",
  44915=>"000000111",
  44916=>"101001111",
  44917=>"011000000",
  44918=>"000001111",
  44919=>"110110001",
  44920=>"001010011",
  44921=>"011011000",
  44922=>"011000011",
  44923=>"000000110",
  44924=>"000110111",
  44925=>"100100000",
  44926=>"000001010",
  44927=>"000000111",
  44928=>"001000110",
  44929=>"100100001",
  44930=>"111000000",
  44931=>"111000001",
  44932=>"111101011",
  44933=>"000100010",
  44934=>"011011101",
  44935=>"000000000",
  44936=>"001001001",
  44937=>"010010010",
  44938=>"010000000",
  44939=>"000000000",
  44940=>"000110001",
  44941=>"101111000",
  44942=>"000110110",
  44943=>"001000001",
  44944=>"011101101",
  44945=>"000111110",
  44946=>"111000001",
  44947=>"100101101",
  44948=>"000110110",
  44949=>"100000100",
  44950=>"000110000",
  44951=>"000000001",
  44952=>"111111111",
  44953=>"111011000",
  44954=>"001111111",
  44955=>"000010000",
  44956=>"110000101",
  44957=>"010110110",
  44958=>"000001111",
  44959=>"101001001",
  44960=>"000000111",
  44961=>"010111110",
  44962=>"000000000",
  44963=>"001000100",
  44964=>"111000000",
  44965=>"101001011",
  44966=>"000000000",
  44967=>"000001111",
  44968=>"111111010",
  44969=>"010000001",
  44970=>"001000000",
  44971=>"001000000",
  44972=>"011000000",
  44973=>"101000000",
  44974=>"100111011",
  44975=>"000110000",
  44976=>"100000110",
  44977=>"111011101",
  44978=>"111010110",
  44979=>"000000100",
  44980=>"010011010",
  44981=>"110100110",
  44982=>"111101000",
  44983=>"000110111",
  44984=>"101011001",
  44985=>"000000100",
  44986=>"000101001",
  44987=>"110011100",
  44988=>"111111111",
  44989=>"111111111",
  44990=>"000100100",
  44991=>"011101111",
  44992=>"000110000",
  44993=>"001000000",
  44994=>"001111011",
  44995=>"001001111",
  44996=>"000000111",
  44997=>"101100001",
  44998=>"110110101",
  44999=>"010111111",
  45000=>"010000101",
  45001=>"111001001",
  45002=>"000000001",
  45003=>"111111110",
  45004=>"000101110",
  45005=>"100000011",
  45006=>"011001000",
  45007=>"001000111",
  45008=>"010001000",
  45009=>"000000001",
  45010=>"000000000",
  45011=>"111100100",
  45012=>"111111111",
  45013=>"101001011",
  45014=>"001001000",
  45015=>"000000000",
  45016=>"001001011",
  45017=>"000000001",
  45018=>"000000011",
  45019=>"011000111",
  45020=>"110111001",
  45021=>"110100110",
  45022=>"111001001",
  45023=>"110111111",
  45024=>"111000001",
  45025=>"011110110",
  45026=>"000110110",
  45027=>"000001001",
  45028=>"000000000",
  45029=>"101000001",
  45030=>"100000000",
  45031=>"011111000",
  45032=>"000101101",
  45033=>"110001000",
  45034=>"011111110",
  45035=>"111000000",
  45036=>"000000001",
  45037=>"111111111",
  45038=>"111001000",
  45039=>"111000001",
  45040=>"110101001",
  45041=>"011110010",
  45042=>"111000000",
  45043=>"101001101",
  45044=>"110110001",
  45045=>"000001111",
  45046=>"100000000",
  45047=>"001001011",
  45048=>"000010111",
  45049=>"101111011",
  45050=>"111001001",
  45051=>"101110000",
  45052=>"111111001",
  45053=>"000010000",
  45054=>"010010011",
  45055=>"111001001",
  45056=>"111000101",
  45057=>"100111111",
  45058=>"000000111",
  45059=>"000011010",
  45060=>"001001111",
  45061=>"101100010",
  45062=>"000100111",
  45063=>"111010001",
  45064=>"100010000",
  45065=>"000111111",
  45066=>"000011011",
  45067=>"010111101",
  45068=>"111000000",
  45069=>"000101111",
  45070=>"100111111",
  45071=>"001010010",
  45072=>"010110000",
  45073=>"000000000",
  45074=>"111110000",
  45075=>"000000000",
  45076=>"101011000",
  45077=>"110000000",
  45078=>"101000010",
  45079=>"010000001",
  45080=>"110111000",
  45081=>"000100000",
  45082=>"000000001",
  45083=>"000111010",
  45084=>"001101000",
  45085=>"111111000",
  45086=>"111000110",
  45087=>"000000111",
  45088=>"000010000",
  45089=>"000011111",
  45090=>"111010001",
  45091=>"111111001",
  45092=>"100001111",
  45093=>"001001000",
  45094=>"000101010",
  45095=>"101001111",
  45096=>"000000010",
  45097=>"010100101",
  45098=>"111000111",
  45099=>"000101011",
  45100=>"111101001",
  45101=>"111111000",
  45102=>"101111111",
  45103=>"011011111",
  45104=>"111001101",
  45105=>"001101011",
  45106=>"111111111",
  45107=>"111010000",
  45108=>"011001111",
  45109=>"111000000",
  45110=>"000000000",
  45111=>"001111111",
  45112=>"110101000",
  45113=>"001000111",
  45114=>"000000110",
  45115=>"101000001",
  45116=>"101001001",
  45117=>"000101101",
  45118=>"000000110",
  45119=>"101100110",
  45120=>"111010000",
  45121=>"010000000",
  45122=>"100000011",
  45123=>"101011101",
  45124=>"101000000",
  45125=>"010000001",
  45126=>"000100111",
  45127=>"111111111",
  45128=>"111011001",
  45129=>"010111010",
  45130=>"111101111",
  45131=>"000000111",
  45132=>"111010111",
  45133=>"011110111",
  45134=>"100101101",
  45135=>"111111110",
  45136=>"000001111",
  45137=>"000010000",
  45138=>"111111111",
  45139=>"100110000",
  45140=>"000100010",
  45141=>"110111111",
  45142=>"000000111",
  45143=>"110111010",
  45144=>"010000000",
  45145=>"000001000",
  45146=>"001011111",
  45147=>"100100101",
  45148=>"111010000",
  45149=>"000001000",
  45150=>"111111000",
  45151=>"011111111",
  45152=>"000000000",
  45153=>"111111111",
  45154=>"100000000",
  45155=>"100100101",
  45156=>"111010000",
  45157=>"000000100",
  45158=>"100111111",
  45159=>"001111111",
  45160=>"101000010",
  45161=>"110000000",
  45162=>"111111100",
  45163=>"110000000",
  45164=>"101000110",
  45165=>"111111000",
  45166=>"111000001",
  45167=>"001111111",
  45168=>"001111111",
  45169=>"000101110",
  45170=>"110000000",
  45171=>"010000001",
  45172=>"111000000",
  45173=>"001000000",
  45174=>"011001111",
  45175=>"000000111",
  45176=>"110111010",
  45177=>"000000111",
  45178=>"111110101",
  45179=>"110111000",
  45180=>"011110100",
  45181=>"111000010",
  45182=>"111111111",
  45183=>"000101111",
  45184=>"111000000",
  45185=>"000111000",
  45186=>"111111000",
  45187=>"111010011",
  45188=>"001110111",
  45189=>"000100000",
  45190=>"000100000",
  45191=>"110100000",
  45192=>"100011111",
  45193=>"000110000",
  45194=>"010010000",
  45195=>"000111101",
  45196=>"000000000",
  45197=>"000111011",
  45198=>"111000000",
  45199=>"000010011",
  45200=>"101111001",
  45201=>"111101010",
  45202=>"000001101",
  45203=>"010111000",
  45204=>"111111010",
  45205=>"100111000",
  45206=>"010001101",
  45207=>"010100100",
  45208=>"010011010",
  45209=>"111010011",
  45210=>"000001000",
  45211=>"100111110",
  45212=>"010011001",
  45213=>"111011000",
  45214=>"010111111",
  45215=>"000000011",
  45216=>"011101111",
  45217=>"110000000",
  45218=>"001111101",
  45219=>"000000000",
  45220=>"111001001",
  45221=>"000000001",
  45222=>"111011001",
  45223=>"100011001",
  45224=>"111111111",
  45225=>"111011001",
  45226=>"111000101",
  45227=>"000000111",
  45228=>"010010111",
  45229=>"000010111",
  45230=>"000001011",
  45231=>"000000011",
  45232=>"101100000",
  45233=>"011000000",
  45234=>"110000000",
  45235=>"001000110",
  45236=>"111111010",
  45237=>"010011111",
  45238=>"111000000",
  45239=>"110000000",
  45240=>"001000100",
  45241=>"001011000",
  45242=>"111111111",
  45243=>"000000100",
  45244=>"011001100",
  45245=>"111000111",
  45246=>"011001001",
  45247=>"010000111",
  45248=>"000100010",
  45249=>"000010110",
  45250=>"111011000",
  45251=>"100100110",
  45252=>"110000111",
  45253=>"110110011",
  45254=>"011000000",
  45255=>"101111100",
  45256=>"111111101",
  45257=>"001000000",
  45258=>"000000000",
  45259=>"110000000",
  45260=>"000010010",
  45261=>"110010001",
  45262=>"000001110",
  45263=>"110011000",
  45264=>"111111010",
  45265=>"011000111",
  45266=>"010111111",
  45267=>"111111111",
  45268=>"100111111",
  45269=>"000100000",
  45270=>"001111111",
  45271=>"010111111",
  45272=>"000000000",
  45273=>"001000000",
  45274=>"101100100",
  45275=>"110110110",
  45276=>"011000100",
  45277=>"000110111",
  45278=>"000000000",
  45279=>"111001100",
  45280=>"000100110",
  45281=>"110111111",
  45282=>"111000000",
  45283=>"000100111",
  45284=>"000000011",
  45285=>"001111010",
  45286=>"111111110",
  45287=>"001000100",
  45288=>"111101101",
  45289=>"010111000",
  45290=>"000110110",
  45291=>"111000111",
  45292=>"110111111",
  45293=>"111011001",
  45294=>"000000010",
  45295=>"111000000",
  45296=>"000001000",
  45297=>"111111110",
  45298=>"001001101",
  45299=>"110111000",
  45300=>"101001011",
  45301=>"000111111",
  45302=>"000000111",
  45303=>"111111000",
  45304=>"111011000",
  45305=>"000101010",
  45306=>"000010001",
  45307=>"001011000",
  45308=>"010000000",
  45309=>"000010000",
  45310=>"110100010",
  45311=>"111111111",
  45312=>"000000001",
  45313=>"110001111",
  45314=>"000000110",
  45315=>"010101001",
  45316=>"100100110",
  45317=>"001000110",
  45318=>"110000111",
  45319=>"111111111",
  45320=>"001001111",
  45321=>"111000011",
  45322=>"001111110",
  45323=>"000000100",
  45324=>"000000000",
  45325=>"000110110",
  45326=>"000000011",
  45327=>"111111000",
  45328=>"111111110",
  45329=>"110111111",
  45330=>"101000000",
  45331=>"011111111",
  45332=>"111111000",
  45333=>"001001011",
  45334=>"010100000",
  45335=>"010011111",
  45336=>"000000011",
  45337=>"011001000",
  45338=>"000100000",
  45339=>"000000000",
  45340=>"000100000",
  45341=>"100100111",
  45342=>"000001111",
  45343=>"010101000",
  45344=>"011111000",
  45345=>"000010000",
  45346=>"011111111",
  45347=>"010011111",
  45348=>"000110010",
  45349=>"101001110",
  45350=>"000110010",
  45351=>"100111110",
  45352=>"011111010",
  45353=>"000001000",
  45354=>"000000000",
  45355=>"000000000",
  45356=>"010011011",
  45357=>"101101000",
  45358=>"111111111",
  45359=>"001000000",
  45360=>"000111000",
  45361=>"111011111",
  45362=>"110111000",
  45363=>"000011111",
  45364=>"111111110",
  45365=>"111101101",
  45366=>"110110010",
  45367=>"001000111",
  45368=>"000001000",
  45369=>"001000000",
  45370=>"100110111",
  45371=>"010110000",
  45372=>"010011001",
  45373=>"010000111",
  45374=>"010000111",
  45375=>"110000000",
  45376=>"111011010",
  45377=>"000011111",
  45378=>"010000111",
  45379=>"101101111",
  45380=>"111110111",
  45381=>"111001000",
  45382=>"001000000",
  45383=>"111000000",
  45384=>"010111111",
  45385=>"010110110",
  45386=>"111111001",
  45387=>"111111111",
  45388=>"000000000",
  45389=>"011011110",
  45390=>"001001001",
  45391=>"000000000",
  45392=>"010000000",
  45393=>"110111110",
  45394=>"111000000",
  45395=>"001001000",
  45396=>"100000111",
  45397=>"111110110",
  45398=>"010011001",
  45399=>"101111000",
  45400=>"000000000",
  45401=>"000000000",
  45402=>"000000100",
  45403=>"011011011",
  45404=>"000000000",
  45405=>"111110000",
  45406=>"000000000",
  45407=>"001100100",
  45408=>"000000000",
  45409=>"010110100",
  45410=>"000110111",
  45411=>"111101000",
  45412=>"001111101",
  45413=>"100000101",
  45414=>"110110110",
  45415=>"001000000",
  45416=>"110001000",
  45417=>"001001111",
  45418=>"100000000",
  45419=>"101000010",
  45420=>"000000000",
  45421=>"101111001",
  45422=>"101000111",
  45423=>"100111111",
  45424=>"110110110",
  45425=>"000000000",
  45426=>"000000100",
  45427=>"000000111",
  45428=>"010110111",
  45429=>"111000111",
  45430=>"100000000",
  45431=>"001101111",
  45432=>"010000110",
  45433=>"000000000",
  45434=>"000111111",
  45435=>"111111101",
  45436=>"011001010",
  45437=>"100000000",
  45438=>"111111011",
  45439=>"100111001",
  45440=>"000000000",
  45441=>"111000000",
  45442=>"000000000",
  45443=>"000001110",
  45444=>"001000111",
  45445=>"000000110",
  45446=>"100110110",
  45447=>"000101001",
  45448=>"011011111",
  45449=>"000010111",
  45450=>"111111111",
  45451=>"001001010",
  45452=>"010000000",
  45453=>"110000111",
  45454=>"001001000",
  45455=>"000000110",
  45456=>"111101101",
  45457=>"000000111",
  45458=>"111111111",
  45459=>"001000110",
  45460=>"100010000",
  45461=>"101000000",
  45462=>"111001001",
  45463=>"110110000",
  45464=>"011101110",
  45465=>"110100010",
  45466=>"000000010",
  45467=>"111000011",
  45468=>"111100000",
  45469=>"111111111",
  45470=>"011111111",
  45471=>"101000001",
  45472=>"000000000",
  45473=>"111100000",
  45474=>"000000100",
  45475=>"000001110",
  45476=>"101001111",
  45477=>"110000000",
  45478=>"011111011",
  45479=>"100001111",
  45480=>"111001000",
  45481=>"000001101",
  45482=>"000000000",
  45483=>"101001000",
  45484=>"011000111",
  45485=>"000000000",
  45486=>"101101100",
  45487=>"011000110",
  45488=>"000000000",
  45489=>"000100101",
  45490=>"010110000",
  45491=>"010000100",
  45492=>"111111111",
  45493=>"000101111",
  45494=>"001000000",
  45495=>"111101111",
  45496=>"101100100",
  45497=>"111111100",
  45498=>"001111101",
  45499=>"011111111",
  45500=>"000110010",
  45501=>"010010000",
  45502=>"110000001",
  45503=>"001000000",
  45504=>"111101100",
  45505=>"001000111",
  45506=>"000111101",
  45507=>"101100110",
  45508=>"001000000",
  45509=>"111101000",
  45510=>"010011000",
  45511=>"111111110",
  45512=>"110000000",
  45513=>"000101111",
  45514=>"001000000",
  45515=>"111111111",
  45516=>"111000101",
  45517=>"100100001",
  45518=>"100101101",
  45519=>"101111111",
  45520=>"000010110",
  45521=>"010010000",
  45522=>"111111000",
  45523=>"111101101",
  45524=>"000000100",
  45525=>"111011111",
  45526=>"101000000",
  45527=>"100000100",
  45528=>"000000001",
  45529=>"100111011",
  45530=>"100000000",
  45531=>"111111110",
  45532=>"000000011",
  45533=>"110111110",
  45534=>"001000000",
  45535=>"001110100",
  45536=>"000000000",
  45537=>"000010111",
  45538=>"111111000",
  45539=>"011111111",
  45540=>"111011111",
  45541=>"111101111",
  45542=>"000000000",
  45543=>"011011011",
  45544=>"111111100",
  45545=>"111011110",
  45546=>"010111111",
  45547=>"101111010",
  45548=>"111111111",
  45549=>"001000000",
  45550=>"010010000",
  45551=>"111111111",
  45552=>"000000000",
  45553=>"011001000",
  45554=>"101000000",
  45555=>"110000000",
  45556=>"001010110",
  45557=>"000100110",
  45558=>"111101000",
  45559=>"000011111",
  45560=>"101111011",
  45561=>"111111111",
  45562=>"000000000",
  45563=>"101000000",
  45564=>"010111011",
  45565=>"000111001",
  45566=>"001011011",
  45567=>"010010011",
  45568=>"000100100",
  45569=>"000000000",
  45570=>"000000001",
  45571=>"000011101",
  45572=>"110100000",
  45573=>"011110000",
  45574=>"111010000",
  45575=>"100100111",
  45576=>"010011001",
  45577=>"111111000",
  45578=>"000000001",
  45579=>"110111111",
  45580=>"000000100",
  45581=>"111111000",
  45582=>"100100000",
  45583=>"111111111",
  45584=>"001000100",
  45585=>"101000101",
  45586=>"001000001",
  45587=>"111111010",
  45588=>"111101111",
  45589=>"001000000",
  45590=>"000011111",
  45591=>"000001000",
  45592=>"010101100",
  45593=>"100100000",
  45594=>"110011000",
  45595=>"000000000",
  45596=>"100000000",
  45597=>"010001000",
  45598=>"111010000",
  45599=>"010010010",
  45600=>"000111001",
  45601=>"111101111",
  45602=>"101101111",
  45603=>"101100110",
  45604=>"010100000",
  45605=>"000011011",
  45606=>"111110000",
  45607=>"111111000",
  45608=>"000000010",
  45609=>"000100111",
  45610=>"111111000",
  45611=>"100011111",
  45612=>"111111100",
  45613=>"000100101",
  45614=>"100000010",
  45615=>"010000111",
  45616=>"111000000",
  45617=>"011011000",
  45618=>"111101101",
  45619=>"111101111",
  45620=>"100000000",
  45621=>"111101111",
  45622=>"000000000",
  45623=>"111111001",
  45624=>"101111111",
  45625=>"111101000",
  45626=>"101110011",
  45627=>"110000011",
  45628=>"111000000",
  45629=>"110111010",
  45630=>"000100000",
  45631=>"001011010",
  45632=>"010101111",
  45633=>"000011001",
  45634=>"000000101",
  45635=>"110011001",
  45636=>"111111011",
  45637=>"010111111",
  45638=>"010011000",
  45639=>"111111001",
  45640=>"011011110",
  45641=>"000000111",
  45642=>"101100110",
  45643=>"111111111",
  45644=>"101111000",
  45645=>"011111101",
  45646=>"110110000",
  45647=>"000000101",
  45648=>"100001001",
  45649=>"000000111",
  45650=>"010010000",
  45651=>"011000000",
  45652=>"000000000",
  45653=>"000100000",
  45654=>"011011000",
  45655=>"000010000",
  45656=>"111111110",
  45657=>"000001001",
  45658=>"110011011",
  45659=>"010110001",
  45660=>"000000011",
  45661=>"001001111",
  45662=>"000000000",
  45663=>"111110000",
  45664=>"010011010",
  45665=>"101000100",
  45666=>"000100100",
  45667=>"111111000",
  45668=>"010010010",
  45669=>"000100100",
  45670=>"000000111",
  45671=>"010000000",
  45672=>"100111111",
  45673=>"111100011",
  45674=>"000000010",
  45675=>"111111101",
  45676=>"101000000",
  45677=>"111000111",
  45678=>"000000111",
  45679=>"111000111",
  45680=>"101101000",
  45681=>"000000111",
  45682=>"000000000",
  45683=>"111111000",
  45684=>"000011111",
  45685=>"000100100",
  45686=>"100000111",
  45687=>"111111111",
  45688=>"111001000",
  45689=>"000011010",
  45690=>"011111110",
  45691=>"000000111",
  45692=>"000000110",
  45693=>"110100000",
  45694=>"000000111",
  45695=>"010110100",
  45696=>"101100100",
  45697=>"000010011",
  45698=>"111000000",
  45699=>"111111001",
  45700=>"111110010",
  45701=>"101101111",
  45702=>"010100110",
  45703=>"110100100",
  45704=>"111100100",
  45705=>"000000000",
  45706=>"000111110",
  45707=>"111000101",
  45708=>"000011111",
  45709=>"010101111",
  45710=>"000100111",
  45711=>"111001110",
  45712=>"100100111",
  45713=>"101111011",
  45714=>"001000010",
  45715=>"111100000",
  45716=>"110000000",
  45717=>"001001101",
  45718=>"111111101",
  45719=>"111101111",
  45720=>"001111010",
  45721=>"000010011",
  45722=>"111111000",
  45723=>"100101100",
  45724=>"011111111",
  45725=>"011111111",
  45726=>"110101101",
  45727=>"110111000",
  45728=>"011010001",
  45729=>"000001100",
  45730=>"111101111",
  45731=>"011001000",
  45732=>"110100100",
  45733=>"011010000",
  45734=>"111110000",
  45735=>"001000100",
  45736=>"111011100",
  45737=>"000011111",
  45738=>"101111111",
  45739=>"101111000",
  45740=>"000000101",
  45741=>"011000001",
  45742=>"100111001",
  45743=>"111000111",
  45744=>"100100111",
  45745=>"110101100",
  45746=>"000000111",
  45747=>"000000100",
  45748=>"111110111",
  45749=>"000010000",
  45750=>"110110110",
  45751=>"000000101",
  45752=>"111111001",
  45753=>"001000001",
  45754=>"000000100",
  45755=>"000100111",
  45756=>"110000011",
  45757=>"000111111",
  45758=>"110110000",
  45759=>"101110111",
  45760=>"000000101",
  45761=>"000000000",
  45762=>"101011111",
  45763=>"111100100",
  45764=>"101100011",
  45765=>"000010111",
  45766=>"111111000",
  45767=>"000000000",
  45768=>"000010000",
  45769=>"000000000",
  45770=>"100000100",
  45771=>"010001111",
  45772=>"000000000",
  45773=>"100100000",
  45774=>"100111010",
  45775=>"000111010",
  45776=>"111011000",
  45777=>"111111110",
  45778=>"110000001",
  45779=>"011101010",
  45780=>"100000001",
  45781=>"000000010",
  45782=>"100111110",
  45783=>"000000011",
  45784=>"000000110",
  45785=>"101100100",
  45786=>"110011100",
  45787=>"101100101",
  45788=>"000100111",
  45789=>"100111111",
  45790=>"111111000",
  45791=>"011111000",
  45792=>"000001010",
  45793=>"000000101",
  45794=>"000010000",
  45795=>"010000000",
  45796=>"100111001",
  45797=>"000100111",
  45798=>"011111111",
  45799=>"011111100",
  45800=>"111101000",
  45801=>"101101010",
  45802=>"001100111",
  45803=>"101101101",
  45804=>"000000100",
  45805=>"010111000",
  45806=>"011010101",
  45807=>"000000000",
  45808=>"111111010",
  45809=>"000011111",
  45810=>"111011000",
  45811=>"011011100",
  45812=>"111110000",
  45813=>"111111010",
  45814=>"101100000",
  45815=>"110101011",
  45816=>"000000111",
  45817=>"000001111",
  45818=>"110100111",
  45819=>"000000000",
  45820=>"010111000",
  45821=>"000000000",
  45822=>"110100110",
  45823=>"000000000",
  45824=>"001001010",
  45825=>"000101110",
  45826=>"000000001",
  45827=>"000000000",
  45828=>"101111111",
  45829=>"000001001",
  45830=>"011111111",
  45831=>"111111111",
  45832=>"000000001",
  45833=>"010110101",
  45834=>"001011011",
  45835=>"001000111",
  45836=>"000000000",
  45837=>"000000000",
  45838=>"000011110",
  45839=>"101111001",
  45840=>"110100111",
  45841=>"000010011",
  45842=>"000001001",
  45843=>"101101100",
  45844=>"101000100",
  45845=>"000111000",
  45846=>"111111110",
  45847=>"111111000",
  45848=>"101001000",
  45849=>"111001001",
  45850=>"000000000",
  45851=>"000000101",
  45852=>"101101111",
  45853=>"101000001",
  45854=>"010010011",
  45855=>"010111110",
  45856=>"111101101",
  45857=>"111111111",
  45858=>"000010111",
  45859=>"111110000",
  45860=>"010001101",
  45861=>"100111010",
  45862=>"110011001",
  45863=>"111110000",
  45864=>"000000000",
  45865=>"000001010",
  45866=>"111111111",
  45867=>"010001101",
  45868=>"000100100",
  45869=>"101010000",
  45870=>"111101111",
  45871=>"011110111",
  45872=>"111000000",
  45873=>"111110110",
  45874=>"001101000",
  45875=>"100000000",
  45876=>"101000111",
  45877=>"111111111",
  45878=>"110111111",
  45879=>"000000000",
  45880=>"111000000",
  45881=>"000000010",
  45882=>"000000000",
  45883=>"101110111",
  45884=>"111001000",
  45885=>"111111000",
  45886=>"001000101",
  45887=>"111111011",
  45888=>"001101111",
  45889=>"010101110",
  45890=>"000000000",
  45891=>"011011100",
  45892=>"111010111",
  45893=>"101000000",
  45894=>"110011001",
  45895=>"101010111",
  45896=>"000011100",
  45897=>"000110101",
  45898=>"100000000",
  45899=>"111110000",
  45900=>"001000110",
  45901=>"000100011",
  45902=>"101001010",
  45903=>"001101100",
  45904=>"001110111",
  45905=>"111111000",
  45906=>"010110011",
  45907=>"011000000",
  45908=>"000000000",
  45909=>"111111100",
  45910=>"101001111",
  45911=>"000010100",
  45912=>"000000011",
  45913=>"001001110",
  45914=>"000011011",
  45915=>"001100100",
  45916=>"111110000",
  45917=>"000000000",
  45918=>"111111111",
  45919=>"110000000",
  45920=>"111111111",
  45921=>"011001000",
  45922=>"000000101",
  45923=>"100010010",
  45924=>"000001100",
  45925=>"000000000",
  45926=>"000000000",
  45927=>"011111111",
  45928=>"101010111",
  45929=>"101001011",
  45930=>"000001111",
  45931=>"100111000",
  45932=>"001101100",
  45933=>"010111111",
  45934=>"000011000",
  45935=>"000000110",
  45936=>"110011011",
  45937=>"000000111",
  45938=>"011011110",
  45939=>"100111000",
  45940=>"111111111",
  45941=>"000000000",
  45942=>"000010101",
  45943=>"000010111",
  45944=>"001010111",
  45945=>"000111111",
  45946=>"001111000",
  45947=>"101101100",
  45948=>"111100000",
  45949=>"110100001",
  45950=>"111111111",
  45951=>"101000000",
  45952=>"110001000",
  45953=>"100100000",
  45954=>"111111110",
  45955=>"000100101",
  45956=>"000101111",
  45957=>"000000000",
  45958=>"110110111",
  45959=>"111110100",
  45960=>"001111111",
  45961=>"110100111",
  45962=>"111110000",
  45963=>"111111111",
  45964=>"010010000",
  45965=>"001000001",
  45966=>"111100011",
  45967=>"000001001",
  45968=>"111111001",
  45969=>"000000111",
  45970=>"110101000",
  45971=>"000000001",
  45972=>"000000100",
  45973=>"000000111",
  45974=>"000010010",
  45975=>"000001011",
  45976=>"011011001",
  45977=>"001000001",
  45978=>"111111010",
  45979=>"100100001",
  45980=>"000000100",
  45981=>"001000111",
  45982=>"111000000",
  45983=>"011111101",
  45984=>"101111100",
  45985=>"100101111",
  45986=>"001000100",
  45987=>"000010001",
  45988=>"010000000",
  45989=>"101001000",
  45990=>"000110000",
  45991=>"001000100",
  45992=>"111111000",
  45993=>"001001000",
  45994=>"000110110",
  45995=>"000000000",
  45996=>"000000001",
  45997=>"000000100",
  45998=>"000101011",
  45999=>"000111110",
  46000=>"000000010",
  46001=>"100000001",
  46002=>"111000000",
  46003=>"000100110",
  46004=>"001011111",
  46005=>"101011101",
  46006=>"011101111",
  46007=>"001000101",
  46008=>"010100000",
  46009=>"011011111",
  46010=>"111111000",
  46011=>"010010101",
  46012=>"010000000",
  46013=>"111010010",
  46014=>"011011111",
  46015=>"000000101",
  46016=>"000010000",
  46017=>"000011001",
  46018=>"101110000",
  46019=>"001001111",
  46020=>"011111000",
  46021=>"001000100",
  46022=>"000000010",
  46023=>"110111011",
  46024=>"100101111",
  46025=>"010111001",
  46026=>"111111111",
  46027=>"101101000",
  46028=>"000000100",
  46029=>"101111101",
  46030=>"101001101",
  46031=>"111111101",
  46032=>"001000111",
  46033=>"001011000",
  46034=>"001101000",
  46035=>"000100101",
  46036=>"010011000",
  46037=>"110100110",
  46038=>"000000010",
  46039=>"000100100",
  46040=>"111110110",
  46041=>"111001100",
  46042=>"111101101",
  46043=>"111010000",
  46044=>"110111101",
  46045=>"000001111",
  46046=>"000101101",
  46047=>"110000000",
  46048=>"000110101",
  46049=>"000000110",
  46050=>"000000111",
  46051=>"111111011",
  46052=>"000010111",
  46053=>"000000101",
  46054=>"101001110",
  46055=>"011111100",
  46056=>"101101000",
  46057=>"011000000",
  46058=>"000110110",
  46059=>"110111010",
  46060=>"100000111",
  46061=>"100101001",
  46062=>"100000000",
  46063=>"111001000",
  46064=>"110101010",
  46065=>"100101001",
  46066=>"010000000",
  46067=>"100101111",
  46068=>"100100100",
  46069=>"000110010",
  46070=>"111111000",
  46071=>"001101111",
  46072=>"111111000",
  46073=>"010000000",
  46074=>"110100111",
  46075=>"101100000",
  46076=>"111110000",
  46077=>"100110011",
  46078=>"001111101",
  46079=>"001000111",
  46080=>"111110101",
  46081=>"000000000",
  46082=>"100000111",
  46083=>"010000000",
  46084=>"100100110",
  46085=>"001000111",
  46086=>"001111001",
  46087=>"000110111",
  46088=>"111001000",
  46089=>"110100111",
  46090=>"110000000",
  46091=>"101100000",
  46092=>"111100111",
  46093=>"000000100",
  46094=>"011110100",
  46095=>"111111000",
  46096=>"000000001",
  46097=>"100100000",
  46098=>"000010111",
  46099=>"000110000",
  46100=>"110110100",
  46101=>"111101111",
  46102=>"000001111",
  46103=>"011111111",
  46104=>"110000000",
  46105=>"111111101",
  46106=>"000101100",
  46107=>"100100111",
  46108=>"000100110",
  46109=>"001010010",
  46110=>"101111000",
  46111=>"111000000",
  46112=>"000111101",
  46113=>"010000001",
  46114=>"001000010",
  46115=>"010010010",
  46116=>"000100011",
  46117=>"010010010",
  46118=>"011011000",
  46119=>"000000000",
  46120=>"111100110",
  46121=>"111101111",
  46122=>"000000110",
  46123=>"100000100",
  46124=>"100100110",
  46125=>"110010011",
  46126=>"010000000",
  46127=>"001011010",
  46128=>"111111000",
  46129=>"110110111",
  46130=>"101111111",
  46131=>"000110101",
  46132=>"111010000",
  46133=>"000000111",
  46134=>"001000000",
  46135=>"010111000",
  46136=>"111001000",
  46137=>"010111001",
  46138=>"101101111",
  46139=>"101000110",
  46140=>"001111001",
  46141=>"111111000",
  46142=>"000000000",
  46143=>"111101001",
  46144=>"000100100",
  46145=>"000000101",
  46146=>"111111000",
  46147=>"000110000",
  46148=>"101111111",
  46149=>"111101011",
  46150=>"001100100",
  46151=>"001100101",
  46152=>"000100101",
  46153=>"010111010",
  46154=>"000000111",
  46155=>"100001001",
  46156=>"001111101",
  46157=>"110110110",
  46158=>"011001111",
  46159=>"101000111",
  46160=>"000000100",
  46161=>"101111100",
  46162=>"100100110",
  46163=>"001100010",
  46164=>"000000110",
  46165=>"110110100",
  46166=>"011011000",
  46167=>"110010000",
  46168=>"000000101",
  46169=>"100000101",
  46170=>"100000010",
  46171=>"010000001",
  46172=>"010111000",
  46173=>"001001000",
  46174=>"010010010",
  46175=>"010001011",
  46176=>"100100111",
  46177=>"001010000",
  46178=>"000000111",
  46179=>"000110100",
  46180=>"111100000",
  46181=>"100100001",
  46182=>"110111110",
  46183=>"110111000",
  46184=>"010010110",
  46185=>"100101111",
  46186=>"010111011",
  46187=>"110110011",
  46188=>"111111111",
  46189=>"100101111",
  46190=>"000100110",
  46191=>"001101111",
  46192=>"010100000",
  46193=>"110001001",
  46194=>"110000000",
  46195=>"001111000",
  46196=>"100111011",
  46197=>"001100111",
  46198=>"110001111",
  46199=>"101000101",
  46200=>"000000110",
  46201=>"000000010",
  46202=>"001111110",
  46203=>"111101011",
  46204=>"110110010",
  46205=>"100000000",
  46206=>"110010111",
  46207=>"000010000",
  46208=>"010000000",
  46209=>"101101010",
  46210=>"000000000",
  46211=>"001000110",
  46212=>"000111111",
  46213=>"010010000",
  46214=>"110100110",
  46215=>"011011000",
  46216=>"111011000",
  46217=>"110010010",
  46218=>"001011010",
  46219=>"000100101",
  46220=>"000000101",
  46221=>"000000001",
  46222=>"011111000",
  46223=>"000000100",
  46224=>"011011011",
  46225=>"000010010",
  46226=>"111000001",
  46227=>"101101111",
  46228=>"010010111",
  46229=>"000000000",
  46230=>"010010000",
  46231=>"111100100",
  46232=>"000000000",
  46233=>"010000110",
  46234=>"111011010",
  46235=>"101000000",
  46236=>"010000111",
  46237=>"101000111",
  46238=>"111010000",
  46239=>"110000111",
  46240=>"101111001",
  46241=>"001001111",
  46242=>"111111000",
  46243=>"111111011",
  46244=>"000000000",
  46245=>"100100100",
  46246=>"001101100",
  46247=>"001001001",
  46248=>"010101111",
  46249=>"000000010",
  46250=>"111101100",
  46251=>"100100111",
  46252=>"000001000",
  46253=>"000010100",
  46254=>"111011001",
  46255=>"100111111",
  46256=>"111000101",
  46257=>"100000001",
  46258=>"111111101",
  46259=>"101110100",
  46260=>"001011001",
  46261=>"111111000",
  46262=>"001000100",
  46263=>"111110010",
  46264=>"001011000",
  46265=>"101100000",
  46266=>"010111111",
  46267=>"000011111",
  46268=>"101101110",
  46269=>"101111111",
  46270=>"001000100",
  46271=>"001100111",
  46272=>"010010000",
  46273=>"000000111",
  46274=>"000111001",
  46275=>"100100100",
  46276=>"010011000",
  46277=>"110100100",
  46278=>"010000000",
  46279=>"000000100",
  46280=>"000000001",
  46281=>"101001111",
  46282=>"111011010",
  46283=>"111100000",
  46284=>"111011111",
  46285=>"101011001",
  46286=>"000000000",
  46287=>"000001000",
  46288=>"000000100",
  46289=>"111111111",
  46290=>"111111111",
  46291=>"111111100",
  46292=>"100000000",
  46293=>"000000000",
  46294=>"000100000",
  46295=>"001111111",
  46296=>"010111011",
  46297=>"000111011",
  46298=>"101101110",
  46299=>"100000111",
  46300=>"000100000",
  46301=>"000000100",
  46302=>"000111100",
  46303=>"010110000",
  46304=>"010010110",
  46305=>"000000111",
  46306=>"001101111",
  46307=>"111000011",
  46308=>"000000100",
  46309=>"101101110",
  46310=>"000000101",
  46311=>"010110110",
  46312=>"000000101",
  46313=>"010111001",
  46314=>"011010010",
  46315=>"111101101",
  46316=>"000000111",
  46317=>"000000111",
  46318=>"000000000",
  46319=>"000000101",
  46320=>"001000000",
  46321=>"011000001",
  46322=>"000000111",
  46323=>"000100100",
  46324=>"010001001",
  46325=>"000010110",
  46326=>"000000000",
  46327=>"100000101",
  46328=>"101000011",
  46329=>"000001010",
  46330=>"111101111",
  46331=>"100110000",
  46332=>"111111000",
  46333=>"011111011",
  46334=>"011011011",
  46335=>"000000000",
  46336=>"011010011",
  46337=>"100100000",
  46338=>"101000111",
  46339=>"000001111",
  46340=>"101001000",
  46341=>"000001010",
  46342=>"111101111",
  46343=>"111111100",
  46344=>"010110110",
  46345=>"111110110",
  46346=>"000100110",
  46347=>"000100010",
  46348=>"000000111",
  46349=>"010010010",
  46350=>"100011011",
  46351=>"101000000",
  46352=>"101100110",
  46353=>"111111111",
  46354=>"101010101",
  46355=>"111101000",
  46356=>"111111111",
  46357=>"010111000",
  46358=>"101101101",
  46359=>"111011001",
  46360=>"000000010",
  46361=>"100100110",
  46362=>"000011001",
  46363=>"010011011",
  46364=>"101001100",
  46365=>"111010101",
  46366=>"010001000",
  46367=>"000010111",
  46368=>"000110010",
  46369=>"000101010",
  46370=>"010111000",
  46371=>"101100101",
  46372=>"010001011",
  46373=>"010000100",
  46374=>"010110010",
  46375=>"011011001",
  46376=>"010111010",
  46377=>"101100010",
  46378=>"001000000",
  46379=>"111100000",
  46380=>"110100111",
  46381=>"000111111",
  46382=>"011010000",
  46383=>"000101001",
  46384=>"110011110",
  46385=>"000001001",
  46386=>"111111100",
  46387=>"110011111",
  46388=>"100000101",
  46389=>"100000000",
  46390=>"011011000",
  46391=>"010000000",
  46392=>"011010010",
  46393=>"101000000",
  46394=>"000111010",
  46395=>"000001101",
  46396=>"011000110",
  46397=>"111111000",
  46398=>"000000010",
  46399=>"001110110",
  46400=>"111111100",
  46401=>"001101110",
  46402=>"111010110",
  46403=>"001000000",
  46404=>"111101101",
  46405=>"001111100",
  46406=>"111000101",
  46407=>"100000000",
  46408=>"000110111",
  46409=>"010010000",
  46410=>"110000101",
  46411=>"110100101",
  46412=>"111111010",
  46413=>"010001010",
  46414=>"000100111",
  46415=>"001101111",
  46416=>"101111000",
  46417=>"010001000",
  46418=>"010000100",
  46419=>"011001101",
  46420=>"101101100",
  46421=>"000000111",
  46422=>"011001010",
  46423=>"100000100",
  46424=>"111111110",
  46425=>"000100110",
  46426=>"001001000",
  46427=>"110100011",
  46428=>"000000000",
  46429=>"000000000",
  46430=>"111001111",
  46431=>"000000001",
  46432=>"101100000",
  46433=>"000000001",
  46434=>"000000000",
  46435=>"101110000",
  46436=>"000000111",
  46437=>"000100010",
  46438=>"011001001",
  46439=>"010010110",
  46440=>"000001101",
  46441=>"111111000",
  46442=>"000000000",
  46443=>"111000000",
  46444=>"010111110",
  46445=>"101111010",
  46446=>"111100100",
  46447=>"000000111",
  46448=>"000001000",
  46449=>"000101111",
  46450=>"011110100",
  46451=>"111000000",
  46452=>"000000000",
  46453=>"011000100",
  46454=>"101110010",
  46455=>"101000000",
  46456=>"001010111",
  46457=>"011100000",
  46458=>"101101101",
  46459=>"000011010",
  46460=>"100100001",
  46461=>"110000000",
  46462=>"111001001",
  46463=>"000010000",
  46464=>"111101100",
  46465=>"100101101",
  46466=>"111000000",
  46467=>"101100010",
  46468=>"011011111",
  46469=>"111001001",
  46470=>"100000001",
  46471=>"011100100",
  46472=>"001011001",
  46473=>"111001000",
  46474=>"111100000",
  46475=>"010000100",
  46476=>"110110011",
  46477=>"111111010",
  46478=>"110000111",
  46479=>"010000000",
  46480=>"011011010",
  46481=>"011001000",
  46482=>"111110001",
  46483=>"010000000",
  46484=>"100010000",
  46485=>"000000010",
  46486=>"101100101",
  46487=>"000001111",
  46488=>"110001010",
  46489=>"011000000",
  46490=>"111111001",
  46491=>"100000010",
  46492=>"111001000",
  46493=>"111001011",
  46494=>"010111110",
  46495=>"101100101",
  46496=>"100110111",
  46497=>"000000000",
  46498=>"011000000",
  46499=>"011000000",
  46500=>"010001011",
  46501=>"011011001",
  46502=>"111111100",
  46503=>"111100101",
  46504=>"100101101",
  46505=>"101100000",
  46506=>"000010000",
  46507=>"001101000",
  46508=>"101100110",
  46509=>"010010010",
  46510=>"110110100",
  46511=>"000001010",
  46512=>"100000010",
  46513=>"110111001",
  46514=>"111011111",
  46515=>"000000100",
  46516=>"111111000",
  46517=>"111000111",
  46518=>"111110100",
  46519=>"010111101",
  46520=>"010110010",
  46521=>"000010101",
  46522=>"010010000",
  46523=>"101000110",
  46524=>"011100000",
  46525=>"111111010",
  46526=>"110011011",
  46527=>"101011100",
  46528=>"100100101",
  46529=>"101000000",
  46530=>"010000000",
  46531=>"001100110",
  46532=>"101101101",
  46533=>"110010001",
  46534=>"011000011",
  46535=>"111001000",
  46536=>"000000110",
  46537=>"111111000",
  46538=>"000101111",
  46539=>"000000101",
  46540=>"011011010",
  46541=>"001000000",
  46542=>"101000000",
  46543=>"000100111",
  46544=>"000010010",
  46545=>"010001110",
  46546=>"010010111",
  46547=>"101101111",
  46548=>"110010010",
  46549=>"111001000",
  46550=>"100111111",
  46551=>"000001111",
  46552=>"000000001",
  46553=>"000001111",
  46554=>"011001111",
  46555=>"101101100",
  46556=>"001101111",
  46557=>"101111011",
  46558=>"111111000",
  46559=>"010111111",
  46560=>"010101100",
  46561=>"001000000",
  46562=>"111111011",
  46563=>"011101111",
  46564=>"110100000",
  46565=>"111111000",
  46566=>"111010000",
  46567=>"001011010",
  46568=>"111000111",
  46569=>"000111111",
  46570=>"001001001",
  46571=>"101100101",
  46572=>"000101101",
  46573=>"101110010",
  46574=>"000110000",
  46575=>"101101000",
  46576=>"111111001",
  46577=>"000110100",
  46578=>"010001101",
  46579=>"001000110",
  46580=>"110110111",
  46581=>"100000000",
  46582=>"000010001",
  46583=>"010000000",
  46584=>"111111111",
  46585=>"110000110",
  46586=>"100111111",
  46587=>"000001101",
  46588=>"001000101",
  46589=>"010110111",
  46590=>"111000010",
  46591=>"001001011",
  46592=>"110100101",
  46593=>"011010000",
  46594=>"001001101",
  46595=>"000000101",
  46596=>"110011010",
  46597=>"110110000",
  46598=>"000000101",
  46599=>"111011101",
  46600=>"000100111",
  46601=>"010010000",
  46602=>"011100100",
  46603=>"111100000",
  46604=>"000111111",
  46605=>"101111011",
  46606=>"100111111",
  46607=>"101001111",
  46608=>"001010111",
  46609=>"000000101",
  46610=>"000010101",
  46611=>"101010000",
  46612=>"000100110",
  46613=>"110111000",
  46614=>"000100010",
  46615=>"101000100",
  46616=>"000001001",
  46617=>"111000110",
  46618=>"101111111",
  46619=>"000101111",
  46620=>"000010111",
  46621=>"100000000",
  46622=>"001000001",
  46623=>"101101100",
  46624=>"001000100",
  46625=>"000101111",
  46626=>"000010000",
  46627=>"010011010",
  46628=>"000100110",
  46629=>"110110110",
  46630=>"011111000",
  46631=>"111000000",
  46632=>"010011010",
  46633=>"110111111",
  46634=>"010100010",
  46635=>"011101111",
  46636=>"111000110",
  46637=>"000000010",
  46638=>"111011110",
  46639=>"010000010",
  46640=>"111000000",
  46641=>"000101111",
  46642=>"000000101",
  46643=>"000010010",
  46644=>"000101000",
  46645=>"011001000",
  46646=>"100110110",
  46647=>"011001011",
  46648=>"111101000",
  46649=>"000010100",
  46650=>"111000000",
  46651=>"010011100",
  46652=>"000000000",
  46653=>"110111000",
  46654=>"001100100",
  46655=>"100100110",
  46656=>"111111110",
  46657=>"111111000",
  46658=>"110000100",
  46659=>"001001000",
  46660=>"000000000",
  46661=>"001001001",
  46662=>"010000010",
  46663=>"111111100",
  46664=>"000000111",
  46665=>"000000011",
  46666=>"000000101",
  46667=>"101101111",
  46668=>"000000100",
  46669=>"100011011",
  46670=>"000100111",
  46671=>"101001111",
  46672=>"000100111",
  46673=>"111010000",
  46674=>"100000000",
  46675=>"000000000",
  46676=>"101000000",
  46677=>"011001111",
  46678=>"001011011",
  46679=>"110010010",
  46680=>"110100111",
  46681=>"000000010",
  46682=>"001110000",
  46683=>"111000000",
  46684=>"000000000",
  46685=>"001001011",
  46686=>"001001011",
  46687=>"001000000",
  46688=>"101000000",
  46689=>"011110110",
  46690=>"000000111",
  46691=>"100011000",
  46692=>"110101000",
  46693=>"110110000",
  46694=>"111111000",
  46695=>"101101000",
  46696=>"000000000",
  46697=>"010010110",
  46698=>"000000110",
  46699=>"000111110",
  46700=>"011111000",
  46701=>"010010000",
  46702=>"011000100",
  46703=>"111111110",
  46704=>"001101011",
  46705=>"111101010",
  46706=>"001001001",
  46707=>"000000001",
  46708=>"010000010",
  46709=>"000000000",
  46710=>"111001111",
  46711=>"101111111",
  46712=>"110111110",
  46713=>"000000100",
  46714=>"000010111",
  46715=>"111110111",
  46716=>"000110111",
  46717=>"010010000",
  46718=>"000000000",
  46719=>"000101111",
  46720=>"111101000",
  46721=>"010001000",
  46722=>"100000111",
  46723=>"000101110",
  46724=>"000010110",
  46725=>"111100100",
  46726=>"111011001",
  46727=>"100000000",
  46728=>"110111011",
  46729=>"101111111",
  46730=>"101010100",
  46731=>"100101100",
  46732=>"000011010",
  46733=>"100101000",
  46734=>"010011111",
  46735=>"001001001",
  46736=>"101100100",
  46737=>"001001001",
  46738=>"000000000",
  46739=>"000000101",
  46740=>"000010110",
  46741=>"010000111",
  46742=>"101110101",
  46743=>"001011010",
  46744=>"010001101",
  46745=>"111100000",
  46746=>"111111100",
  46747=>"000000011",
  46748=>"100000011",
  46749=>"001000000",
  46750=>"000100011",
  46751=>"011000000",
  46752=>"101000011",
  46753=>"101101011",
  46754=>"000010100",
  46755=>"111001000",
  46756=>"000100000",
  46757=>"111000100",
  46758=>"000000000",
  46759=>"000000000",
  46760=>"000000110",
  46761=>"000110111",
  46762=>"111111110",
  46763=>"100000100",
  46764=>"010110110",
  46765=>"000001111",
  46766=>"000100110",
  46767=>"111000111",
  46768=>"011000000",
  46769=>"100000001",
  46770=>"111011111",
  46771=>"000000010",
  46772=>"011011000",
  46773=>"000010010",
  46774=>"110101000",
  46775=>"000011000",
  46776=>"000000001",
  46777=>"000010111",
  46778=>"101000010",
  46779=>"000100111",
  46780=>"111010000",
  46781=>"111111000",
  46782=>"001011011",
  46783=>"101111010",
  46784=>"101000101",
  46785=>"111000000",
  46786=>"100110011",
  46787=>"101111010",
  46788=>"000010000",
  46789=>"001000000",
  46790=>"000000010",
  46791=>"010010001",
  46792=>"001010000",
  46793=>"111101001",
  46794=>"111111000",
  46795=>"101111110",
  46796=>"110010000",
  46797=>"000011111",
  46798=>"101111011",
  46799=>"000111010",
  46800=>"111111010",
  46801=>"110100110",
  46802=>"101000100",
  46803=>"100111111",
  46804=>"010010001",
  46805=>"101111101",
  46806=>"010000111",
  46807=>"101010011",
  46808=>"001000000",
  46809=>"000000110",
  46810=>"101000111",
  46811=>"010000000",
  46812=>"001111001",
  46813=>"111111000",
  46814=>"111101000",
  46815=>"001010110",
  46816=>"101101101",
  46817=>"100100111",
  46818=>"010111110",
  46819=>"000110111",
  46820=>"101000001",
  46821=>"110100000",
  46822=>"111100101",
  46823=>"001011011",
  46824=>"011000000",
  46825=>"010011110",
  46826=>"110000001",
  46827=>"000010000",
  46828=>"011111000",
  46829=>"111111000",
  46830=>"111111000",
  46831=>"110000000",
  46832=>"001110000",
  46833=>"001000111",
  46834=>"011000000",
  46835=>"100000110",
  46836=>"101001011",
  46837=>"101111111",
  46838=>"000010000",
  46839=>"011100101",
  46840=>"001000000",
  46841=>"101000000",
  46842=>"110001111",
  46843=>"000101111",
  46844=>"010010111",
  46845=>"111101001",
  46846=>"011110000",
  46847=>"001000101",
  46848=>"111110111",
  46849=>"011000000",
  46850=>"101000000",
  46851=>"000100111",
  46852=>"100011011",
  46853=>"001011111",
  46854=>"000011111",
  46855=>"111111101",
  46856=>"000011010",
  46857=>"001000101",
  46858=>"001000100",
  46859=>"101100000",
  46860=>"000011111",
  46861=>"000110010",
  46862=>"101100110",
  46863=>"000000100",
  46864=>"111000100",
  46865=>"010010000",
  46866=>"101000000",
  46867=>"111111000",
  46868=>"011000000",
  46869=>"111001010",
  46870=>"001110110",
  46871=>"001011010",
  46872=>"111101101",
  46873=>"000000001",
  46874=>"000011010",
  46875=>"101000000",
  46876=>"101100000",
  46877=>"000001000",
  46878=>"000111101",
  46879=>"000010010",
  46880=>"010000000",
  46881=>"100111111",
  46882=>"000000111",
  46883=>"000111111",
  46884=>"110110110",
  46885=>"111001011",
  46886=>"000011110",
  46887=>"000000110",
  46888=>"011011011",
  46889=>"000000111",
  46890=>"100100000",
  46891=>"010000001",
  46892=>"011000100",
  46893=>"100100010",
  46894=>"000000111",
  46895=>"000001001",
  46896=>"001000111",
  46897=>"011011001",
  46898=>"100110000",
  46899=>"111111111",
  46900=>"111001101",
  46901=>"111101101",
  46902=>"110110011",
  46903=>"111100000",
  46904=>"000000011",
  46905=>"101100000",
  46906=>"000001100",
  46907=>"110000111",
  46908=>"000100000",
  46909=>"111111011",
  46910=>"000000000",
  46911=>"001011100",
  46912=>"100000111",
  46913=>"001000100",
  46914=>"001000000",
  46915=>"101111111",
  46916=>"000101001",
  46917=>"000000000",
  46918=>"111001000",
  46919=>"000011010",
  46920=>"000100111",
  46921=>"111100000",
  46922=>"001101100",
  46923=>"101000000",
  46924=>"111100101",
  46925=>"011011011",
  46926=>"100100000",
  46927=>"000000000",
  46928=>"100110110",
  46929=>"110111111",
  46930=>"000011010",
  46931=>"000011001",
  46932=>"111000000",
  46933=>"011110110",
  46934=>"011011011",
  46935=>"101000000",
  46936=>"000010100",
  46937=>"000001001",
  46938=>"111100001",
  46939=>"001011011",
  46940=>"100000000",
  46941=>"011010000",
  46942=>"100111011",
  46943=>"011101101",
  46944=>"000000000",
  46945=>"111110111",
  46946=>"111100000",
  46947=>"110110000",
  46948=>"110000010",
  46949=>"001000100",
  46950=>"111000000",
  46951=>"110101101",
  46952=>"010000101",
  46953=>"111111001",
  46954=>"100111111",
  46955=>"000001110",
  46956=>"011001000",
  46957=>"111010010",
  46958=>"001100111",
  46959=>"001000100",
  46960=>"111100001",
  46961=>"000000011",
  46962=>"001011101",
  46963=>"000111111",
  46964=>"000100110",
  46965=>"111000100",
  46966=>"101000000",
  46967=>"100000010",
  46968=>"000000000",
  46969=>"010000001",
  46970=>"010000100",
  46971=>"111111011",
  46972=>"011111100",
  46973=>"001010000",
  46974=>"111010000",
  46975=>"111101101",
  46976=>"000000000",
  46977=>"111111110",
  46978=>"101000000",
  46979=>"100000111",
  46980=>"010111111",
  46981=>"101000000",
  46982=>"111100110",
  46983=>"111000001",
  46984=>"000111000",
  46985=>"111000000",
  46986=>"011110000",
  46987=>"001011110",
  46988=>"000000010",
  46989=>"111101001",
  46990=>"111101000",
  46991=>"011000101",
  46992=>"110100111",
  46993=>"000000110",
  46994=>"110000011",
  46995=>"101101111",
  46996=>"010010010",
  46997=>"000111111",
  46998=>"001000000",
  46999=>"000000011",
  47000=>"111101000",
  47001=>"000101010",
  47002=>"000111011",
  47003=>"101011000",
  47004=>"011100100",
  47005=>"111100100",
  47006=>"000100100",
  47007=>"111100100",
  47008=>"000001000",
  47009=>"010000000",
  47010=>"111001101",
  47011=>"010000000",
  47012=>"010011111",
  47013=>"000000001",
  47014=>"000110110",
  47015=>"111111101",
  47016=>"000111010",
  47017=>"010000000",
  47018=>"001110011",
  47019=>"111000100",
  47020=>"000000010",
  47021=>"000010010",
  47022=>"111101000",
  47023=>"101010111",
  47024=>"000000100",
  47025=>"000110000",
  47026=>"000100111",
  47027=>"000100100",
  47028=>"110001001",
  47029=>"000001101",
  47030=>"000000100",
  47031=>"011111000",
  47032=>"000001001",
  47033=>"100111111",
  47034=>"111101000",
  47035=>"100111101",
  47036=>"110111000",
  47037=>"000010111",
  47038=>"000110011",
  47039=>"000100111",
  47040=>"101000000",
  47041=>"111000111",
  47042=>"000001000",
  47043=>"101110111",
  47044=>"110000000",
  47045=>"101000100",
  47046=>"111111111",
  47047=>"111111011",
  47048=>"011001000",
  47049=>"100101000",
  47050=>"000011100",
  47051=>"000000000",
  47052=>"111100100",
  47053=>"100101101",
  47054=>"101101101",
  47055=>"000111111",
  47056=>"100111011",
  47057=>"010100110",
  47058=>"011000000",
  47059=>"000101010",
  47060=>"111000000",
  47061=>"110011011",
  47062=>"000100000",
  47063=>"000000011",
  47064=>"111000000",
  47065=>"111111101",
  47066=>"000011111",
  47067=>"011101101",
  47068=>"001011011",
  47069=>"000011011",
  47070=>"000000101",
  47071=>"101111111",
  47072=>"000000000",
  47073=>"101000111",
  47074=>"000111111",
  47075=>"111101001",
  47076=>"111000101",
  47077=>"111000101",
  47078=>"000000111",
  47079=>"110011000",
  47080=>"111111001",
  47081=>"111111111",
  47082=>"001100000",
  47083=>"000000000",
  47084=>"010111111",
  47085=>"000111111",
  47086=>"010000000",
  47087=>"001000010",
  47088=>"110111000",
  47089=>"000010001",
  47090=>"000000111",
  47091=>"100110111",
  47092=>"011011100",
  47093=>"111000000",
  47094=>"000000100",
  47095=>"011001000",
  47096=>"001111111",
  47097=>"111111001",
  47098=>"001000000",
  47099=>"110110000",
  47100=>"111110010",
  47101=>"111111100",
  47102=>"101111001",
  47103=>"111100100",
  47104=>"001001001",
  47105=>"100101000",
  47106=>"101000000",
  47107=>"010101101",
  47108=>"111000001",
  47109=>"011101101",
  47110=>"111101000",
  47111=>"110111110",
  47112=>"011000101",
  47113=>"110011000",
  47114=>"111000100",
  47115=>"000111111",
  47116=>"111110111",
  47117=>"100110010",
  47118=>"100000100",
  47119=>"000000111",
  47120=>"000110011",
  47121=>"000000000",
  47122=>"000000000",
  47123=>"111001100",
  47124=>"111000000",
  47125=>"000000111",
  47126=>"001000000",
  47127=>"001010010",
  47128=>"111000000",
  47129=>"000110110",
  47130=>"000101111",
  47131=>"000000000",
  47132=>"001000000",
  47133=>"000000101",
  47134=>"110111101",
  47135=>"101000111",
  47136=>"101101000",
  47137=>"011110001",
  47138=>"101010010",
  47139=>"000000110",
  47140=>"111111110",
  47141=>"010001000",
  47142=>"000010111",
  47143=>"000010111",
  47144=>"110010111",
  47145=>"000110010",
  47146=>"000110111",
  47147=>"010000000",
  47148=>"000011010",
  47149=>"000011111",
  47150=>"000110111",
  47151=>"000101100",
  47152=>"110111000",
  47153=>"111101001",
  47154=>"000111000",
  47155=>"111101000",
  47156=>"110000011",
  47157=>"000101001",
  47158=>"010110111",
  47159=>"000000110",
  47160=>"110111100",
  47161=>"111000001",
  47162=>"000000111",
  47163=>"000000000",
  47164=>"000110011",
  47165=>"111011111",
  47166=>"000000101",
  47167=>"100101110",
  47168=>"111000100",
  47169=>"001101000",
  47170=>"101111100",
  47171=>"000000011",
  47172=>"000000110",
  47173=>"000000001",
  47174=>"000000000",
  47175=>"111000000",
  47176=>"000111111",
  47177=>"010000000",
  47178=>"111001100",
  47179=>"111111101",
  47180=>"111111000",
  47181=>"100001111",
  47182=>"101001110",
  47183=>"111110111",
  47184=>"111001111",
  47185=>"111111000",
  47186=>"100111000",
  47187=>"000111000",
  47188=>"000000100",
  47189=>"000110111",
  47190=>"111111111",
  47191=>"000111010",
  47192=>"110000010",
  47193=>"000000001",
  47194=>"110000000",
  47195=>"000111101",
  47196=>"000000000",
  47197=>"000000000",
  47198=>"000011011",
  47199=>"111000000",
  47200=>"000011111",
  47201=>"010000000",
  47202=>"111000000",
  47203=>"011011000",
  47204=>"001000001",
  47205=>"100111010",
  47206=>"000000111",
  47207=>"001000000",
  47208=>"011101101",
  47209=>"111111111",
  47210=>"101111111",
  47211=>"000101111",
  47212=>"000111111",
  47213=>"111000010",
  47214=>"111100000",
  47215=>"001101000",
  47216=>"000110100",
  47217=>"000000111",
  47218=>"000010111",
  47219=>"011000000",
  47220=>"001001000",
  47221=>"010001100",
  47222=>"000000111",
  47223=>"000001000",
  47224=>"110111000",
  47225=>"011000100",
  47226=>"010000001",
  47227=>"101000001",
  47228=>"000000001",
  47229=>"000110000",
  47230=>"000111111",
  47231=>"111000011",
  47232=>"011111101",
  47233=>"111101000",
  47234=>"000011011",
  47235=>"000000111",
  47236=>"111110111",
  47237=>"101111000",
  47238=>"100111100",
  47239=>"111000100",
  47240=>"100100001",
  47241=>"000000001",
  47242=>"111110001",
  47243=>"101111011",
  47244=>"111010000",
  47245=>"111101000",
  47246=>"100000000",
  47247=>"111000001",
  47248=>"011001100",
  47249=>"000000000",
  47250=>"000111001",
  47251=>"000111101",
  47252=>"111000110",
  47253=>"000111000",
  47254=>"111111000",
  47255=>"010000001",
  47256=>"110111111",
  47257=>"110100000",
  47258=>"000110111",
  47259=>"101110000",
  47260=>"111111110",
  47261=>"000010010",
  47262=>"111111000",
  47263=>"100101111",
  47264=>"011001100",
  47265=>"011000000",
  47266=>"000101111",
  47267=>"111000000",
  47268=>"000111101",
  47269=>"010000001",
  47270=>"000000111",
  47271=>"010011111",
  47272=>"000000010",
  47273=>"000000100",
  47274=>"100000010",
  47275=>"101001001",
  47276=>"001001010",
  47277=>"011110111",
  47278=>"000000111",
  47279=>"111111111",
  47280=>"000000000",
  47281=>"111000011",
  47282=>"000111011",
  47283=>"101000100",
  47284=>"000000001",
  47285=>"101111010",
  47286=>"000001000",
  47287=>"101111011",
  47288=>"001011010",
  47289=>"011001001",
  47290=>"011000000",
  47291=>"010111110",
  47292=>"010101101",
  47293=>"111011011",
  47294=>"000000001",
  47295=>"011101000",
  47296=>"010110111",
  47297=>"101111000",
  47298=>"111111111",
  47299=>"100101111",
  47300=>"000110111",
  47301=>"001011001",
  47302=>"010111101",
  47303=>"111000000",
  47304=>"011111011",
  47305=>"000000000",
  47306=>"101000000",
  47307=>"111101100",
  47308=>"000010011",
  47309=>"100000110",
  47310=>"111000101",
  47311=>"111101000",
  47312=>"100000111",
  47313=>"101000100",
  47314=>"011000001",
  47315=>"000000000",
  47316=>"000010110",
  47317=>"111001111",
  47318=>"111101111",
  47319=>"000111011",
  47320=>"000111111",
  47321=>"011000111",
  47322=>"101000000",
  47323=>"111111000",
  47324=>"000110000",
  47325=>"110001010",
  47326=>"010001011",
  47327=>"100110111",
  47328=>"111000000",
  47329=>"111001111",
  47330=>"111111111",
  47331=>"001000100",
  47332=>"111000101",
  47333=>"110000000",
  47334=>"000110000",
  47335=>"000000000",
  47336=>"100111111",
  47337=>"011000101",
  47338=>"001000011",
  47339=>"111001000",
  47340=>"000010011",
  47341=>"010111111",
  47342=>"111000001",
  47343=>"000010111",
  47344=>"000111101",
  47345=>"110011111",
  47346=>"000111111",
  47347=>"000000110",
  47348=>"011110110",
  47349=>"111101000",
  47350=>"101000000",
  47351=>"010111111",
  47352=>"000110010",
  47353=>"010111101",
  47354=>"001000000",
  47355=>"001001111",
  47356=>"000010111",
  47357=>"111100000",
  47358=>"100100100",
  47359=>"010110110",
  47360=>"001001101",
  47361=>"111111000",
  47362=>"000000101",
  47363=>"000001000",
  47364=>"000011011",
  47365=>"000000110",
  47366=>"000110100",
  47367=>"000110110",
  47368=>"000110000",
  47369=>"011001101",
  47370=>"010010010",
  47371=>"101111000",
  47372=>"100111110",
  47373=>"101100000",
  47374=>"000111011",
  47375=>"101100000",
  47376=>"110111111",
  47377=>"111000111",
  47378=>"100000000",
  47379=>"000000010",
  47380=>"110000100",
  47381=>"111000000",
  47382=>"000010011",
  47383=>"101000111",
  47384=>"001000000",
  47385=>"111011000",
  47386=>"000000010",
  47387=>"001111111",
  47388=>"101110000",
  47389=>"100000000",
  47390=>"111000011",
  47391=>"011001000",
  47392=>"010011111",
  47393=>"000000110",
  47394=>"111000010",
  47395=>"111100011",
  47396=>"100111011",
  47397=>"101101010",
  47398=>"111010000",
  47399=>"000100100",
  47400=>"111000000",
  47401=>"000111100",
  47402=>"000000000",
  47403=>"101111010",
  47404=>"100111111",
  47405=>"111001111",
  47406=>"000100011",
  47407=>"000100001",
  47408=>"111000000",
  47409=>"001100100",
  47410=>"111010001",
  47411=>"000100110",
  47412=>"101001111",
  47413=>"111100111",
  47414=>"000000011",
  47415=>"011110000",
  47416=>"111000110",
  47417=>"000100110",
  47418=>"100000000",
  47419=>"111111111",
  47420=>"011111110",
  47421=>"111111101",
  47422=>"000000101",
  47423=>"110110111",
  47424=>"100100111",
  47425=>"000110110",
  47426=>"001000011",
  47427=>"001110100",
  47428=>"000001000",
  47429=>"100110100",
  47430=>"000100110",
  47431=>"000101101",
  47432=>"111001101",
  47433=>"101011111",
  47434=>"000110110",
  47435=>"101111111",
  47436=>"000000011",
  47437=>"011011110",
  47438=>"000001011",
  47439=>"101001110",
  47440=>"000001000",
  47441=>"111111111",
  47442=>"111010111",
  47443=>"001001000",
  47444=>"110000000",
  47445=>"110100110",
  47446=>"001001110",
  47447=>"111011101",
  47448=>"000001000",
  47449=>"000100110",
  47450=>"011101100",
  47451=>"011000000",
  47452=>"010111000",
  47453=>"000001001",
  47454=>"111011000",
  47455=>"111000000",
  47456=>"000000010",
  47457=>"111000111",
  47458=>"000000111",
  47459=>"100011111",
  47460=>"000110101",
  47461=>"000000101",
  47462=>"000111100",
  47463=>"110000000",
  47464=>"110011100",
  47465=>"111000111",
  47466=>"000000111",
  47467=>"000000110",
  47468=>"010010111",
  47469=>"111111000",
  47470=>"000000000",
  47471=>"001111110",
  47472=>"110001011",
  47473=>"010000000",
  47474=>"001100110",
  47475=>"010000000",
  47476=>"000000010",
  47477=>"001000000",
  47478=>"000100000",
  47479=>"000010000",
  47480=>"000110000",
  47481=>"011111010",
  47482=>"110111001",
  47483=>"111111101",
  47484=>"101101101",
  47485=>"100100000",
  47486=>"110000000",
  47487=>"111000000",
  47488=>"000000000",
  47489=>"010000010",
  47490=>"010010000",
  47491=>"011110110",
  47492=>"101101111",
  47493=>"110011100",
  47494=>"001100110",
  47495=>"011101100",
  47496=>"011111110",
  47497=>"101111110",
  47498=>"011011001",
  47499=>"101100000",
  47500=>"111000000",
  47501=>"110000000",
  47502=>"111110000",
  47503=>"000101000",
  47504=>"001001011",
  47505=>"000111111",
  47506=>"111001000",
  47507=>"000110101",
  47508=>"011001111",
  47509=>"010000101",
  47510=>"010111010",
  47511=>"011010100",
  47512=>"110010000",
  47513=>"111111101",
  47514=>"111011001",
  47515=>"000000000",
  47516=>"000001010",
  47517=>"100110010",
  47518=>"000000111",
  47519=>"000101111",
  47520=>"000010011",
  47521=>"010111111",
  47522=>"000111101",
  47523=>"011111000",
  47524=>"100110111",
  47525=>"100110010",
  47526=>"110110000",
  47527=>"000111100",
  47528=>"010010011",
  47529=>"000000010",
  47530=>"111000000",
  47531=>"000000000",
  47532=>"010111111",
  47533=>"000000111",
  47534=>"100100111",
  47535=>"011010000",
  47536=>"110110000",
  47537=>"011011011",
  47538=>"000001000",
  47539=>"100100001",
  47540=>"111111010",
  47541=>"010010000",
  47542=>"010011100",
  47543=>"001001000",
  47544=>"110111100",
  47545=>"000111010",
  47546=>"010000000",
  47547=>"011011110",
  47548=>"010001000",
  47549=>"000000000",
  47550=>"011010011",
  47551=>"110000000",
  47552=>"001101011",
  47553=>"010010011",
  47554=>"111110000",
  47555=>"001001110",
  47556=>"000101000",
  47557=>"100101101",
  47558=>"110000000",
  47559=>"000001101",
  47560=>"000000111",
  47561=>"000111010",
  47562=>"010110000",
  47563=>"111110010",
  47564=>"000011010",
  47565=>"000100000",
  47566=>"010000000",
  47567=>"111110111",
  47568=>"001111111",
  47569=>"000111111",
  47570=>"111101110",
  47571=>"101000000",
  47572=>"011000000",
  47573=>"110111100",
  47574=>"000000111",
  47575=>"000011111",
  47576=>"111000000",
  47577=>"011100000",
  47578=>"000000110",
  47579=>"111000000",
  47580=>"010110110",
  47581=>"111100000",
  47582=>"111010000",
  47583=>"010001101",
  47584=>"000111111",
  47585=>"110100101",
  47586=>"111011000",
  47587=>"100110111",
  47588=>"000000000",
  47589=>"110011111",
  47590=>"000100111",
  47591=>"010011011",
  47592=>"000000001",
  47593=>"010011000",
  47594=>"111011011",
  47595=>"010010000",
  47596=>"111010000",
  47597=>"000001000",
  47598=>"111001000",
  47599=>"011000000",
  47600=>"110100000",
  47601=>"011001111",
  47602=>"001000000",
  47603=>"000010001",
  47604=>"110110111",
  47605=>"001011010",
  47606=>"001000000",
  47607=>"111111000",
  47608=>"010011000",
  47609=>"000000000",
  47610=>"111101100",
  47611=>"000101111",
  47612=>"010111101",
  47613=>"111000000",
  47614=>"010111111",
  47615=>"000111111",
  47616=>"100100110",
  47617=>"000000110",
  47618=>"011000111",
  47619=>"001000100",
  47620=>"001000001",
  47621=>"111010000",
  47622=>"111001000",
  47623=>"110010111",
  47624=>"001011011",
  47625=>"000110010",
  47626=>"001100100",
  47627=>"101111010",
  47628=>"111000000",
  47629=>"010011000",
  47630=>"110001001",
  47631=>"111000001",
  47632=>"000111101",
  47633=>"000111100",
  47634=>"111000001",
  47635=>"000101111",
  47636=>"001110111",
  47637=>"001000110",
  47638=>"111010001",
  47639=>"111111111",
  47640=>"110000000",
  47641=>"000001111",
  47642=>"000100110",
  47643=>"000100000",
  47644=>"100000010",
  47645=>"111000000",
  47646=>"111111011",
  47647=>"010101000",
  47648=>"011000000",
  47649=>"000010000",
  47650=>"111100000",
  47651=>"000001000",
  47652=>"010000001",
  47653=>"001100110",
  47654=>"101100111",
  47655=>"000110010",
  47656=>"010000000",
  47657=>"010100010",
  47658=>"000101111",
  47659=>"000010110",
  47660=>"010110001",
  47661=>"000000110",
  47662=>"101111001",
  47663=>"010101111",
  47664=>"111110000",
  47665=>"111100000",
  47666=>"000001101",
  47667=>"111111110",
  47668=>"011001100",
  47669=>"000000000",
  47670=>"001001000",
  47671=>"000010000",
  47672=>"111111010",
  47673=>"110010111",
  47674=>"111000101",
  47675=>"000001111",
  47676=>"011001001",
  47677=>"000010000",
  47678=>"000000011",
  47679=>"001011111",
  47680=>"111111111",
  47681=>"100100100",
  47682=>"001001111",
  47683=>"001000101",
  47684=>"100010110",
  47685=>"010011001",
  47686=>"111111000",
  47687=>"011111100",
  47688=>"100010001",
  47689=>"000111110",
  47690=>"000110000",
  47691=>"001011101",
  47692=>"111111100",
  47693=>"001001000",
  47694=>"010000100",
  47695=>"100111111",
  47696=>"111101000",
  47697=>"001000000",
  47698=>"000111000",
  47699=>"111111000",
  47700=>"000000000",
  47701=>"010001101",
  47702=>"110101101",
  47703=>"010111111",
  47704=>"001011111",
  47705=>"111001001",
  47706=>"010100100",
  47707=>"100110110",
  47708=>"000011011",
  47709=>"110000001",
  47710=>"110000111",
  47711=>"011001000",
  47712=>"000101111",
  47713=>"000000110",
  47714=>"101001111",
  47715=>"110110001",
  47716=>"111000000",
  47717=>"011110001",
  47718=>"000110110",
  47719=>"111001000",
  47720=>"110111000",
  47721=>"000111111",
  47722=>"110010101",
  47723=>"111001110",
  47724=>"000101101",
  47725=>"100001011",
  47726=>"111111000",
  47727=>"101000000",
  47728=>"111011000",
  47729=>"101110110",
  47730=>"100110000",
  47731=>"111101111",
  47732=>"111010000",
  47733=>"110001000",
  47734=>"000000110",
  47735=>"000101111",
  47736=>"110100100",
  47737=>"111111110",
  47738=>"010000010",
  47739=>"110000000",
  47740=>"110110100",
  47741=>"011011000",
  47742=>"001111010",
  47743=>"111101101",
  47744=>"111111000",
  47745=>"110010000",
  47746=>"000101111",
  47747=>"000111100",
  47748=>"111111010",
  47749=>"110101100",
  47750=>"000001111",
  47751=>"000011101",
  47752=>"110100000",
  47753=>"010000000",
  47754=>"111101000",
  47755=>"100101000",
  47756=>"110010000",
  47757=>"111000001",
  47758=>"101111000",
  47759=>"001001111",
  47760=>"111000100",
  47761=>"111001000",
  47762=>"000010111",
  47763=>"111111001",
  47764=>"111111001",
  47765=>"110000110",
  47766=>"110111111",
  47767=>"010001001",
  47768=>"000101111",
  47769=>"110000111",
  47770=>"111010111",
  47771=>"110000101",
  47772=>"110011011",
  47773=>"000110110",
  47774=>"101111100",
  47775=>"111110110",
  47776=>"110001001",
  47777=>"000101000",
  47778=>"001011000",
  47779=>"000111111",
  47780=>"111110011",
  47781=>"011001001",
  47782=>"011011111",
  47783=>"000101001",
  47784=>"000111101",
  47785=>"000100111",
  47786=>"111110001",
  47787=>"111010010",
  47788=>"111001000",
  47789=>"111100111",
  47790=>"011001000",
  47791=>"000111111",
  47792=>"110000000",
  47793=>"110111000",
  47794=>"010000101",
  47795=>"000000100",
  47796=>"110100000",
  47797=>"110111101",
  47798=>"000000000",
  47799=>"111001011",
  47800=>"100100000",
  47801=>"110110111",
  47802=>"100000000",
  47803=>"111111000",
  47804=>"101000000",
  47805=>"000111111",
  47806=>"100110110",
  47807=>"101000000",
  47808=>"111001100",
  47809=>"000111111",
  47810=>"111110110",
  47811=>"110100000",
  47812=>"000000001",
  47813=>"111010010",
  47814=>"111100011",
  47815=>"100110111",
  47816=>"111111001",
  47817=>"010000000",
  47818=>"111111111",
  47819=>"000111111",
  47820=>"101111111",
  47821=>"001011001",
  47822=>"111111000",
  47823=>"000000000",
  47824=>"000000111",
  47825=>"111110101",
  47826=>"010010010",
  47827=>"111100100",
  47828=>"101110010",
  47829=>"011011100",
  47830=>"111111111",
  47831=>"000011110",
  47832=>"000101111",
  47833=>"111101100",
  47834=>"011001101",
  47835=>"111101000",
  47836=>"110110101",
  47837=>"111000111",
  47838=>"101101010",
  47839=>"100111110",
  47840=>"000001101",
  47841=>"111011000",
  47842=>"111000101",
  47843=>"111011000",
  47844=>"000000100",
  47845=>"000111010",
  47846=>"111111111",
  47847=>"100100001",
  47848=>"010111111",
  47849=>"110000000",
  47850=>"100000011",
  47851=>"000101111",
  47852=>"111101001",
  47853=>"111001101",
  47854=>"000000000",
  47855=>"010000000",
  47856=>"111101000",
  47857=>"111011111",
  47858=>"100110000",
  47859=>"010010101",
  47860=>"011011001",
  47861=>"010000000",
  47862=>"100100011",
  47863=>"011010000",
  47864=>"000010101",
  47865=>"001001100",
  47866=>"111110000",
  47867=>"010110101",
  47868=>"111110111",
  47869=>"000000111",
  47870=>"011000000",
  47871=>"000111010",
  47872=>"111101100",
  47873=>"001101100",
  47874=>"001000000",
  47875=>"111001001",
  47876=>"010001000",
  47877=>"000000001",
  47878=>"111111000",
  47879=>"000010110",
  47880=>"111110000",
  47881=>"000010000",
  47882=>"001001000",
  47883=>"101000100",
  47884=>"111000101",
  47885=>"110110001",
  47886=>"001011000",
  47887=>"001101110",
  47888=>"010000010",
  47889=>"000000001",
  47890=>"000000011",
  47891=>"110111110",
  47892=>"111111100",
  47893=>"000001001",
  47894=>"111101101",
  47895=>"101000011",
  47896=>"100111000",
  47897=>"111111000",
  47898=>"010000000",
  47899=>"000100101",
  47900=>"000111111",
  47901=>"000001101",
  47902=>"110000111",
  47903=>"101001000",
  47904=>"000111000",
  47905=>"111101111",
  47906=>"111100000",
  47907=>"111111010",
  47908=>"011011000",
  47909=>"100101100",
  47910=>"110010000",
  47911=>"100010010",
  47912=>"001001100",
  47913=>"110010000",
  47914=>"001000010",
  47915=>"001000111",
  47916=>"111111100",
  47917=>"000010110",
  47918=>"111010101",
  47919=>"001000111",
  47920=>"001001110",
  47921=>"101000000",
  47922=>"000000000",
  47923=>"001001101",
  47924=>"000000111",
  47925=>"101000000",
  47926=>"100110101",
  47927=>"000000111",
  47928=>"010011110",
  47929=>"100000000",
  47930=>"010000000",
  47931=>"101111000",
  47932=>"100100011",
  47933=>"011111101",
  47934=>"000000100",
  47935=>"011111000",
  47936=>"101001000",
  47937=>"010111101",
  47938=>"111111111",
  47939=>"000100110",
  47940=>"100111101",
  47941=>"010000010",
  47942=>"111100000",
  47943=>"110010110",
  47944=>"111010110",
  47945=>"000101111",
  47946=>"000000001",
  47947=>"110100000",
  47948=>"010110000",
  47949=>"011101000",
  47950=>"001100000",
  47951=>"001111111",
  47952=>"101001000",
  47953=>"001011111",
  47954=>"111101111",
  47955=>"011001101",
  47956=>"001000110",
  47957=>"000000010",
  47958=>"100111110",
  47959=>"111111000",
  47960=>"010000110",
  47961=>"110110010",
  47962=>"100100000",
  47963=>"110110000",
  47964=>"000000000",
  47965=>"001000000",
  47966=>"010110110",
  47967=>"000001000",
  47968=>"110111000",
  47969=>"011001111",
  47970=>"010000000",
  47971=>"111001000",
  47972=>"001111000",
  47973=>"001011101",
  47974=>"000111010",
  47975=>"000000000",
  47976=>"111111000",
  47977=>"000000010",
  47978=>"110010111",
  47979=>"111001011",
  47980=>"000111000",
  47981=>"000000111",
  47982=>"111100110",
  47983=>"000110110",
  47984=>"101100100",
  47985=>"111101101",
  47986=>"011011101",
  47987=>"001001000",
  47988=>"010000100",
  47989=>"000000000",
  47990=>"111110111",
  47991=>"111000000",
  47992=>"000000110",
  47993=>"010111010",
  47994=>"111111111",
  47995=>"011000111",
  47996=>"110110100",
  47997=>"100100100",
  47998=>"011100010",
  47999=>"001000000",
  48000=>"111110110",
  48001=>"111001000",
  48002=>"110000111",
  48003=>"111101110",
  48004=>"100000011",
  48005=>"111110110",
  48006=>"001000011",
  48007=>"011011000",
  48008=>"101111000",
  48009=>"000001101",
  48010=>"000000000",
  48011=>"111111111",
  48012=>"001000101",
  48013=>"101000001",
  48014=>"001010110",
  48015=>"001001000",
  48016=>"111100000",
  48017=>"001001001",
  48018=>"110111000",
  48019=>"000000111",
  48020=>"011000100",
  48021=>"111110110",
  48022=>"110110110",
  48023=>"011011011",
  48024=>"001011101",
  48025=>"000111111",
  48026=>"010111000",
  48027=>"100000110",
  48028=>"010111000",
  48029=>"000110111",
  48030=>"000010111",
  48031=>"111111101",
  48032=>"111110010",
  48033=>"111000111",
  48034=>"111110110",
  48035=>"000000000",
  48036=>"010001011",
  48037=>"011111100",
  48038=>"011110101",
  48039=>"010111010",
  48040=>"000001111",
  48041=>"000110111",
  48042=>"001000000",
  48043=>"000010001",
  48044=>"111000110",
  48045=>"110010000",
  48046=>"100101100",
  48047=>"001000000",
  48048=>"001000000",
  48049=>"110100000",
  48050=>"011010000",
  48051=>"000110000",
  48052=>"101111111",
  48053=>"000001101",
  48054=>"100001000",
  48055=>"101110111",
  48056=>"001011000",
  48057=>"110110101",
  48058=>"110000000",
  48059=>"110110000",
  48060=>"100000010",
  48061=>"101111111",
  48062=>"110110000",
  48063=>"000000101",
  48064=>"110100000",
  48065=>"001001100",
  48066=>"010000111",
  48067=>"111101000",
  48068=>"000010000",
  48069=>"000001011",
  48070=>"000011000",
  48071=>"010000000",
  48072=>"101111010",
  48073=>"000000000",
  48074=>"001000000",
  48075=>"000111111",
  48076=>"000111111",
  48077=>"111011001",
  48078=>"101111101",
  48079=>"110111100",
  48080=>"001000111",
  48081=>"010110100",
  48082=>"111111000",
  48083=>"000000111",
  48084=>"000010111",
  48085=>"011001110",
  48086=>"110000111",
  48087=>"110000000",
  48088=>"110000111",
  48089=>"000000001",
  48090=>"111111000",
  48091=>"000000101",
  48092=>"000001100",
  48093=>"101000000",
  48094=>"000000000",
  48095=>"000001010",
  48096=>"000000001",
  48097=>"101001111",
  48098=>"001000111",
  48099=>"111011100",
  48100=>"111101100",
  48101=>"111010000",
  48102=>"111100001",
  48103=>"011011011",
  48104=>"000001000",
  48105=>"000000111",
  48106=>"001000101",
  48107=>"111000001",
  48108=>"000000001",
  48109=>"000000000",
  48110=>"010000000",
  48111=>"101100100",
  48112=>"101101001",
  48113=>"010000010",
  48114=>"110010100",
  48115=>"011011110",
  48116=>"111111001",
  48117=>"010011000",
  48118=>"000010010",
  48119=>"101000110",
  48120=>"000111111",
  48121=>"010010110",
  48122=>"111000001",
  48123=>"110010000",
  48124=>"101111010",
  48125=>"000000110",
  48126=>"100111000",
  48127=>"001001111",
  48128=>"100000000",
  48129=>"101000000",
  48130=>"000000000",
  48131=>"001000111",
  48132=>"000011011",
  48133=>"001011111",
  48134=>"111100100",
  48135=>"111000100",
  48136=>"000000011",
  48137=>"001000000",
  48138=>"100010011",
  48139=>"100100110",
  48140=>"010011010",
  48141=>"001011000",
  48142=>"100100110",
  48143=>"111101011",
  48144=>"111010001",
  48145=>"001011111",
  48146=>"101001101",
  48147=>"011110000",
  48148=>"011001000",
  48149=>"100111010",
  48150=>"000111010",
  48151=>"110111111",
  48152=>"111101000",
  48153=>"110000000",
  48154=>"100000000",
  48155=>"000010010",
  48156=>"100000000",
  48157=>"100100111",
  48158=>"000100111",
  48159=>"000000100",
  48160=>"111101111",
  48161=>"000010100",
  48162=>"100101111",
  48163=>"000100001",
  48164=>"010010000",
  48165=>"100001000",
  48166=>"111100000",
  48167=>"001110101",
  48168=>"011000000",
  48169=>"001000011",
  48170=>"101100000",
  48171=>"000010111",
  48172=>"000011001",
  48173=>"101010010",
  48174=>"010010111",
  48175=>"000111101",
  48176=>"101111111",
  48177=>"011001000",
  48178=>"111111101",
  48179=>"110100000",
  48180=>"000010000",
  48181=>"111111111",
  48182=>"101111100",
  48183=>"000100101",
  48184=>"000111100",
  48185=>"101101101",
  48186=>"111111101",
  48187=>"000110000",
  48188=>"000001001",
  48189=>"101111101",
  48190=>"000000111",
  48191=>"001000010",
  48192=>"100111111",
  48193=>"001100110",
  48194=>"000000011",
  48195=>"100100000",
  48196=>"000010000",
  48197=>"000101110",
  48198=>"010000000",
  48199=>"001000111",
  48200=>"101010001",
  48201=>"001000000",
  48202=>"101101100",
  48203=>"111100101",
  48204=>"000100101",
  48205=>"111011001",
  48206=>"101110100",
  48207=>"010000000",
  48208=>"111000000",
  48209=>"111000100",
  48210=>"000000101",
  48211=>"000000001",
  48212=>"000000001",
  48213=>"011001101",
  48214=>"000100010",
  48215=>"111100100",
  48216=>"000000101",
  48217=>"000000101",
  48218=>"000000000",
  48219=>"000110010",
  48220=>"010000000",
  48221=>"000010000",
  48222=>"010111000",
  48223=>"100100100",
  48224=>"100100001",
  48225=>"001000000",
  48226=>"000011100",
  48227=>"001011001",
  48228=>"011000111",
  48229=>"001111111",
  48230=>"110011100",
  48231=>"100000011",
  48232=>"110101000",
  48233=>"011111111",
  48234=>"111111100",
  48235=>"001100100",
  48236=>"000101111",
  48237=>"000101110",
  48238=>"000000000",
  48239=>"100000100",
  48240=>"000110110",
  48241=>"000011100",
  48242=>"010011011",
  48243=>"111101111",
  48244=>"011000000",
  48245=>"101111010",
  48246=>"000111111",
  48247=>"000100011",
  48248=>"000001000",
  48249=>"011011101",
  48250=>"111111111",
  48251=>"111111101",
  48252=>"011001000",
  48253=>"000001000",
  48254=>"111111110",
  48255=>"111100110",
  48256=>"100101110",
  48257=>"000000000",
  48258=>"000011000",
  48259=>"100100111",
  48260=>"000010000",
  48261=>"111111111",
  48262=>"000100100",
  48263=>"010000000",
  48264=>"001001100",
  48265=>"000000110",
  48266=>"111101000",
  48267=>"000011111",
  48268=>"111100000",
  48269=>"111101111",
  48270=>"000000010",
  48271=>"111000001",
  48272=>"101110001",
  48273=>"010111101",
  48274=>"000100100",
  48275=>"010000000",
  48276=>"111000100",
  48277=>"111010000",
  48278=>"100000000",
  48279=>"110010001",
  48280=>"101001110",
  48281=>"111000000",
  48282=>"000011001",
  48283=>"000010011",
  48284=>"111100000",
  48285=>"000000000",
  48286=>"001000011",
  48287=>"000100101",
  48288=>"010100110",
  48289=>"001000101",
  48290=>"100001111",
  48291=>"000000101",
  48292=>"000000011",
  48293=>"110101101",
  48294=>"100000110",
  48295=>"000111111",
  48296=>"100111000",
  48297=>"000000110",
  48298=>"000011011",
  48299=>"000000010",
  48300=>"010100111",
  48301=>"111000001",
  48302=>"100100100",
  48303=>"111111111",
  48304=>"110011011",
  48305=>"111110001",
  48306=>"000000010",
  48307=>"000000001",
  48308=>"001001011",
  48309=>"101111000",
  48310=>"000000100",
  48311=>"000011111",
  48312=>"000000000",
  48313=>"010000000",
  48314=>"111011010",
  48315=>"101111111",
  48316=>"110100000",
  48317=>"011111111",
  48318=>"010000000",
  48319=>"001111111",
  48320=>"111000000",
  48321=>"101100000",
  48322=>"111001000",
  48323=>"110000000",
  48324=>"100100111",
  48325=>"011001111",
  48326=>"000011000",
  48327=>"111011101",
  48328=>"010100101",
  48329=>"000100111",
  48330=>"000000100",
  48331=>"000100000",
  48332=>"111100011",
  48333=>"110000100",
  48334=>"000010011",
  48335=>"011000010",
  48336=>"100111111",
  48337=>"101110110",
  48338=>"100000100",
  48339=>"111111111",
  48340=>"000000000",
  48341=>"011011011",
  48342=>"000000000",
  48343=>"001000001",
  48344=>"100100000",
  48345=>"000100000",
  48346=>"110001101",
  48347=>"011111111",
  48348=>"110111110",
  48349=>"111011011",
  48350=>"101101000",
  48351=>"000100111",
  48352=>"100000000",
  48353=>"001011011",
  48354=>"011010011",
  48355=>"010100101",
  48356=>"001000000",
  48357=>"000011010",
  48358=>"111111111",
  48359=>"000101100",
  48360=>"010111101",
  48361=>"111111000",
  48362=>"001001000",
  48363=>"001000000",
  48364=>"100000000",
  48365=>"000100100",
  48366=>"101010100",
  48367=>"000000111",
  48368=>"000000101",
  48369=>"010100011",
  48370=>"100000111",
  48371=>"100100000",
  48372=>"001001100",
  48373=>"111011000",
  48374=>"000000101",
  48375=>"000010010",
  48376=>"011111000",
  48377=>"010111011",
  48378=>"111111110",
  48379=>"000000111",
  48380=>"100100000",
  48381=>"000111110",
  48382=>"111111111",
  48383=>"100000100",
  48384=>"010000010",
  48385=>"000011111",
  48386=>"000000000",
  48387=>"000110111",
  48388=>"111101000",
  48389=>"111000010",
  48390=>"111111111",
  48391=>"111101101",
  48392=>"000101111",
  48393=>"000000100",
  48394=>"000100000",
  48395=>"101000100",
  48396=>"110000000",
  48397=>"111011011",
  48398=>"010100100",
  48399=>"111010000",
  48400=>"100011010",
  48401=>"000000110",
  48402=>"000111000",
  48403=>"011000011",
  48404=>"010010000",
  48405=>"000000111",
  48406=>"000011111",
  48407=>"000111111",
  48408=>"111000100",
  48409=>"111010000",
  48410=>"000000111",
  48411=>"000111111",
  48412=>"101111111",
  48413=>"000000011",
  48414=>"010000011",
  48415=>"010011111",
  48416=>"111000010",
  48417=>"010011000",
  48418=>"000111101",
  48419=>"010010000",
  48420=>"000111111",
  48421=>"000001011",
  48422=>"000100111",
  48423=>"000100000",
  48424=>"011111100",
  48425=>"000100000",
  48426=>"100110000",
  48427=>"111101001",
  48428=>"111011010",
  48429=>"100100000",
  48430=>"000100010",
  48431=>"000000101",
  48432=>"101100000",
  48433=>"000000011",
  48434=>"000000000",
  48435=>"111111100",
  48436=>"000000010",
  48437=>"001100100",
  48438=>"011011011",
  48439=>"100000100",
  48440=>"111010000",
  48441=>"011111011",
  48442=>"000000000",
  48443=>"110111000",
  48444=>"111011001",
  48445=>"011111000",
  48446=>"100100001",
  48447=>"101101110",
  48448=>"111101000",
  48449=>"100111111",
  48450=>"111100001",
  48451=>"111100000",
  48452=>"111111000",
  48453=>"000100100",
  48454=>"111111011",
  48455=>"010111111",
  48456=>"000111001",
  48457=>"111110111",
  48458=>"000000000",
  48459=>"000100001",
  48460=>"000000000",
  48461=>"000111111",
  48462=>"111111010",
  48463=>"000000000",
  48464=>"010010011",
  48465=>"111111110",
  48466=>"111001111",
  48467=>"001000000",
  48468=>"100100111",
  48469=>"101111111",
  48470=>"001111110",
  48471=>"101100111",
  48472=>"000000001",
  48473=>"011001000",
  48474=>"101111111",
  48475=>"011111111",
  48476=>"000011010",
  48477=>"000000000",
  48478=>"001111010",
  48479=>"100101100",
  48480=>"111001010",
  48481=>"111000000",
  48482=>"101100111",
  48483=>"100110110",
  48484=>"000010010",
  48485=>"000000001",
  48486=>"000011011",
  48487=>"100000000",
  48488=>"111111000",
  48489=>"000000001",
  48490=>"010101111",
  48491=>"111101000",
  48492=>"000000000",
  48493=>"000100110",
  48494=>"010000000",
  48495=>"000000011",
  48496=>"111111111",
  48497=>"010000000",
  48498=>"111110011",
  48499=>"100000010",
  48500=>"000000101",
  48501=>"100100000",
  48502=>"111011111",
  48503=>"110100111",
  48504=>"110000000",
  48505=>"010110110",
  48506=>"000111111",
  48507=>"100100101",
  48508=>"010001001",
  48509=>"100000011",
  48510=>"110011000",
  48511=>"101100100",
  48512=>"011010000",
  48513=>"111000000",
  48514=>"100011111",
  48515=>"000000100",
  48516=>"111100111",
  48517=>"010100000",
  48518=>"111110111",
  48519=>"011010010",
  48520=>"111001011",
  48521=>"001000000",
  48522=>"111100101",
  48523=>"100100101",
  48524=>"011011000",
  48525=>"000000010",
  48526=>"101000000",
  48527=>"100000001",
  48528=>"110111110",
  48529=>"001011111",
  48530=>"011011000",
  48531=>"011101010",
  48532=>"111001100",
  48533=>"100000100",
  48534=>"000010011",
  48535=>"100000000",
  48536=>"000010000",
  48537=>"111001001",
  48538=>"100110000",
  48539=>"100100100",
  48540=>"111011011",
  48541=>"111101000",
  48542=>"111011111",
  48543=>"100100001",
  48544=>"100111011",
  48545=>"000111010",
  48546=>"010111111",
  48547=>"110100100",
  48548=>"000000100",
  48549=>"111010000",
  48550=>"001111011",
  48551=>"000000011",
  48552=>"010011111",
  48553=>"000000000",
  48554=>"100000100",
  48555=>"100000111",
  48556=>"000011000",
  48557=>"101000110",
  48558=>"100110010",
  48559=>"111110100",
  48560=>"001010000",
  48561=>"100111100",
  48562=>"000100000",
  48563=>"000010001",
  48564=>"000000000",
  48565=>"011111000",
  48566=>"011011000",
  48567=>"011000110",
  48568=>"011010110",
  48569=>"110111001",
  48570=>"111111010",
  48571=>"010111111",
  48572=>"111101000",
  48573=>"111111110",
  48574=>"001001101",
  48575=>"010000001",
  48576=>"000000000",
  48577=>"000000000",
  48578=>"011001000",
  48579=>"000111111",
  48580=>"000100100",
  48581=>"010110111",
  48582=>"010111011",
  48583=>"000000011",
  48584=>"101000000",
  48585=>"000000000",
  48586=>"111011000",
  48587=>"011011111",
  48588=>"000000101",
  48589=>"000010011",
  48590=>"000011011",
  48591=>"000100111",
  48592=>"110000010",
  48593=>"100010110",
  48594=>"111100111",
  48595=>"011000000",
  48596=>"111101110",
  48597=>"000100000",
  48598=>"000100110",
  48599=>"100000111",
  48600=>"000000000",
  48601=>"000000000",
  48602=>"000010111",
  48603=>"100000000",
  48604=>"100110111",
  48605=>"100010111",
  48606=>"111011000",
  48607=>"111010010",
  48608=>"011011011",
  48609=>"101100011",
  48610=>"111110110",
  48611=>"101111111",
  48612=>"100100100",
  48613=>"000101110",
  48614=>"111000011",
  48615=>"000110110",
  48616=>"011000000",
  48617=>"000001111",
  48618=>"001000000",
  48619=>"010010100",
  48620=>"000111101",
  48621=>"111011001",
  48622=>"000100111",
  48623=>"000000000",
  48624=>"100100100",
  48625=>"000101111",
  48626=>"000101111",
  48627=>"110000011",
  48628=>"110111001",
  48629=>"111100111",
  48630=>"010000100",
  48631=>"000100001",
  48632=>"011111110",
  48633=>"111100000",
  48634=>"010000000",
  48635=>"000000001",
  48636=>"001000010",
  48637=>"000100000",
  48638=>"000111001",
  48639=>"101000000",
  48640=>"110110000",
  48641=>"000000001",
  48642=>"000000000",
  48643=>"010000000",
  48644=>"000111101",
  48645=>"011001001",
  48646=>"111000000",
  48647=>"110101001",
  48648=>"101111000",
  48649=>"011000000",
  48650=>"110011011",
  48651=>"000001111",
  48652=>"000000000",
  48653=>"110111101",
  48654=>"011100100",
  48655=>"000010000",
  48656=>"111000001",
  48657=>"000000000",
  48658=>"100111000",
  48659=>"010000001",
  48660=>"000110010",
  48661=>"011000111",
  48662=>"000000111",
  48663=>"011111101",
  48664=>"010000000",
  48665=>"000001111",
  48666=>"111111100",
  48667=>"000000000",
  48668=>"010000000",
  48669=>"111111101",
  48670=>"001011100",
  48671=>"011111000",
  48672=>"000010000",
  48673=>"000000000",
  48674=>"101010101",
  48675=>"101000010",
  48676=>"111110111",
  48677=>"011011011",
  48678=>"011111110",
  48679=>"000110000",
  48680=>"000000001",
  48681=>"000111101",
  48682=>"100111001",
  48683=>"000000000",
  48684=>"111110000",
  48685=>"010000000",
  48686=>"111101101",
  48687=>"000000000",
  48688=>"010111100",
  48689=>"110110111",
  48690=>"100111101",
  48691=>"111111101",
  48692=>"111111000",
  48693=>"010110000",
  48694=>"000100100",
  48695=>"111000001",
  48696=>"101011100",
  48697=>"110000110",
  48698=>"000111010",
  48699=>"000100111",
  48700=>"111010000",
  48701=>"111010001",
  48702=>"000000000",
  48703=>"000101110",
  48704=>"101000000",
  48705=>"001111101",
  48706=>"110001001",
  48707=>"000000001",
  48708=>"000110110",
  48709=>"000000000",
  48710=>"010111000",
  48711=>"000111111",
  48712=>"010110110",
  48713=>"000000010",
  48714=>"000001000",
  48715=>"000000000",
  48716=>"101111000",
  48717=>"100101111",
  48718=>"001111111",
  48719=>"101101101",
  48720=>"111000000",
  48721=>"001000111",
  48722=>"000100101",
  48723=>"000100000",
  48724=>"010111111",
  48725=>"011011011",
  48726=>"100100010",
  48727=>"000010111",
  48728=>"000111011",
  48729=>"011011110",
  48730=>"100000000",
  48731=>"010011001",
  48732=>"111110111",
  48733=>"000110100",
  48734=>"000010010",
  48735=>"000000000",
  48736=>"111111111",
  48737=>"110010000",
  48738=>"111001111",
  48739=>"001000011",
  48740=>"000000110",
  48741=>"111011000",
  48742=>"110000000",
  48743=>"111111000",
  48744=>"010110111",
  48745=>"011110111",
  48746=>"111110000",
  48747=>"110111111",
  48748=>"000000011",
  48749=>"111111001",
  48750=>"000000000",
  48751=>"000000000",
  48752=>"100110110",
  48753=>"000111100",
  48754=>"100000001",
  48755=>"110000000",
  48756=>"011000001",
  48757=>"111111110",
  48758=>"000110100",
  48759=>"111100000",
  48760=>"000111111",
  48761=>"000010110",
  48762=>"001010001",
  48763=>"010110110",
  48764=>"001000100",
  48765=>"111011111",
  48766=>"000011101",
  48767=>"000000000",
  48768=>"101001010",
  48769=>"000000001",
  48770=>"111111110",
  48771=>"111000110",
  48772=>"101001000",
  48773=>"100000000",
  48774=>"100100110",
  48775=>"110000000",
  48776=>"000000111",
  48777=>"011000000",
  48778=>"111011011",
  48779=>"000101110",
  48780=>"000101001",
  48781=>"111111111",
  48782=>"000001110",
  48783=>"110000110",
  48784=>"111110000",
  48785=>"010000000",
  48786=>"111110000",
  48787=>"001001000",
  48788=>"010100000",
  48789=>"101000000",
  48790=>"111111111",
  48791=>"010010000",
  48792=>"010111111",
  48793=>"011111101",
  48794=>"011010111",
  48795=>"101101000",
  48796=>"111010000",
  48797=>"000000100",
  48798=>"101111111",
  48799=>"101001000",
  48800=>"010110110",
  48801=>"000111101",
  48802=>"110111000",
  48803=>"101000000",
  48804=>"111001111",
  48805=>"100000110",
  48806=>"000000000",
  48807=>"000111000",
  48808=>"000000000",
  48809=>"000111111",
  48810=>"111001011",
  48811=>"101000000",
  48812=>"101001000",
  48813=>"111000011",
  48814=>"101110010",
  48815=>"111000000",
  48816=>"000000000",
  48817=>"111100000",
  48818=>"000010111",
  48819=>"101101011",
  48820=>"010111111",
  48821=>"010010000",
  48822=>"010111111",
  48823=>"111111000",
  48824=>"110001110",
  48825=>"001001000",
  48826=>"010000101",
  48827=>"101111111",
  48828=>"111010110",
  48829=>"001001111",
  48830=>"100110011",
  48831=>"110111010",
  48832=>"000001111",
  48833=>"111000001",
  48834=>"001000110",
  48835=>"111000101",
  48836=>"000110111",
  48837=>"111001011",
  48838=>"000010001",
  48839=>"000111111",
  48840=>"000100101",
  48841=>"000000010",
  48842=>"000000111",
  48843=>"000110110",
  48844=>"110111001",
  48845=>"100000011",
  48846=>"000011011",
  48847=>"111110010",
  48848=>"111111001",
  48849=>"111011110",
  48850=>"000000010",
  48851=>"111111011",
  48852=>"000000000",
  48853=>"011011001",
  48854=>"000000110",
  48855=>"110011111",
  48856=>"110111000",
  48857=>"111110000",
  48858=>"000001111",
  48859=>"000011000",
  48860=>"000100010",
  48861=>"111111101",
  48862=>"000111111",
  48863=>"111000000",
  48864=>"101010010",
  48865=>"100000000",
  48866=>"111110000",
  48867=>"000111011",
  48868=>"110110101",
  48869=>"010011000",
  48870=>"111111001",
  48871=>"101001111",
  48872=>"111000111",
  48873=>"001111110",
  48874=>"011111100",
  48875=>"001001111",
  48876=>"111101111",
  48877=>"011111101",
  48878=>"011000011",
  48879=>"000000000",
  48880=>"000000000",
  48881=>"011110100",
  48882=>"101101000",
  48883=>"100110000",
  48884=>"111001000",
  48885=>"010000000",
  48886=>"010111111",
  48887=>"111000101",
  48888=>"000110110",
  48889=>"000000001",
  48890=>"000000100",
  48891=>"010010010",
  48892=>"111000111",
  48893=>"011111000",
  48894=>"011011111",
  48895=>"111101001",
  48896=>"000001000",
  48897=>"011011010",
  48898=>"100001110",
  48899=>"111100110",
  48900=>"111100100",
  48901=>"111111011",
  48902=>"000000110",
  48903=>"001110110",
  48904=>"111110111",
  48905=>"011011000",
  48906=>"000000110",
  48907=>"110110100",
  48908=>"011111111",
  48909=>"111011000",
  48910=>"111100000",
  48911=>"100111101",
  48912=>"001010010",
  48913=>"100011111",
  48914=>"110100001",
  48915=>"100011011",
  48916=>"100100001",
  48917=>"000011011",
  48918=>"010011011",
  48919=>"111100100",
  48920=>"000001100",
  48921=>"011001111",
  48922=>"011011010",
  48923=>"011001011",
  48924=>"001110011",
  48925=>"000000010",
  48926=>"011011000",
  48927=>"000000100",
  48928=>"100100001",
  48929=>"000010100",
  48930=>"110010001",
  48931=>"000011011",
  48932=>"110110100",
  48933=>"100101101",
  48934=>"011011010",
  48935=>"111010111",
  48936=>"100111100",
  48937=>"100100100",
  48938=>"011111011",
  48939=>"011000001",
  48940=>"001000001",
  48941=>"111010111",
  48942=>"011010101",
  48943=>"100000100",
  48944=>"011010001",
  48945=>"100100100",
  48946=>"001111101",
  48947=>"011111001",
  48948=>"000101001",
  48949=>"001011000",
  48950=>"011011010",
  48951=>"011010011",
  48952=>"011001000",
  48953=>"001011000",
  48954=>"100100100",
  48955=>"011011111",
  48956=>"100001101",
  48957=>"100100101",
  48958=>"001011011",
  48959=>"111111101",
  48960=>"001000011",
  48961=>"111011011",
  48962=>"110111011",
  48963=>"000011110",
  48964=>"101011011",
  48965=>"110000000",
  48966=>"000111111",
  48967=>"110000111",
  48968=>"110111111",
  48969=>"100110111",
  48970=>"101100011",
  48971=>"001000111",
  48972=>"111011011",
  48973=>"101100100",
  48974=>"100100101",
  48975=>"100100111",
  48976=>"110000110",
  48977=>"000100100",
  48978=>"010111111",
  48979=>"001000011",
  48980=>"110000000",
  48981=>"001111101",
  48982=>"100100100",
  48983=>"000011000",
  48984=>"111001000",
  48985=>"111110011",
  48986=>"101101101",
  48987=>"000000111",
  48988=>"011011011",
  48989=>"001000000",
  48990=>"011010011",
  48991=>"011010011",
  48992=>"011011011",
  48993=>"011011011",
  48994=>"100001011",
  48995=>"111111000",
  48996=>"100100101",
  48997=>"001100101",
  48998=>"000111000",
  48999=>"101000000",
  49000=>"011011000",
  49001=>"010011001",
  49002=>"110110111",
  49003=>"110010101",
  49004=>"111111101",
  49005=>"100100101",
  49006=>"000000001",
  49007=>"000000011",
  49008=>"001111110",
  49009=>"011011111",
  49010=>"000011011",
  49011=>"110100111",
  49012=>"011010111",
  49013=>"000000011",
  49014=>"011011010",
  49015=>"011111011",
  49016=>"111011000",
  49017=>"110001111",
  49018=>"100100100",
  49019=>"001100100",
  49020=>"111111101",
  49021=>"110100000",
  49022=>"000000101",
  49023=>"011011110",
  49024=>"110000000",
  49025=>"111100100",
  49026=>"011011011",
  49027=>"011001101",
  49028=>"111100110",
  49029=>"111010101",
  49030=>"101100101",
  49031=>"101011000",
  49032=>"101100100",
  49033=>"101100111",
  49034=>"111101111",
  49035=>"111000011",
  49036=>"110111110",
  49037=>"001100100",
  49038=>"111100101",
  49039=>"001001010",
  49040=>"110000100",
  49041=>"110110011",
  49042=>"000011110",
  49043=>"011011000",
  49044=>"110110110",
  49045=>"001011011",
  49046=>"111001011",
  49047=>"111100100",
  49048=>"000111100",
  49049=>"110000000",
  49050=>"100101100",
  49051=>"000001001",
  49052=>"011101011",
  49053=>"000001001",
  49054=>"011011011",
  49055=>"100100001",
  49056=>"100000000",
  49057=>"011000000",
  49058=>"100111100",
  49059=>"100101011",
  49060=>"101100101",
  49061=>"100000001",
  49062=>"100100100",
  49063=>"011011011",
  49064=>"011011011",
  49065=>"001011111",
  49066=>"100100100",
  49067=>"000011001",
  49068=>"100100001",
  49069=>"010110110",
  49070=>"110111101",
  49071=>"000010111",
  49072=>"010010000",
  49073=>"000011011",
  49074=>"100100100",
  49075=>"100101101",
  49076=>"100110101",
  49077=>"111110110",
  49078=>"011010111",
  49079=>"100100000",
  49080=>"001011011",
  49081=>"001101101",
  49082=>"111011101",
  49083=>"101100110",
  49084=>"100000001",
  49085=>"100110111",
  49086=>"001011000",
  49087=>"011010110",
  49088=>"110111010",
  49089=>"011011011",
  49090=>"011011111",
  49091=>"111101111",
  49092=>"000000100",
  49093=>"111100000",
  49094=>"011000000",
  49095=>"100000111",
  49096=>"101001000",
  49097=>"011011100",
  49098=>"111011000",
  49099=>"001001011",
  49100=>"011011010",
  49101=>"000011001",
  49102=>"011010000",
  49103=>"110111100",
  49104=>"100100100",
  49105=>"100100111",
  49106=>"011111100",
  49107=>"100111101",
  49108=>"000111000",
  49109=>"101101111",
  49110=>"110011001",
  49111=>"111111001",
  49112=>"010110111",
  49113=>"000011011",
  49114=>"101100111",
  49115=>"100101111",
  49116=>"111100111",
  49117=>"001000110",
  49118=>"011011111",
  49119=>"110000110",
  49120=>"100010011",
  49121=>"110100111",
  49122=>"000000100",
  49123=>"110100111",
  49124=>"010010011",
  49125=>"110111110",
  49126=>"110100011",
  49127=>"000001010",
  49128=>"001001111",
  49129=>"011011111",
  49130=>"001001001",
  49131=>"101101000",
  49132=>"000011010",
  49133=>"000000111",
  49134=>"000000000",
  49135=>"100100001",
  49136=>"111001001",
  49137=>"000000011",
  49138=>"011010000",
  49139=>"100100111",
  49140=>"111110000",
  49141=>"001001001",
  49142=>"101001001",
  49143=>"001001001",
  49144=>"001011010",
  49145=>"110100100",
  49146=>"011100100",
  49147=>"111011011",
  49148=>"001001101",
  49149=>"110111111",
  49150=>"011100001",
  49151=>"111100101",
  49152=>"100010111",
  49153=>"000000001",
  49154=>"111001001",
  49155=>"001000110",
  49156=>"101000011",
  49157=>"100110111",
  49158=>"111101000",
  49159=>"000101000",
  49160=>"000010111",
  49161=>"111001110",
  49162=>"001000100",
  49163=>"110100000",
  49164=>"110000000",
  49165=>"010101001",
  49166=>"001000010",
  49167=>"000110111",
  49168=>"110110000",
  49169=>"111101000",
  49170=>"111111000",
  49171=>"111111100",
  49172=>"111111111",
  49173=>"101000000",
  49174=>"000110111",
  49175=>"111111000",
  49176=>"111001000",
  49177=>"001110100",
  49178=>"000110111",
  49179=>"010000011",
  49180=>"111001101",
  49181=>"101111001",
  49182=>"111111111",
  49183=>"101110110",
  49184=>"000011111",
  49185=>"100110111",
  49186=>"000101100",
  49187=>"000100110",
  49188=>"100011001",
  49189=>"011111110",
  49190=>"110000000",
  49191=>"101000111",
  49192=>"001110110",
  49193=>"000010110",
  49194=>"011101000",
  49195=>"000111110",
  49196=>"000110101",
  49197=>"101010000",
  49198=>"000110001",
  49199=>"001111001",
  49200=>"111001010",
  49201=>"000011011",
  49202=>"101111000",
  49203=>"010111001",
  49204=>"111011101",
  49205=>"111001100",
  49206=>"000000110",
  49207=>"011001001",
  49208=>"011111111",
  49209=>"111001001",
  49210=>"111101100",
  49211=>"000001101",
  49212=>"000100010",
  49213=>"111111011",
  49214=>"100000000",
  49215=>"000001111",
  49216=>"000101000",
  49217=>"000011100",
  49218=>"000001001",
  49219=>"100110111",
  49220=>"010111111",
  49221=>"100000001",
  49222=>"111001000",
  49223=>"000010110",
  49224=>"100001110",
  49225=>"000111111",
  49226=>"111001001",
  49227=>"110101000",
  49228=>"000110010",
  49229=>"000100100",
  49230=>"000000100",
  49231=>"001011101",
  49232=>"111001010",
  49233=>"010111101",
  49234=>"111101001",
  49235=>"000000001",
  49236=>"111001000",
  49237=>"101111110",
  49238=>"111000001",
  49239=>"111111000",
  49240=>"111011100",
  49241=>"100100100",
  49242=>"111000000",
  49243=>"100000011",
  49244=>"001011000",
  49245=>"001001011",
  49246=>"101110111",
  49247=>"001111111",
  49248=>"000111111",
  49249=>"000000111",
  49250=>"110101001",
  49251=>"111000000",
  49252=>"000000101",
  49253=>"011101110",
  49254=>"100000001",
  49255=>"111110010",
  49256=>"000010011",
  49257=>"111111000",
  49258=>"011111101",
  49259=>"000111111",
  49260=>"000000010",
  49261=>"111101000",
  49262=>"111000000",
  49263=>"101000101",
  49264=>"000000010",
  49265=>"001111001",
  49266=>"000010011",
  49267=>"110111000",
  49268=>"010110101",
  49269=>"111101100",
  49270=>"000000000",
  49271=>"000101111",
  49272=>"111111000",
  49273=>"111101000",
  49274=>"100000110",
  49275=>"101101111",
  49276=>"100111110",
  49277=>"000100100",
  49278=>"100110111",
  49279=>"100000110",
  49280=>"100000000",
  49281=>"010111100",
  49282=>"000110000",
  49283=>"000000000",
  49284=>"000111111",
  49285=>"111001001",
  49286=>"100110110",
  49287=>"100000100",
  49288=>"000000001",
  49289=>"111001001",
  49290=>"110000100",
  49291=>"110110110",
  49292=>"000000110",
  49293=>"101000100",
  49294=>"110000000",
  49295=>"111001001",
  49296=>"010010011",
  49297=>"000000111",
  49298=>"000011110",
  49299=>"000000000",
  49300=>"011001011",
  49301=>"101111000",
  49302=>"111111111",
  49303=>"000011011",
  49304=>"101110010",
  49305=>"000010010",
  49306=>"111001001",
  49307=>"101001001",
  49308=>"110111101",
  49309=>"111101000",
  49310=>"111000001",
  49311=>"111101000",
  49312=>"011000100",
  49313=>"010111000",
  49314=>"000010110",
  49315=>"101111010",
  49316=>"111010010",
  49317=>"010001000",
  49318=>"000110110",
  49319=>"000000111",
  49320=>"000110111",
  49321=>"000111101",
  49322=>"111101000",
  49323=>"111101001",
  49324=>"000000000",
  49325=>"000110111",
  49326=>"111100100",
  49327=>"111101001",
  49328=>"010111111",
  49329=>"010011101",
  49330=>"110110110",
  49331=>"001100110",
  49332=>"000011111",
  49333=>"110100000",
  49334=>"000000100",
  49335=>"111000111",
  49336=>"000010111",
  49337=>"000000111",
  49338=>"000010000",
  49339=>"000001000",
  49340=>"110111101",
  49341=>"111111111",
  49342=>"000110110",
  49343=>"000000000",
  49344=>"111101101",
  49345=>"010111000",
  49346=>"000111011",
  49347=>"111000011",
  49348=>"111111101",
  49349=>"000000001",
  49350=>"000000111",
  49351=>"111001000",
  49352=>"010010000",
  49353=>"011000010",
  49354=>"001111110",
  49355=>"111001000",
  49356=>"000011011",
  49357=>"100111111",
  49358=>"111101101",
  49359=>"000000011",
  49360=>"111000000",
  49361=>"000000110",
  49362=>"001100110",
  49363=>"010110111",
  49364=>"111000000",
  49365=>"110100110",
  49366=>"110110111",
  49367=>"010000001",
  49368=>"000111101",
  49369=>"000000110",
  49370=>"100110000",
  49371=>"111001000",
  49372=>"000011101",
  49373=>"001011111",
  49374=>"110000000",
  49375=>"111101001",
  49376=>"001111111",
  49377=>"111001100",
  49378=>"001010000",
  49379=>"011011011",
  49380=>"111111000",
  49381=>"000010110",
  49382=>"000001001",
  49383=>"010101100",
  49384=>"000010000",
  49385=>"000101010",
  49386=>"000001001",
  49387=>"010111100",
  49388=>"000110111",
  49389=>"000000000",
  49390=>"000001001",
  49391=>"111011110",
  49392=>"110110111",
  49393=>"000000100",
  49394=>"111010011",
  49395=>"000100100",
  49396=>"000010110",
  49397=>"111001000",
  49398=>"000000100",
  49399=>"000100000",
  49400=>"000111111",
  49401=>"000111001",
  49402=>"010110000",
  49403=>"100010111",
  49404=>"111001000",
  49405=>"000110111",
  49406=>"101110110",
  49407=>"111001000",
  49408=>"110100110",
  49409=>"000100100",
  49410=>"010010000",
  49411=>"000000000",
  49412=>"110110100",
  49413=>"000000000",
  49414=>"111001101",
  49415=>"010110100",
  49416=>"000000000",
  49417=>"000000101",
  49418=>"101111010",
  49419=>"101100111",
  49420=>"000100100",
  49421=>"011101000",
  49422=>"100000000",
  49423=>"000000000",
  49424=>"010000000",
  49425=>"111000011",
  49426=>"011010111",
  49427=>"001000000",
  49428=>"000011000",
  49429=>"111111011",
  49430=>"010001000",
  49431=>"110110111",
  49432=>"111000100",
  49433=>"111011110",
  49434=>"111111111",
  49435=>"000000000",
  49436=>"000111011",
  49437=>"000101111",
  49438=>"001001011",
  49439=>"010000000",
  49440=>"001000000",
  49441=>"110111111",
  49442=>"000000101",
  49443=>"000000000",
  49444=>"010111110",
  49445=>"001011011",
  49446=>"111001000",
  49447=>"101101111",
  49448=>"111111111",
  49449=>"000101100",
  49450=>"000000000",
  49451=>"000000100",
  49452=>"110110110",
  49453=>"110100001",
  49454=>"111100010",
  49455=>"110111111",
  49456=>"110111111",
  49457=>"010110000",
  49458=>"000100111",
  49459=>"011111011",
  49460=>"111111111",
  49461=>"000000000",
  49462=>"111011001",
  49463=>"101001000",
  49464=>"010111100",
  49465=>"001101101",
  49466=>"000000100",
  49467=>"110111010",
  49468=>"111001001",
  49469=>"111111111",
  49470=>"010100000",
  49471=>"000100001",
  49472=>"000000100",
  49473=>"001001111",
  49474=>"111111000",
  49475=>"100100000",
  49476=>"101101000",
  49477=>"000000111",
  49478=>"000000000",
  49479=>"000000100",
  49480=>"000000100",
  49481=>"000000000",
  49482=>"010111111",
  49483=>"110111011",
  49484=>"000000000",
  49485=>"000100010",
  49486=>"110010010",
  49487=>"010000010",
  49488=>"101011010",
  49489=>"010111111",
  49490=>"001101010",
  49491=>"001000000",
  49492=>"000000000",
  49493=>"010100111",
  49494=>"011111101",
  49495=>"001001111",
  49496=>"001000000",
  49497=>"111111110",
  49498=>"011010000",
  49499=>"111111110",
  49500=>"111111111",
  49501=>"011000000",
  49502=>"111011010",
  49503=>"111000000",
  49504=>"000000000",
  49505=>"001101011",
  49506=>"000000000",
  49507=>"110111000",
  49508=>"000111010",
  49509=>"000000000",
  49510=>"101110000",
  49511=>"000011000",
  49512=>"000111000",
  49513=>"000011111",
  49514=>"001000100",
  49515=>"110111011",
  49516=>"110010011",
  49517=>"010111111",
  49518=>"000111000",
  49519=>"000100100",
  49520=>"111111111",
  49521=>"000010001",
  49522=>"110110100",
  49523=>"000101010",
  49524=>"000100011",
  49525=>"000000100",
  49526=>"111111000",
  49527=>"000101101",
  49528=>"000000000",
  49529=>"100000000",
  49530=>"100110111",
  49531=>"111000111",
  49532=>"010111001",
  49533=>"100000001",
  49534=>"111110011",
  49535=>"000000000",
  49536=>"000100000",
  49537=>"001111010",
  49538=>"000000111",
  49539=>"110111111",
  49540=>"011000000",
  49541=>"000000000",
  49542=>"110110110",
  49543=>"110000000",
  49544=>"000011011",
  49545=>"111111111",
  49546=>"100001001",
  49547=>"000111111",
  49548=>"010011001",
  49549=>"100111001",
  49550=>"110010011",
  49551=>"000000000",
  49552=>"000111101",
  49553=>"111111011",
  49554=>"000000100",
  49555=>"011000001",
  49556=>"110100100",
  49557=>"000000000",
  49558=>"101100100",
  49559=>"000000010",
  49560=>"100100101",
  49561=>"010110001",
  49562=>"000000000",
  49563=>"000000000",
  49564=>"001111111",
  49565=>"110000000",
  49566=>"000000111",
  49567=>"101000000",
  49568=>"100110111",
  49569=>"010000110",
  49570=>"001000000",
  49571=>"000000000",
  49572=>"111101001",
  49573=>"100100010",
  49574=>"111011100",
  49575=>"010011011",
  49576=>"110111110",
  49577=>"100010100",
  49578=>"000000010",
  49579=>"000001100",
  49580=>"111001111",
  49581=>"100000000",
  49582=>"001111111",
  49583=>"001111001",
  49584=>"111100000",
  49585=>"000110011",
  49586=>"101100101",
  49587=>"000100000",
  49588=>"001011110",
  49589=>"001000000",
  49590=>"100000100",
  49591=>"111101100",
  49592=>"110000100",
  49593=>"010000000",
  49594=>"111001111",
  49595=>"100000010",
  49596=>"000111011",
  49597=>"100010110",
  49598=>"000000000",
  49599=>"011011111",
  49600=>"011111011",
  49601=>"111111111",
  49602=>"101111111",
  49603=>"000111110",
  49604=>"000111111",
  49605=>"111010010",
  49606=>"000000100",
  49607=>"111011011",
  49608=>"100001111",
  49609=>"100101101",
  49610=>"111100100",
  49611=>"101000001",
  49612=>"000010000",
  49613=>"001111100",
  49614=>"111111010",
  49615=>"110010011",
  49616=>"011000100",
  49617=>"100000000",
  49618=>"001110000",
  49619=>"000000000",
  49620=>"111111111",
  49621=>"001101110",
  49622=>"101000000",
  49623=>"000000111",
  49624=>"011011011",
  49625=>"000101011",
  49626=>"100110111",
  49627=>"000000101",
  49628=>"010010011",
  49629=>"000000101",
  49630=>"111110011",
  49631=>"101001000",
  49632=>"110111111",
  49633=>"000011011",
  49634=>"000000001",
  49635=>"011010000",
  49636=>"101000011",
  49637=>"000000000",
  49638=>"100000000",
  49639=>"110110110",
  49640=>"000101000",
  49641=>"000111011",
  49642=>"011011011",
  49643=>"111100110",
  49644=>"000000000",
  49645=>"000000110",
  49646=>"001001111",
  49647=>"110000000",
  49648=>"101000110",
  49649=>"100100010",
  49650=>"101100100",
  49651=>"110000000",
  49652=>"001001011",
  49653=>"010111011",
  49654=>"000000000",
  49655=>"110111011",
  49656=>"010010010",
  49657=>"011111101",
  49658=>"000011000",
  49659=>"000000000",
  49660=>"000000000",
  49661=>"101000101",
  49662=>"010010000",
  49663=>"111110000",
  49664=>"010000001",
  49665=>"011010001",
  49666=>"111100111",
  49667=>"000000000",
  49668=>"000000000",
  49669=>"100100001",
  49670=>"001110111",
  49671=>"000101000",
  49672=>"000001110",
  49673=>"111111111",
  49674=>"111110100",
  49675=>"000000001",
  49676=>"000000000",
  49677=>"010010000",
  49678=>"110110000",
  49679=>"111101000",
  49680=>"001111111",
  49681=>"000111000",
  49682=>"111111111",
  49683=>"000000100",
  49684=>"000011011",
  49685=>"000000000",
  49686=>"000010000",
  49687=>"111111000",
  49688=>"000001000",
  49689=>"011010110",
  49690=>"001001101",
  49691=>"111111101",
  49692=>"111110011",
  49693=>"000011000",
  49694=>"000111000",
  49695=>"010000000",
  49696=>"000100101",
  49697=>"000000000",
  49698=>"101000000",
  49699=>"111000110",
  49700=>"011110101",
  49701=>"010110100",
  49702=>"100000000",
  49703=>"101110111",
  49704=>"001010000",
  49705=>"000011010",
  49706=>"111111111",
  49707=>"100111101",
  49708=>"000011011",
  49709=>"010010000",
  49710=>"110111001",
  49711=>"111111111",
  49712=>"000111010",
  49713=>"111110110",
  49714=>"011001001",
  49715=>"111111101",
  49716=>"010000100",
  49717=>"000000110",
  49718=>"111010000",
  49719=>"111110111",
  49720=>"111111111",
  49721=>"111111010",
  49722=>"111111011",
  49723=>"111100101",
  49724=>"010011011",
  49725=>"111111111",
  49726=>"000000000",
  49727=>"010100000",
  49728=>"111010000",
  49729=>"101111001",
  49730=>"011000000",
  49731=>"000000000",
  49732=>"101111000",
  49733=>"101000000",
  49734=>"111100001",
  49735=>"111111111",
  49736=>"011111110",
  49737=>"101111111",
  49738=>"111001111",
  49739=>"010000000",
  49740=>"111110101",
  49741=>"111111011",
  49742=>"101000110",
  49743=>"001100011",
  49744=>"000000000",
  49745=>"111111111",
  49746=>"000000010",
  49747=>"010111000",
  49748=>"010010110",
  49749=>"111111000",
  49750=>"111111111",
  49751=>"101000101",
  49752=>"111011001",
  49753=>"111000000",
  49754=>"110110010",
  49755=>"000111110",
  49756=>"111111100",
  49757=>"111100100",
  49758=>"011111111",
  49759=>"000000000",
  49760=>"110111111",
  49761=>"111000000",
  49762=>"111101100",
  49763=>"011111010",
  49764=>"000110010",
  49765=>"010000000",
  49766=>"111011111",
  49767=>"000100101",
  49768=>"000010010",
  49769=>"110010000",
  49770=>"011110000",
  49771=>"110100001",
  49772=>"010111010",
  49773=>"111110010",
  49774=>"000010100",
  49775=>"000111001",
  49776=>"110110001",
  49777=>"000110110",
  49778=>"100111000",
  49779=>"010011011",
  49780=>"100111111",
  49781=>"000000011",
  49782=>"111000000",
  49783=>"111011111",
  49784=>"101100011",
  49785=>"111111010",
  49786=>"010111111",
  49787=>"001101001",
  49788=>"101100111",
  49789=>"111011000",
  49790=>"100101111",
  49791=>"111011010",
  49792=>"010101001",
  49793=>"000000000",
  49794=>"011111000",
  49795=>"000001011",
  49796=>"000000000",
  49797=>"010011011",
  49798=>"100111000",
  49799=>"000010110",
  49800=>"011011000",
  49801=>"101111001",
  49802=>"100110011",
  49803=>"111000001",
  49804=>"000010111",
  49805=>"000001001",
  49806=>"101101111",
  49807=>"000011011",
  49808=>"010111100",
  49809=>"110100000",
  49810=>"001110111",
  49811=>"110010000",
  49812=>"000101100",
  49813=>"100000000",
  49814=>"000000000",
  49815=>"101100100",
  49816=>"110110011",
  49817=>"010111101",
  49818=>"111110000",
  49819=>"111001000",
  49820=>"000110100",
  49821=>"111111111",
  49822=>"101010111",
  49823=>"000010000",
  49824=>"011111011",
  49825=>"000111000",
  49826=>"111111001",
  49827=>"000100010",
  49828=>"110110000",
  49829=>"000010000",
  49830=>"101011001",
  49831=>"000111000",
  49832=>"011010111",
  49833=>"010000001",
  49834=>"111011101",
  49835=>"100111100",
  49836=>"011111101",
  49837=>"111100111",
  49838=>"110111100",
  49839=>"000010000",
  49840=>"111101111",
  49841=>"000010001",
  49842=>"111111111",
  49843=>"111001011",
  49844=>"000100100",
  49845=>"111111010",
  49846=>"000000010",
  49847=>"111110101",
  49848=>"011011110",
  49849=>"000110100",
  49850=>"111111110",
  49851=>"000000111",
  49852=>"000110001",
  49853=>"111111111",
  49854=>"000010011",
  49855=>"010110111",
  49856=>"011111010",
  49857=>"000100111",
  49858=>"111011001",
  49859=>"111100000",
  49860=>"101000111",
  49861=>"111001001",
  49862=>"111101001",
  49863=>"111111111",
  49864=>"011011000",
  49865=>"000000000",
  49866=>"001000111",
  49867=>"010001110",
  49868=>"000000000",
  49869=>"001011110",
  49870=>"010100111",
  49871=>"000000101",
  49872=>"111111110",
  49873=>"000010010",
  49874=>"000000000",
  49875=>"110101011",
  49876=>"011011100",
  49877=>"101000000",
  49878=>"111111000",
  49879=>"000000111",
  49880=>"000000010",
  49881=>"110011110",
  49882=>"110110111",
  49883=>"110111110",
  49884=>"000111100",
  49885=>"110111111",
  49886=>"000111111",
  49887=>"110111110",
  49888=>"110000011",
  49889=>"110010000",
  49890=>"111010100",
  49891=>"100010000",
  49892=>"000000000",
  49893=>"000000000",
  49894=>"101100000",
  49895=>"010011000",
  49896=>"000000000",
  49897=>"000110010",
  49898=>"111011000",
  49899=>"010001000",
  49900=>"111000100",
  49901=>"010001100",
  49902=>"111111111",
  49903=>"011111111",
  49904=>"000000000",
  49905=>"101100001",
  49906=>"100111101",
  49907=>"011011110",
  49908=>"011011000",
  49909=>"111110000",
  49910=>"111111111",
  49911=>"001000101",
  49912=>"000111111",
  49913=>"011110011",
  49914=>"111111111",
  49915=>"100000000",
  49916=>"111111111",
  49917=>"011001000",
  49918=>"111111100",
  49919=>"001110110",
  49920=>"011010000",
  49921=>"000000010",
  49922=>"110111111",
  49923=>"010010000",
  49924=>"100110110",
  49925=>"000110111",
  49926=>"010111000",
  49927=>"111000000",
  49928=>"000000000",
  49929=>"000000000",
  49930=>"000000000",
  49931=>"010010000",
  49932=>"000111000",
  49933=>"000010000",
  49934=>"101101101",
  49935=>"111111111",
  49936=>"000000000",
  49937=>"011110000",
  49938=>"010100100",
  49939=>"000000000",
  49940=>"100001000",
  49941=>"011111011",
  49942=>"111111111",
  49943=>"111000000",
  49944=>"000100000",
  49945=>"001111111",
  49946=>"101000000",
  49947=>"111110111",
  49948=>"011111101",
  49949=>"010011011",
  49950=>"111110100",
  49951=>"010100000",
  49952=>"011110000",
  49953=>"000110000",
  49954=>"111100100",
  49955=>"111000000",
  49956=>"011001011",
  49957=>"111111001",
  49958=>"011011000",
  49959=>"101000110",
  49960=>"000000000",
  49961=>"000000001",
  49962=>"000010110",
  49963=>"111100111",
  49964=>"100011000",
  49965=>"100010000",
  49966=>"111101111",
  49967=>"111110111",
  49968=>"000000000",
  49969=>"100100100",
  49970=>"011000011",
  49971=>"111111101",
  49972=>"000000110",
  49973=>"000111000",
  49974=>"001011011",
  49975=>"010000101",
  49976=>"111111000",
  49977=>"111001101",
  49978=>"000001000",
  49979=>"000000000",
  49980=>"111110101",
  49981=>"101111111",
  49982=>"010000000",
  49983=>"000100000",
  49984=>"110000100",
  49985=>"110010110",
  49986=>"011100000",
  49987=>"001100110",
  49988=>"010111111",
  49989=>"000001111",
  49990=>"010010010",
  49991=>"000101111",
  49992=>"010000000",
  49993=>"101000001",
  49994=>"000000111",
  49995=>"000000000",
  49996=>"101000101",
  49997=>"110111111",
  49998=>"101111001",
  49999=>"111111111",
  50000=>"111111011",
  50001=>"000110111",
  50002=>"010111010",
  50003=>"001111001",
  50004=>"000100100",
  50005=>"001010010",
  50006=>"110100111",
  50007=>"100000000",
  50008=>"000000000",
  50009=>"110110100",
  50010=>"001011001",
  50011=>"100100000",
  50012=>"010011000",
  50013=>"011001001",
  50014=>"111111111",
  50015=>"100001011",
  50016=>"000000110",
  50017=>"111000111",
  50018=>"000000000",
  50019=>"011011110",
  50020=>"010111101",
  50021=>"100100000",
  50022=>"000110000",
  50023=>"110110000",
  50024=>"010111000",
  50025=>"111101100",
  50026=>"111100000",
  50027=>"000000000",
  50028=>"111100101",
  50029=>"000000000",
  50030=>"010111011",
  50031=>"111111111",
  50032=>"000110110",
  50033=>"111011000",
  50034=>"100110000",
  50035=>"111000111",
  50036=>"000000111",
  50037=>"111010101",
  50038=>"111111000",
  50039=>"000100110",
  50040=>"110110100",
  50041=>"111011000",
  50042=>"000100001",
  50043=>"111111111",
  50044=>"110110111",
  50045=>"100100000",
  50046=>"000000001",
  50047=>"001011011",
  50048=>"100111111",
  50049=>"111110100",
  50050=>"000000001",
  50051=>"100111111",
  50052=>"111111100",
  50053=>"000000000",
  50054=>"110100100",
  50055=>"110010111",
  50056=>"001011111",
  50057=>"000101111",
  50058=>"000000000",
  50059=>"111111111",
  50060=>"000011111",
  50061=>"000111010",
  50062=>"111111111",
  50063=>"111000001",
  50064=>"010100100",
  50065=>"110110110",
  50066=>"100000000",
  50067=>"111100011",
  50068=>"111001100",
  50069=>"010111111",
  50070=>"000111110",
  50071=>"000000001",
  50072=>"011011011",
  50073=>"111011101",
  50074=>"110111011",
  50075=>"000000000",
  50076=>"000011001",
  50077=>"010111111",
  50078=>"000000000",
  50079=>"101000111",
  50080=>"110110100",
  50081=>"111110011",
  50082=>"111111010",
  50083=>"100101111",
  50084=>"000000000",
  50085=>"101011000",
  50086=>"101001001",
  50087=>"000011011",
  50088=>"110100111",
  50089=>"111111000",
  50090=>"000000000",
  50091=>"011101111",
  50092=>"110100000",
  50093=>"111111111",
  50094=>"111111011",
  50095=>"000001101",
  50096=>"111100111",
  50097=>"001000100",
  50098=>"111001111",
  50099=>"110110010",
  50100=>"000101000",
  50101=>"011100000",
  50102=>"111110110",
  50103=>"010111110",
  50104=>"000011100",
  50105=>"101101001",
  50106=>"000000010",
  50107=>"010110111",
  50108=>"111111111",
  50109=>"111111111",
  50110=>"000000000",
  50111=>"111111111",
  50112=>"010010000",
  50113=>"000000110",
  50114=>"111000001",
  50115=>"001001001",
  50116=>"000000001",
  50117=>"000111011",
  50118=>"110100001",
  50119=>"000000100",
  50120=>"111001111",
  50121=>"001000000",
  50122=>"011111010",
  50123=>"010111110",
  50124=>"100110111",
  50125=>"001011011",
  50126=>"110000000",
  50127=>"100000000",
  50128=>"111100100",
  50129=>"000100100",
  50130=>"101101111",
  50131=>"000101111",
  50132=>"101000101",
  50133=>"110110000",
  50134=>"110110000",
  50135=>"100000000",
  50136=>"100000000",
  50137=>"011111011",
  50138=>"101000001",
  50139=>"101100100",
  50140=>"101110101",
  50141=>"000001000",
  50142=>"000011111",
  50143=>"110011000",
  50144=>"000000001",
  50145=>"011111101",
  50146=>"000000000",
  50147=>"001101101",
  50148=>"101000000",
  50149=>"010110110",
  50150=>"000110010",
  50151=>"100110010",
  50152=>"000100000",
  50153=>"011100110",
  50154=>"111111000",
  50155=>"111000000",
  50156=>"000010000",
  50157=>"101000001",
  50158=>"111111111",
  50159=>"101000000",
  50160=>"000000000",
  50161=>"110011111",
  50162=>"111000000",
  50163=>"110111010",
  50164=>"111000001",
  50165=>"001111101",
  50166=>"000000010",
  50167=>"111101100",
  50168=>"111111110",
  50169=>"001111000",
  50170=>"000111111",
  50171=>"111100001",
  50172=>"111111111",
  50173=>"010111010",
  50174=>"010100000",
  50175=>"110100110",
  50176=>"000000111",
  50177=>"000000100",
  50178=>"101000100",
  50179=>"000000000",
  50180=>"100100100",
  50181=>"111000000",
  50182=>"101001111",
  50183=>"100100000",
  50184=>"000000111",
  50185=>"110000101",
  50186=>"000001001",
  50187=>"010011000",
  50188=>"001010010",
  50189=>"111101000",
  50190=>"100100010",
  50191=>"101011111",
  50192=>"101000100",
  50193=>"111000101",
  50194=>"010101100",
  50195=>"000100000",
  50196=>"001110111",
  50197=>"111011101",
  50198=>"000000110",
  50199=>"101101001",
  50200=>"111100000",
  50201=>"000000000",
  50202=>"001101111",
  50203=>"111111111",
  50204=>"111011100",
  50205=>"000100101",
  50206=>"100101101",
  50207=>"000111111",
  50208=>"100101111",
  50209=>"011111000",
  50210=>"100010111",
  50211=>"000011110",
  50212=>"010111011",
  50213=>"001100001",
  50214=>"101000111",
  50215=>"000000011",
  50216=>"000011111",
  50217=>"001110111",
  50218=>"100101101",
  50219=>"110011110",
  50220=>"011000110",
  50221=>"111010010",
  50222=>"011101101",
  50223=>"010111101",
  50224=>"011110111",
  50225=>"000011010",
  50226=>"010000010",
  50227=>"110111111",
  50228=>"111000000",
  50229=>"101010111",
  50230=>"110100000",
  50231=>"011000100",
  50232=>"111111100",
  50233=>"101000000",
  50234=>"011010011",
  50235=>"100011011",
  50236=>"100000100",
  50237=>"111111111",
  50238=>"000100000",
  50239=>"000011001",
  50240=>"000000111",
  50241=>"001001011",
  50242=>"101111111",
  50243=>"000100101",
  50244=>"000011011",
  50245=>"101000000",
  50246=>"101101101",
  50247=>"111111000",
  50248=>"111100000",
  50249=>"110101101",
  50250=>"000000000",
  50251=>"111111101",
  50252=>"011100101",
  50253=>"000101110",
  50254=>"000100011",
  50255=>"111111100",
  50256=>"111000000",
  50257=>"011010000",
  50258=>"011010000",
  50259=>"010011001",
  50260=>"111000001",
  50261=>"001111100",
  50262=>"101000010",
  50263=>"111000100",
  50264=>"011111011",
  50265=>"011001000",
  50266=>"100100110",
  50267=>"000011011",
  50268=>"000101010",
  50269=>"100001001",
  50270=>"111011111",
  50271=>"100000111",
  50272=>"000010101",
  50273=>"010101000",
  50274=>"111000100",
  50275=>"001001001",
  50276=>"000011010",
  50277=>"011000000",
  50278=>"010101011",
  50279=>"100010011",
  50280=>"000010010",
  50281=>"111000000",
  50282=>"010111101",
  50283=>"111000010",
  50284=>"000100111",
  50285=>"111101111",
  50286=>"010000101",
  50287=>"111010000",
  50288=>"001000110",
  50289=>"111000000",
  50290=>"011001000",
  50291=>"100001011",
  50292=>"111001000",
  50293=>"011000100",
  50294=>"111000000",
  50295=>"000000111",
  50296=>"011000101",
  50297=>"111010100",
  50298=>"000111111",
  50299=>"000110001",
  50300=>"000110000",
  50301=>"000000100",
  50302=>"000010000",
  50303=>"101101000",
  50304=>"001101101",
  50305=>"111101101",
  50306=>"001000110",
  50307=>"000000000",
  50308=>"010011001",
  50309=>"000001111",
  50310=>"100111100",
  50311=>"100000001",
  50312=>"110111011",
  50313=>"000000010",
  50314=>"000100100",
  50315=>"100010000",
  50316=>"000110111",
  50317=>"000100010",
  50318=>"000101010",
  50319=>"001000000",
  50320=>"010100010",
  50321=>"000110011",
  50322=>"011001000",
  50323=>"111101000",
  50324=>"000100111",
  50325=>"111000000",
  50326=>"111110111",
  50327=>"000001011",
  50328=>"111110010",
  50329=>"000000000",
  50330=>"000000000",
  50331=>"001011100",
  50332=>"100100111",
  50333=>"010101111",
  50334=>"101111000",
  50335=>"110110100",
  50336=>"001101010",
  50337=>"011000101",
  50338=>"000000101",
  50339=>"001000111",
  50340=>"010000101",
  50341=>"100000011",
  50342=>"000110110",
  50343=>"110101111",
  50344=>"111100000",
  50345=>"100000110",
  50346=>"101111101",
  50347=>"111100000",
  50348=>"000001010",
  50349=>"001101000",
  50350=>"110001001",
  50351=>"000010010",
  50352=>"000011100",
  50353=>"010011101",
  50354=>"000000010",
  50355=>"010010110",
  50356=>"101011011",
  50357=>"011111010",
  50358=>"001000001",
  50359=>"000000000",
  50360=>"001000001",
  50361=>"000001001",
  50362=>"000000001",
  50363=>"010111011",
  50364=>"010010011",
  50365=>"101000110",
  50366=>"001100010",
  50367=>"011010111",
  50368=>"111000001",
  50369=>"100000100",
  50370=>"111000100",
  50371=>"101101111",
  50372=>"100000100",
  50373=>"110110011",
  50374=>"110110110",
  50375=>"010000111",
  50376=>"110000000",
  50377=>"101010111",
  50378=>"100100111",
  50379=>"111011111",
  50380=>"000100100",
  50381=>"000001000",
  50382=>"000000000",
  50383=>"100010011",
  50384=>"111010000",
  50385=>"100100111",
  50386=>"000000010",
  50387=>"000101111",
  50388=>"101111111",
  50389=>"110110000",
  50390=>"111111100",
  50391=>"101100100",
  50392=>"010010000",
  50393=>"010010111",
  50394=>"000100001",
  50395=>"111100101",
  50396=>"000010001",
  50397=>"101001101",
  50398=>"000011111",
  50399=>"111101101",
  50400=>"011110110",
  50401=>"111101000",
  50402=>"101011011",
  50403=>"000001011",
  50404=>"100000101",
  50405=>"000111010",
  50406=>"000010011",
  50407=>"011100100",
  50408=>"110101101",
  50409=>"000000111",
  50410=>"000100100",
  50411=>"011100000",
  50412=>"000010010",
  50413=>"010010001",
  50414=>"100000000",
  50415=>"100100101",
  50416=>"010111010",
  50417=>"011011100",
  50418=>"000000101",
  50419=>"000110110",
  50420=>"001101100",
  50421=>"001001000",
  50422=>"100101101",
  50423=>"100001111",
  50424=>"111000000",
  50425=>"111110101",
  50426=>"011111101",
  50427=>"101111111",
  50428=>"111101111",
  50429=>"000011011",
  50430=>"000100011",
  50431=>"111100100",
  50432=>"001100010",
  50433=>"001011000",
  50434=>"100000110",
  50435=>"001010111",
  50436=>"000000010",
  50437=>"100000000",
  50438=>"001001010",
  50439=>"111000001",
  50440=>"010100110",
  50441=>"110010100",
  50442=>"001011001",
  50443=>"100110100",
  50444=>"110100100",
  50445=>"000000000",
  50446=>"100001101",
  50447=>"001010000",
  50448=>"010000000",
  50449=>"111111000",
  50450=>"000100001",
  50451=>"100100110",
  50452=>"011001001",
  50453=>"011110110",
  50454=>"011101000",
  50455=>"100111000",
  50456=>"001000000",
  50457=>"000000011",
  50458=>"100001001",
  50459=>"110111111",
  50460=>"111011011",
  50461=>"011000000",
  50462=>"110110111",
  50463=>"100111011",
  50464=>"100100110",
  50465=>"111101001",
  50466=>"001001000",
  50467=>"011111101",
  50468=>"010001000",
  50469=>"001000100",
  50470=>"000100000",
  50471=>"111010011",
  50472=>"111110100",
  50473=>"011011001",
  50474=>"000000010",
  50475=>"000111011",
  50476=>"000001011",
  50477=>"011111100",
  50478=>"111001101",
  50479=>"100101000",
  50480=>"111110100",
  50481=>"011001011",
  50482=>"111000111",
  50483=>"100001010",
  50484=>"010001000",
  50485=>"010010000",
  50486=>"010011010",
  50487=>"110001100",
  50488=>"100100111",
  50489=>"110100000",
  50490=>"000110111",
  50491=>"111110111",
  50492=>"010110100",
  50493=>"111011001",
  50494=>"001000000",
  50495=>"000111110",
  50496=>"110110111",
  50497=>"001001011",
  50498=>"100100100",
  50499=>"100110010",
  50500=>"000011000",
  50501=>"100110101",
  50502=>"011111110",
  50503=>"011100100",
  50504=>"011101010",
  50505=>"011010110",
  50506=>"111110110",
  50507=>"011100110",
  50508=>"111101110",
  50509=>"111011000",
  50510=>"000110111",
  50511=>"000101000",
  50512=>"100011011",
  50513=>"011101011",
  50514=>"001100000",
  50515=>"111010000",
  50516=>"010011001",
  50517=>"011000011",
  50518=>"001001001",
  50519=>"110110101",
  50520=>"000111011",
  50521=>"011011111",
  50522=>"010001001",
  50523=>"001011111",
  50524=>"010000100",
  50525=>"000001000",
  50526=>"111110111",
  50527=>"111111010",
  50528=>"111011010",
  50529=>"001001100",
  50530=>"000100111",
  50531=>"001011011",
  50532=>"100100111",
  50533=>"111111111",
  50534=>"110100111",
  50535=>"100000000",
  50536=>"000110111",
  50537=>"110000101",
  50538=>"011110100",
  50539=>"010010000",
  50540=>"111101001",
  50541=>"001001000",
  50542=>"000001000",
  50543=>"011111000",
  50544=>"010001001",
  50545=>"111110001",
  50546=>"110000001",
  50547=>"011010000",
  50548=>"000001000",
  50549=>"110100110",
  50550=>"000011010",
  50551=>"000000111",
  50552=>"100100100",
  50553=>"011011001",
  50554=>"100101011",
  50555=>"010100110",
  50556=>"001001000",
  50557=>"110100110",
  50558=>"100110110",
  50559=>"110110110",
  50560=>"111110000",
  50561=>"100100011",
  50562=>"011011111",
  50563=>"001001011",
  50564=>"011100001",
  50565=>"001000000",
  50566=>"011111000",
  50567=>"100000011",
  50568=>"000001111",
  50569=>"100110001",
  50570=>"000010000",
  50571=>"100111001",
  50572=>"010110010",
  50573=>"110110010",
  50574=>"000010111",
  50575=>"000000000",
  50576=>"001001000",
  50577=>"000110100",
  50578=>"000110110",
  50579=>"000110000",
  50580=>"001101101",
  50581=>"010100100",
  50582=>"011011111",
  50583=>"100110010",
  50584=>"110111111",
  50585=>"010100000",
  50586=>"000100110",
  50587=>"000110100",
  50588=>"111100000",
  50589=>"000111010",
  50590=>"001101111",
  50591=>"111100110",
  50592=>"011100011",
  50593=>"010000011",
  50594=>"100100111",
  50595=>"000100101",
  50596=>"001010011",
  50597=>"110011110",
  50598=>"000100001",
  50599=>"010000000",
  50600=>"001011000",
  50601=>"000110110",
  50602=>"000100110",
  50603=>"110111011",
  50604=>"111000011",
  50605=>"110000101",
  50606=>"000011011",
  50607=>"000100110",
  50608=>"100110100",
  50609=>"110110001",
  50610=>"001111011",
  50611=>"110100000",
  50612=>"101001000",
  50613=>"000001000",
  50614=>"001001001",
  50615=>"110001000",
  50616=>"011000000",
  50617=>"001100010",
  50618=>"011100100",
  50619=>"100100100",
  50620=>"000000111",
  50621=>"011111001",
  50622=>"100100111",
  50623=>"111110000",
  50624=>"100000100",
  50625=>"001011000",
  50626=>"001110000",
  50627=>"111001001",
  50628=>"000000101",
  50629=>"001001110",
  50630=>"111100000",
  50631=>"000100110",
  50632=>"110100110",
  50633=>"100001001",
  50634=>"100111011",
  50635=>"000110010",
  50636=>"110110111",
  50637=>"111101100",
  50638=>"000011001",
  50639=>"000100110",
  50640=>"100011001",
  50641=>"010011001",
  50642=>"000100000",
  50643=>"111011000",
  50644=>"010001001",
  50645=>"000011101",
  50646=>"001001001",
  50647=>"100011000",
  50648=>"111000011",
  50649=>"000000000",
  50650=>"000110101",
  50651=>"110100100",
  50652=>"011010111",
  50653=>"100100100",
  50654=>"011001000",
  50655=>"000100010",
  50656=>"100100100",
  50657=>"111011001",
  50658=>"010110110",
  50659=>"010010110",
  50660=>"110000000",
  50661=>"011010011",
  50662=>"000000000",
  50663=>"000011011",
  50664=>"110010000",
  50665=>"000001001",
  50666=>"111011011",
  50667=>"010110110",
  50668=>"100100100",
  50669=>"111001001",
  50670=>"110100100",
  50671=>"011100100",
  50672=>"100100110",
  50673=>"011011000",
  50674=>"111110110",
  50675=>"011011001",
  50676=>"101111100",
  50677=>"100011001",
  50678=>"000000100",
  50679=>"000000000",
  50680=>"000100010",
  50681=>"111100110",
  50682=>"111111110",
  50683=>"111111001",
  50684=>"010110000",
  50685=>"011000010",
  50686=>"001011111",
  50687=>"011011110",
  50688=>"101111110",
  50689=>"000000000",
  50690=>"101001000",
  50691=>"000000001",
  50692=>"000100110",
  50693=>"111101111",
  50694=>"101110110",
  50695=>"100100000",
  50696=>"101001000",
  50697=>"001000000",
  50698=>"011111011",
  50699=>"001011111",
  50700=>"001100111",
  50701=>"111100101",
  50702=>"110000110",
  50703=>"111111010",
  50704=>"000000010",
  50705=>"000000000",
  50706=>"001101101",
  50707=>"010110111",
  50708=>"010110101",
  50709=>"111000111",
  50710=>"001101000",
  50711=>"111111000",
  50712=>"010000010",
  50713=>"000000000",
  50714=>"100101111",
  50715=>"000000101",
  50716=>"100010000",
  50717=>"011110101",
  50718=>"111101000",
  50719=>"000000111",
  50720=>"110001000",
  50721=>"000010000",
  50722=>"000101111",
  50723=>"000000111",
  50724=>"011100111",
  50725=>"111001111",
  50726=>"000000011",
  50727=>"000110000",
  50728=>"011010011",
  50729=>"100111111",
  50730=>"110010010",
  50731=>"000010000",
  50732=>"011100001",
  50733=>"111100111",
  50734=>"111111111",
  50735=>"110000111",
  50736=>"111101001",
  50737=>"100111010",
  50738=>"000001000",
  50739=>"111111111",
  50740=>"000011111",
  50741=>"001000011",
  50742=>"000000011",
  50743=>"000110100",
  50744=>"111101001",
  50745=>"001001111",
  50746=>"001111101",
  50747=>"010000110",
  50748=>"000011111",
  50749=>"011110110",
  50750=>"101000000",
  50751=>"101001100",
  50752=>"100000000",
  50753=>"000010101",
  50754=>"101101000",
  50755=>"001101101",
  50756=>"100111111",
  50757=>"101101001",
  50758=>"111010010",
  50759=>"111101111",
  50760=>"110001100",
  50761=>"000100000",
  50762=>"000101101",
  50763=>"111010110",
  50764=>"101101111",
  50765=>"111111111",
  50766=>"000011010",
  50767=>"100100001",
  50768=>"000000010",
  50769=>"111010000",
  50770=>"010010111",
  50771=>"011001000",
  50772=>"000000110",
  50773=>"001001000",
  50774=>"010010111",
  50775=>"000000000",
  50776=>"101111011",
  50777=>"000101111",
  50778=>"100001011",
  50779=>"000001111",
  50780=>"110111010",
  50781=>"100000001",
  50782=>"110010111",
  50783=>"100100111",
  50784=>"100101111",
  50785=>"001000100",
  50786=>"111000111",
  50787=>"011100100",
  50788=>"011111110",
  50789=>"111010010",
  50790=>"001001111",
  50791=>"101111111",
  50792=>"000101111",
  50793=>"111110001",
  50794=>"101110010",
  50795=>"001111010",
  50796=>"010000101",
  50797=>"111111100",
  50798=>"001100100",
  50799=>"111111100",
  50800=>"100100100",
  50801=>"000110010",
  50802=>"100000000",
  50803=>"111100000",
  50804=>"110111110",
  50805=>"101000101",
  50806=>"111011000",
  50807=>"000001111",
  50808=>"000000101",
  50809=>"000111111",
  50810=>"111111111",
  50811=>"111101000",
  50812=>"000001000",
  50813=>"111101000",
  50814=>"101111111",
  50815=>"001001101",
  50816=>"010010001",
  50817=>"100100101",
  50818=>"000110111",
  50819=>"000010010",
  50820=>"111000110",
  50821=>"010110111",
  50822=>"110110101",
  50823=>"000100000",
  50824=>"001001001",
  50825=>"000010110",
  50826=>"111010000",
  50827=>"000011000",
  50828=>"000001000",
  50829=>"101101111",
  50830=>"000010000",
  50831=>"000000011",
  50832=>"001111111",
  50833=>"111101110",
  50834=>"111010000",
  50835=>"100000001",
  50836=>"000000010",
  50837=>"000111111",
  50838=>"110110010",
  50839=>"100100110",
  50840=>"001001001",
  50841=>"000000000",
  50842=>"110111011",
  50843=>"100000000",
  50844=>"101111000",
  50845=>"000000000",
  50846=>"010111000",
  50847=>"001101000",
  50848=>"001000000",
  50849=>"010001000",
  50850=>"000000000",
  50851=>"000000000",
  50852=>"111111011",
  50853=>"111111111",
  50854=>"001111001",
  50855=>"000100001",
  50856=>"011011011",
  50857=>"111001000",
  50858=>"111000000",
  50859=>"000000100",
  50860=>"000001000",
  50861=>"001001111",
  50862=>"011011010",
  50863=>"001000110",
  50864=>"000100101",
  50865=>"000001011",
  50866=>"000001100",
  50867=>"000101011",
  50868=>"111111011",
  50869=>"011011011",
  50870=>"011100111",
  50871=>"111011000",
  50872=>"000110111",
  50873=>"000001000",
  50874=>"110111111",
  50875=>"110100111",
  50876=>"010000111",
  50877=>"100001000",
  50878=>"100000000",
  50879=>"000000000",
  50880=>"111000100",
  50881=>"000011010",
  50882=>"110111111",
  50883=>"001100110",
  50884=>"111111111",
  50885=>"111110001",
  50886=>"111111000",
  50887=>"111111000",
  50888=>"000110011",
  50889=>"000000101",
  50890=>"000111011",
  50891=>"000010000",
  50892=>"000110111",
  50893=>"000100000",
  50894=>"000000010",
  50895=>"100100000",
  50896=>"000011111",
  50897=>"011001001",
  50898=>"100000010",
  50899=>"111111111",
  50900=>"000000111",
  50901=>"000000100",
  50902=>"101100101",
  50903=>"010110000",
  50904=>"011011001",
  50905=>"000111111",
  50906=>"000001000",
  50907=>"111011000",
  50908=>"001000000",
  50909=>"000101110",
  50910=>"100101011",
  50911=>"110110000",
  50912=>"000000101",
  50913=>"111000000",
  50914=>"111110111",
  50915=>"100100100",
  50916=>"000000000",
  50917=>"010111110",
  50918=>"101011010",
  50919=>"010010110",
  50920=>"000111111",
  50921=>"010111110",
  50922=>"110011000",
  50923=>"100000010",
  50924=>"000101111",
  50925=>"111011011",
  50926=>"101001000",
  50927=>"100001111",
  50928=>"000000011",
  50929=>"111011101",
  50930=>"001100101",
  50931=>"101101101",
  50932=>"011011111",
  50933=>"000101111",
  50934=>"101011111",
  50935=>"001001101",
  50936=>"010000000",
  50937=>"110111101",
  50938=>"101101111",
  50939=>"010111111",
  50940=>"111111011",
  50941=>"001111110",
  50942=>"100011110",
  50943=>"000000000",
  50944=>"100000110",
  50945=>"000000000",
  50946=>"100111111",
  50947=>"100000000",
  50948=>"001100100",
  50949=>"011000011",
  50950=>"111111111",
  50951=>"001101101",
  50952=>"000100100",
  50953=>"000111000",
  50954=>"001001011",
  50955=>"001101111",
  50956=>"010000000",
  50957=>"110000000",
  50958=>"110100100",
  50959=>"111111111",
  50960=>"011000111",
  50961=>"101111111",
  50962=>"011011011",
  50963=>"000000000",
  50964=>"000000000",
  50965=>"001010111",
  50966=>"110011111",
  50967=>"111111000",
  50968=>"001000000",
  50969=>"010000010",
  50970=>"100100101",
  50971=>"111111111",
  50972=>"000001100",
  50973=>"101111011",
  50974=>"000010011",
  50975=>"101101000",
  50976=>"000011010",
  50977=>"111000111",
  50978=>"110111101",
  50979=>"001111111",
  50980=>"011011010",
  50981=>"001000010",
  50982=>"000010010",
  50983=>"111111011",
  50984=>"011000000",
  50985=>"100100100",
  50986=>"010000110",
  50987=>"000011010",
  50988=>"111011011",
  50989=>"000000001",
  50990=>"000111111",
  50991=>"110111111",
  50992=>"111111000",
  50993=>"110110111",
  50994=>"010001101",
  50995=>"010011011",
  50996=>"111111111",
  50997=>"111100110",
  50998=>"011111111",
  50999=>"111101101",
  51000=>"000000000",
  51001=>"001111100",
  51002=>"111111111",
  51003=>"111111111",
  51004=>"001011101",
  51005=>"111111000",
  51006=>"000000000",
  51007=>"010100101",
  51008=>"111100111",
  51009=>"010010010",
  51010=>"001010000",
  51011=>"000000100",
  51012=>"111000011",
  51013=>"000000100",
  51014=>"110000000",
  51015=>"100111111",
  51016=>"000000000",
  51017=>"101000111",
  51018=>"100101001",
  51019=>"110000000",
  51020=>"000111111",
  51021=>"100100100",
  51022=>"001001011",
  51023=>"000000101",
  51024=>"000111011",
  51025=>"111111111",
  51026=>"101000100",
  51027=>"001100111",
  51028=>"000100000",
  51029=>"111101111",
  51030=>"111011001",
  51031=>"000100110",
  51032=>"001111111",
  51033=>"110110110",
  51034=>"111101100",
  51035=>"011011111",
  51036=>"001111100",
  51037=>"000110110",
  51038=>"011000111",
  51039=>"000100011",
  51040=>"000000000",
  51041=>"000000000",
  51042=>"010000010",
  51043=>"111011000",
  51044=>"101011111",
  51045=>"111000100",
  51046=>"000000000",
  51047=>"101100000",
  51048=>"111000000",
  51049=>"010010111",
  51050=>"000000010",
  51051=>"000100001",
  51052=>"001000000",
  51053=>"011111111",
  51054=>"101000100",
  51055=>"111000101",
  51056=>"100100100",
  51057=>"010010000",
  51058=>"110011011",
  51059=>"111111001",
  51060=>"000100000",
  51061=>"001111001",
  51062=>"001000100",
  51063=>"111111111",
  51064=>"001000111",
  51065=>"000111010",
  51066=>"110100001",
  51067=>"111111111",
  51068=>"100011111",
  51069=>"010001111",
  51070=>"110001111",
  51071=>"000000000",
  51072=>"010000001",
  51073=>"100100000",
  51074=>"010110111",
  51075=>"111111101",
  51076=>"101000000",
  51077=>"111000100",
  51078=>"110010000",
  51079=>"101110110",
  51080=>"001000001",
  51081=>"001100010",
  51082=>"111000010",
  51083=>"100010010",
  51084=>"000000000",
  51085=>"010001011",
  51086=>"000111111",
  51087=>"001001101",
  51088=>"111011000",
  51089=>"111000000",
  51090=>"011000100",
  51091=>"111000000",
  51092=>"000000000",
  51093=>"111001101",
  51094=>"011111111",
  51095=>"001001000",
  51096=>"110101100",
  51097=>"100001111",
  51098=>"111111101",
  51099=>"101000000",
  51100=>"000110100",
  51101=>"010000111",
  51102=>"001000111",
  51103=>"000011000",
  51104=>"100111111",
  51105=>"011111011",
  51106=>"111000000",
  51107=>"110111101",
  51108=>"111000000",
  51109=>"110110110",
  51110=>"000001001",
  51111=>"011001100",
  51112=>"000000010",
  51113=>"111111001",
  51114=>"010001100",
  51115=>"001101111",
  51116=>"111000001",
  51117=>"000000000",
  51118=>"001101111",
  51119=>"001000000",
  51120=>"001101101",
  51121=>"000001100",
  51122=>"010011011",
  51123=>"000011011",
  51124=>"111000001",
  51125=>"000100001",
  51126=>"011011010",
  51127=>"111000000",
  51128=>"110110110",
  51129=>"001000100",
  51130=>"000000000",
  51131=>"000101100",
  51132=>"000110111",
  51133=>"001011011",
  51134=>"110010101",
  51135=>"000111000",
  51136=>"000000111",
  51137=>"000011000",
  51138=>"000000000",
  51139=>"100110110",
  51140=>"111111110",
  51141=>"000000001",
  51142=>"111111000",
  51143=>"000100111",
  51144=>"101111111",
  51145=>"000101100",
  51146=>"000000000",
  51147=>"010010111",
  51148=>"000000111",
  51149=>"011110110",
  51150=>"111111000",
  51151=>"010011111",
  51152=>"011000000",
  51153=>"011000000",
  51154=>"111000100",
  51155=>"111101110",
  51156=>"000111111",
  51157=>"010000000",
  51158=>"001111111",
  51159=>"000000000",
  51160=>"011000000",
  51161=>"111000000",
  51162=>"000010111",
  51163=>"011100000",
  51164=>"111111001",
  51165=>"111011000",
  51166=>"111100000",
  51167=>"101000000",
  51168=>"000000000",
  51169=>"111000011",
  51170=>"111001011",
  51171=>"000111111",
  51172=>"000101100",
  51173=>"100100111",
  51174=>"000000000",
  51175=>"100111111",
  51176=>"011000111",
  51177=>"000001101",
  51178=>"100111011",
  51179=>"000000000",
  51180=>"000100100",
  51181=>"011001101",
  51182=>"001000000",
  51183=>"010000111",
  51184=>"000111100",
  51185=>"000100000",
  51186=>"111000000",
  51187=>"111010000",
  51188=>"011000001",
  51189=>"111111110",
  51190=>"000010101",
  51191=>"111110011",
  51192=>"000000000",
  51193=>"111101101",
  51194=>"000101100",
  51195=>"111010010",
  51196=>"000011111",
  51197=>"100100010",
  51198=>"101001111",
  51199=>"000000001",
  51200=>"011001011",
  51201=>"000101101",
  51202=>"001001000",
  51203=>"000001000",
  51204=>"001000101",
  51205=>"111110000",
  51206=>"010111111",
  51207=>"001110110",
  51208=>"110111110",
  51209=>"111111111",
  51210=>"001000000",
  51211=>"010000000",
  51212=>"000010111",
  51213=>"110111101",
  51214=>"010101001",
  51215=>"000001100",
  51216=>"000000001",
  51217=>"111111110",
  51218=>"100111001",
  51219=>"010100000",
  51220=>"110010101",
  51221=>"111101111",
  51222=>"000001001",
  51223=>"000001001",
  51224=>"100111111",
  51225=>"001000101",
  51226=>"010000000",
  51227=>"000111111",
  51228=>"111000000",
  51229=>"000101010",
  51230=>"010100010",
  51231=>"000111111",
  51232=>"111000000",
  51233=>"110000111",
  51234=>"001001110",
  51235=>"000110000",
  51236=>"000010011",
  51237=>"111000100",
  51238=>"000000000",
  51239=>"011100110",
  51240=>"011001000",
  51241=>"110110000",
  51242=>"110000000",
  51243=>"000000000",
  51244=>"111001001",
  51245=>"001001100",
  51246=>"111000111",
  51247=>"100111100",
  51248=>"000000001",
  51249=>"011111100",
  51250=>"000000111",
  51251=>"000000000",
  51252=>"000010110",
  51253=>"100011010",
  51254=>"000000000",
  51255=>"000101101",
  51256=>"000010011",
  51257=>"001101111",
  51258=>"001101101",
  51259=>"010110100",
  51260=>"110111011",
  51261=>"111111111",
  51262=>"000000100",
  51263=>"011111010",
  51264=>"000010111",
  51265=>"000101111",
  51266=>"101101101",
  51267=>"011001001",
  51268=>"111101000",
  51269=>"110110110",
  51270=>"000000011",
  51271=>"111010000",
  51272=>"000111101",
  51273=>"111000101",
  51274=>"001000111",
  51275=>"111110010",
  51276=>"111111100",
  51277=>"110110111",
  51278=>"110110011",
  51279=>"011111111",
  51280=>"000000010",
  51281=>"000111111",
  51282=>"010111001",
  51283=>"011011111",
  51284=>"101101001",
  51285=>"110111110",
  51286=>"011111001",
  51287=>"001000000",
  51288=>"111111001",
  51289=>"100000100",
  51290=>"100111100",
  51291=>"111010011",
  51292=>"000101101",
  51293=>"010010000",
  51294=>"101111011",
  51295=>"100001111",
  51296=>"110111101",
  51297=>"000001001",
  51298=>"001000000",
  51299=>"011011001",
  51300=>"001010111",
  51301=>"100000111",
  51302=>"000000000",
  51303=>"110111100",
  51304=>"111001000",
  51305=>"111000000",
  51306=>"101001101",
  51307=>"100000110",
  51308=>"110111111",
  51309=>"000000000",
  51310=>"110010000",
  51311=>"111010000",
  51312=>"110000101",
  51313=>"000000000",
  51314=>"001001000",
  51315=>"101010000",
  51316=>"110011000",
  51317=>"111000001",
  51318=>"011111111",
  51319=>"111110110",
  51320=>"000001000",
  51321=>"101000111",
  51322=>"000100000",
  51323=>"001101001",
  51324=>"110000001",
  51325=>"100100100",
  51326=>"001000111",
  51327=>"110000000",
  51328=>"101111110",
  51329=>"000000000",
  51330=>"111111111",
  51331=>"000101111",
  51332=>"110111111",
  51333=>"000100111",
  51334=>"111001011",
  51335=>"000000100",
  51336=>"100000000",
  51337=>"001101111",
  51338=>"101001110",
  51339=>"010000000",
  51340=>"110000000",
  51341=>"010001000",
  51342=>"000010010",
  51343=>"001000001",
  51344=>"101000100",
  51345=>"000000111",
  51346=>"010100010",
  51347=>"000000110",
  51348=>"000010010",
  51349=>"111000000",
  51350=>"010000101",
  51351=>"010011011",
  51352=>"111010000",
  51353=>"101001110",
  51354=>"001101001",
  51355=>"000000011",
  51356=>"000100000",
  51357=>"000000110",
  51358=>"100101101",
  51359=>"010000000",
  51360=>"001100101",
  51361=>"001000000",
  51362=>"011101111",
  51363=>"000000000",
  51364=>"111000000",
  51365=>"001111111",
  51366=>"110110000",
  51367=>"110000001",
  51368=>"010000001",
  51369=>"000101010",
  51370=>"110111000",
  51371=>"011000000",
  51372=>"111111110",
  51373=>"001001000",
  51374=>"100000100",
  51375=>"001001111",
  51376=>"111001110",
  51377=>"100011011",
  51378=>"111111000",
  51379=>"001010000",
  51380=>"001100111",
  51381=>"110010000",
  51382=>"000100111",
  51383=>"110110000",
  51384=>"011011110",
  51385=>"000000110",
  51386=>"111000000",
  51387=>"001111111",
  51388=>"100110111",
  51389=>"111110000",
  51390=>"110110011",
  51391=>"000000000",
  51392=>"001001111",
  51393=>"000111000",
  51394=>"100101111",
  51395=>"000010001",
  51396=>"101101000",
  51397=>"001001001",
  51398=>"001010010",
  51399=>"110101001",
  51400=>"111101011",
  51401=>"000111111",
  51402=>"001100110",
  51403=>"111110110",
  51404=>"011100110",
  51405=>"011000000",
  51406=>"000000000",
  51407=>"110110111",
  51408=>"000000000",
  51409=>"110100001",
  51410=>"011010000",
  51411=>"001111100",
  51412=>"000010000",
  51413=>"001100100",
  51414=>"110000000",
  51415=>"101111111",
  51416=>"100111101",
  51417=>"000000000",
  51418=>"000100111",
  51419=>"101000000",
  51420=>"100010001",
  51421=>"010111110",
  51422=>"110111010",
  51423=>"001001000",
  51424=>"101110010",
  51425=>"101001111",
  51426=>"000000000",
  51427=>"001110110",
  51428=>"111001000",
  51429=>"110010000",
  51430=>"110010101",
  51431=>"111111111",
  51432=>"000000000",
  51433=>"000000000",
  51434=>"111100000",
  51435=>"000000000",
  51436=>"000000000",
  51437=>"010001010",
  51438=>"001000001",
  51439=>"011110000",
  51440=>"111110000",
  51441=>"000000000",
  51442=>"101000011",
  51443=>"100111011",
  51444=>"110100110",
  51445=>"100100000",
  51446=>"000001000",
  51447=>"001001010",
  51448=>"000000000",
  51449=>"101101001",
  51450=>"111111111",
  51451=>"000111111",
  51452=>"001101111",
  51453=>"011000000",
  51454=>"010100100",
  51455=>"000001111",
  51456=>"011010100",
  51457=>"110110110",
  51458=>"111000000",
  51459=>"110110001",
  51460=>"000111111",
  51461=>"100000100",
  51462=>"111111000",
  51463=>"110100110",
  51464=>"111001111",
  51465=>"110000000",
  51466=>"000000100",
  51467=>"100111111",
  51468=>"100000000",
  51469=>"000111111",
  51470=>"000000000",
  51471=>"110100000",
  51472=>"110110110",
  51473=>"111111110",
  51474=>"111011011",
  51475=>"000110101",
  51476=>"111110111",
  51477=>"110111000",
  51478=>"010001001",
  51479=>"110010110",
  51480=>"001110101",
  51481=>"110100111",
  51482=>"010111000",
  51483=>"111011010",
  51484=>"101110111",
  51485=>"010010111",
  51486=>"111000010",
  51487=>"100101001",
  51488=>"100000100",
  51489=>"010110111",
  51490=>"101001000",
  51491=>"101111010",
  51492=>"001000001",
  51493=>"000010010",
  51494=>"111001001",
  51495=>"110110110",
  51496=>"100000000",
  51497=>"001111110",
  51498=>"110100000",
  51499=>"101111111",
  51500=>"000011001",
  51501=>"111001000",
  51502=>"101111000",
  51503=>"111110110",
  51504=>"110000001",
  51505=>"000011111",
  51506=>"011110010",
  51507=>"011010001",
  51508=>"111010000",
  51509=>"000000110",
  51510=>"000100110",
  51511=>"000000110",
  51512=>"110000110",
  51513=>"010110100",
  51514=>"101000000",
  51515=>"000000000",
  51516=>"100000011",
  51517=>"000101001",
  51518=>"000000000",
  51519=>"111001001",
  51520=>"111010110",
  51521=>"111111110",
  51522=>"111111001",
  51523=>"011011000",
  51524=>"000110000",
  51525=>"110000011",
  51526=>"000001111",
  51527=>"111011000",
  51528=>"100100100",
  51529=>"111001110",
  51530=>"000000001",
  51531=>"001000000",
  51532=>"111000000",
  51533=>"000000000",
  51534=>"001111101",
  51535=>"000000110",
  51536=>"000001101",
  51537=>"110010000",
  51538=>"110101010",
  51539=>"011001101",
  51540=>"111100000",
  51541=>"111000000",
  51542=>"011011111",
  51543=>"110111000",
  51544=>"000010010",
  51545=>"000001001",
  51546=>"000110111",
  51547=>"011000001",
  51548=>"011111111",
  51549=>"011011001",
  51550=>"111110010",
  51551=>"100100000",
  51552=>"100110111",
  51553=>"111110000",
  51554=>"111000000",
  51555=>"000011011",
  51556=>"000001101",
  51557=>"111111111",
  51558=>"100100110",
  51559=>"110001001",
  51560=>"100000001",
  51561=>"110000000",
  51562=>"101000000",
  51563=>"000011110",
  51564=>"000000010",
  51565=>"000110110",
  51566=>"000111001",
  51567=>"110000100",
  51568=>"101100101",
  51569=>"000111000",
  51570=>"000001111",
  51571=>"111010011",
  51572=>"110110000",
  51573=>"001000001",
  51574=>"001101000",
  51575=>"111000000",
  51576=>"111110100",
  51577=>"111110110",
  51578=>"011110101",
  51579=>"111000000",
  51580=>"100000011",
  51581=>"100000000",
  51582=>"110110011",
  51583=>"001001000",
  51584=>"000110110",
  51585=>"111000000",
  51586=>"111000010",
  51587=>"010010000",
  51588=>"000000111",
  51589=>"111001011",
  51590=>"000111001",
  51591=>"000110110",
  51592=>"001100001",
  51593=>"000010110",
  51594=>"000000001",
  51595=>"010000010",
  51596=>"101110000",
  51597=>"110000000",
  51598=>"011111000",
  51599=>"000000000",
  51600=>"111001001",
  51601=>"001011000",
  51602=>"001010000",
  51603=>"000000111",
  51604=>"001000110",
  51605=>"110111110",
  51606=>"000000010",
  51607=>"100001010",
  51608=>"110100000",
  51609=>"110000000",
  51610=>"111000000",
  51611=>"110111000",
  51612=>"000001001",
  51613=>"111000000",
  51614=>"011101000",
  51615=>"010111010",
  51616=>"000110001",
  51617=>"111111110",
  51618=>"101101000",
  51619=>"110011001",
  51620=>"111110110",
  51621=>"000100111",
  51622=>"111111001",
  51623=>"111111000",
  51624=>"000010000",
  51625=>"010000001",
  51626=>"111111001",
  51627=>"000110010",
  51628=>"001000111",
  51629=>"101001000",
  51630=>"100110111",
  51631=>"010001111",
  51632=>"101110110",
  51633=>"000100111",
  51634=>"110000000",
  51635=>"001001000",
  51636=>"101001000",
  51637=>"000000001",
  51638=>"010000111",
  51639=>"000000000",
  51640=>"001010000",
  51641=>"000001100",
  51642=>"101111000",
  51643=>"010010011",
  51644=>"111111001",
  51645=>"110111101",
  51646=>"111000000",
  51647=>"010010110",
  51648=>"001001111",
  51649=>"000001111",
  51650=>"110111111",
  51651=>"111001000",
  51652=>"000000010",
  51653=>"000001101",
  51654=>"010000000",
  51655=>"101001000",
  51656=>"110000000",
  51657=>"001100111",
  51658=>"000111111",
  51659=>"000110110",
  51660=>"111111000",
  51661=>"011100100",
  51662=>"000010111",
  51663=>"110010111",
  51664=>"000000000",
  51665=>"000101111",
  51666=>"000111101",
  51667=>"001111011",
  51668=>"101001000",
  51669=>"000111111",
  51670=>"011111000",
  51671=>"110110110",
  51672=>"000100110",
  51673=>"000110111",
  51674=>"011010000",
  51675=>"000000011",
  51676=>"010000001",
  51677=>"111000000",
  51678=>"010010111",
  51679=>"010110110",
  51680=>"111011111",
  51681=>"110001111",
  51682=>"111000000",
  51683=>"001100010",
  51684=>"111010000",
  51685=>"001001100",
  51686=>"100110100",
  51687=>"011111111",
  51688=>"111110000",
  51689=>"000010100",
  51690=>"001001100",
  51691=>"111111000",
  51692=>"000100000",
  51693=>"000110111",
  51694=>"010010010",
  51695=>"001101100",
  51696=>"111000110",
  51697=>"000111011",
  51698=>"111011001",
  51699=>"000001011",
  51700=>"100110010",
  51701=>"000000111",
  51702=>"000000000",
  51703=>"111111110",
  51704=>"000110110",
  51705=>"110001011",
  51706=>"111000111",
  51707=>"001001111",
  51708=>"111001000",
  51709=>"000010000",
  51710=>"000000000",
  51711=>"101001001",
  51712=>"010011001",
  51713=>"110111111",
  51714=>"111000101",
  51715=>"000010000",
  51716=>"001100110",
  51717=>"111010000",
  51718=>"101111111",
  51719=>"000100000",
  51720=>"000100110",
  51721=>"000101100",
  51722=>"000000011",
  51723=>"110111000",
  51724=>"000000100",
  51725=>"011000100",
  51726=>"001011010",
  51727=>"111011001",
  51728=>"111111000",
  51729=>"100101101",
  51730=>"010111100",
  51731=>"111111000",
  51732=>"101110110",
  51733=>"000001011",
  51734=>"111011011",
  51735=>"011111000",
  51736=>"010011000",
  51737=>"010010000",
  51738=>"000111011",
  51739=>"000111111",
  51740=>"111000010",
  51741=>"000111111",
  51742=>"111000000",
  51743=>"000010010",
  51744=>"010010110",
  51745=>"000010000",
  51746=>"000000001",
  51747=>"000011111",
  51748=>"000010010",
  51749=>"011111010",
  51750=>"000100000",
  51751=>"111011111",
  51752=>"001011111",
  51753=>"000000000",
  51754=>"110111110",
  51755=>"111100100",
  51756=>"100111100",
  51757=>"101010000",
  51758=>"011010000",
  51759=>"111111100",
  51760=>"111101100",
  51761=>"101011001",
  51762=>"101110001",
  51763=>"111111000",
  51764=>"111000111",
  51765=>"000101010",
  51766=>"001110100",
  51767=>"010111010",
  51768=>"111101001",
  51769=>"000000000",
  51770=>"010011010",
  51771=>"101111101",
  51772=>"110110100",
  51773=>"101011011",
  51774=>"111111101",
  51775=>"010111111",
  51776=>"111101000",
  51777=>"111011000",
  51778=>"111000000",
  51779=>"111111011",
  51780=>"110111010",
  51781=>"000111011",
  51782=>"111000010",
  51783=>"111111010",
  51784=>"000110100",
  51785=>"000111000",
  51786=>"000111000",
  51787=>"000010000",
  51788=>"111000000",
  51789=>"000011000",
  51790=>"000100010",
  51791=>"111000111",
  51792=>"010111111",
  51793=>"000111111",
  51794=>"011111010",
  51795=>"111011001",
  51796=>"101111010",
  51797=>"111011011",
  51798=>"100111011",
  51799=>"111101111",
  51800=>"110110100",
  51801=>"011011011",
  51802=>"000011011",
  51803=>"110111000",
  51804=>"111110000",
  51805=>"100111011",
  51806=>"110000100",
  51807=>"111101110",
  51808=>"100111111",
  51809=>"010010011",
  51810=>"111101111",
  51811=>"110100110",
  51812=>"000010000",
  51813=>"001010011",
  51814=>"000000000",
  51815=>"000111000",
  51816=>"110111010",
  51817=>"111111101",
  51818=>"000011110",
  51819=>"110101000",
  51820=>"000000100",
  51821=>"000111000",
  51822=>"110111000",
  51823=>"011111111",
  51824=>"100110111",
  51825=>"000000111",
  51826=>"110011001",
  51827=>"100001101",
  51828=>"110010010",
  51829=>"011110000",
  51830=>"101101100",
  51831=>"110111101",
  51832=>"111111110",
  51833=>"000111110",
  51834=>"001000010",
  51835=>"000000000",
  51836=>"100110110",
  51837=>"011110100",
  51838=>"101100111",
  51839=>"010000111",
  51840=>"111110000",
  51841=>"111100000",
  51842=>"010111111",
  51843=>"000011011",
  51844=>"100000000",
  51845=>"110110100",
  51846=>"111111000",
  51847=>"010111011",
  51848=>"001011011",
  51849=>"000001010",
  51850=>"000011000",
  51851=>"111111000",
  51852=>"101010011",
  51853=>"111101010",
  51854=>"110101111",
  51855=>"101001010",
  51856=>"100010011",
  51857=>"111111010",
  51858=>"010010000",
  51859=>"111111110",
  51860=>"011111111",
  51861=>"111101101",
  51862=>"101001001",
  51863=>"000110010",
  51864=>"000001000",
  51865=>"111111001",
  51866=>"011111000",
  51867=>"111000111",
  51868=>"000010000",
  51869=>"111001110",
  51870=>"111111101",
  51871=>"000000000",
  51872=>"000011000",
  51873=>"101111111",
  51874=>"010111101",
  51875=>"000100010",
  51876=>"100101100",
  51877=>"100110100",
  51878=>"001111000",
  51879=>"011100000",
  51880=>"101100101",
  51881=>"000110111",
  51882=>"100100100",
  51883=>"111000111",
  51884=>"111111001",
  51885=>"111011101",
  51886=>"011110111",
  51887=>"000000000",
  51888=>"011011111",
  51889=>"011011000",
  51890=>"110011000",
  51891=>"101110110",
  51892=>"000011000",
  51893=>"101111000",
  51894=>"000011011",
  51895=>"010010001",
  51896=>"011011001",
  51897=>"000011010",
  51898=>"010111111",
  51899=>"100110010",
  51900=>"111010101",
  51901=>"111001101",
  51902=>"000011011",
  51903=>"010001001",
  51904=>"010000010",
  51905=>"111111111",
  51906=>"111111000",
  51907=>"101111111",
  51908=>"000000001",
  51909=>"111111110",
  51910=>"011111110",
  51911=>"111111111",
  51912=>"000111010",
  51913=>"101111010",
  51914=>"111111011",
  51915=>"101101111",
  51916=>"111011011",
  51917=>"011011110",
  51918=>"111010111",
  51919=>"010111010",
  51920=>"101000001",
  51921=>"000010000",
  51922=>"000010010",
  51923=>"000011111",
  51924=>"111000111",
  51925=>"110110110",
  51926=>"101000000",
  51927=>"010111101",
  51928=>"000000000",
  51929=>"000111010",
  51930=>"000110000",
  51931=>"111000111",
  51932=>"111110110",
  51933=>"000000000",
  51934=>"000010000",
  51935=>"000011100",
  51936=>"111000010",
  51937=>"101100111",
  51938=>"000000101",
  51939=>"000001111",
  51940=>"101101000",
  51941=>"110110010",
  51942=>"111111111",
  51943=>"100110110",
  51944=>"110011000",
  51945=>"110111101",
  51946=>"011001100",
  51947=>"000000111",
  51948=>"000100110",
  51949=>"010111010",
  51950=>"111111111",
  51951=>"000110001",
  51952=>"111111000",
  51953=>"010110110",
  51954=>"011000001",
  51955=>"000110100",
  51956=>"000011011",
  51957=>"010000011",
  51958=>"111010010",
  51959=>"111111010",
  51960=>"011100000",
  51961=>"011010000",
  51962=>"000000000",
  51963=>"000111111",
  51964=>"011011000",
  51965=>"110110100",
  51966=>"000011001",
  51967=>"101000101",
  51968=>"100110011",
  51969=>"111011000",
  51970=>"001000001",
  51971=>"010011000",
  51972=>"111110110",
  51973=>"101101000",
  51974=>"000100101",
  51975=>"000011011",
  51976=>"111110110",
  51977=>"000111010",
  51978=>"100100110",
  51979=>"000000000",
  51980=>"111111111",
  51981=>"000000000",
  51982=>"011010000",
  51983=>"000000100",
  51984=>"000100111",
  51985=>"110100000",
  51986=>"001000000",
  51987=>"111110111",
  51988=>"000000000",
  51989=>"000100000",
  51990=>"000011111",
  51991=>"111111010",
  51992=>"111111010",
  51993=>"011000001",
  51994=>"001000000",
  51995=>"010100110",
  51996=>"100000100",
  51997=>"101000101",
  51998=>"001000111",
  51999=>"011111011",
  52000=>"100111000",
  52001=>"000010110",
  52002=>"100000000",
  52003=>"011000000",
  52004=>"011010100",
  52005=>"100101100",
  52006=>"000010010",
  52007=>"111000111",
  52008=>"000010001",
  52009=>"000000010",
  52010=>"111000111",
  52011=>"000111111",
  52012=>"010010011",
  52013=>"010010000",
  52014=>"100111111",
  52015=>"000000000",
  52016=>"100010010",
  52017=>"101111111",
  52018=>"110000011",
  52019=>"000010011",
  52020=>"110100101",
  52021=>"010100000",
  52022=>"000111110",
  52023=>"000110000",
  52024=>"010011010",
  52025=>"111101000",
  52026=>"000110000",
  52027=>"000100010",
  52028=>"000001110",
  52029=>"111111101",
  52030=>"000000110",
  52031=>"001101011",
  52032=>"111011000",
  52033=>"000000000",
  52034=>"010111000",
  52035=>"110111110",
  52036=>"000000000",
  52037=>"011001000",
  52038=>"111000010",
  52039=>"011100000",
  52040=>"001010111",
  52041=>"111001111",
  52042=>"011000010",
  52043=>"101000000",
  52044=>"111100111",
  52045=>"111111111",
  52046=>"111111111",
  52047=>"110111111",
  52048=>"001001011",
  52049=>"111111111",
  52050=>"000000110",
  52051=>"000011001",
  52052=>"000001100",
  52053=>"000011100",
  52054=>"100110110",
  52055=>"011000111",
  52056=>"111001111",
  52057=>"111111001",
  52058=>"001001001",
  52059=>"001000000",
  52060=>"000000000",
  52061=>"101111001",
  52062=>"000000000",
  52063=>"011111100",
  52064=>"111111101",
  52065=>"100000000",
  52066=>"011101111",
  52067=>"000000000",
  52068=>"010011011",
  52069=>"000001000",
  52070=>"000000000",
  52071=>"111111110",
  52072=>"100010000",
  52073=>"000100000",
  52074=>"000010110",
  52075=>"100000100",
  52076=>"111100000",
  52077=>"000100100",
  52078=>"000000111",
  52079=>"100100111",
  52080=>"100000000",
  52081=>"100100010",
  52082=>"000110010",
  52083=>"011110100",
  52084=>"100000011",
  52085=>"111000000",
  52086=>"111010000",
  52087=>"010000000",
  52088=>"111111000",
  52089=>"010111010",
  52090=>"000100010",
  52091=>"110011011",
  52092=>"110001001",
  52093=>"000011010",
  52094=>"100100001",
  52095=>"011101101",
  52096=>"000111000",
  52097=>"100111110",
  52098=>"000010000",
  52099=>"111111111",
  52100=>"000000000",
  52101=>"000010000",
  52102=>"101110011",
  52103=>"001000010",
  52104=>"011110000",
  52105=>"010101100",
  52106=>"011000010",
  52107=>"000111011",
  52108=>"000000000",
  52109=>"111100000",
  52110=>"110110000",
  52111=>"100000000",
  52112=>"110110111",
  52113=>"000010000",
  52114=>"000000010",
  52115=>"100000110",
  52116=>"111000000",
  52117=>"100111111",
  52118=>"111110100",
  52119=>"011111011",
  52120=>"000100000",
  52121=>"011111010",
  52122=>"101101111",
  52123=>"111110000",
  52124=>"000000011",
  52125=>"010111111",
  52126=>"100011010",
  52127=>"110111110",
  52128=>"011011011",
  52129=>"000110000",
  52130=>"111110111",
  52131=>"100111111",
  52132=>"000110010",
  52133=>"100110110",
  52134=>"011000011",
  52135=>"111100110",
  52136=>"110110100",
  52137=>"111111101",
  52138=>"010011010",
  52139=>"111111100",
  52140=>"101101100",
  52141=>"011101111",
  52142=>"100011010",
  52143=>"001111111",
  52144=>"100000001",
  52145=>"100111111",
  52146=>"000011011",
  52147=>"110111111",
  52148=>"111011101",
  52149=>"111010000",
  52150=>"001000000",
  52151=>"001100000",
  52152=>"100110100",
  52153=>"101010100",
  52154=>"110000000",
  52155=>"111000000",
  52156=>"011000000",
  52157=>"010101111",
  52158=>"110110010",
  52159=>"000000000",
  52160=>"000111111",
  52161=>"010111010",
  52162=>"100110100",
  52163=>"000000101",
  52164=>"000000100",
  52165=>"000110111",
  52166=>"001111000",
  52167=>"000000000",
  52168=>"111101000",
  52169=>"001000000",
  52170=>"111100001",
  52171=>"000100010",
  52172=>"010010010",
  52173=>"001100100",
  52174=>"100111000",
  52175=>"101111111",
  52176=>"000010000",
  52177=>"110111010",
  52178=>"111011001",
  52179=>"111111011",
  52180=>"011011011",
  52181=>"110111000",
  52182=>"010010010",
  52183=>"111111110",
  52184=>"010111111",
  52185=>"000000000",
  52186=>"000110111",
  52187=>"000000000",
  52188=>"010110000",
  52189=>"111001011",
  52190=>"000000000",
  52191=>"111001111",
  52192=>"000000101",
  52193=>"000011000",
  52194=>"000101111",
  52195=>"111011111",
  52196=>"011010010",
  52197=>"000000000",
  52198=>"111000100",
  52199=>"110111110",
  52200=>"111100011",
  52201=>"001001011",
  52202=>"101000000",
  52203=>"111110111",
  52204=>"000100101",
  52205=>"111101111",
  52206=>"001101000",
  52207=>"000010000",
  52208=>"111111001",
  52209=>"110011011",
  52210=>"100111010",
  52211=>"100110000",
  52212=>"000011111",
  52213=>"000000001",
  52214=>"101011000",
  52215=>"111010100",
  52216=>"000000000",
  52217=>"000000110",
  52218=>"111111111",
  52219=>"000100100",
  52220=>"100111111",
  52221=>"000001000",
  52222=>"111111011",
  52223=>"111000000",
  52224=>"111110111",
  52225=>"000000001",
  52226=>"111101000",
  52227=>"111111001",
  52228=>"111010000",
  52229=>"011011000",
  52230=>"000101100",
  52231=>"000111000",
  52232=>"111111000",
  52233=>"000000101",
  52234=>"110100000",
  52235=>"110111110",
  52236=>"111111101",
  52237=>"111111110",
  52238=>"111111000",
  52239=>"000011111",
  52240=>"111011000",
  52241=>"111101001",
  52242=>"111111101",
  52243=>"100101001",
  52244=>"111111000",
  52245=>"111111000",
  52246=>"000000111",
  52247=>"100001111",
  52248=>"111111001",
  52249=>"110000010",
  52250=>"111111101",
  52251=>"000000101",
  52252=>"000000000",
  52253=>"010111101",
  52254=>"111010110",
  52255=>"111000001",
  52256=>"011111111",
  52257=>"110010000",
  52258=>"000100110",
  52259=>"000000000",
  52260=>"000010010",
  52261=>"001001111",
  52262=>"111111000",
  52263=>"000000110",
  52264=>"111111001",
  52265=>"000111110",
  52266=>"000000111",
  52267=>"000000000",
  52268=>"000000110",
  52269=>"100101001",
  52270=>"000010100",
  52271=>"111001000",
  52272=>"000010111",
  52273=>"000010111",
  52274=>"010111000",
  52275=>"000010111",
  52276=>"100001111",
  52277=>"011101111",
  52278=>"011111111",
  52279=>"101010111",
  52280=>"101000101",
  52281=>"111100000",
  52282=>"000111111",
  52283=>"110101000",
  52284=>"000010011",
  52285=>"000111111",
  52286=>"011000000",
  52287=>"000000011",
  52288=>"111100000",
  52289=>"000010010",
  52290=>"101111000",
  52291=>"100101100",
  52292=>"010111111",
  52293=>"000011001",
  52294=>"010000111",
  52295=>"000000001",
  52296=>"010101010",
  52297=>"010011000",
  52298=>"111111101",
  52299=>"101111111",
  52300=>"000010000",
  52301=>"011000001",
  52302=>"010011011",
  52303=>"000111111",
  52304=>"111101101",
  52305=>"011011111",
  52306=>"000001111",
  52307=>"000110111",
  52308=>"011111000",
  52309=>"000010110",
  52310=>"100010001",
  52311=>"111111110",
  52312=>"100100000",
  52313=>"000000001",
  52314=>"001000000",
  52315=>"100000010",
  52316=>"101101000",
  52317=>"011110000",
  52318=>"111111010",
  52319=>"001001011",
  52320=>"001000011",
  52321=>"000111101",
  52322=>"111111000",
  52323=>"110110011",
  52324=>"100111000",
  52325=>"000101111",
  52326=>"000100100",
  52327=>"000000000",
  52328=>"110010101",
  52329=>"111111111",
  52330=>"000000111",
  52331=>"000000011",
  52332=>"000111001",
  52333=>"101000000",
  52334=>"111111000",
  52335=>"000000111",
  52336=>"000001000",
  52337=>"000000000",
  52338=>"110111110",
  52339=>"011111101",
  52340=>"000000000",
  52341=>"111101000",
  52342=>"000001111",
  52343=>"000001000",
  52344=>"001101111",
  52345=>"000000110",
  52346=>"000001000",
  52347=>"111110001",
  52348=>"010011001",
  52349=>"000011111",
  52350=>"111111110",
  52351=>"001000000",
  52352=>"000010010",
  52353=>"100011111",
  52354=>"000000111",
  52355=>"000111100",
  52356=>"101101100",
  52357=>"111101111",
  52358=>"000000111",
  52359=>"010110000",
  52360=>"000010000",
  52361=>"001101000",
  52362=>"111111000",
  52363=>"010111111",
  52364=>"111111000",
  52365=>"111001111",
  52366=>"000000001",
  52367=>"111111000",
  52368=>"110110100",
  52369=>"111101101",
  52370=>"000000111",
  52371=>"000110110",
  52372=>"111010000",
  52373=>"111000000",
  52374=>"111000110",
  52375=>"010110100",
  52376=>"000000011",
  52377=>"000000111",
  52378=>"111111010",
  52379=>"111111000",
  52380=>"000001000",
  52381=>"000110001",
  52382=>"000000111",
  52383=>"000111001",
  52384=>"010100010",
  52385=>"111000010",
  52386=>"011000110",
  52387=>"000000000",
  52388=>"110000000",
  52389=>"001011000",
  52390=>"000000010",
  52391=>"000001000",
  52392=>"111000000",
  52393=>"111101101",
  52394=>"111111000",
  52395=>"101111000",
  52396=>"001000000",
  52397=>"010111000",
  52398=>"111010111",
  52399=>"011010001",
  52400=>"000000001",
  52401=>"111001001",
  52402=>"100100001",
  52403=>"000000000",
  52404=>"001110111",
  52405=>"011101111",
  52406=>"111101100",
  52407=>"000001011",
  52408=>"000000000",
  52409=>"000000000",
  52410=>"000000101",
  52411=>"000010111",
  52412=>"111111100",
  52413=>"111010000",
  52414=>"011011000",
  52415=>"010111101",
  52416=>"111111000",
  52417=>"001000111",
  52418=>"101111011",
  52419=>"000110011",
  52420=>"000000010",
  52421=>"110001000",
  52422=>"000000000",
  52423=>"110110010",
  52424=>"000100011",
  52425=>"111100100",
  52426=>"110001000",
  52427=>"111000000",
  52428=>"010000000",
  52429=>"000110100",
  52430=>"000000100",
  52431=>"111110000",
  52432=>"001010111",
  52433=>"011011001",
  52434=>"111111000",
  52435=>"000011111",
  52436=>"111001000",
  52437=>"101110110",
  52438=>"111111000",
  52439=>"001110111",
  52440=>"000111111",
  52441=>"111111000",
  52442=>"000001000",
  52443=>"011111101",
  52444=>"000111111",
  52445=>"001100110",
  52446=>"001100001",
  52447=>"111110111",
  52448=>"111111000",
  52449=>"111101001",
  52450=>"010010111",
  52451=>"111111000",
  52452=>"111011001",
  52453=>"111000000",
  52454=>"001111011",
  52455=>"000010110",
  52456=>"010010111",
  52457=>"000000101",
  52458=>"011001001",
  52459=>"101001001",
  52460=>"101101010",
  52461=>"000000010",
  52462=>"010111000",
  52463=>"000110000",
  52464=>"000000111",
  52465=>"110010000",
  52466=>"000000000",
  52467=>"000111111",
  52468=>"001011110",
  52469=>"111110000",
  52470=>"000000100",
  52471=>"010111000",
  52472=>"111011111",
  52473=>"110000111",
  52474=>"000010000",
  52475=>"111110001",
  52476=>"100000111",
  52477=>"000000101",
  52478=>"010000111",
  52479=>"000000000",
  52480=>"000111110",
  52481=>"000100000",
  52482=>"001100100",
  52483=>"000110000",
  52484=>"000011110",
  52485=>"001010110",
  52486=>"110100010",
  52487=>"000000011",
  52488=>"110100100",
  52489=>"000000010",
  52490=>"111111010",
  52491=>"000011000",
  52492=>"100100011",
  52493=>"010111010",
  52494=>"000101001",
  52495=>"100000100",
  52496=>"111100001",
  52497=>"111110100",
  52498=>"101100101",
  52499=>"100000000",
  52500=>"101001100",
  52501=>"000011111",
  52502=>"111110000",
  52503=>"000011010",
  52504=>"011111100",
  52505=>"011010011",
  52506=>"001100100",
  52507=>"000100000",
  52508=>"101011111",
  52509=>"111011010",
  52510=>"011111111",
  52511=>"000000010",
  52512=>"000100000",
  52513=>"000000000",
  52514=>"111001111",
  52515=>"111111011",
  52516=>"000001000",
  52517=>"010000101",
  52518=>"101000100",
  52519=>"000111101",
  52520=>"111101111",
  52521=>"001000101",
  52522=>"000000100",
  52523=>"111100100",
  52524=>"100110001",
  52525=>"111111101",
  52526=>"100101111",
  52527=>"010111000",
  52528=>"000010000",
  52529=>"011011010",
  52530=>"011101011",
  52531=>"000111111",
  52532=>"000101111",
  52533=>"100010101",
  52534=>"010100000",
  52535=>"010011011",
  52536=>"111100111",
  52537=>"101111101",
  52538=>"111100000",
  52539=>"010011011",
  52540=>"001011001",
  52541=>"111111111",
  52542=>"000000000",
  52543=>"110111011",
  52544=>"010100100",
  52545=>"111011100",
  52546=>"101000000",
  52547=>"111000101",
  52548=>"111000010",
  52549=>"000000100",
  52550=>"000011010",
  52551=>"110001001",
  52552=>"100100110",
  52553=>"010011010",
  52554=>"001000100",
  52555=>"000011011",
  52556=>"101100111",
  52557=>"110000110",
  52558=>"100110111",
  52559=>"110010111",
  52560=>"011000000",
  52561=>"011010000",
  52562=>"000010111",
  52563=>"001001000",
  52564=>"111101000",
  52565=>"010000000",
  52566=>"100110010",
  52567=>"011111111",
  52568=>"000001100",
  52569=>"000100110",
  52570=>"000110110",
  52571=>"001011000",
  52572=>"100100100",
  52573=>"001001001",
  52574=>"111111100",
  52575=>"000111011",
  52576=>"111100100",
  52577=>"001000100",
  52578=>"111000001",
  52579=>"010111011",
  52580=>"000000000",
  52581=>"000100110",
  52582=>"000000000",
  52583=>"000000010",
  52584=>"100111010",
  52585=>"001001111",
  52586=>"111000100",
  52587=>"110001111",
  52588=>"111000000",
  52589=>"011111111",
  52590=>"000011010",
  52591=>"000000010",
  52592=>"001011011",
  52593=>"011000000",
  52594=>"100001110",
  52595=>"100100000",
  52596=>"011111000",
  52597=>"100101111",
  52598=>"100010111",
  52599=>"111000110",
  52600=>"011100110",
  52601=>"100000110",
  52602=>"010010000",
  52603=>"101111000",
  52604=>"110111011",
  52605=>"100111110",
  52606=>"110000000",
  52607=>"100011011",
  52608=>"011010000",
  52609=>"000000001",
  52610=>"010011000",
  52611=>"000011010",
  52612=>"011011001",
  52613=>"000011011",
  52614=>"101101000",
  52615=>"001101111",
  52616=>"000110000",
  52617=>"110111010",
  52618=>"000111000",
  52619=>"100111111",
  52620=>"000101100",
  52621=>"101000100",
  52622=>"100111111",
  52623=>"110101001",
  52624=>"101110110",
  52625=>"011000000",
  52626=>"000011011",
  52627=>"110010101",
  52628=>"000000000",
  52629=>"001101101",
  52630=>"111100100",
  52631=>"111100110",
  52632=>"010000000",
  52633=>"101101011",
  52634=>"111000000",
  52635=>"111011111",
  52636=>"000011011",
  52637=>"100111111",
  52638=>"011111110",
  52639=>"111101010",
  52640=>"101011110",
  52641=>"111110100",
  52642=>"000101111",
  52643=>"110111110",
  52644=>"000010100",
  52645=>"100110110",
  52646=>"110001101",
  52647=>"110100000",
  52648=>"000000000",
  52649=>"111111100",
  52650=>"111100000",
  52651=>"000101100",
  52652=>"000001000",
  52653=>"000001011",
  52654=>"110011000",
  52655=>"111001100",
  52656=>"111100100",
  52657=>"001011001",
  52658=>"101100101",
  52659=>"100100111",
  52660=>"100011001",
  52661=>"000000100",
  52662=>"111100100",
  52663=>"001100001",
  52664=>"111010010",
  52665=>"000011011",
  52666=>"101011000",
  52667=>"000111100",
  52668=>"111011011",
  52669=>"111111111",
  52670=>"000000011",
  52671=>"001000101",
  52672=>"111101111",
  52673=>"000000111",
  52674=>"011011000",
  52675=>"000000100",
  52676=>"000011100",
  52677=>"110110110",
  52678=>"000011011",
  52679=>"111101111",
  52680=>"111111000",
  52681=>"000000000",
  52682=>"000110100",
  52683=>"000011011",
  52684=>"101101110",
  52685=>"001111110",
  52686=>"000100101",
  52687=>"010001001",
  52688=>"111111100",
  52689=>"111011011",
  52690=>"011010010",
  52691=>"111111000",
  52692=>"010100010",
  52693=>"000100100",
  52694=>"000000000",
  52695=>"010011000",
  52696=>"010111011",
  52697=>"010111100",
  52698=>"110110111",
  52699=>"010100100",
  52700=>"100001000",
  52701=>"110100000",
  52702=>"111101111",
  52703=>"100000000",
  52704=>"100100000",
  52705=>"111111001",
  52706=>"001011101",
  52707=>"001011000",
  52708=>"111010000",
  52709=>"000010100",
  52710=>"101010010",
  52711=>"010111100",
  52712=>"111000101",
  52713=>"010101001",
  52714=>"101000011",
  52715=>"111101101",
  52716=>"000000111",
  52717=>"000000000",
  52718=>"111100010",
  52719=>"011100100",
  52720=>"100100111",
  52721=>"100011001",
  52722=>"101011111",
  52723=>"110101100",
  52724=>"000001011",
  52725=>"000101000",
  52726=>"100000101",
  52727=>"111111000",
  52728=>"000001000",
  52729=>"111000010",
  52730=>"010000000",
  52731=>"011011101",
  52732=>"000000000",
  52733=>"000011011",
  52734=>"001001000",
  52735=>"000011011",
  52736=>"011000000",
  52737=>"000010000",
  52738=>"101101111",
  52739=>"000100111",
  52740=>"100011010",
  52741=>"011000010",
  52742=>"011111010",
  52743=>"000011110",
  52744=>"000000000",
  52745=>"000000101",
  52746=>"001011001",
  52747=>"100111000",
  52748=>"001000110",
  52749=>"101111101",
  52750=>"011111100",
  52751=>"110001111",
  52752=>"010101111",
  52753=>"101111000",
  52754=>"101111111",
  52755=>"000010100",
  52756=>"000000010",
  52757=>"010010000",
  52758=>"000000111",
  52759=>"000111100",
  52760=>"111100111",
  52761=>"001001000",
  52762=>"100100110",
  52763=>"111000100",
  52764=>"000000000",
  52765=>"101000101",
  52766=>"010000101",
  52767=>"100111000",
  52768=>"010010111",
  52769=>"110110111",
  52770=>"111010000",
  52771=>"000000000",
  52772=>"000111001",
  52773=>"011000000",
  52774=>"010111000",
  52775=>"001010000",
  52776=>"000000111",
  52777=>"011110101",
  52778=>"010010100",
  52779=>"111101111",
  52780=>"001000001",
  52781=>"101000111",
  52782=>"011000101",
  52783=>"100000111",
  52784=>"010101000",
  52785=>"110001000",
  52786=>"000000101",
  52787=>"000000000",
  52788=>"111110101",
  52789=>"010001000",
  52790=>"011011010",
  52791=>"000000001",
  52792=>"111000010",
  52793=>"000000101",
  52794=>"000001010",
  52795=>"111000101",
  52796=>"000001000",
  52797=>"111010110",
  52798=>"000000111",
  52799=>"110000100",
  52800=>"100000001",
  52801=>"011000101",
  52802=>"001111111",
  52803=>"001001000",
  52804=>"000000000",
  52805=>"100000011",
  52806=>"010011000",
  52807=>"111111111",
  52808=>"100101001",
  52809=>"101000110",
  52810=>"001000110",
  52811=>"100101001",
  52812=>"000000100",
  52813=>"101100100",
  52814=>"001110000",
  52815=>"101000000",
  52816=>"111111111",
  52817=>"101111111",
  52818=>"011000111",
  52819=>"011000010",
  52820=>"101000101",
  52821=>"110111111",
  52822=>"001111101",
  52823=>"000011001",
  52824=>"001011111",
  52825=>"000011010",
  52826=>"100111000",
  52827=>"011111100",
  52828=>"010000000",
  52829=>"001101111",
  52830=>"111000101",
  52831=>"100100001",
  52832=>"111001010",
  52833=>"111000111",
  52834=>"000000111",
  52835=>"011001011",
  52836=>"101111011",
  52837=>"011011110",
  52838=>"111101001",
  52839=>"000000000",
  52840=>"110100101",
  52841=>"011011111",
  52842=>"111011000",
  52843=>"011111001",
  52844=>"111000111",
  52845=>"111011100",
  52846=>"001000101",
  52847=>"000111010",
  52848=>"100000110",
  52849=>"100010010",
  52850=>"110010010",
  52851=>"101000000",
  52852=>"011010000",
  52853=>"000100010",
  52854=>"010010000",
  52855=>"100101101",
  52856=>"000000111",
  52857=>"000111110",
  52858=>"110110001",
  52859=>"101111111",
  52860=>"111010011",
  52861=>"101000111",
  52862=>"010111111",
  52863=>"100000101",
  52864=>"111010001",
  52865=>"000000100",
  52866=>"000000000",
  52867=>"000010100",
  52868=>"111100000",
  52869=>"100000000",
  52870=>"110100100",
  52871=>"010111111",
  52872=>"111100101",
  52873=>"110000000",
  52874=>"011010011",
  52875=>"000111111",
  52876=>"010000000",
  52877=>"010101111",
  52878=>"111101111",
  52879=>"000001111",
  52880=>"111100000",
  52881=>"010110000",
  52882=>"111110000",
  52883=>"010010011",
  52884=>"101111011",
  52885=>"000010110",
  52886=>"000100111",
  52887=>"100100000",
  52888=>"010010111",
  52889=>"001000001",
  52890=>"100111101",
  52891=>"000000111",
  52892=>"110000100",
  52893=>"111101111",
  52894=>"111111000",
  52895=>"100101000",
  52896=>"111111100",
  52897=>"000000101",
  52898=>"101111011",
  52899=>"111111100",
  52900=>"101110000",
  52901=>"100111001",
  52902=>"011000000",
  52903=>"010001000",
  52904=>"000000010",
  52905=>"111101111",
  52906=>"000000000",
  52907=>"000010010",
  52908=>"000000000",
  52909=>"000001011",
  52910=>"010001011",
  52911=>"010000000",
  52912=>"101001111",
  52913=>"011110100",
  52914=>"101101111",
  52915=>"100110001",
  52916=>"111111111",
  52917=>"011000010",
  52918=>"110001001",
  52919=>"011011000",
  52920=>"011000110",
  52921=>"110111010",
  52922=>"111000000",
  52923=>"110000000",
  52924=>"011001101",
  52925=>"111011000",
  52926=>"000000011",
  52927=>"000000000",
  52928=>"111001001",
  52929=>"010101101",
  52930=>"111111000",
  52931=>"111011010",
  52932=>"000111000",
  52933=>"101111101",
  52934=>"010011000",
  52935=>"011000111",
  52936=>"000111111",
  52937=>"101100100",
  52938=>"111111111",
  52939=>"000110000",
  52940=>"011011101",
  52941=>"100010110",
  52942=>"101111110",
  52943=>"110101111",
  52944=>"001110101",
  52945=>"111011110",
  52946=>"000000010",
  52947=>"110111000",
  52948=>"000100110",
  52949=>"000001101",
  52950=>"000000011",
  52951=>"010100111",
  52952=>"010000000",
  52953=>"000010010",
  52954=>"001101000",
  52955=>"101001111",
  52956=>"010000011",
  52957=>"100101101",
  52958=>"101111000",
  52959=>"011101010",
  52960=>"110101101",
  52961=>"001001010",
  52962=>"111101000",
  52963=>"111111000",
  52964=>"010101101",
  52965=>"100010000",
  52966=>"100111111",
  52967=>"010110100",
  52968=>"111110111",
  52969=>"111000011",
  52970=>"000110100",
  52971=>"110110000",
  52972=>"000110000",
  52973=>"010010000",
  52974=>"101000000",
  52975=>"000001010",
  52976=>"000110010",
  52977=>"011111100",
  52978=>"010000000",
  52979=>"001000110",
  52980=>"110011011",
  52981=>"111000000",
  52982=>"000010110",
  52983=>"001000110",
  52984=>"111000000",
  52985=>"011101111",
  52986=>"101000000",
  52987=>"111111110",
  52988=>"010101111",
  52989=>"000010000",
  52990=>"001001000",
  52991=>"010000001",
  52992=>"001000100",
  52993=>"000111111",
  52994=>"000000111",
  52995=>"000000001",
  52996=>"101000000",
  52997=>"000000110",
  52998=>"111001000",
  52999=>"010000001",
  53000=>"000000010",
  53001=>"111000000",
  53002=>"110001100",
  53003=>"000101101",
  53004=>"000010111",
  53005=>"111101000",
  53006=>"000000000",
  53007=>"011101111",
  53008=>"111100000",
  53009=>"011010011",
  53010=>"000000111",
  53011=>"000010000",
  53012=>"111111111",
  53013=>"101101111",
  53014=>"011110000",
  53015=>"111111100",
  53016=>"111000101",
  53017=>"001001000",
  53018=>"011000000",
  53019=>"000010110",
  53020=>"111110000",
  53021=>"000000000",
  53022=>"000010110",
  53023=>"000000001",
  53024=>"011001001",
  53025=>"000111100",
  53026=>"100101001",
  53027=>"000000010",
  53028=>"000000011",
  53029=>"010100001",
  53030=>"000010010",
  53031=>"010101001",
  53032=>"000010011",
  53033=>"111111010",
  53034=>"010010000",
  53035=>"100000101",
  53036=>"001011011",
  53037=>"011110110",
  53038=>"001010111",
  53039=>"100001101",
  53040=>"111010000",
  53041=>"000010110",
  53042=>"101011000",
  53043=>"101000000",
  53044=>"111101000",
  53045=>"001101000",
  53046=>"111100000",
  53047=>"001101100",
  53048=>"000111111",
  53049=>"000000111",
  53050=>"000010011",
  53051=>"110110011",
  53052=>"011101001",
  53053=>"111111110",
  53054=>"000111101",
  53055=>"111000000",
  53056=>"111000011",
  53057=>"111111101",
  53058=>"000000010",
  53059=>"011001000",
  53060=>"000110111",
  53061=>"101111000",
  53062=>"001000001",
  53063=>"001000111",
  53064=>"111111100",
  53065=>"011000000",
  53066=>"001100000",
  53067=>"001111000",
  53068=>"000000111",
  53069=>"000000110",
  53070=>"000000011",
  53071=>"101000110",
  53072=>"101101000",
  53073=>"000101000",
  53074=>"110111111",
  53075=>"001000000",
  53076=>"111001001",
  53077=>"101100000",
  53078=>"100001000",
  53079=>"111000000",
  53080=>"111111111",
  53081=>"000110110",
  53082=>"001100110",
  53083=>"000011011",
  53084=>"000111110",
  53085=>"000110110",
  53086=>"101101111",
  53087=>"110100001",
  53088=>"111000000",
  53089=>"111101000",
  53090=>"000000111",
  53091=>"000011001",
  53092=>"000000001",
  53093=>"011111001",
  53094=>"111101000",
  53095=>"000001111",
  53096=>"000010000",
  53097=>"001111000",
  53098=>"001111111",
  53099=>"100001101",
  53100=>"110000111",
  53101=>"111111000",
  53102=>"001011111",
  53103=>"001010000",
  53104=>"001000111",
  53105=>"000111111",
  53106=>"010001100",
  53107=>"111101000",
  53108=>"010010110",
  53109=>"000001001",
  53110=>"011010000",
  53111=>"101001000",
  53112=>"000000010",
  53113=>"000110111",
  53114=>"000010111",
  53115=>"110010010",
  53116=>"001001001",
  53117=>"000000000",
  53118=>"001111111",
  53119=>"000001101",
  53120=>"111011000",
  53121=>"000110000",
  53122=>"111001011",
  53123=>"111100111",
  53124=>"000010111",
  53125=>"111101000",
  53126=>"110011000",
  53127=>"110100000",
  53128=>"100000010",
  53129=>"001000101",
  53130=>"111101000",
  53131=>"001001111",
  53132=>"000101011",
  53133=>"011011101",
  53134=>"000000011",
  53135=>"000001000",
  53136=>"000000110",
  53137=>"000000111",
  53138=>"101111001",
  53139=>"000101111",
  53140=>"111111000",
  53141=>"010010000",
  53142=>"100001000",
  53143=>"000010000",
  53144=>"110010011",
  53145=>"000111111",
  53146=>"010100000",
  53147=>"000000000",
  53148=>"000100001",
  53149=>"000000000",
  53150=>"001111101",
  53151=>"000000010",
  53152=>"101001111",
  53153=>"111111100",
  53154=>"000001001",
  53155=>"000100110",
  53156=>"000110111",
  53157=>"001110110",
  53158=>"001000001",
  53159=>"011001001",
  53160=>"111111000",
  53161=>"011001000",
  53162=>"000111111",
  53163=>"000010111",
  53164=>"111111111",
  53165=>"000101111",
  53166=>"100101100",
  53167=>"111000000",
  53168=>"001001110",
  53169=>"000101100",
  53170=>"000000000",
  53171=>"000001011",
  53172=>"100110000",
  53173=>"000000000",
  53174=>"000000000",
  53175=>"000000011",
  53176=>"110100100",
  53177=>"111011001",
  53178=>"110100001",
  53179=>"000000111",
  53180=>"011111110",
  53181=>"000000001",
  53182=>"001000010",
  53183=>"111111010",
  53184=>"000000100",
  53185=>"000000111",
  53186=>"111111000",
  53187=>"000000010",
  53188=>"100000001",
  53189=>"100100110",
  53190=>"000011011",
  53191=>"000000011",
  53192=>"101101101",
  53193=>"000111011",
  53194=>"101000000",
  53195=>"000001110",
  53196=>"000000000",
  53197=>"110100100",
  53198=>"111100100",
  53199=>"010111101",
  53200=>"000100101",
  53201=>"011111100",
  53202=>"001100000",
  53203=>"000000101",
  53204=>"000001111",
  53205=>"110111001",
  53206=>"011000011",
  53207=>"110000000",
  53208=>"000111111",
  53209=>"000000000",
  53210=>"001011011",
  53211=>"011000000",
  53212=>"100011100",
  53213=>"001111110",
  53214=>"000000000",
  53215=>"110000010",
  53216=>"000010010",
  53217=>"000011011",
  53218=>"001001101",
  53219=>"011111111",
  53220=>"000000001",
  53221=>"000000100",
  53222=>"001000111",
  53223=>"000001011",
  53224=>"000000010",
  53225=>"111111100",
  53226=>"110101101",
  53227=>"111001000",
  53228=>"000111000",
  53229=>"000000100",
  53230=>"000000000",
  53231=>"000110111",
  53232=>"111101100",
  53233=>"000011011",
  53234=>"111000000",
  53235=>"001011011",
  53236=>"100100000",
  53237=>"000101111",
  53238=>"000100000",
  53239=>"000000110",
  53240=>"000010000",
  53241=>"000010000",
  53242=>"000000110",
  53243=>"111111100",
  53244=>"000100001",
  53245=>"000000000",
  53246=>"001000110",
  53247=>"100000000",
  53248=>"101100110",
  53249=>"110111101",
  53250=>"100000100",
  53251=>"000001000",
  53252=>"001011011",
  53253=>"111001001",
  53254=>"000000111",
  53255=>"111111101",
  53256=>"000000001",
  53257=>"110000000",
  53258=>"011111011",
  53259=>"110100101",
  53260=>"000000010",
  53261=>"000001111",
  53262=>"111110100",
  53263=>"000000110",
  53264=>"010000000",
  53265=>"011010000",
  53266=>"000111111",
  53267=>"000111101",
  53268=>"101111111",
  53269=>"101100000",
  53270=>"111011111",
  53271=>"101101000",
  53272=>"000110111",
  53273=>"001000010",
  53274=>"000000000",
  53275=>"111000000",
  53276=>"000111101",
  53277=>"011101000",
  53278=>"000101000",
  53279=>"011011000",
  53280=>"010111111",
  53281=>"100000000",
  53282=>"001111111",
  53283=>"101001111",
  53284=>"000110111",
  53285=>"000001001",
  53286=>"000011000",
  53287=>"100000110",
  53288=>"010000000",
  53289=>"000010000",
  53290=>"000001001",
  53291=>"101000100",
  53292=>"000111111",
  53293=>"111011011",
  53294=>"100101001",
  53295=>"000011110",
  53296=>"111000000",
  53297=>"011001111",
  53298=>"000010100",
  53299=>"010010000",
  53300=>"000010111",
  53301=>"111011001",
  53302=>"110100100",
  53303=>"111100000",
  53304=>"101111111",
  53305=>"111010110",
  53306=>"101000111",
  53307=>"101100101",
  53308=>"001001111",
  53309=>"111000101",
  53310=>"001000000",
  53311=>"000111001",
  53312=>"111111111",
  53313=>"000111101",
  53314=>"011000000",
  53315=>"100010001",
  53316=>"000001111",
  53317=>"000100000",
  53318=>"110100111",
  53319=>"000000110",
  53320=>"011010010",
  53321=>"111101101",
  53322=>"100000001",
  53323=>"001000000",
  53324=>"010100111",
  53325=>"011011010",
  53326=>"110110011",
  53327=>"001101100",
  53328=>"011101000",
  53329=>"101111111",
  53330=>"111100000",
  53331=>"110111000",
  53332=>"000000100",
  53333=>"010000000",
  53334=>"110111111",
  53335=>"000010000",
  53336=>"000011001",
  53337=>"110001011",
  53338=>"111001000",
  53339=>"000000011",
  53340=>"111000010",
  53341=>"101111110",
  53342=>"111111111",
  53343=>"100000001",
  53344=>"000000000",
  53345=>"110111100",
  53346=>"111101101",
  53347=>"001111010",
  53348=>"111000011",
  53349=>"111101111",
  53350=>"101110011",
  53351=>"010010101",
  53352=>"000010010",
  53353=>"101111111",
  53354=>"110111111",
  53355=>"000000000",
  53356=>"100111111",
  53357=>"111111000",
  53358=>"000100111",
  53359=>"000111111",
  53360=>"011111110",
  53361=>"101001000",
  53362=>"001001001",
  53363=>"000000000",
  53364=>"000101111",
  53365=>"100111111",
  53366=>"010111001",
  53367=>"000111111",
  53368=>"000010111",
  53369=>"000011111",
  53370=>"111000000",
  53371=>"110111111",
  53372=>"000000011",
  53373=>"000011011",
  53374=>"100100000",
  53375=>"100100100",
  53376=>"110101111",
  53377=>"000000100",
  53378=>"111101011",
  53379=>"101111111",
  53380=>"010111000",
  53381=>"111111110",
  53382=>"000110001",
  53383=>"011000000",
  53384=>"110100111",
  53385=>"110100000",
  53386=>"100011001",
  53387=>"000100000",
  53388=>"011100000",
  53389=>"000000010",
  53390=>"100000000",
  53391=>"111000001",
  53392=>"000010100",
  53393=>"000101101",
  53394=>"000000000",
  53395=>"000000000",
  53396=>"110110000",
  53397=>"111101001",
  53398=>"001010111",
  53399=>"010000000",
  53400=>"001000001",
  53401=>"000111111",
  53402=>"111000000",
  53403=>"110000010",
  53404=>"111000010",
  53405=>"000000000",
  53406=>"100111111",
  53407=>"111101101",
  53408=>"011001111",
  53409=>"010000000",
  53410=>"101000000",
  53411=>"000010111",
  53412=>"101001000",
  53413=>"010000100",
  53414=>"100001101",
  53415=>"011001111",
  53416=>"000000000",
  53417=>"100010001",
  53418=>"100100011",
  53419=>"000000000",
  53420=>"100111111",
  53421=>"111101111",
  53422=>"011010001",
  53423=>"111000000",
  53424=>"000000000",
  53425=>"110100100",
  53426=>"000010000",
  53427=>"000000011",
  53428=>"000111111",
  53429=>"111111010",
  53430=>"000001011",
  53431=>"000000000",
  53432=>"100110111",
  53433=>"011001000",
  53434=>"000001000",
  53435=>"000000000",
  53436=>"111101111",
  53437=>"000000101",
  53438=>"100000001",
  53439=>"011101111",
  53440=>"010100101",
  53441=>"111000000",
  53442=>"000111001",
  53443=>"111101101",
  53444=>"101001111",
  53445=>"111001001",
  53446=>"100011010",
  53447=>"111000001",
  53448=>"111101000",
  53449=>"100000000",
  53450=>"111111110",
  53451=>"110010000",
  53452=>"111111111",
  53453=>"111100100",
  53454=>"010100101",
  53455=>"000011111",
  53456=>"011011100",
  53457=>"111111110",
  53458=>"000000000",
  53459=>"000000010",
  53460=>"101100111",
  53461=>"001000001",
  53462=>"010011111",
  53463=>"010110010",
  53464=>"101111000",
  53465=>"010011000",
  53466=>"110100111",
  53467=>"101001000",
  53468=>"100110110",
  53469=>"000010011",
  53470=>"001001001",
  53471=>"000111011",
  53472=>"000111000",
  53473=>"111111000",
  53474=>"010110111",
  53475=>"010000000",
  53476=>"000000111",
  53477=>"001111111",
  53478=>"000000000",
  53479=>"000011111",
  53480=>"000000000",
  53481=>"011111101",
  53482=>"000110110",
  53483=>"011100000",
  53484=>"000000000",
  53485=>"000000111",
  53486=>"000000010",
  53487=>"111000111",
  53488=>"100100111",
  53489=>"110100000",
  53490=>"101100101",
  53491=>"011011111",
  53492=>"010011011",
  53493=>"111111000",
  53494=>"000000010",
  53495=>"111000000",
  53496=>"000000011",
  53497=>"111111111",
  53498=>"010010110",
  53499=>"111111111",
  53500=>"101111111",
  53501=>"010000000",
  53502=>"111000110",
  53503=>"111110100",
  53504=>"110010000",
  53505=>"000010111",
  53506=>"001001001",
  53507=>"111001000",
  53508=>"000010001",
  53509=>"100001111",
  53510=>"001001001",
  53511=>"000011000",
  53512=>"110100110",
  53513=>"000000010",
  53514=>"001000000",
  53515=>"000000001",
  53516=>"001001011",
  53517=>"100110110",
  53518=>"000100010",
  53519=>"110110001",
  53520=>"100110000",
  53521=>"110000110",
  53522=>"000001111",
  53523=>"000100110",
  53524=>"110110001",
  53525=>"000001001",
  53526=>"100110111",
  53527=>"110000110",
  53528=>"000000000",
  53529=>"100111110",
  53530=>"000000000",
  53531=>"101001000",
  53532=>"010110001",
  53533=>"001001110",
  53534=>"110110100",
  53535=>"011011000",
  53536=>"110110010",
  53537=>"010110001",
  53538=>"111001000",
  53539=>"110011100",
  53540=>"100100000",
  53541=>"110111001",
  53542=>"110110000",
  53543=>"001000100",
  53544=>"010110000",
  53545=>"110110010",
  53546=>"100110110",
  53547=>"000000111",
  53548=>"001110111",
  53549=>"101100110",
  53550=>"110110111",
  53551=>"110001001",
  53552=>"111111000",
  53553=>"100111100",
  53554=>"111010110",
  53555=>"111011110",
  53556=>"110000000",
  53557=>"001001111",
  53558=>"100001011",
  53559=>"000001001",
  53560=>"110000010",
  53561=>"001110110",
  53562=>"000001101",
  53563=>"111001001",
  53564=>"100100100",
  53565=>"111111001",
  53566=>"000000000",
  53567=>"110110111",
  53568=>"110110001",
  53569=>"110110000",
  53570=>"110111000",
  53571=>"111100000",
  53572=>"011111111",
  53573=>"110110100",
  53574=>"000000110",
  53575=>"111100000",
  53576=>"110011111",
  53577=>"110110010",
  53578=>"010000011",
  53579=>"010000010",
  53580=>"110100010",
  53581=>"000011000",
  53582=>"001101100",
  53583=>"001000110",
  53584=>"011011010",
  53585=>"100111110",
  53586=>"001001111",
  53587=>"111001100",
  53588=>"011000110",
  53589=>"010110110",
  53590=>"011010000",
  53591=>"101101000",
  53592=>"000001001",
  53593=>"110100111",
  53594=>"101101001",
  53595=>"011100110",
  53596=>"000000000",
  53597=>"000011010",
  53598=>"110100000",
  53599=>"110110110",
  53600=>"110110110",
  53601=>"110110110",
  53602=>"001001001",
  53603=>"110111000",
  53604=>"010110000",
  53605=>"100000110",
  53606=>"110110000",
  53607=>"001000010",
  53608=>"110110110",
  53609=>"111001001",
  53610=>"100010110",
  53611=>"111110101",
  53612=>"010110000",
  53613=>"001000001",
  53614=>"111001101",
  53615=>"000000000",
  53616=>"000100110",
  53617=>"110000001",
  53618=>"010100110",
  53619=>"111111110",
  53620=>"010111010",
  53621=>"000000000",
  53622=>"010010000",
  53623=>"110111000",
  53624=>"001000110",
  53625=>"111001000",
  53626=>"001001000",
  53627=>"000000001",
  53628=>"000110110",
  53629=>"110100100",
  53630=>"001101111",
  53631=>"110000100",
  53632=>"011100000",
  53633=>"110001000",
  53634=>"110000110",
  53635=>"010111100",
  53636=>"000000110",
  53637=>"111000101",
  53638=>"010110010",
  53639=>"000110001",
  53640=>"111011010",
  53641=>"111111111",
  53642=>"001110011",
  53643=>"111000000",
  53644=>"000000001",
  53645=>"001011111",
  53646=>"100000000",
  53647=>"011000000",
  53648=>"010010000",
  53649=>"111111001",
  53650=>"001001000",
  53651=>"111000001",
  53652=>"000110100",
  53653=>"000000110",
  53654=>"110110000",
  53655=>"000010000",
  53656=>"000001000",
  53657=>"001111110",
  53658=>"001001110",
  53659=>"100000001",
  53660=>"001001110",
  53661=>"000110110",
  53662=>"001110110",
  53663=>"101001001",
  53664=>"001011111",
  53665=>"100110110",
  53666=>"110100000",
  53667=>"010000111",
  53668=>"111110000",
  53669=>"000011000",
  53670=>"011011011",
  53671=>"000010000",
  53672=>"001101110",
  53673=>"000000110",
  53674=>"001001111",
  53675=>"001010010",
  53676=>"110111101",
  53677=>"110110110",
  53678=>"000011011",
  53679=>"001001111",
  53680=>"110110000",
  53681=>"011011000",
  53682=>"111000000",
  53683=>"011000000",
  53684=>"110100110",
  53685=>"111111111",
  53686=>"000000101",
  53687=>"000010101",
  53688=>"011010011",
  53689=>"001110110",
  53690=>"010110010",
  53691=>"111110110",
  53692=>"001100000",
  53693=>"111001111",
  53694=>"000000100",
  53695=>"101001011",
  53696=>"100001101",
  53697=>"001001111",
  53698=>"111000001",
  53699=>"100100100",
  53700=>"101000000",
  53701=>"100000001",
  53702=>"010011000",
  53703=>"000110101",
  53704=>"100110110",
  53705=>"000111000",
  53706=>"010111111",
  53707=>"000000000",
  53708=>"000110111",
  53709=>"000110110",
  53710=>"111001000",
  53711=>"100110010",
  53712=>"111001011",
  53713=>"100110100",
  53714=>"110011110",
  53715=>"011010111",
  53716=>"100100101",
  53717=>"010001000",
  53718=>"000110000",
  53719=>"000110110",
  53720=>"001001111",
  53721=>"000000000",
  53722=>"000100000",
  53723=>"001001001",
  53724=>"011100100",
  53725=>"001110111",
  53726=>"010000000",
  53727=>"110000010",
  53728=>"001000001",
  53729=>"100000001",
  53730=>"001001101",
  53731=>"011011000",
  53732=>"001001000",
  53733=>"001001111",
  53734=>"110000011",
  53735=>"010111110",
  53736=>"000000111",
  53737=>"011111110",
  53738=>"010000001",
  53739=>"000001000",
  53740=>"001001011",
  53741=>"001001111",
  53742=>"000001000",
  53743=>"000001000",
  53744=>"001001111",
  53745=>"011001000",
  53746=>"000101110",
  53747=>"000010110",
  53748=>"110101011",
  53749=>"011001001",
  53750=>"011001010",
  53751=>"110000110",
  53752=>"101101111",
  53753=>"001000111",
  53754=>"111001101",
  53755=>"011001000",
  53756=>"110110000",
  53757=>"001001001",
  53758=>"100101000",
  53759=>"000000000",
  53760=>"111101110",
  53761=>"000010001",
  53762=>"100100101",
  53763=>"000101101",
  53764=>"110111100",
  53765=>"100000001",
  53766=>"100100100",
  53767=>"111111011",
  53768=>"111000100",
  53769=>"000000010",
  53770=>"010011000",
  53771=>"000011011",
  53772=>"000000111",
  53773=>"101000110",
  53774=>"101011111",
  53775=>"011111000",
  53776=>"011011000",
  53777=>"000111101",
  53778=>"111100000",
  53779=>"000010111",
  53780=>"000100001",
  53781=>"011011000",
  53782=>"100100000",
  53783=>"000111110",
  53784=>"110100000",
  53785=>"011111010",
  53786=>"101111010",
  53787=>"101100111",
  53788=>"100100001",
  53789=>"101100000",
  53790=>"111101101",
  53791=>"000100000",
  53792=>"101101011",
  53793=>"100100000",
  53794=>"011011111",
  53795=>"000100100",
  53796=>"110111100",
  53797=>"010000110",
  53798=>"111111010",
  53799=>"100100000",
  53800=>"110111111",
  53801=>"000000000",
  53802=>"000000110",
  53803=>"101110111",
  53804=>"101011111",
  53805=>"000000011",
  53806=>"011011000",
  53807=>"111001000",
  53808=>"011000000",
  53809=>"100111111",
  53810=>"000110010",
  53811=>"010011011",
  53812=>"011011000",
  53813=>"101101011",
  53814=>"001011011",
  53815=>"101100011",
  53816=>"011100001",
  53817=>"101100000",
  53818=>"010011100",
  53819=>"111100111",
  53820=>"001111001",
  53821=>"011100010",
  53822=>"000000000",
  53823=>"110111011",
  53824=>"111101000",
  53825=>"000000010",
  53826=>"111011000",
  53827=>"001001101",
  53828=>"000100101",
  53829=>"000100011",
  53830=>"011011011",
  53831=>"100000101",
  53832=>"000000110",
  53833=>"101100111",
  53834=>"101100100",
  53835=>"011011001",
  53836=>"101100111",
  53837=>"001001001",
  53838=>"001101110",
  53839=>"100111110",
  53840=>"000000111",
  53841=>"111110100",
  53842=>"110111100",
  53843=>"100000100",
  53844=>"000100000",
  53845=>"011011101",
  53846=>"001011111",
  53847=>"111111000",
  53848=>"101100100",
  53849=>"000100110",
  53850=>"000111000",
  53851=>"011011000",
  53852=>"010011010",
  53853=>"100101000",
  53854=>"111110111",
  53855=>"100110000",
  53856=>"000000111",
  53857=>"000011000",
  53858=>"000000001",
  53859=>"100101111",
  53860=>"100111110",
  53861=>"100101110",
  53862=>"111111110",
  53863=>"100000000",
  53864=>"011111000",
  53865=>"100111011",
  53866=>"001000110",
  53867=>"010010000",
  53868=>"011000000",
  53869=>"011011000",
  53870=>"010011010",
  53871=>"001000100",
  53872=>"111111001",
  53873=>"011111100",
  53874=>"011011000",
  53875=>"100000000",
  53876=>"010111111",
  53877=>"100100111",
  53878=>"101010010",
  53879=>"000000111",
  53880=>"001100111",
  53881=>"000000000",
  53882=>"001100010",
  53883=>"000000100",
  53884=>"111010100",
  53885=>"001000100",
  53886=>"110011010",
  53887=>"101100101",
  53888=>"101000111",
  53889=>"111001000",
  53890=>"011000111",
  53891=>"000100000",
  53892=>"100111011",
  53893=>"000000110",
  53894=>"111111101",
  53895=>"001011000",
  53896=>"110111101",
  53897=>"011111010",
  53898=>"011011011",
  53899=>"000000111",
  53900=>"100000000",
  53901=>"111001011",
  53902=>"001000000",
  53903=>"000001000",
  53904=>"001101011",
  53905=>"101111111",
  53906=>"100000100",
  53907=>"000100100",
  53908=>"010010011",
  53909=>"101011001",
  53910=>"011011010",
  53911=>"110110100",
  53912=>"011111111",
  53913=>"111011010",
  53914=>"000011111",
  53915=>"000000000",
  53916=>"100111111",
  53917=>"010010011",
  53918=>"010000000",
  53919=>"100100111",
  53920=>"100101100",
  53921=>"111101111",
  53922=>"011100100",
  53923=>"101000111",
  53924=>"011011000",
  53925=>"111010001",
  53926=>"111001011",
  53927=>"111000000",
  53928=>"000000011",
  53929=>"000000100",
  53930=>"000000111",
  53931=>"100101011",
  53932=>"110111110",
  53933=>"100100011",
  53934=>"001000011",
  53935=>"000010011",
  53936=>"000000111",
  53937=>"000000011",
  53938=>"100111000",
  53939=>"000001001",
  53940=>"001101010",
  53941=>"010011001",
  53942=>"101110111",
  53943=>"100111111",
  53944=>"101011010",
  53945=>"000011010",
  53946=>"111010000",
  53947=>"001011011",
  53948=>"000000010",
  53949=>"011000110",
  53950=>"101001111",
  53951=>"000000000",
  53952=>"011011000",
  53953=>"111100000",
  53954=>"011000111",
  53955=>"011100000",
  53956=>"110100111",
  53957=>"110100001",
  53958=>"111000011",
  53959=>"111011100",
  53960=>"010011011",
  53961=>"001100100",
  53962=>"001011111",
  53963=>"001111101",
  53964=>"111111011",
  53965=>"001011111",
  53966=>"010011110",
  53967=>"000011111",
  53968=>"011001011",
  53969=>"000001001",
  53970=>"011111000",
  53971=>"111111111",
  53972=>"001000110",
  53973=>"111111100",
  53974=>"100100101",
  53975=>"011011011",
  53976=>"100100111",
  53977=>"100110010",
  53978=>"001000001",
  53979=>"111111111",
  53980=>"100100101",
  53981=>"110001001",
  53982=>"001100110",
  53983=>"000000011",
  53984=>"000011000",
  53985=>"000100100",
  53986=>"000100000",
  53987=>"111111100",
  53988=>"000000000",
  53989=>"011000011",
  53990=>"100000110",
  53991=>"000000100",
  53992=>"100100000",
  53993=>"000110011",
  53994=>"010011010",
  53995=>"111111100",
  53996=>"101100100",
  53997=>"111100111",
  53998=>"101000110",
  53999=>"000000000",
  54000=>"100000011",
  54001=>"101110100",
  54002=>"000100000",
  54003=>"000000101",
  54004=>"110110011",
  54005=>"001111100",
  54006=>"000001111",
  54007=>"000000100",
  54008=>"001011110",
  54009=>"111001000",
  54010=>"011111111",
  54011=>"111011010",
  54012=>"011011000",
  54013=>"100100000",
  54014=>"011110110",
  54015=>"010011101",
  54016=>"100000110",
  54017=>"111000000",
  54018=>"011010000",
  54019=>"101101001",
  54020=>"000011011",
  54021=>"111101001",
  54022=>"100000001",
  54023=>"001111011",
  54024=>"000000000",
  54025=>"000000001",
  54026=>"000111111",
  54027=>"101101111",
  54028=>"000001001",
  54029=>"001000111",
  54030=>"100111001",
  54031=>"110111111",
  54032=>"101110111",
  54033=>"110010010",
  54034=>"111110000",
  54035=>"000101010",
  54036=>"000000000",
  54037=>"111110110",
  54038=>"011011111",
  54039=>"000100111",
  54040=>"010000000",
  54041=>"111110000",
  54042=>"110000000",
  54043=>"100111011",
  54044=>"101000000",
  54045=>"001001101",
  54046=>"111111000",
  54047=>"000000001",
  54048=>"000000000",
  54049=>"111101000",
  54050=>"000000000",
  54051=>"111001001",
  54052=>"000000111",
  54053=>"001001011",
  54054=>"000000101",
  54055=>"010001000",
  54056=>"000001000",
  54057=>"000000101",
  54058=>"100110110",
  54059=>"000000000",
  54060=>"011111111",
  54061=>"111110101",
  54062=>"010011011",
  54063=>"000000000",
  54064=>"000000000",
  54065=>"110110111",
  54066=>"011000001",
  54067=>"111011010",
  54068=>"001000100",
  54069=>"000001110",
  54070=>"011001001",
  54071=>"000000000",
  54072=>"111011011",
  54073=>"101000101",
  54074=>"000000000",
  54075=>"000000000",
  54076=>"000000001",
  54077=>"110111000",
  54078=>"000000000",
  54079=>"000001001",
  54080=>"110110101",
  54081=>"110010110",
  54082=>"110111000",
  54083=>"111111000",
  54084=>"100111111",
  54085=>"000001111",
  54086=>"000101000",
  54087=>"110000110",
  54088=>"001011101",
  54089=>"111111111",
  54090=>"111001011",
  54091=>"011111111",
  54092=>"111011001",
  54093=>"101100011",
  54094=>"011111000",
  54095=>"010011111",
  54096=>"011010111",
  54097=>"111010010",
  54098=>"000001101",
  54099=>"000000101",
  54100=>"101101111",
  54101=>"001111111",
  54102=>"000011000",
  54103=>"000111111",
  54104=>"111111110",
  54105=>"100100110",
  54106=>"100101100",
  54107=>"110111111",
  54108=>"111111011",
  54109=>"000000000",
  54110=>"010110010",
  54111=>"011010010",
  54112=>"000000001",
  54113=>"010111111",
  54114=>"000000001",
  54115=>"001111001",
  54116=>"011001001",
  54117=>"001011010",
  54118=>"001001101",
  54119=>"000000001",
  54120=>"000100111",
  54121=>"000000001",
  54122=>"001101000",
  54123=>"010101110",
  54124=>"000000000",
  54125=>"110111110",
  54126=>"001000001",
  54127=>"111011000",
  54128=>"011111101",
  54129=>"000001000",
  54130=>"111000110",
  54131=>"000000010",
  54132=>"000101111",
  54133=>"100000101",
  54134=>"000111110",
  54135=>"000000001",
  54136=>"100000000",
  54137=>"010010000",
  54138=>"010000111",
  54139=>"111101101",
  54140=>"010000001",
  54141=>"000000000",
  54142=>"000000011",
  54143=>"011111111",
  54144=>"010101010",
  54145=>"111111010",
  54146=>"000000000",
  54147=>"000111101",
  54148=>"101000000",
  54149=>"001001111",
  54150=>"000000011",
  54151=>"110010001",
  54152=>"111111001",
  54153=>"000000100",
  54154=>"011111111",
  54155=>"101101111",
  54156=>"001001001",
  54157=>"111111111",
  54158=>"111111010",
  54159=>"001000101",
  54160=>"001000100",
  54161=>"101111101",
  54162=>"001100111",
  54163=>"111000101",
  54164=>"111001011",
  54165=>"010000000",
  54166=>"111111111",
  54167=>"001001111",
  54168=>"101111111",
  54169=>"000000000",
  54170=>"111111111",
  54171=>"000000000",
  54172=>"101001111",
  54173=>"111111111",
  54174=>"111111111",
  54175=>"000001111",
  54176=>"101111011",
  54177=>"111111011",
  54178=>"101000001",
  54179=>"101111100",
  54180=>"000111110",
  54181=>"001101111",
  54182=>"010101001",
  54183=>"111011110",
  54184=>"111111111",
  54185=>"111001001",
  54186=>"100001001",
  54187=>"111101001",
  54188=>"000000000",
  54189=>"111001011",
  54190=>"010111011",
  54191=>"000111111",
  54192=>"101000000",
  54193=>"011110100",
  54194=>"001000000",
  54195=>"111001001",
  54196=>"110111111",
  54197=>"000000000",
  54198=>"000000100",
  54199=>"101000000",
  54200=>"100000010",
  54201=>"011010100",
  54202=>"101001000",
  54203=>"111010000",
  54204=>"000001011",
  54205=>"111110010",
  54206=>"000000100",
  54207=>"000000001",
  54208=>"010010010",
  54209=>"000110111",
  54210=>"010111111",
  54211=>"110001000",
  54212=>"101001111",
  54213=>"110110011",
  54214=>"000101000",
  54215=>"010111011",
  54216=>"100100101",
  54217=>"100110011",
  54218=>"000000011",
  54219=>"000001111",
  54220=>"100000100",
  54221=>"010000000",
  54222=>"000000000",
  54223=>"000000101",
  54224=>"110100111",
  54225=>"110111111",
  54226=>"111010000",
  54227=>"001001000",
  54228=>"001000001",
  54229=>"000000010",
  54230=>"111111010",
  54231=>"110110110",
  54232=>"000000111",
  54233=>"000001100",
  54234=>"110011111",
  54235=>"101101111",
  54236=>"110111001",
  54237=>"110001000",
  54238=>"011100010",
  54239=>"011000010",
  54240=>"000000101",
  54241=>"101001111",
  54242=>"111111111",
  54243=>"011111111",
  54244=>"000000001",
  54245=>"001001011",
  54246=>"000000111",
  54247=>"000110110",
  54248=>"001000101",
  54249=>"011010000",
  54250=>"000101100",
  54251=>"000000111",
  54252=>"001000000",
  54253=>"001101111",
  54254=>"110110000",
  54255=>"001000001",
  54256=>"011001000",
  54257=>"011111100",
  54258=>"001001000",
  54259=>"001011111",
  54260=>"001011011",
  54261=>"010111000",
  54262=>"010000110",
  54263=>"000000111",
  54264=>"000000111",
  54265=>"101111111",
  54266=>"000010000",
  54267=>"011010010",
  54268=>"111111111",
  54269=>"111101111",
  54270=>"100100100",
  54271=>"010011000",
  54272=>"101101101",
  54273=>"000011010",
  54274=>"111001011",
  54275=>"111011010",
  54276=>"100111110",
  54277=>"011001101",
  54278=>"100100000",
  54279=>"000100100",
  54280=>"110100010",
  54281=>"000000000",
  54282=>"001101100",
  54283=>"111011001",
  54284=>"000110110",
  54285=>"110011000",
  54286=>"100100100",
  54287=>"100100000",
  54288=>"110101100",
  54289=>"100000100",
  54290=>"110000111",
  54291=>"000001001",
  54292=>"011001011",
  54293=>"111001001",
  54294=>"111001111",
  54295=>"000100100",
  54296=>"110000000",
  54297=>"011001100",
  54298=>"000001001",
  54299=>"111001000",
  54300=>"001000100",
  54301=>"000000010",
  54302=>"011011010",
  54303=>"001111100",
  54304=>"011111111",
  54305=>"000001111",
  54306=>"000001001",
  54307=>"100110110",
  54308=>"011111110",
  54309=>"011001110",
  54310=>"011011011",
  54311=>"000110110",
  54312=>"111011001",
  54313=>"011011011",
  54314=>"111110010",
  54315=>"011001000",
  54316=>"000110101",
  54317=>"100010001",
  54318=>"011011000",
  54319=>"001000101",
  54320=>"010000000",
  54321=>"111001001",
  54322=>"000011011",
  54323=>"000111110",
  54324=>"110001100",
  54325=>"100100011",
  54326=>"101001001",
  54327=>"110110000",
  54328=>"001001011",
  54329=>"000000110",
  54330=>"010001011",
  54331=>"010100000",
  54332=>"000000000",
  54333=>"111110100",
  54334=>"000001001",
  54335=>"100110001",
  54336=>"000000111",
  54337=>"011111011",
  54338=>"111011100",
  54339=>"111101100",
  54340=>"001000000",
  54341=>"011111001",
  54342=>"100110110",
  54343=>"111110111",
  54344=>"100111010",
  54345=>"110000000",
  54346=>"101001110",
  54347=>"100110100",
  54348=>"011001001",
  54349=>"000000000",
  54350=>"010010111",
  54351=>"000111101",
  54352=>"101001001",
  54353=>"110001110",
  54354=>"001100101",
  54355=>"000101000",
  54356=>"011001011",
  54357=>"111101111",
  54358=>"000000000",
  54359=>"011111110",
  54360=>"111011111",
  54361=>"001101001",
  54362=>"010100011",
  54363=>"001001000",
  54364=>"110110110",
  54365=>"001000100",
  54366=>"001001111",
  54367=>"100011001",
  54368=>"011111111",
  54369=>"111011001",
  54370=>"001001011",
  54371=>"101100000",
  54372=>"001000000",
  54373=>"101111111",
  54374=>"111011000",
  54375=>"010110010",
  54376=>"011001001",
  54377=>"000000110",
  54378=>"110000000",
  54379=>"110110111",
  54380=>"001110111",
  54381=>"000100100",
  54382=>"111001001",
  54383=>"001001000",
  54384=>"111111111",
  54385=>"010010010",
  54386=>"101001011",
  54387=>"100111100",
  54388=>"110100000",
  54389=>"110010000",
  54390=>"000011001",
  54391=>"011001011",
  54392=>"011010011",
  54393=>"101000100",
  54394=>"001000001",
  54395=>"000000101",
  54396=>"000001110",
  54397=>"010000000",
  54398=>"110001001",
  54399=>"101110100",
  54400=>"011100000",
  54401=>"111000011",
  54402=>"111101110",
  54403=>"011111000",
  54404=>"000001111",
  54405=>"011011001",
  54406=>"011011010",
  54407=>"000100110",
  54408=>"000100100",
  54409=>"110100110",
  54410=>"011000001",
  54411=>"001110100",
  54412=>"111001000",
  54413=>"100000000",
  54414=>"000110100",
  54415=>"000000100",
  54416=>"011111001",
  54417=>"111011010",
  54418=>"010010111",
  54419=>"110001110",
  54420=>"010000010",
  54421=>"111001111",
  54422=>"000000101",
  54423=>"000000000",
  54424=>"110011100",
  54425=>"011011011",
  54426=>"001001001",
  54427=>"010001011",
  54428=>"111010000",
  54429=>"110101100",
  54430=>"111000000",
  54431=>"011100000",
  54432=>"001111111",
  54433=>"111110011",
  54434=>"001111110",
  54435=>"110000001",
  54436=>"011011111",
  54437=>"000100000",
  54438=>"000111000",
  54439=>"000101111",
  54440=>"111000000",
  54441=>"110010001",
  54442=>"001001011",
  54443=>"111011011",
  54444=>"000111111",
  54445=>"100100100",
  54446=>"001001111",
  54447=>"011110000",
  54448=>"110000001",
  54449=>"011111010",
  54450=>"000011000",
  54451=>"000011100",
  54452=>"111111111",
  54453=>"110101111",
  54454=>"011011001",
  54455=>"011011110",
  54456=>"000111111",
  54457=>"000000000",
  54458=>"111010000",
  54459=>"111111000",
  54460=>"000111110",
  54461=>"111001000",
  54462=>"011111111",
  54463=>"100000000",
  54464=>"111000000",
  54465=>"000000100",
  54466=>"010011000",
  54467=>"000000100",
  54468=>"000110100",
  54469=>"100001010",
  54470=>"000100110",
  54471=>"110000010",
  54472=>"000110111",
  54473=>"011010000",
  54474=>"110111111",
  54475=>"011001011",
  54476=>"111111000",
  54477=>"100100101",
  54478=>"100000001",
  54479=>"000000111",
  54480=>"101001000",
  54481=>"110111111",
  54482=>"100000100",
  54483=>"101111111",
  54484=>"110000100",
  54485=>"001001001",
  54486=>"011000100",
  54487=>"110000000",
  54488=>"100110100",
  54489=>"010010010",
  54490=>"000000001",
  54491=>"101101110",
  54492=>"111011111",
  54493=>"001011001",
  54494=>"001010110",
  54495=>"011011110",
  54496=>"011010101",
  54497=>"001000000",
  54498=>"111000000",
  54499=>"001111011",
  54500=>"110000100",
  54501=>"000100100",
  54502=>"110111100",
  54503=>"110110110",
  54504=>"001001001",
  54505=>"011001001",
  54506=>"010000010",
  54507=>"111111001",
  54508=>"110000000",
  54509=>"110000000",
  54510=>"100000100",
  54511=>"100110100",
  54512=>"100000001",
  54513=>"000101101",
  54514=>"111011000",
  54515=>"100000000",
  54516=>"101100000",
  54517=>"001011111",
  54518=>"000110110",
  54519=>"000001001",
  54520=>"111011001",
  54521=>"100011000",
  54522=>"111001111",
  54523=>"000010101",
  54524=>"001001111",
  54525=>"000100100",
  54526=>"000110100",
  54527=>"110110110",
  54528=>"111000000",
  54529=>"000101101",
  54530=>"000110111",
  54531=>"010100111",
  54532=>"111111111",
  54533=>"111111101",
  54534=>"111111000",
  54535=>"000000110",
  54536=>"111110000",
  54537=>"000000111",
  54538=>"000000100",
  54539=>"111111000",
  54540=>"000111111",
  54541=>"111111111",
  54542=>"100000010",
  54543=>"101110011",
  54544=>"111101111",
  54545=>"001000101",
  54546=>"100101001",
  54547=>"101000011",
  54548=>"011111000",
  54549=>"010010001",
  54550=>"111001100",
  54551=>"001000011",
  54552=>"001000000",
  54553=>"101111111",
  54554=>"101010010",
  54555=>"010101100",
  54556=>"101101000",
  54557=>"000010100",
  54558=>"101111000",
  54559=>"100100010",
  54560=>"111101111",
  54561=>"011111001",
  54562=>"000000010",
  54563=>"000010111",
  54564=>"000000011",
  54565=>"011111001",
  54566=>"000100111",
  54567=>"011111011",
  54568=>"010010001",
  54569=>"110100111",
  54570=>"111000100",
  54571=>"000100100",
  54572=>"000000000",
  54573=>"010100110",
  54574=>"101000100",
  54575=>"110001001",
  54576=>"000000101",
  54577=>"011101111",
  54578=>"011001000",
  54579=>"111010000",
  54580=>"111100000",
  54581=>"110111110",
  54582=>"101000100",
  54583=>"111010001",
  54584=>"111000010",
  54585=>"000010010",
  54586=>"000000000",
  54587=>"000000000",
  54588=>"001001010",
  54589=>"111111000",
  54590=>"100000000",
  54591=>"111111001",
  54592=>"100100110",
  54593=>"101101111",
  54594=>"001101111",
  54595=>"110110111",
  54596=>"101111001",
  54597=>"000100000",
  54598=>"101001110",
  54599=>"011000010",
  54600=>"101001001",
  54601=>"011111101",
  54602=>"000000000",
  54603=>"111101101",
  54604=>"000010111",
  54605=>"000001111",
  54606=>"010101111",
  54607=>"000000110",
  54608=>"101000001",
  54609=>"011000000",
  54610=>"111111101",
  54611=>"110100101",
  54612=>"111000000",
  54613=>"111011101",
  54614=>"001000001",
  54615=>"000000000",
  54616=>"111110101",
  54617=>"010001111",
  54618=>"000010110",
  54619=>"100100110",
  54620=>"111111111",
  54621=>"001001001",
  54622=>"110011110",
  54623=>"011011001",
  54624=>"010011111",
  54625=>"111011000",
  54626=>"000011111",
  54627=>"001000001",
  54628=>"100100110",
  54629=>"100101111",
  54630=>"010010000",
  54631=>"010010111",
  54632=>"111000000",
  54633=>"111000000",
  54634=>"010000111",
  54635=>"110111010",
  54636=>"111011110",
  54637=>"000000101",
  54638=>"000000111",
  54639=>"001001000",
  54640=>"110101100",
  54641=>"111000000",
  54642=>"101000001",
  54643=>"010111100",
  54644=>"001000000",
  54645=>"000000000",
  54646=>"000000000",
  54647=>"101110111",
  54648=>"001010000",
  54649=>"101101110",
  54650=>"010101111",
  54651=>"010101001",
  54652=>"001101010",
  54653=>"001000100",
  54654=>"011010001",
  54655=>"111111000",
  54656=>"000010110",
  54657=>"101100100",
  54658=>"110111001",
  54659=>"100111111",
  54660=>"010000000",
  54661=>"110101111",
  54662=>"100110110",
  54663=>"000000011",
  54664=>"001111001",
  54665=>"001001000",
  54666=>"111100110",
  54667=>"000001000",
  54668=>"011010011",
  54669=>"100000011",
  54670=>"000111011",
  54671=>"000000000",
  54672=>"111100110",
  54673=>"111101001",
  54674=>"000110000",
  54675=>"111101000",
  54676=>"111001000",
  54677=>"111000000",
  54678=>"111011110",
  54679=>"000011000",
  54680=>"001000010",
  54681=>"100000001",
  54682=>"110010111",
  54683=>"111111000",
  54684=>"000001101",
  54685=>"000000011",
  54686=>"010000111",
  54687=>"001000100",
  54688=>"011110111",
  54689=>"001110001",
  54690=>"011011010",
  54691=>"111000000",
  54692=>"111010000",
  54693=>"000001111",
  54694=>"000110011",
  54695=>"001011000",
  54696=>"111011010",
  54697=>"000111100",
  54698=>"011000111",
  54699=>"111000000",
  54700=>"111010011",
  54701=>"100000000",
  54702=>"001001100",
  54703=>"010111111",
  54704=>"011111101",
  54705=>"011100101",
  54706=>"001001001",
  54707=>"000100100",
  54708=>"001100110",
  54709=>"000011111",
  54710=>"000010111",
  54711=>"000111111",
  54712=>"110000100",
  54713=>"011100100",
  54714=>"111111001",
  54715=>"011000000",
  54716=>"000010100",
  54717=>"111111111",
  54718=>"001011000",
  54719=>"011000000",
  54720=>"001001011",
  54721=>"110000000",
  54722=>"101000111",
  54723=>"111100100",
  54724=>"000110010",
  54725=>"110100001",
  54726=>"110101101",
  54727=>"000010000",
  54728=>"010000111",
  54729=>"000000010",
  54730=>"101111111",
  54731=>"101101111",
  54732=>"011011011",
  54733=>"110001000",
  54734=>"101000000",
  54735=>"111111011",
  54736=>"100111000",
  54737=>"110111010",
  54738=>"010011110",
  54739=>"101101101",
  54740=>"010101101",
  54741=>"100100100",
  54742=>"101001000",
  54743=>"011001001",
  54744=>"000000000",
  54745=>"000111010",
  54746=>"000101111",
  54747=>"000000100",
  54748=>"111001100",
  54749=>"111010010",
  54750=>"000011000",
  54751=>"110011001",
  54752=>"000000000",
  54753=>"111000000",
  54754=>"000011111",
  54755=>"011001101",
  54756=>"001001001",
  54757=>"111001011",
  54758=>"111111010",
  54759=>"110000011",
  54760=>"011101001",
  54761=>"111011000",
  54762=>"000001001",
  54763=>"010000000",
  54764=>"000000000",
  54765=>"000010111",
  54766=>"000000000",
  54767=>"000100001",
  54768=>"111011000",
  54769=>"011001100",
  54770=>"000000000",
  54771=>"110101101",
  54772=>"011000101",
  54773=>"000000011",
  54774=>"000000000",
  54775=>"101000001",
  54776=>"000000000",
  54777=>"001000000",
  54778=>"001100101",
  54779=>"000101111",
  54780=>"110001011",
  54781=>"000000000",
  54782=>"110111111",
  54783=>"000000000",
  54784=>"000101111",
  54785=>"111111100",
  54786=>"110000110",
  54787=>"111001000",
  54788=>"000110011",
  54789=>"011001001",
  54790=>"011101101",
  54791=>"000000000",
  54792=>"100001011",
  54793=>"000000100",
  54794=>"111000100",
  54795=>"000000000",
  54796=>"000001001",
  54797=>"110110110",
  54798=>"111000000",
  54799=>"111011111",
  54800=>"111000010",
  54801=>"111001010",
  54802=>"001001000",
  54803=>"111111000",
  54804=>"101000010",
  54805=>"111110100",
  54806=>"001111110",
  54807=>"111011111",
  54808=>"101000110",
  54809=>"100111001",
  54810=>"101100101",
  54811=>"000111011",
  54812=>"110110111",
  54813=>"110110000",
  54814=>"000000011",
  54815=>"111101111",
  54816=>"000000110",
  54817=>"000100011",
  54818=>"101111110",
  54819=>"101111101",
  54820=>"101101100",
  54821=>"011111100",
  54822=>"011011110",
  54823=>"000000000",
  54824=>"111110111",
  54825=>"000110110",
  54826=>"111000101",
  54827=>"101111001",
  54828=>"010000000",
  54829=>"000000000",
  54830=>"100001001",
  54831=>"110011011",
  54832=>"111100000",
  54833=>"000001001",
  54834=>"111011010",
  54835=>"110110000",
  54836=>"010111111",
  54837=>"000010001",
  54838=>"010110101",
  54839=>"000101111",
  54840=>"000000000",
  54841=>"001001100",
  54842=>"111001000",
  54843=>"101110000",
  54844=>"100110000",
  54845=>"101111111",
  54846=>"001001100",
  54847=>"100010001",
  54848=>"111011111",
  54849=>"111111000",
  54850=>"000000000",
  54851=>"010110111",
  54852=>"101000000",
  54853=>"111101001",
  54854=>"010001101",
  54855=>"110110011",
  54856=>"000000000",
  54857=>"001111011",
  54858=>"001100100",
  54859=>"111001111",
  54860=>"100000000",
  54861=>"011010011",
  54862=>"101001110",
  54863=>"110010000",
  54864=>"101110111",
  54865=>"110111111",
  54866=>"110101000",
  54867=>"111011000",
  54868=>"000110010",
  54869=>"010000100",
  54870=>"111110111",
  54871=>"000100110",
  54872=>"110101111",
  54873=>"111001000",
  54874=>"000001001",
  54875=>"010000000",
  54876=>"111001000",
  54877=>"111000100",
  54878=>"111110010",
  54879=>"000111111",
  54880=>"111111111",
  54881=>"001000001",
  54882=>"111000000",
  54883=>"001111110",
  54884=>"000000010",
  54885=>"001110010",
  54886=>"110100010",
  54887=>"100110110",
  54888=>"001111110",
  54889=>"111101000",
  54890=>"000000000",
  54891=>"111110010",
  54892=>"111000000",
  54893=>"011000001",
  54894=>"000001101",
  54895=>"101111001",
  54896=>"111010100",
  54897=>"000000000",
  54898=>"010011111",
  54899=>"001001000",
  54900=>"111001101",
  54901=>"111001101",
  54902=>"000100000",
  54903=>"010010010",
  54904=>"110110100",
  54905=>"000111000",
  54906=>"101000011",
  54907=>"111001101",
  54908=>"001000000",
  54909=>"101111001",
  54910=>"111010110",
  54911=>"111000111",
  54912=>"100110111",
  54913=>"111100110",
  54914=>"111111111",
  54915=>"101000010",
  54916=>"111101000",
  54917=>"111000001",
  54918=>"110111001",
  54919=>"000000010",
  54920=>"011011011",
  54921=>"111000110",
  54922=>"111100111",
  54923=>"101110000",
  54924=>"000110111",
  54925=>"000000111",
  54926=>"111001000",
  54927=>"110001001",
  54928=>"001101101",
  54929=>"000101110",
  54930=>"111101101",
  54931=>"010110010",
  54932=>"000000100",
  54933=>"001000000",
  54934=>"111111000",
  54935=>"110001000",
  54936=>"010000000",
  54937=>"111011000",
  54938=>"111010000",
  54939=>"000000000",
  54940=>"000001001",
  54941=>"000000000",
  54942=>"000000110",
  54943=>"111100000",
  54944=>"000000011",
  54945=>"000111111",
  54946=>"111001010",
  54947=>"001000000",
  54948=>"000000111",
  54949=>"001000110",
  54950=>"111111010",
  54951=>"000000000",
  54952=>"101101010",
  54953=>"000101101",
  54954=>"101000111",
  54955=>"111011011",
  54956=>"110111111",
  54957=>"110000000",
  54958=>"010111110",
  54959=>"111001001",
  54960=>"001000111",
  54961=>"111101100",
  54962=>"111000001",
  54963=>"001001001",
  54964=>"111000110",
  54965=>"010111110",
  54966=>"001111111",
  54967=>"000011000",
  54968=>"001011001",
  54969=>"001000000",
  54970=>"010111111",
  54971=>"110101110",
  54972=>"111110001",
  54973=>"111001001",
  54974=>"011000100",
  54975=>"000101011",
  54976=>"000110111",
  54977=>"101000001",
  54978=>"110111111",
  54979=>"101111101",
  54980=>"010000001",
  54981=>"000000110",
  54982=>"000000100",
  54983=>"000110101",
  54984=>"110000000",
  54985=>"001111111",
  54986=>"111101111",
  54987=>"111000010",
  54988=>"000000010",
  54989=>"000000010",
  54990=>"000101011",
  54991=>"111001101",
  54992=>"111111110",
  54993=>"011001111",
  54994=>"111001000",
  54995=>"111111111",
  54996=>"111111100",
  54997=>"001011111",
  54998=>"000001011",
  54999=>"001001010",
  55000=>"010011000",
  55001=>"111000001",
  55002=>"001011101",
  55003=>"111000000",
  55004=>"100111110",
  55005=>"101101001",
  55006=>"010100101",
  55007=>"000110000",
  55008=>"000000000",
  55009=>"000000010",
  55010=>"010110111",
  55011=>"111000001",
  55012=>"000010110",
  55013=>"111001111",
  55014=>"001000001",
  55015=>"000111111",
  55016=>"110101101",
  55017=>"111111111",
  55018=>"110000001",
  55019=>"000101001",
  55020=>"101000000",
  55021=>"000010000",
  55022=>"111000001",
  55023=>"110000011",
  55024=>"010111010",
  55025=>"000000001",
  55026=>"000000000",
  55027=>"111100001",
  55028=>"000001001",
  55029=>"101000110",
  55030=>"000000001",
  55031=>"010010000",
  55032=>"000000000",
  55033=>"001101110",
  55034=>"111110111",
  55035=>"000000001",
  55036=>"000111101",
  55037=>"011100001",
  55038=>"000100000",
  55039=>"110000000",
  55040=>"110100110",
  55041=>"110110110",
  55042=>"001001011",
  55043=>"110100000",
  55044=>"010110110",
  55045=>"100110100",
  55046=>"001001011",
  55047=>"000001010",
  55048=>"100100110",
  55049=>"001001000",
  55050=>"001001111",
  55051=>"000000000",
  55052=>"110011011",
  55053=>"100001000",
  55054=>"111001001",
  55055=>"001010001",
  55056=>"000110100",
  55057=>"000001100",
  55058=>"000000011",
  55059=>"111000000",
  55060=>"000001011",
  55061=>"001011110",
  55062=>"100100110",
  55063=>"100000000",
  55064=>"011011111",
  55065=>"100000100",
  55066=>"100110100",
  55067=>"011011111",
  55068=>"000011110",
  55069=>"010010011",
  55070=>"011011111",
  55071=>"011000111",
  55072=>"111000100",
  55073=>"100100101",
  55074=>"110011011",
  55075=>"110110000",
  55076=>"111111101",
  55077=>"001001011",
  55078=>"110110000",
  55079=>"011011001",
  55080=>"100100000",
  55081=>"000100100",
  55082=>"011000000",
  55083=>"100110100",
  55084=>"110111101",
  55085=>"001011111",
  55086=>"100100111",
  55087=>"110011110",
  55088=>"000110110",
  55089=>"101100001",
  55090=>"001111110",
  55091=>"011011001",
  55092=>"011001011",
  55093=>"101010000",
  55094=>"001101110",
  55095=>"011101000",
  55096=>"011001001",
  55097=>"011001011",
  55098=>"000001100",
  55099=>"000011000",
  55100=>"001011111",
  55101=>"101101000",
  55102=>"100001001",
  55103=>"100100110",
  55104=>"000000111",
  55105=>"000111001",
  55106=>"111111000",
  55107=>"000110010",
  55108=>"100100100",
  55109=>"111011010",
  55110=>"011011001",
  55111=>"100101001",
  55112=>"110010111",
  55113=>"101001001",
  55114=>"001011111",
  55115=>"011011111",
  55116=>"110000100",
  55117=>"100000010",
  55118=>"110010001",
  55119=>"011011101",
  55120=>"100100001",
  55121=>"100110110",
  55122=>"100001001",
  55123=>"010000000",
  55124=>"001001001",
  55125=>"001011101",
  55126=>"111111101",
  55127=>"000001111",
  55128=>"011001001",
  55129=>"011001001",
  55130=>"011011111",
  55131=>"110101010",
  55132=>"100100000",
  55133=>"000110100",
  55134=>"101111111",
  55135=>"000100000",
  55136=>"100100100",
  55137=>"100100110",
  55138=>"000001011",
  55139=>"011011110",
  55140=>"011001011",
  55141=>"001001001",
  55142=>"011011011",
  55143=>"101101001",
  55144=>"100101100",
  55145=>"110011111",
  55146=>"100111100",
  55147=>"100111010",
  55148=>"100100010",
  55149=>"001100111",
  55150=>"000001100",
  55151=>"000011111",
  55152=>"110010011",
  55153=>"010000101",
  55154=>"110011001",
  55155=>"110110110",
  55156=>"111111100",
  55157=>"011011110",
  55158=>"111010101",
  55159=>"100101011",
  55160=>"000000100",
  55161=>"111110111",
  55162=>"000001000",
  55163=>"110101100",
  55164=>"001001011",
  55165=>"100000000",
  55166=>"111101101",
  55167=>"000011111",
  55168=>"110110110",
  55169=>"000000100",
  55170=>"100000111",
  55171=>"110010001",
  55172=>"000011111",
  55173=>"000000000",
  55174=>"100110111",
  55175=>"000000000",
  55176=>"000000000",
  55177=>"011011111",
  55178=>"000000001",
  55179=>"110000000",
  55180=>"000100100",
  55181=>"011000111",
  55182=>"001011011",
  55183=>"011001000",
  55184=>"011001010",
  55185=>"111011110",
  55186=>"001001100",
  55187=>"010011011",
  55188=>"000010000",
  55189=>"011111111",
  55190=>"001001101",
  55191=>"110110100",
  55192=>"110001011",
  55193=>"000100110",
  55194=>"011011000",
  55195=>"000100100",
  55196=>"011000000",
  55197=>"011011110",
  55198=>"101000101",
  55199=>"011001011",
  55200=>"110110001",
  55201=>"000101100",
  55202=>"100011001",
  55203=>"011010100",
  55204=>"100011100",
  55205=>"100000000",
  55206=>"110100000",
  55207=>"111100000",
  55208=>"000010111",
  55209=>"010100000",
  55210=>"011001110",
  55211=>"001101011",
  55212=>"100100000",
  55213=>"100100111",
  55214=>"001011111",
  55215=>"101100001",
  55216=>"010110001",
  55217=>"111110111",
  55218=>"000011110",
  55219=>"001001111",
  55220=>"111111100",
  55221=>"111011000",
  55222=>"100111000",
  55223=>"110001011",
  55224=>"110100100",
  55225=>"100010000",
  55226=>"100000000",
  55227=>"111000001",
  55228=>"100000000",
  55229=>"100100110",
  55230=>"100100000",
  55231=>"111111110",
  55232=>"001001111",
  55233=>"001000001",
  55234=>"001111100",
  55235=>"010000000",
  55236=>"001010010",
  55237=>"111111111",
  55238=>"111000000",
  55239=>"000100111",
  55240=>"110000001",
  55241=>"111110000",
  55242=>"100010110",
  55243=>"011011110",
  55244=>"001001011",
  55245=>"101000001",
  55246=>"001001001",
  55247=>"100100000",
  55248=>"011001001",
  55249=>"000100000",
  55250=>"100010001",
  55251=>"100110110",
  55252=>"011000111",
  55253=>"001000100",
  55254=>"111000011",
  55255=>"000111101",
  55256=>"011001011",
  55257=>"110010100",
  55258=>"000000001",
  55259=>"001001010",
  55260=>"001010111",
  55261=>"100110100",
  55262=>"110110100",
  55263=>"001001011",
  55264=>"100100101",
  55265=>"011011011",
  55266=>"000000011",
  55267=>"111110100",
  55268=>"000000000",
  55269=>"110110110",
  55270=>"100100100",
  55271=>"100011111",
  55272=>"100100110",
  55273=>"111010110",
  55274=>"001001011",
  55275=>"100010011",
  55276=>"110110100",
  55277=>"100100000",
  55278=>"000010100",
  55279=>"110110010",
  55280=>"110110100",
  55281=>"010010000",
  55282=>"101011010",
  55283=>"100100010",
  55284=>"110001001",
  55285=>"011001001",
  55286=>"010000100",
  55287=>"000100010",
  55288=>"001001111",
  55289=>"010011100",
  55290=>"100000010",
  55291=>"011110010",
  55292=>"001001011",
  55293=>"100110000",
  55294=>"011111011",
  55295=>"001001011",
  55296=>"011011000",
  55297=>"111111111",
  55298=>"101000101",
  55299=>"101100111",
  55300=>"111111100",
  55301=>"011101011",
  55302=>"111100111",
  55303=>"100000000",
  55304=>"000110110",
  55305=>"001000101",
  55306=>"111000111",
  55307=>"110101111",
  55308=>"000111011",
  55309=>"011111000",
  55310=>"110001011",
  55311=>"000000000",
  55312=>"010011111",
  55313=>"001000101",
  55314=>"100101101",
  55315=>"001111111",
  55316=>"111001111",
  55317=>"000110000",
  55318=>"000000001",
  55319=>"111000000",
  55320=>"110100100",
  55321=>"000111110",
  55322=>"011100010",
  55323=>"000001011",
  55324=>"000000000",
  55325=>"110110010",
  55326=>"110011111",
  55327=>"000110000",
  55328=>"001000001",
  55329=>"111111111",
  55330=>"100100111",
  55331=>"111110000",
  55332=>"110101100",
  55333=>"110100000",
  55334=>"110111011",
  55335=>"111010101",
  55336=>"111011000",
  55337=>"000000000",
  55338=>"111100100",
  55339=>"000001110",
  55340=>"000000100",
  55341=>"111111111",
  55342=>"111001101",
  55343=>"000111011",
  55344=>"111100000",
  55345=>"111111101",
  55346=>"011111111",
  55347=>"111101101",
  55348=>"011101011",
  55349=>"110111111",
  55350=>"101101110",
  55351=>"010111000",
  55352=>"111000000",
  55353=>"000110000",
  55354=>"000100100",
  55355=>"000000001",
  55356=>"110100000",
  55357=>"111111000",
  55358=>"000000101",
  55359=>"111110000",
  55360=>"001000010",
  55361=>"111111010",
  55362=>"110111011",
  55363=>"010101000",
  55364=>"011001000",
  55365=>"000000000",
  55366=>"000110110",
  55367=>"100000000",
  55368=>"111111111",
  55369=>"111001011",
  55370=>"001000001",
  55371=>"111000000",
  55372=>"111100100",
  55373=>"111101101",
  55374=>"011111001",
  55375=>"000000000",
  55376=>"100101111",
  55377=>"110111010",
  55378=>"000000000",
  55379=>"011001000",
  55380=>"111000000",
  55381=>"111110101",
  55382=>"111100111",
  55383=>"011111000",
  55384=>"111101001",
  55385=>"010000100",
  55386=>"011100000",
  55387=>"010000111",
  55388=>"000000000",
  55389=>"011001011",
  55390=>"011000001",
  55391=>"110001011",
  55392=>"000101000",
  55393=>"111111011",
  55394=>"001000000",
  55395=>"110111100",
  55396=>"100100000",
  55397=>"010011001",
  55398=>"110110000",
  55399=>"110110110",
  55400=>"111000101",
  55401=>"111110111",
  55402=>"010101100",
  55403=>"000110000",
  55404=>"111001001",
  55405=>"000000100",
  55406=>"011011011",
  55407=>"000000111",
  55408=>"011111111",
  55409=>"010000000",
  55410=>"011001001",
  55411=>"010110000",
  55412=>"111000000",
  55413=>"000001000",
  55414=>"000110111",
  55415=>"000001111",
  55416=>"000000000",
  55417=>"000000000",
  55418=>"000010111",
  55419=>"000101100",
  55420=>"110100110",
  55421=>"100100100",
  55422=>"111110001",
  55423=>"101101101",
  55424=>"111000000",
  55425=>"111000110",
  55426=>"000111011",
  55427=>"000000010",
  55428=>"110110101",
  55429=>"111100001",
  55430=>"111011001",
  55431=>"001011000",
  55432=>"111111111",
  55433=>"111001011",
  55434=>"010000000",
  55435=>"110110000",
  55436=>"111111010",
  55437=>"011000001",
  55438=>"111111111",
  55439=>"000000000",
  55440=>"111100110",
  55441=>"011111000",
  55442=>"101110000",
  55443=>"111110111",
  55444=>"001111111",
  55445=>"000000100",
  55446=>"110111111",
  55447=>"000011000",
  55448=>"010010011",
  55449=>"000110100",
  55450=>"101111111",
  55451=>"000000001",
  55452=>"000000010",
  55453=>"100001101",
  55454=>"101101111",
  55455=>"000000000",
  55456=>"111110110",
  55457=>"000000000",
  55458=>"111010010",
  55459=>"010111101",
  55460=>"110010110",
  55461=>"110110010",
  55462=>"000000111",
  55463=>"000111000",
  55464=>"110000111",
  55465=>"001111101",
  55466=>"101001001",
  55467=>"000000001",
  55468=>"000000010",
  55469=>"011010111",
  55470=>"010000000",
  55471=>"000001110",
  55472=>"101111001",
  55473=>"111111101",
  55474=>"001000100",
  55475=>"100100111",
  55476=>"000011000",
  55477=>"100000101",
  55478=>"000000001",
  55479=>"000000000",
  55480=>"011011000",
  55481=>"000111111",
  55482=>"000101000",
  55483=>"111101111",
  55484=>"111010010",
  55485=>"111001000",
  55486=>"001111111",
  55487=>"010111111",
  55488=>"000010000",
  55489=>"111111010",
  55490=>"111111101",
  55491=>"110001110",
  55492=>"000111000",
  55493=>"110110111",
  55494=>"111101000",
  55495=>"000000000",
  55496=>"000111111",
  55497=>"000000000",
  55498=>"110111101",
  55499=>"110001101",
  55500=>"010000001",
  55501=>"001010111",
  55502=>"000000110",
  55503=>"000001010",
  55504=>"000010000",
  55505=>"000101000",
  55506=>"001110010",
  55507=>"110101000",
  55508=>"101000111",
  55509=>"110111110",
  55510=>"111111010",
  55511=>"111000000",
  55512=>"000000000",
  55513=>"000001101",
  55514=>"000110011",
  55515=>"111100110",
  55516=>"010000100",
  55517=>"101010110",
  55518=>"000001111",
  55519=>"100110100",
  55520=>"111010010",
  55521=>"001000100",
  55522=>"111110000",
  55523=>"011101000",
  55524=>"000000100",
  55525=>"010111111",
  55526=>"000000001",
  55527=>"100100011",
  55528=>"110001000",
  55529=>"100010110",
  55530=>"111101010",
  55531=>"000000000",
  55532=>"111111011",
  55533=>"110111111",
  55534=>"001000000",
  55535=>"111001010",
  55536=>"111111010",
  55537=>"100010010",
  55538=>"000000111",
  55539=>"000100110",
  55540=>"100101010",
  55541=>"111000111",
  55542=>"000000001",
  55543=>"000000100",
  55544=>"001000010",
  55545=>"111111000",
  55546=>"111001000",
  55547=>"100110111",
  55548=>"000000011",
  55549=>"000000000",
  55550=>"011111011",
  55551=>"010101001",
  55552=>"101111100",
  55553=>"000000111",
  55554=>"000100000",
  55555=>"001001011",
  55556=>"101110110",
  55557=>"101011001",
  55558=>"111111111",
  55559=>"000000011",
  55560=>"100110000",
  55561=>"001000011",
  55562=>"000000100",
  55563=>"000000000",
  55564=>"101111111",
  55565=>"000001000",
  55566=>"100100000",
  55567=>"111011101",
  55568=>"001000010",
  55569=>"000000110",
  55570=>"000000110",
  55571=>"000000111",
  55572=>"111111101",
  55573=>"010110111",
  55574=>"011111000",
  55575=>"010000000",
  55576=>"101000111",
  55577=>"111101101",
  55578=>"101001111",
  55579=>"011000000",
  55580=>"110001111",
  55581=>"111110111",
  55582=>"100100011",
  55583=>"110001101",
  55584=>"100000000",
  55585=>"001001111",
  55586=>"000111111",
  55587=>"111111110",
  55588=>"110000110",
  55589=>"001111011",
  55590=>"001000111",
  55591=>"111000000",
  55592=>"110111101",
  55593=>"001111111",
  55594=>"000101000",
  55595=>"111001000",
  55596=>"100110111",
  55597=>"101000110",
  55598=>"000000111",
  55599=>"110111101",
  55600=>"000100001",
  55601=>"111100010",
  55602=>"000111011",
  55603=>"100011001",
  55604=>"000100000",
  55605=>"110000010",
  55606=>"100110100",
  55607=>"100111111",
  55608=>"101001101",
  55609=>"100000000",
  55610=>"101001000",
  55611=>"111111100",
  55612=>"110100111",
  55613=>"010111010",
  55614=>"000000011",
  55615=>"001100110",
  55616=>"111100010",
  55617=>"001100111",
  55618=>"000100111",
  55619=>"100000000",
  55620=>"000001001",
  55621=>"000101000",
  55622=>"111110000",
  55623=>"101000000",
  55624=>"011100111",
  55625=>"000000010",
  55626=>"000000000",
  55627=>"000001111",
  55628=>"000000100",
  55629=>"000100011",
  55630=>"110111110",
  55631=>"000000011",
  55632=>"000011111",
  55633=>"111010000",
  55634=>"101100000",
  55635=>"000010000",
  55636=>"000001000",
  55637=>"011011111",
  55638=>"011110110",
  55639=>"001000000",
  55640=>"000110111",
  55641=>"001011010",
  55642=>"000001011",
  55643=>"000000011",
  55644=>"100101101",
  55645=>"001100000",
  55646=>"111111000",
  55647=>"001000100",
  55648=>"000101101",
  55649=>"000000111",
  55650=>"000000101",
  55651=>"000110110",
  55652=>"100001001",
  55653=>"010101101",
  55654=>"101111010",
  55655=>"011111111",
  55656=>"000000001",
  55657=>"101000000",
  55658=>"111000000",
  55659=>"000000001",
  55660=>"100101101",
  55661=>"000000100",
  55662=>"100000000",
  55663=>"011011111",
  55664=>"100001101",
  55665=>"001101101",
  55666=>"000001001",
  55667=>"001000100",
  55668=>"100110111",
  55669=>"000000001",
  55670=>"000100111",
  55671=>"011111010",
  55672=>"010101100",
  55673=>"101111010",
  55674=>"000100111",
  55675=>"111010010",
  55676=>"100001101",
  55677=>"001001010",
  55678=>"011010010",
  55679=>"000000000",
  55680=>"101000100",
  55681=>"000000011",
  55682=>"110110000",
  55683=>"111010110",
  55684=>"010010010",
  55685=>"110000111",
  55686=>"000001100",
  55687=>"001100101",
  55688=>"001001101",
  55689=>"111110101",
  55690=>"100100100",
  55691=>"111100010",
  55692=>"111001000",
  55693=>"010011111",
  55694=>"000000001",
  55695=>"000000110",
  55696=>"100111011",
  55697=>"000000110",
  55698=>"100101001",
  55699=>"000000010",
  55700=>"000000100",
  55701=>"100000000",
  55702=>"101101000",
  55703=>"000110110",
  55704=>"101110000",
  55705=>"111111011",
  55706=>"011100000",
  55707=>"010000000",
  55708=>"100111111",
  55709=>"100000111",
  55710=>"100001111",
  55711=>"000001111",
  55712=>"111100101",
  55713=>"000000001",
  55714=>"111101000",
  55715=>"100101111",
  55716=>"111100100",
  55717=>"100100111",
  55718=>"000111001",
  55719=>"110001011",
  55720=>"111000000",
  55721=>"000001100",
  55722=>"100100000",
  55723=>"000100111",
  55724=>"010010011",
  55725=>"000000101",
  55726=>"000110110",
  55727=>"111111111",
  55728=>"111000100",
  55729=>"000101110",
  55730=>"001011000",
  55731=>"000101000",
  55732=>"011011111",
  55733=>"111011000",
  55734=>"011111111",
  55735=>"101101101",
  55736=>"011000111",
  55737=>"010000011",
  55738=>"010011001",
  55739=>"100101101",
  55740=>"101111101",
  55741=>"000101111",
  55742=>"111001010",
  55743=>"000000000",
  55744=>"100010110",
  55745=>"000000010",
  55746=>"000111011",
  55747=>"101110110",
  55748=>"010100001",
  55749=>"110011011",
  55750=>"000011000",
  55751=>"101100000",
  55752=>"111101001",
  55753=>"010111000",
  55754=>"111111010",
  55755=>"000100100",
  55756=>"000010001",
  55757=>"000000110",
  55758=>"000111010",
  55759=>"000111100",
  55760=>"000010110",
  55761=>"111011111",
  55762=>"000110111",
  55763=>"111011010",
  55764=>"010000100",
  55765=>"000111100",
  55766=>"001001000",
  55767=>"111001111",
  55768=>"111010000",
  55769=>"000110001",
  55770=>"101111100",
  55771=>"100000111",
  55772=>"110011110",
  55773=>"001011011",
  55774=>"001111110",
  55775=>"000111001",
  55776=>"010010000",
  55777=>"100101011",
  55778=>"111011000",
  55779=>"001100101",
  55780=>"000100000",
  55781=>"111111111",
  55782=>"111100110",
  55783=>"000011011",
  55784=>"111101101",
  55785=>"111110111",
  55786=>"000001001",
  55787=>"101111101",
  55788=>"010000000",
  55789=>"000000000",
  55790=>"111001000",
  55791=>"111101011",
  55792=>"111111110",
  55793=>"011110110",
  55794=>"000100000",
  55795=>"110110000",
  55796=>"000010011",
  55797=>"101000110",
  55798=>"000000111",
  55799=>"000010010",
  55800=>"001000000",
  55801=>"101000010",
  55802=>"111111011",
  55803=>"010011101",
  55804=>"111101000",
  55805=>"011011111",
  55806=>"111111110",
  55807=>"000000010",
  55808=>"010111111",
  55809=>"110000000",
  55810=>"111010000",
  55811=>"000000001",
  55812=>"010110101",
  55813=>"000110000",
  55814=>"101110110",
  55815=>"000000111",
  55816=>"001110101",
  55817=>"110100000",
  55818=>"001110111",
  55819=>"000100110",
  55820=>"110000000",
  55821=>"000001100",
  55822=>"100001011",
  55823=>"110000111",
  55824=>"110101111",
  55825=>"000000111",
  55826=>"111111111",
  55827=>"000111111",
  55828=>"000000000",
  55829=>"110111000",
  55830=>"000100010",
  55831=>"000000111",
  55832=>"010000001",
  55833=>"111010001",
  55834=>"000101111",
  55835=>"111110100",
  55836=>"001101111",
  55837=>"000010010",
  55838=>"111001111",
  55839=>"101101000",
  55840=>"010010000",
  55841=>"000000111",
  55842=>"000010000",
  55843=>"100000000",
  55844=>"011000000",
  55845=>"000000011",
  55846=>"111100000",
  55847=>"000011000",
  55848=>"011000000",
  55849=>"100111111",
  55850=>"101000111",
  55851=>"011000000",
  55852=>"001000111",
  55853=>"101010000",
  55854=>"000001000",
  55855=>"000011010",
  55856=>"000111111",
  55857=>"101110100",
  55858=>"001111111",
  55859=>"000100111",
  55860=>"011001010",
  55861=>"000001111",
  55862=>"100001011",
  55863=>"010011111",
  55864=>"010000001",
  55865=>"111101101",
  55866=>"000000000",
  55867=>"001001110",
  55868=>"001001001",
  55869=>"011011001",
  55870=>"000000000",
  55871=>"101100010",
  55872=>"101101111",
  55873=>"110010010",
  55874=>"000110010",
  55875=>"011111100",
  55876=>"000010000",
  55877=>"011111000",
  55878=>"111110101",
  55879=>"010010011",
  55880=>"001001001",
  55881=>"111101101",
  55882=>"001000000",
  55883=>"010101011",
  55884=>"011111000",
  55885=>"101101000",
  55886=>"001011001",
  55887=>"011111011",
  55888=>"101111000",
  55889=>"111111111",
  55890=>"000010111",
  55891=>"001100100",
  55892=>"111101001",
  55893=>"000000110",
  55894=>"101101110",
  55895=>"000000111",
  55896=>"110011111",
  55897=>"100000100",
  55898=>"100100000",
  55899=>"011001110",
  55900=>"101000000",
  55901=>"101101000",
  55902=>"111111111",
  55903=>"100001011",
  55904=>"111111111",
  55905=>"111111111",
  55906=>"000000000",
  55907=>"001101100",
  55908=>"111111000",
  55909=>"011011111",
  55910=>"110010111",
  55911=>"111111000",
  55912=>"100000011",
  55913=>"010000111",
  55914=>"001001111",
  55915=>"100111000",
  55916=>"000000000",
  55917=>"001100111",
  55918=>"000000000",
  55919=>"000000111",
  55920=>"110111010",
  55921=>"000000111",
  55922=>"010000110",
  55923=>"010010011",
  55924=>"000000011",
  55925=>"001000000",
  55926=>"111000111",
  55927=>"100000000",
  55928=>"000000100",
  55929=>"001001000",
  55930=>"000111111",
  55931=>"000000000",
  55932=>"001001111",
  55933=>"101011000",
  55934=>"011111010",
  55935=>"111101000",
  55936=>"100000111",
  55937=>"011111111",
  55938=>"001000000",
  55939=>"001001000",
  55940=>"000000111",
  55941=>"111110010",
  55942=>"000000110",
  55943=>"110001001",
  55944=>"110111011",
  55945=>"000000111",
  55946=>"101111011",
  55947=>"111010000",
  55948=>"110010000",
  55949=>"111011101",
  55950=>"111011000",
  55951=>"111000001",
  55952=>"001111110",
  55953=>"001111111",
  55954=>"111000001",
  55955=>"111111111",
  55956=>"000001101",
  55957=>"000000111",
  55958=>"110111000",
  55959=>"001001011",
  55960=>"000100111",
  55961=>"100010000",
  55962=>"001011101",
  55963=>"001100001",
  55964=>"111110111",
  55965=>"111111111",
  55966=>"000100111",
  55967=>"010110101",
  55968=>"001111100",
  55969=>"110011111",
  55970=>"111111010",
  55971=>"111011000",
  55972=>"110001111",
  55973=>"111010001",
  55974=>"100110101",
  55975=>"001000010",
  55976=>"000000111",
  55977=>"010000000",
  55978=>"110000000",
  55979=>"000111111",
  55980=>"000000000",
  55981=>"101101111",
  55982=>"101101000",
  55983=>"110110000",
  55984=>"111111100",
  55985=>"001101100",
  55986=>"001000000",
  55987=>"011100100",
  55988=>"111011010",
  55989=>"000000111",
  55990=>"011011000",
  55991=>"101101001",
  55992=>"000100000",
  55993=>"011101100",
  55994=>"101010010",
  55995=>"110111101",
  55996=>"111111000",
  55997=>"011010111",
  55998=>"100011111",
  55999=>"000000000",
  56000=>"100111000",
  56001=>"100111000",
  56002=>"000000011",
  56003=>"100011011",
  56004=>"000111000",
  56005=>"100000001",
  56006=>"000010111",
  56007=>"110000000",
  56008=>"111111000",
  56009=>"011010000",
  56010=>"010010000",
  56011=>"000001111",
  56012=>"000110100",
  56013=>"000001001",
  56014=>"010001000",
  56015=>"011011001",
  56016=>"111001010",
  56017=>"110100000",
  56018=>"111010000",
  56019=>"011010111",
  56020=>"111111000",
  56021=>"011001000",
  56022=>"111111000",
  56023=>"000000001",
  56024=>"111110000",
  56025=>"001001111",
  56026=>"110010000",
  56027=>"000000100",
  56028=>"000011111",
  56029=>"111000101",
  56030=>"111010101",
  56031=>"101111111",
  56032=>"110110000",
  56033=>"000001111",
  56034=>"111111011",
  56035=>"111011000",
  56036=>"111001000",
  56037=>"011000000",
  56038=>"111000111",
  56039=>"011011001",
  56040=>"000101111",
  56041=>"111000000",
  56042=>"111101111",
  56043=>"010110111",
  56044=>"000110111",
  56045=>"010101011",
  56046=>"001000000",
  56047=>"101101111",
  56048=>"001001111",
  56049=>"001010000",
  56050=>"000000000",
  56051=>"001000000",
  56052=>"110010011",
  56053=>"101011000",
  56054=>"011000000",
  56055=>"011111011",
  56056=>"000000111",
  56057=>"101001111",
  56058=>"111100000",
  56059=>"110001000",
  56060=>"000110111",
  56061=>"000011000",
  56062=>"101111111",
  56063=>"000000101",
  56064=>"000010000",
  56065=>"000000110",
  56066=>"101111111",
  56067=>"110000000",
  56068=>"000011001",
  56069=>"110110000",
  56070=>"111001111",
  56071=>"111010110",
  56072=>"000000110",
  56073=>"111000000",
  56074=>"010000000",
  56075=>"110110010",
  56076=>"000111111",
  56077=>"001001001",
  56078=>"000000011",
  56079=>"000110010",
  56080=>"000000100",
  56081=>"111111000",
  56082=>"001010001",
  56083=>"010000011",
  56084=>"001001111",
  56085=>"011111111",
  56086=>"000001011",
  56087=>"010001111",
  56088=>"111001000",
  56089=>"101111000",
  56090=>"000111111",
  56091=>"010000011",
  56092=>"101110111",
  56093=>"000101000",
  56094=>"000000000",
  56095=>"111101101",
  56096=>"000110000",
  56097=>"100000010",
  56098=>"000000010",
  56099=>"000110111",
  56100=>"001001100",
  56101=>"000000000",
  56102=>"000110111",
  56103=>"001001111",
  56104=>"111000010",
  56105=>"110010001",
  56106=>"111000001",
  56107=>"101000000",
  56108=>"101111011",
  56109=>"011001110",
  56110=>"111111101",
  56111=>"000001000",
  56112=>"111101000",
  56113=>"011011000",
  56114=>"010010101",
  56115=>"100110111",
  56116=>"001000000",
  56117=>"100110110",
  56118=>"000100001",
  56119=>"010001101",
  56120=>"001000010",
  56121=>"111000000",
  56122=>"111101101",
  56123=>"111000010",
  56124=>"011010100",
  56125=>"111001010",
  56126=>"000111110",
  56127=>"010110110",
  56128=>"001110111",
  56129=>"000100000",
  56130=>"111110010",
  56131=>"011011000",
  56132=>"001000000",
  56133=>"001000000",
  56134=>"000000001",
  56135=>"111111100",
  56136=>"111100000",
  56137=>"010010010",
  56138=>"110000000",
  56139=>"101101000",
  56140=>"000101001",
  56141=>"100001011",
  56142=>"010111000",
  56143=>"101001111",
  56144=>"001000000",
  56145=>"011011111",
  56146=>"000000000",
  56147=>"011000100",
  56148=>"000010000",
  56149=>"010011111",
  56150=>"011011001",
  56151=>"111110000",
  56152=>"011110101",
  56153=>"110110011",
  56154=>"001111110",
  56155=>"100111110",
  56156=>"000001111",
  56157=>"001001001",
  56158=>"000001111",
  56159=>"110100000",
  56160=>"010000111",
  56161=>"000000000",
  56162=>"110000000",
  56163=>"100001011",
  56164=>"111010000",
  56165=>"111000100",
  56166=>"101000000",
  56167=>"111001001",
  56168=>"111111101",
  56169=>"000100000",
  56170=>"111000000",
  56171=>"001001000",
  56172=>"111111101",
  56173=>"010000001",
  56174=>"000101101",
  56175=>"110000010",
  56176=>"111011111",
  56177=>"100000001",
  56178=>"000000100",
  56179=>"000110010",
  56180=>"111000000",
  56181=>"111000000",
  56182=>"000010010",
  56183=>"000100111",
  56184=>"011011000",
  56185=>"111111000",
  56186=>"111111111",
  56187=>"000111000",
  56188=>"101100001",
  56189=>"110100000",
  56190=>"000001010",
  56191=>"000001101",
  56192=>"000110110",
  56193=>"110111010",
  56194=>"000100111",
  56195=>"010000110",
  56196=>"001010111",
  56197=>"001001101",
  56198=>"001000001",
  56199=>"000010001",
  56200=>"110111100",
  56201=>"000101000",
  56202=>"000100000",
  56203=>"111100000",
  56204=>"111101101",
  56205=>"000111111",
  56206=>"111111111",
  56207=>"110000000",
  56208=>"001100001",
  56209=>"111110111",
  56210=>"001000101",
  56211=>"111100010",
  56212=>"001011110",
  56213=>"111010110",
  56214=>"001111111",
  56215=>"000111110",
  56216=>"110101000",
  56217=>"000000111",
  56218=>"000000110",
  56219=>"000000000",
  56220=>"111000101",
  56221=>"110111000",
  56222=>"110011011",
  56223=>"111010000",
  56224=>"100110111",
  56225=>"001000000",
  56226=>"110111001",
  56227=>"010111001",
  56228=>"111110110",
  56229=>"000111111",
  56230=>"101110101",
  56231=>"111111011",
  56232=>"111100111",
  56233=>"000010010",
  56234=>"111110110",
  56235=>"111110010",
  56236=>"101110110",
  56237=>"110111110",
  56238=>"111110010",
  56239=>"111011111",
  56240=>"111110101",
  56241=>"011011000",
  56242=>"000001000",
  56243=>"001001001",
  56244=>"010010111",
  56245=>"000111111",
  56246=>"000000010",
  56247=>"000110110",
  56248=>"110000110",
  56249=>"000100100",
  56250=>"000000110",
  56251=>"111001010",
  56252=>"010000111",
  56253=>"111111110",
  56254=>"000011011",
  56255=>"000000000",
  56256=>"000000000",
  56257=>"000100000",
  56258=>"110010111",
  56259=>"001111100",
  56260=>"100001101",
  56261=>"111001001",
  56262=>"110111010",
  56263=>"011000000",
  56264=>"000010000",
  56265=>"000000110",
  56266=>"000000110",
  56267=>"101000001",
  56268=>"111010100",
  56269=>"001001100",
  56270=>"110111110",
  56271=>"010101000",
  56272=>"000110110",
  56273=>"000110100",
  56274=>"111000000",
  56275=>"000110111",
  56276=>"001011111",
  56277=>"100100100",
  56278=>"000000101",
  56279=>"101001101",
  56280=>"101001001",
  56281=>"000000110",
  56282=>"001111110",
  56283=>"111001000",
  56284=>"001000000",
  56285=>"111110110",
  56286=>"000110111",
  56287=>"111001001",
  56288=>"000010110",
  56289=>"000000100",
  56290=>"101111111",
  56291=>"001111101",
  56292=>"100101000",
  56293=>"111111000",
  56294=>"011111111",
  56295=>"111011111",
  56296=>"011010010",
  56297=>"000000001",
  56298=>"010000001",
  56299=>"000000111",
  56300=>"111111111",
  56301=>"110110100",
  56302=>"000010000",
  56303=>"000100110",
  56304=>"000000111",
  56305=>"111000101",
  56306=>"111000000",
  56307=>"000001111",
  56308=>"100000011",
  56309=>"000000000",
  56310=>"110101000",
  56311=>"110000000",
  56312=>"000000110",
  56313=>"011111101",
  56314=>"000000010",
  56315=>"000000011",
  56316=>"100111111",
  56317=>"101000000",
  56318=>"010111111",
  56319=>"111100001",
  56320=>"000100100",
  56321=>"100000001",
  56322=>"000000001",
  56323=>"000001000",
  56324=>"111111000",
  56325=>"111111111",
  56326=>"001001111",
  56327=>"111010000",
  56328=>"010011000",
  56329=>"111101001",
  56330=>"000010111",
  56331=>"000000000",
  56332=>"000000111",
  56333=>"110111110",
  56334=>"011011011",
  56335=>"001000000",
  56336=>"111110010",
  56337=>"001000111",
  56338=>"000100100",
  56339=>"101001000",
  56340=>"011101111",
  56341=>"100100000",
  56342=>"101000001",
  56343=>"001001001",
  56344=>"001000111",
  56345=>"110111111",
  56346=>"110111000",
  56347=>"011000000",
  56348=>"000010000",
  56349=>"000001101",
  56350=>"011111111",
  56351=>"110000000",
  56352=>"001001011",
  56353=>"110110110",
  56354=>"110100010",
  56355=>"110010110",
  56356=>"101100000",
  56357=>"001011011",
  56358=>"010110010",
  56359=>"000000000",
  56360=>"010111110",
  56361=>"000000100",
  56362=>"000001101",
  56363=>"000000010",
  56364=>"101100101",
  56365=>"001010111",
  56366=>"000101111",
  56367=>"101001001",
  56368=>"110111110",
  56369=>"001100111",
  56370=>"001111110",
  56371=>"001111110",
  56372=>"000000001",
  56373=>"001100011",
  56374=>"000000001",
  56375=>"000000100",
  56376=>"011000001",
  56377=>"001000001",
  56378=>"101101110",
  56379=>"000001111",
  56380=>"100010100",
  56381=>"001111010",
  56382=>"000000000",
  56383=>"011111000",
  56384=>"111111111",
  56385=>"101101111",
  56386=>"101000111",
  56387=>"110111111",
  56388=>"000001101",
  56389=>"001110110",
  56390=>"011011000",
  56391=>"101101010",
  56392=>"101000110",
  56393=>"110010000",
  56394=>"001000111",
  56395=>"000001110",
  56396=>"110000000",
  56397=>"111100010",
  56398=>"000011001",
  56399=>"001000010",
  56400=>"100000000",
  56401=>"000011111",
  56402=>"001000101",
  56403=>"101100000",
  56404=>"101000111",
  56405=>"011110010",
  56406=>"011011011",
  56407=>"111111000",
  56408=>"101101111",
  56409=>"101100101",
  56410=>"111010000",
  56411=>"111001001",
  56412=>"000110000",
  56413=>"000000011",
  56414=>"101011001",
  56415=>"011111110",
  56416=>"001000000",
  56417=>"001111110",
  56418=>"000000001",
  56419=>"001000000",
  56420=>"100110100",
  56421=>"111110111",
  56422=>"001011110",
  56423=>"111101000",
  56424=>"111110010",
  56425=>"001001011",
  56426=>"000101111",
  56427=>"110110111",
  56428=>"101000011",
  56429=>"101111111",
  56430=>"100100100",
  56431=>"000000111",
  56432=>"111100000",
  56433=>"000111101",
  56434=>"011000100",
  56435=>"001001110",
  56436=>"001101111",
  56437=>"000000011",
  56438=>"110110000",
  56439=>"111111000",
  56440=>"000010111",
  56441=>"111010010",
  56442=>"000111101",
  56443=>"000001010",
  56444=>"011011001",
  56445=>"101000000",
  56446=>"111110000",
  56447=>"110110110",
  56448=>"001001111",
  56449=>"001010011",
  56450=>"001010101",
  56451=>"000101110",
  56452=>"101000111",
  56453=>"111101110",
  56454=>"010100111",
  56455=>"110110110",
  56456=>"011011101",
  56457=>"001011111",
  56458=>"000000111",
  56459=>"101001111",
  56460=>"010000000",
  56461=>"001110111",
  56462=>"101000000",
  56463=>"000000000",
  56464=>"001001111",
  56465=>"111110000",
  56466=>"110000000",
  56467=>"101000110",
  56468=>"111010000",
  56469=>"111101001",
  56470=>"100001111",
  56471=>"011011111",
  56472=>"111111110",
  56473=>"010110010",
  56474=>"001111110",
  56475=>"101100110",
  56476=>"001101100",
  56477=>"001000111",
  56478=>"000111101",
  56479=>"001001111",
  56480=>"100100010",
  56481=>"000010000",
  56482=>"000001111",
  56483=>"001101000",
  56484=>"000000000",
  56485=>"111100100",
  56486=>"110110110",
  56487=>"000000110",
  56488=>"111101111",
  56489=>"110110110",
  56490=>"010000101",
  56491=>"000000001",
  56492=>"011111110",
  56493=>"110010000",
  56494=>"101111011",
  56495=>"001000110",
  56496=>"110110000",
  56497=>"001001011",
  56498=>"000100111",
  56499=>"000101101",
  56500=>"111111111",
  56501=>"000000001",
  56502=>"000000010",
  56503=>"101111101",
  56504=>"011010011",
  56505=>"011101010",
  56506=>"010000110",
  56507=>"110110100",
  56508=>"001001010",
  56509=>"111110000",
  56510=>"001000000",
  56511=>"000101101",
  56512=>"000000001",
  56513=>"101001000",
  56514=>"010111010",
  56515=>"110110001",
  56516=>"000101111",
  56517=>"001101111",
  56518=>"111000000",
  56519=>"010010000",
  56520=>"110000000",
  56521=>"111110010",
  56522=>"001001111",
  56523=>"001000000",
  56524=>"000000000",
  56525=>"111000000",
  56526=>"101000000",
  56527=>"110110000",
  56528=>"111011000",
  56529=>"110100110",
  56530=>"110110000",
  56531=>"100000000",
  56532=>"111000000",
  56533=>"000000111",
  56534=>"001100101",
  56535=>"111111101",
  56536=>"011110111",
  56537=>"000000000",
  56538=>"011001000",
  56539=>"001001101",
  56540=>"001001101",
  56541=>"011001111",
  56542=>"000000110",
  56543=>"111101101",
  56544=>"010010000",
  56545=>"000001101",
  56546=>"001001111",
  56547=>"100101111",
  56548=>"001000000",
  56549=>"000001011",
  56550=>"111001111",
  56551=>"011100100",
  56552=>"000101111",
  56553=>"000000000",
  56554=>"001100111",
  56555=>"001001001",
  56556=>"110000000",
  56557=>"000111000",
  56558=>"000000000",
  56559=>"100110111",
  56560=>"000000111",
  56561=>"001101111",
  56562=>"101001111",
  56563=>"001011100",
  56564=>"110101000",
  56565=>"111001100",
  56566=>"000000000",
  56567=>"101011110",
  56568=>"010110010",
  56569=>"001001010",
  56570=>"000000000",
  56571=>"111001001",
  56572=>"000111111",
  56573=>"100101101",
  56574=>"110110011",
  56575=>"000010110",
  56576=>"011011100",
  56577=>"001001100",
  56578=>"111101101",
  56579=>"110010000",
  56580=>"100110110",
  56581=>"111000010",
  56582=>"000010000",
  56583=>"100010010",
  56584=>"001011100",
  56585=>"101100100",
  56586=>"000110110",
  56587=>"111101111",
  56588=>"000000000",
  56589=>"010111111",
  56590=>"111100010",
  56591=>"111011001",
  56592=>"011100100",
  56593=>"111000000",
  56594=>"101100101",
  56595=>"000000000",
  56596=>"111100000",
  56597=>"110000000",
  56598=>"111101101",
  56599=>"111111101",
  56600=>"101000111",
  56601=>"001010010",
  56602=>"000111101",
  56603=>"000001001",
  56604=>"111011000",
  56605=>"000000000",
  56606=>"111101001",
  56607=>"011111010",
  56608=>"101001000",
  56609=>"000111111",
  56610=>"100000011",
  56611=>"000010011",
  56612=>"001001001",
  56613=>"110010010",
  56614=>"111111000",
  56615=>"000010000",
  56616=>"111111111",
  56617=>"111111100",
  56618=>"101111111",
  56619=>"101000000",
  56620=>"011111011",
  56621=>"010010010",
  56622=>"110000100",
  56623=>"110110111",
  56624=>"111001000",
  56625=>"101100100",
  56626=>"101010010",
  56627=>"001010111",
  56628=>"000000001",
  56629=>"000100000",
  56630=>"010110100",
  56631=>"000000010",
  56632=>"100000011",
  56633=>"000011010",
  56634=>"000001001",
  56635=>"101101000",
  56636=>"100110010",
  56637=>"000111000",
  56638=>"000101100",
  56639=>"111111100",
  56640=>"111101000",
  56641=>"111111000",
  56642=>"000011111",
  56643=>"011101000",
  56644=>"010111011",
  56645=>"011000101",
  56646=>"000100111",
  56647=>"011011010",
  56648=>"000000010",
  56649=>"000000000",
  56650=>"000110100",
  56651=>"000010111",
  56652=>"111000001",
  56653=>"000110100",
  56654=>"101101001",
  56655=>"110111010",
  56656=>"010010011",
  56657=>"111101111",
  56658=>"010010000",
  56659=>"011000000",
  56660=>"000110000",
  56661=>"101000100",
  56662=>"000110100",
  56663=>"100100100",
  56664=>"000111011",
  56665=>"000111000",
  56666=>"000001000",
  56667=>"000101111",
  56668=>"000000000",
  56669=>"010101101",
  56670=>"111000000",
  56671=>"100000001",
  56672=>"111111010",
  56673=>"000000000",
  56674=>"100100101",
  56675=>"111110100",
  56676=>"100111100",
  56677=>"000110100",
  56678=>"011010010",
  56679=>"111000000",
  56680=>"111101111",
  56681=>"111111110",
  56682=>"101000111",
  56683=>"111010100",
  56684=>"000001010",
  56685=>"111111111",
  56686=>"000100000",
  56687=>"110110101",
  56688=>"110101010",
  56689=>"111101000",
  56690=>"011101001",
  56691=>"100010100",
  56692=>"110111001",
  56693=>"111100101",
  56694=>"000000111",
  56695=>"111100000",
  56696=>"111000000",
  56697=>"000111111",
  56698=>"101000011",
  56699=>"100100110",
  56700=>"100110000",
  56701=>"010010000",
  56702=>"101100010",
  56703=>"111100111",
  56704=>"000010000",
  56705=>"111100100",
  56706=>"110110101",
  56707=>"010111111",
  56708=>"000010010",
  56709=>"111111000",
  56710=>"110010001",
  56711=>"000100000",
  56712=>"001110110",
  56713=>"000100010",
  56714=>"111111111",
  56715=>"111100111",
  56716=>"101100101",
  56717=>"111000001",
  56718=>"000010001",
  56719=>"000000000",
  56720=>"011111100",
  56721=>"000000000",
  56722=>"101101100",
  56723=>"000000000",
  56724=>"000101110",
  56725=>"101100101",
  56726=>"010111000",
  56727=>"100100100",
  56728=>"100010010",
  56729=>"111111011",
  56730=>"111111000",
  56731=>"111000100",
  56732=>"000010011",
  56733=>"100101000",
  56734=>"011011010",
  56735=>"010111101",
  56736=>"100101001",
  56737=>"101100101",
  56738=>"111111000",
  56739=>"000000011",
  56740=>"001101000",
  56741=>"000111001",
  56742=>"111000001",
  56743=>"000010010",
  56744=>"011000000",
  56745=>"000101110",
  56746=>"111110111",
  56747=>"000111101",
  56748=>"010101111",
  56749=>"000000011",
  56750=>"000110100",
  56751=>"000000110",
  56752=>"011000010",
  56753=>"000001000",
  56754=>"111101101",
  56755=>"001001010",
  56756=>"111011000",
  56757=>"001010000",
  56758=>"000100111",
  56759=>"000001000",
  56760=>"000010010",
  56761=>"000000010",
  56762=>"010111111",
  56763=>"000010010",
  56764=>"110111111",
  56765=>"111101111",
  56766=>"111001001",
  56767=>"101101010",
  56768=>"000000000",
  56769=>"000000111",
  56770=>"111111100",
  56771=>"110001001",
  56772=>"001111011",
  56773=>"011001111",
  56774=>"000011011",
  56775=>"101100111",
  56776=>"101010100",
  56777=>"111101100",
  56778=>"111001111",
  56779=>"101000000",
  56780=>"111100000",
  56781=>"001001010",
  56782=>"100000000",
  56783=>"111111111",
  56784=>"010000000",
  56785=>"000011001",
  56786=>"000010111",
  56787=>"111111000",
  56788=>"100100001",
  56789=>"100000010",
  56790=>"010111110",
  56791=>"010111010",
  56792=>"111001000",
  56793=>"100010011",
  56794=>"011011010",
  56795=>"101100111",
  56796=>"111111001",
  56797=>"100011000",
  56798=>"000111111",
  56799=>"000000000",
  56800=>"101000101",
  56801=>"011000000",
  56802=>"111000001",
  56803=>"001001111",
  56804=>"101000000",
  56805=>"111000010",
  56806=>"101111101",
  56807=>"000010101",
  56808=>"000000000",
  56809=>"000010000",
  56810=>"100001101",
  56811=>"000000111",
  56812=>"111000000",
  56813=>"111000001",
  56814=>"000000000",
  56815=>"000110100",
  56816=>"000000000",
  56817=>"010100111",
  56818=>"111101000",
  56819=>"000011001",
  56820=>"000010001",
  56821=>"000000111",
  56822=>"000000010",
  56823=>"000000011",
  56824=>"111001000",
  56825=>"000010011",
  56826=>"010001111",
  56827=>"000111010",
  56828=>"011111111",
  56829=>"111100000",
  56830=>"010011011",
  56831=>"111111111",
  56832=>"001111111",
  56833=>"001000100",
  56834=>"001010000",
  56835=>"111011001",
  56836=>"000100111",
  56837=>"000001000",
  56838=>"101000000",
  56839=>"111011111",
  56840=>"111001001",
  56841=>"001010110",
  56842=>"000110110",
  56843=>"000000000",
  56844=>"001101101",
  56845=>"111000000",
  56846=>"011111010",
  56847=>"100110010",
  56848=>"111001000",
  56849=>"111000000",
  56850=>"110001000",
  56851=>"110110000",
  56852=>"011111111",
  56853=>"111111001",
  56854=>"001011001",
  56855=>"111000101",
  56856=>"001000000",
  56857=>"111001001",
  56858=>"001000000",
  56859=>"000110110",
  56860=>"000001000",
  56861=>"000111110",
  56862=>"010110001",
  56863=>"111001000",
  56864=>"001010000",
  56865=>"011000001",
  56866=>"000000110",
  56867=>"000000100",
  56868=>"100100001",
  56869=>"110100100",
  56870=>"011111000",
  56871=>"000000000",
  56872=>"000110110",
  56873=>"000000110",
  56874=>"001001001",
  56875=>"010111010",
  56876=>"010111111",
  56877=>"001111010",
  56878=>"011111111",
  56879=>"101000000",
  56880=>"000000110",
  56881=>"000101101",
  56882=>"100000111",
  56883=>"110110111",
  56884=>"001110110",
  56885=>"100110111",
  56886=>"010111001",
  56887=>"111001001",
  56888=>"110000001",
  56889=>"111001001",
  56890=>"101001000",
  56891=>"111110110",
  56892=>"101111110",
  56893=>"011011111",
  56894=>"001000000",
  56895=>"000101100",
  56896=>"110101000",
  56897=>"100100111",
  56898=>"111001000",
  56899=>"111001000",
  56900=>"001001000",
  56901=>"001000000",
  56902=>"000000101",
  56903=>"000000100",
  56904=>"001001000",
  56905=>"111000000",
  56906=>"111001001",
  56907=>"111001001",
  56908=>"111011000",
  56909=>"001100100",
  56910=>"001111111",
  56911=>"110110110",
  56912=>"111100000",
  56913=>"110111111",
  56914=>"111101110",
  56915=>"010000000",
  56916=>"110000000",
  56917=>"001110110",
  56918=>"001011001",
  56919=>"011000000",
  56920=>"111001000",
  56921=>"011100100",
  56922=>"011111111",
  56923=>"111111010",
  56924=>"001001001",
  56925=>"000000000",
  56926=>"000110100",
  56927=>"101000001",
  56928=>"001011000",
  56929=>"110001000",
  56930=>"000001111",
  56931=>"101101100",
  56932=>"111111001",
  56933=>"011000000",
  56934=>"000001001",
  56935=>"000110110",
  56936=>"111010100",
  56937=>"110010000",
  56938=>"000000110",
  56939=>"001001000",
  56940=>"000010110",
  56941=>"110110110",
  56942=>"111011011",
  56943=>"000000000",
  56944=>"000110110",
  56945=>"001000111",
  56946=>"110011000",
  56947=>"010110010",
  56948=>"000000000",
  56949=>"011001000",
  56950=>"011001000",
  56951=>"001110000",
  56952=>"010000000",
  56953=>"111110100",
  56954=>"000110110",
  56955=>"000000000",
  56956=>"011011110",
  56957=>"111100000",
  56958=>"011000001",
  56959=>"111100000",
  56960=>"100000000",
  56961=>"111001000",
  56962=>"000110110",
  56963=>"000000111",
  56964=>"110111001",
  56965=>"000110111",
  56966=>"001111110",
  56967=>"111101100",
  56968=>"011011011",
  56969=>"000110110",
  56970=>"111110000",
  56971=>"000101100",
  56972=>"111101110",
  56973=>"100110110",
  56974=>"001110110",
  56975=>"110101000",
  56976=>"111001000",
  56977=>"101101100",
  56978=>"001000000",
  56979=>"100111101",
  56980=>"110110110",
  56981=>"110000000",
  56982=>"101111100",
  56983=>"000001111",
  56984=>"000110110",
  56985=>"100001101",
  56986=>"000110111",
  56987=>"000000000",
  56988=>"111111001",
  56989=>"000110110",
  56990=>"111111111",
  56991=>"111001001",
  56992=>"001000001",
  56993=>"000000001",
  56994=>"001001000",
  56995=>"111000001",
  56996=>"000001010",
  56997=>"011010000",
  56998=>"001110111",
  56999=>"000110110",
  57000=>"000010110",
  57001=>"000101001",
  57002=>"000000000",
  57003=>"111010001",
  57004=>"000000000",
  57005=>"111101000",
  57006=>"100100000",
  57007=>"100001000",
  57008=>"010001001",
  57009=>"111001011",
  57010=>"110001000",
  57011=>"000001100",
  57012=>"001111111",
  57013=>"110000000",
  57014=>"010000000",
  57015=>"000110110",
  57016=>"100111110",
  57017=>"110111110",
  57018=>"000110111",
  57019=>"101000111",
  57020=>"100111111",
  57021=>"000110111",
  57022=>"000000000",
  57023=>"001000000",
  57024=>"111001000",
  57025=>"000000001",
  57026=>"110111000",
  57027=>"001011011",
  57028=>"110110111",
  57029=>"011101110",
  57030=>"111000100",
  57031=>"111001000",
  57032=>"111001111",
  57033=>"111001000",
  57034=>"111111110",
  57035=>"111001001",
  57036=>"111001000",
  57037=>"100100110",
  57038=>"010000111",
  57039=>"110001111",
  57040=>"011001000",
  57041=>"011101010",
  57042=>"111000011",
  57043=>"111111010",
  57044=>"111001001",
  57045=>"010001000",
  57046=>"111001000",
  57047=>"011000110",
  57048=>"111001000",
  57049=>"100000000",
  57050=>"001000000",
  57051=>"100100110",
  57052=>"100001000",
  57053=>"000110110",
  57054=>"101001000",
  57055=>"001110111",
  57056=>"111001000",
  57057=>"111001001",
  57058=>"100101111",
  57059=>"111001001",
  57060=>"111001000",
  57061=>"001011111",
  57062=>"000011011",
  57063=>"110110010",
  57064=>"000111000",
  57065=>"000010000",
  57066=>"000110110",
  57067=>"001001101",
  57068=>"111001000",
  57069=>"110001001",
  57070=>"000001001",
  57071=>"000110010",
  57072=>"000110110",
  57073=>"001010010",
  57074=>"000000000",
  57075=>"010010000",
  57076=>"000110111",
  57077=>"001001111",
  57078=>"110100100",
  57079=>"000110110",
  57080=>"000001001",
  57081=>"110111100",
  57082=>"001110110",
  57083=>"111111000",
  57084=>"000100101",
  57085=>"000110011",
  57086=>"000111111",
  57087=>"111001001",
  57088=>"000000000",
  57089=>"001011111",
  57090=>"000010001",
  57091=>"001000100",
  57092=>"110111110",
  57093=>"110101100",
  57094=>"000000000",
  57095=>"011111001",
  57096=>"111101100",
  57097=>"011000011",
  57098=>"111110100",
  57099=>"100001110",
  57100=>"101011111",
  57101=>"000000110",
  57102=>"110001000",
  57103=>"000011000",
  57104=>"111011011",
  57105=>"001000000",
  57106=>"100000000",
  57107=>"000000010",
  57108=>"110111111",
  57109=>"000100110",
  57110=>"110010010",
  57111=>"111000001",
  57112=>"010000000",
  57113=>"111111011",
  57114=>"100100110",
  57115=>"111110100",
  57116=>"000100111",
  57117=>"000110100",
  57118=>"110010001",
  57119=>"100101111",
  57120=>"000100000",
  57121=>"000000100",
  57122=>"100001101",
  57123=>"111101100",
  57124=>"100101100",
  57125=>"100001101",
  57126=>"111000000",
  57127=>"100010110",
  57128=>"001000110",
  57129=>"100101111",
  57130=>"010000000",
  57131=>"011011011",
  57132=>"100100000",
  57133=>"111001001",
  57134=>"000001001",
  57135=>"110111111",
  57136=>"000000000",
  57137=>"100100111",
  57138=>"000011011",
  57139=>"000001011",
  57140=>"001111110",
  57141=>"010100000",
  57142=>"110100101",
  57143=>"011010010",
  57144=>"100001001",
  57145=>"100110000",
  57146=>"000000011",
  57147=>"000011000",
  57148=>"111011011",
  57149=>"100100100",
  57150=>"010010000",
  57151=>"110111111",
  57152=>"011011011",
  57153=>"100110001",
  57154=>"001101101",
  57155=>"001010110",
  57156=>"000010000",
  57157=>"000010010",
  57158=>"000111111",
  57159=>"010111000",
  57160=>"100111111",
  57161=>"100100100",
  57162=>"011110100",
  57163=>"011011111",
  57164=>"110110011",
  57165=>"110011011",
  57166=>"000000000",
  57167=>"101111111",
  57168=>"100100110",
  57169=>"100000000",
  57170=>"101001011",
  57171=>"000010110",
  57172=>"110000000",
  57173=>"000110111",
  57174=>"100111111",
  57175=>"100000000",
  57176=>"000001000",
  57177=>"100110111",
  57178=>"100001111",
  57179=>"001001001",
  57180=>"001010011",
  57181=>"000001001",
  57182=>"111010011",
  57183=>"110100100",
  57184=>"110100100",
  57185=>"101110110",
  57186=>"110111000",
  57187=>"000001001",
  57188=>"000000100",
  57189=>"101001101",
  57190=>"000101111",
  57191=>"000011011",
  57192=>"011110100",
  57193=>"100000001",
  57194=>"101001000",
  57195=>"011111011",
  57196=>"111000110",
  57197=>"111000101",
  57198=>"010001001",
  57199=>"111000000",
  57200=>"100110101",
  57201=>"111111001",
  57202=>"001011110",
  57203=>"100110101",
  57204=>"110011110",
  57205=>"000101111",
  57206=>"000000000",
  57207=>"101001011",
  57208=>"011000001",
  57209=>"100000000",
  57210=>"000010010",
  57211=>"000011010",
  57212=>"111011011",
  57213=>"100100000",
  57214=>"011011011",
  57215=>"110110100",
  57216=>"111000000",
  57217=>"111000000",
  57218=>"011000000",
  57219=>"101100000",
  57220=>"100100011",
  57221=>"100100110",
  57222=>"000010100",
  57223=>"000000000",
  57224=>"100110100",
  57225=>"000100100",
  57226=>"011001101",
  57227=>"011011000",
  57228=>"111101011",
  57229=>"010001101",
  57230=>"111111100",
  57231=>"001000100",
  57232=>"100110101",
  57233=>"100011011",
  57234=>"010001111",
  57235=>"001001001",
  57236=>"000000110",
  57237=>"111000011",
  57238=>"110000001",
  57239=>"101101111",
  57240=>"111100100",
  57241=>"111011001",
  57242=>"000000011",
  57243=>"011000110",
  57244=>"101100000",
  57245=>"010010011",
  57246=>"000000001",
  57247=>"101001011",
  57248=>"000001101",
  57249=>"000111011",
  57250=>"000001101",
  57251=>"101110011",
  57252=>"010000000",
  57253=>"111111011",
  57254=>"111100000",
  57255=>"110111110",
  57256=>"011111111",
  57257=>"011000100",
  57258=>"000100100",
  57259=>"011000110",
  57260=>"000110100",
  57261=>"100100111",
  57262=>"110110110",
  57263=>"001010111",
  57264=>"001001100",
  57265=>"000011111",
  57266=>"001011000",
  57267=>"000001101",
  57268=>"000100100",
  57269=>"001001001",
  57270=>"000111110",
  57271=>"000111110",
  57272=>"100100110",
  57273=>"111001111",
  57274=>"101011011",
  57275=>"100011011",
  57276=>"110110111",
  57277=>"101100100",
  57278=>"000000100",
  57279=>"111010110",
  57280=>"101011011",
  57281=>"111011011",
  57282=>"011110100",
  57283=>"000110110",
  57284=>"011011110",
  57285=>"110110000",
  57286=>"111000000",
  57287=>"011011011",
  57288=>"110111011",
  57289=>"100100100",
  57290=>"001111011",
  57291=>"001000011",
  57292=>"010110100",
  57293=>"010110000",
  57294=>"000001011",
  57295=>"111011001",
  57296=>"100100000",
  57297=>"000001000",
  57298=>"001101001",
  57299=>"010010100",
  57300=>"011011111",
  57301=>"100100101",
  57302=>"111100101",
  57303=>"111000011",
  57304=>"011111001",
  57305=>"011110110",
  57306=>"000111111",
  57307=>"000000111",
  57308=>"100011000",
  57309=>"010100100",
  57310=>"111100110",
  57311=>"111001111",
  57312=>"001100100",
  57313=>"101011111",
  57314=>"001011011",
  57315=>"100101110",
  57316=>"000100111",
  57317=>"110100100",
  57318=>"110100100",
  57319=>"001001001",
  57320=>"101101110",
  57321=>"011011111",
  57322=>"110010010",
  57323=>"100111000",
  57324=>"001000000",
  57325=>"100111110",
  57326=>"000000000",
  57327=>"100100100",
  57328=>"011000111",
  57329=>"000001110",
  57330=>"111000010",
  57331=>"001011001",
  57332=>"110100001",
  57333=>"000101000",
  57334=>"000011001",
  57335=>"011010010",
  57336=>"011011011",
  57337=>"110100100",
  57338=>"110011011",
  57339=>"011010011",
  57340=>"110111100",
  57341=>"011011011",
  57342=>"100011100",
  57343=>"000001000",
  57344=>"100100111",
  57345=>"110011111",
  57346=>"110000100",
  57347=>"011011011",
  57348=>"101011011",
  57349=>"001100111",
  57350=>"110000100",
  57351=>"000111011",
  57352=>"100101001",
  57353=>"000000000",
  57354=>"100110111",
  57355=>"111101101",
  57356=>"111100100",
  57357=>"110100111",
  57358=>"110111111",
  57359=>"011111111",
  57360=>"100100110",
  57361=>"010011111",
  57362=>"101011111",
  57363=>"011011001",
  57364=>"001111101",
  57365=>"101000100",
  57366=>"000010001",
  57367=>"101111111",
  57368=>"101011111",
  57369=>"111100000",
  57370=>"101111111",
  57371=>"111111101",
  57372=>"100000000",
  57373=>"011111011",
  57374=>"000000111",
  57375=>"101100100",
  57376=>"010100101",
  57377=>"111111111",
  57378=>"011011001",
  57379=>"111000000",
  57380=>"110111111",
  57381=>"000000011",
  57382=>"100011010",
  57383=>"111111101",
  57384=>"001000000",
  57385=>"000111001",
  57386=>"100000000",
  57387=>"000000000",
  57388=>"111111111",
  57389=>"111111101",
  57390=>"000000010",
  57391=>"010110110",
  57392=>"111110011",
  57393=>"111110111",
  57394=>"111011100",
  57395=>"010111001",
  57396=>"111111011",
  57397=>"011011100",
  57398=>"100110100",
  57399=>"001011011",
  57400=>"000111100",
  57401=>"000001111",
  57402=>"000101101",
  57403=>"110010001",
  57404=>"111000000",
  57405=>"111011111",
  57406=>"000000100",
  57407=>"010011111",
  57408=>"001011000",
  57409=>"000000100",
  57410=>"011110111",
  57411=>"110100111",
  57412=>"000000000",
  57413=>"001111000",
  57414=>"000000000",
  57415=>"000000000",
  57416=>"110011101",
  57417=>"010001000",
  57418=>"010010010",
  57419=>"000000111",
  57420=>"010111111",
  57421=>"001111111",
  57422=>"100111111",
  57423=>"101000101",
  57424=>"000000111",
  57425=>"111111100",
  57426=>"001100101",
  57427=>"000110110",
  57428=>"000000111",
  57429=>"011111001",
  57430=>"000110111",
  57431=>"111000000",
  57432=>"100000000",
  57433=>"011011001",
  57434=>"000000111",
  57435=>"110010110",
  57436=>"000111111",
  57437=>"000110100",
  57438=>"000111010",
  57439=>"111000001",
  57440=>"000000001",
  57441=>"111000000",
  57442=>"111000000",
  57443=>"001110100",
  57444=>"000001000",
  57445=>"000000000",
  57446=>"101111101",
  57447=>"001000000",
  57448=>"010010101",
  57449=>"000111011",
  57450=>"010010010",
  57451=>"101100101",
  57452=>"000010111",
  57453=>"010011011",
  57454=>"100100101",
  57455=>"101010111",
  57456=>"011101101",
  57457=>"010000000",
  57458=>"100111101",
  57459=>"010010000",
  57460=>"010010010",
  57461=>"110101101",
  57462=>"001001000",
  57463=>"111001000",
  57464=>"000000110",
  57465=>"000101001",
  57466=>"010000000",
  57467=>"111110100",
  57468=>"011011011",
  57469=>"000001011",
  57470=>"001001101",
  57471=>"100100101",
  57472=>"110100110",
  57473=>"000000000",
  57474=>"010011111",
  57475=>"111111011",
  57476=>"101110111",
  57477=>"000101000",
  57478=>"000000100",
  57479=>"111100100",
  57480=>"100100000",
  57481=>"111111101",
  57482=>"000011111",
  57483=>"001001011",
  57484=>"110000000",
  57485=>"000100101",
  57486=>"001000000",
  57487=>"001000000",
  57488=>"010011011",
  57489=>"000111111",
  57490=>"000111100",
  57491=>"110001000",
  57492=>"001001111",
  57493=>"111001000",
  57494=>"000010110",
  57495=>"111110100",
  57496=>"000101000",
  57497=>"011001000",
  57498=>"100000000",
  57499=>"000100100",
  57500=>"110100100",
  57501=>"111100000",
  57502=>"000100110",
  57503=>"100100100",
  57504=>"000001111",
  57505=>"111111111",
  57506=>"000000001",
  57507=>"110000111",
  57508=>"111111010",
  57509=>"100110100",
  57510=>"101001000",
  57511=>"100000101",
  57512=>"000011010",
  57513=>"001111001",
  57514=>"110101101",
  57515=>"101101111",
  57516=>"001011111",
  57517=>"000111010",
  57518=>"010000100",
  57519=>"101100101",
  57520=>"111100000",
  57521=>"100110100",
  57522=>"111010000",
  57523=>"011000000",
  57524=>"101111111",
  57525=>"011010011",
  57526=>"000001001",
  57527=>"101000000",
  57528=>"110100100",
  57529=>"110011111",
  57530=>"010111011",
  57531=>"110110100",
  57532=>"111101000",
  57533=>"101000000",
  57534=>"100100100",
  57535=>"111010110",
  57536=>"000000011",
  57537=>"000011000",
  57538=>"000100101",
  57539=>"001100110",
  57540=>"011010001",
  57541=>"111111101",
  57542=>"000011011",
  57543=>"111000110",
  57544=>"111101101",
  57545=>"000000000",
  57546=>"110110100",
  57547=>"000100000",
  57548=>"100000100",
  57549=>"111110100",
  57550=>"100011011",
  57551=>"110111010",
  57552=>"111111111",
  57553=>"000111111",
  57554=>"111110000",
  57555=>"011000111",
  57556=>"011101101",
  57557=>"000111111",
  57558=>"000010101",
  57559=>"000000111",
  57560=>"000000000",
  57561=>"111000000",
  57562=>"011100000",
  57563=>"000000011",
  57564=>"000111110",
  57565=>"000101000",
  57566=>"000000000",
  57567=>"010111111",
  57568=>"111100100",
  57569=>"011100110",
  57570=>"111000100",
  57571=>"011011111",
  57572=>"100000000",
  57573=>"010010011",
  57574=>"111100000",
  57575=>"001000010",
  57576=>"111100100",
  57577=>"000000000",
  57578=>"100111111",
  57579=>"100010111",
  57580=>"111000000",
  57581=>"000000111",
  57582=>"001000011",
  57583=>"000000000",
  57584=>"100100101",
  57585=>"000011100",
  57586=>"001000101",
  57587=>"110111110",
  57588=>"011010011",
  57589=>"101111011",
  57590=>"000000111",
  57591=>"111000000",
  57592=>"111000000",
  57593=>"010100111",
  57594=>"110100111",
  57595=>"000101010",
  57596=>"111011110",
  57597=>"000000000",
  57598=>"000111110",
  57599=>"011000000",
  57600=>"001000000",
  57601=>"000000101",
  57602=>"001110000",
  57603=>"111110000",
  57604=>"000001011",
  57605=>"000000000",
  57606=>"111101011",
  57607=>"101001000",
  57608=>"111001011",
  57609=>"101001001",
  57610=>"011011110",
  57611=>"000001101",
  57612=>"111001111",
  57613=>"111111011",
  57614=>"001000011",
  57615=>"111111110",
  57616=>"001001000",
  57617=>"000000000",
  57618=>"000000000",
  57619=>"010001011",
  57620=>"001000000",
  57621=>"001100100",
  57622=>"000100111",
  57623=>"100111111",
  57624=>"100000011",
  57625=>"111110000",
  57626=>"001000000",
  57627=>"000000000",
  57628=>"000101101",
  57629=>"101111111",
  57630=>"010000011",
  57631=>"111111000",
  57632=>"101111010",
  57633=>"000000011",
  57634=>"000011111",
  57635=>"110111111",
  57636=>"100100111",
  57637=>"011000000",
  57638=>"000111010",
  57639=>"010101001",
  57640=>"010010000",
  57641=>"010000001",
  57642=>"010000001",
  57643=>"100000101",
  57644=>"010000110",
  57645=>"000111111",
  57646=>"000111111",
  57647=>"000000011",
  57648=>"010010011",
  57649=>"001011100",
  57650=>"000010101",
  57651=>"110010000",
  57652=>"000000000",
  57653=>"110110100",
  57654=>"001001011",
  57655=>"010101111",
  57656=>"010000010",
  57657=>"000000000",
  57658=>"000000101",
  57659=>"000111111",
  57660=>"110000100",
  57661=>"111101000",
  57662=>"100000000",
  57663=>"011001001",
  57664=>"011000000",
  57665=>"000000000",
  57666=>"111111111",
  57667=>"110001000",
  57668=>"000010010",
  57669=>"010000000",
  57670=>"111111111",
  57671=>"110000000",
  57672=>"000001100",
  57673=>"010010000",
  57674=>"000001000",
  57675=>"010001001",
  57676=>"010011010",
  57677=>"111111101",
  57678=>"110100000",
  57679=>"000000011",
  57680=>"000001111",
  57681=>"110111000",
  57682=>"000001000",
  57683=>"000100111",
  57684=>"010110111",
  57685=>"010001010",
  57686=>"011011111",
  57687=>"111110010",
  57688=>"111110111",
  57689=>"001101001",
  57690=>"110000011",
  57691=>"001000000",
  57692=>"111010000",
  57693=>"001001001",
  57694=>"111111010",
  57695=>"110100000",
  57696=>"010011000",
  57697=>"110010000",
  57698=>"000000000",
  57699=>"111111101",
  57700=>"100000101",
  57701=>"100100101",
  57702=>"110111001",
  57703=>"111001010",
  57704=>"110111110",
  57705=>"000000000",
  57706=>"110101101",
  57707=>"000101000",
  57708=>"000000010",
  57709=>"000010111",
  57710=>"110011000",
  57711=>"010000010",
  57712=>"111111110",
  57713=>"000000000",
  57714=>"100100100",
  57715=>"111111010",
  57716=>"000011111",
  57717=>"000000000",
  57718=>"110110010",
  57719=>"111000000",
  57720=>"000110010",
  57721=>"000000111",
  57722=>"000111111",
  57723=>"000000111",
  57724=>"110110100",
  57725=>"100001011",
  57726=>"000111111",
  57727=>"100111100",
  57728=>"001100100",
  57729=>"111000000",
  57730=>"010000100",
  57731=>"111100101",
  57732=>"000000000",
  57733=>"111111111",
  57734=>"000000000",
  57735=>"111011010",
  57736=>"101001011",
  57737=>"000010111",
  57738=>"000000001",
  57739=>"010000000",
  57740=>"111111000",
  57741=>"000100000",
  57742=>"000000111",
  57743=>"001000000",
  57744=>"011111111",
  57745=>"010110000",
  57746=>"010111011",
  57747=>"101001011",
  57748=>"111111111",
  57749=>"011011111",
  57750=>"011011000",
  57751=>"000000100",
  57752=>"110000000",
  57753=>"010010010",
  57754=>"011111000",
  57755=>"001101111",
  57756=>"010111111",
  57757=>"010000000",
  57758=>"100010111",
  57759=>"000100101",
  57760=>"100100001",
  57761=>"000000011",
  57762=>"111111001",
  57763=>"000000101",
  57764=>"000000001",
  57765=>"011100100",
  57766=>"110110101",
  57767=>"010010111",
  57768=>"110110111",
  57769=>"010101111",
  57770=>"000000001",
  57771=>"010000000",
  57772=>"111000000",
  57773=>"111111000",
  57774=>"000011001",
  57775=>"111111110",
  57776=>"101000000",
  57777=>"001001111",
  57778=>"101110000",
  57779=>"000000100",
  57780=>"101100111",
  57781=>"111111111",
  57782=>"111110000",
  57783=>"111111100",
  57784=>"011001001",
  57785=>"110110111",
  57786=>"101111100",
  57787=>"011111111",
  57788=>"111000000",
  57789=>"111111011",
  57790=>"100100110",
  57791=>"000000000",
  57792=>"010111000",
  57793=>"010010000",
  57794=>"110101111",
  57795=>"001101100",
  57796=>"000010111",
  57797=>"000001110",
  57798=>"111100000",
  57799=>"110100000",
  57800=>"111111010",
  57801=>"111111011",
  57802=>"001000010",
  57803=>"111110111",
  57804=>"010010010",
  57805=>"011011001",
  57806=>"000111010",
  57807=>"011101110",
  57808=>"011111000",
  57809=>"000001011",
  57810=>"110010010",
  57811=>"010101011",
  57812=>"010000000",
  57813=>"000000111",
  57814=>"111110111",
  57815=>"000001111",
  57816=>"001011010",
  57817=>"110101110",
  57818=>"000001000",
  57819=>"011010011",
  57820=>"011011000",
  57821=>"010000111",
  57822=>"011110010",
  57823=>"111000010",
  57824=>"000000000",
  57825=>"000001101",
  57826=>"111110010",
  57827=>"000001101",
  57828=>"010111000",
  57829=>"000000111",
  57830=>"100111111",
  57831=>"001101101",
  57832=>"110100000",
  57833=>"110010000",
  57834=>"100100111",
  57835=>"111111100",
  57836=>"001000100",
  57837=>"111111110",
  57838=>"000000000",
  57839=>"001000010",
  57840=>"100011010",
  57841=>"101110010",
  57842=>"000000000",
  57843=>"001001111",
  57844=>"100100110",
  57845=>"000000111",
  57846=>"110001000",
  57847=>"001111011",
  57848=>"010110111",
  57849=>"001011111",
  57850=>"000100000",
  57851=>"111011000",
  57852=>"001111111",
  57853=>"000000000",
  57854=>"100100111",
  57855=>"100000101",
  57856=>"111101111",
  57857=>"000000111",
  57858=>"000000110",
  57859=>"111111000",
  57860=>"101000001",
  57861=>"110000000",
  57862=>"010111000",
  57863=>"000111111",
  57864=>"010000000",
  57865=>"010010110",
  57866=>"001011011",
  57867=>"000001110",
  57868=>"000000000",
  57869=>"011001001",
  57870=>"000010011",
  57871=>"100000111",
  57872=>"111111000",
  57873=>"111110010",
  57874=>"100100111",
  57875=>"101000100",
  57876=>"010011111",
  57877=>"000110110",
  57878=>"100101101",
  57879=>"101000000",
  57880=>"001000000",
  57881=>"111101101",
  57882=>"101000000",
  57883=>"010000000",
  57884=>"100100101",
  57885=>"011111101",
  57886=>"111111010",
  57887=>"110111001",
  57888=>"001000001",
  57889=>"001001001",
  57890=>"000000100",
  57891=>"000110111",
  57892=>"001000000",
  57893=>"100000010",
  57894=>"000010110",
  57895=>"100000000",
  57896=>"011111101",
  57897=>"100001001",
  57898=>"000111011",
  57899=>"110000000",
  57900=>"111000000",
  57901=>"111111101",
  57902=>"000010000",
  57903=>"110111111",
  57904=>"011110000",
  57905=>"101000100",
  57906=>"101000111",
  57907=>"000100111",
  57908=>"000000111",
  57909=>"101000101",
  57910=>"000111111",
  57911=>"111111111",
  57912=>"001101000",
  57913=>"111111111",
  57914=>"000000000",
  57915=>"000000000",
  57916=>"100001000",
  57917=>"111111111",
  57918=>"000000000",
  57919=>"110110100",
  57920=>"000000000",
  57921=>"110000010",
  57922=>"011011111",
  57923=>"011011011",
  57924=>"011000001",
  57925=>"111001101",
  57926=>"100110111",
  57927=>"100111111",
  57928=>"111101111",
  57929=>"010111000",
  57930=>"101011111",
  57931=>"000000001",
  57932=>"101000010",
  57933=>"100100000",
  57934=>"011000001",
  57935=>"000101000",
  57936=>"010110110",
  57937=>"111111101",
  57938=>"000000110",
  57939=>"011001100",
  57940=>"000000000",
  57941=>"110100000",
  57942=>"111011001",
  57943=>"000111110",
  57944=>"001000000",
  57945=>"000100100",
  57946=>"001001001",
  57947=>"011001000",
  57948=>"000110000",
  57949=>"111001001",
  57950=>"010010111",
  57951=>"110110111",
  57952=>"101100100",
  57953=>"000000000",
  57954=>"111000000",
  57955=>"100100000",
  57956=>"100110100",
  57957=>"111000110",
  57958=>"111101111",
  57959=>"110111010",
  57960=>"000011111",
  57961=>"101111111",
  57962=>"011001100",
  57963=>"010100111",
  57964=>"101111110",
  57965=>"000111000",
  57966=>"000110110",
  57967=>"011001000",
  57968=>"100101001",
  57969=>"000001000",
  57970=>"000100100",
  57971=>"111111010",
  57972=>"000100100",
  57973=>"001000101",
  57974=>"111111111",
  57975=>"000000000",
  57976=>"000000001",
  57977=>"000010011",
  57978=>"000000101",
  57979=>"010100000",
  57980=>"000110100",
  57981=>"111101010",
  57982=>"000010100",
  57983=>"000000001",
  57984=>"000000010",
  57985=>"111101100",
  57986=>"111111101",
  57987=>"111111101",
  57988=>"000101111",
  57989=>"110111001",
  57990=>"001000000",
  57991=>"000000000",
  57992=>"001011001",
  57993=>"000010000",
  57994=>"111111000",
  57995=>"011111110",
  57996=>"001010000",
  57997=>"010111111",
  57998=>"110111111",
  57999=>"000001000",
  58000=>"111001001",
  58001=>"101010111",
  58002=>"101000001",
  58003=>"000111111",
  58004=>"000100001",
  58005=>"000111010",
  58006=>"110111111",
  58007=>"100000000",
  58008=>"011101110",
  58009=>"001001000",
  58010=>"000111111",
  58011=>"010111000",
  58012=>"111101100",
  58013=>"001110111",
  58014=>"110111001",
  58015=>"101100111",
  58016=>"001111101",
  58017=>"111000000",
  58018=>"010111111",
  58019=>"110001000",
  58020=>"101011111",
  58021=>"100000000",
  58022=>"001000001",
  58023=>"111010000",
  58024=>"011011000",
  58025=>"000111110",
  58026=>"111101100",
  58027=>"001000000",
  58028=>"111101101",
  58029=>"010010010",
  58030=>"010010011",
  58031=>"010110110",
  58032=>"101111111",
  58033=>"101001100",
  58034=>"011001001",
  58035=>"001100100",
  58036=>"011010100",
  58037=>"111111000",
  58038=>"101000000",
  58039=>"000101101",
  58040=>"111110000",
  58041=>"010000000",
  58042=>"110111101",
  58043=>"010101111",
  58044=>"100111110",
  58045=>"111000100",
  58046=>"101001101",
  58047=>"011110110",
  58048=>"000110010",
  58049=>"111000000",
  58050=>"111111110",
  58051=>"000000110",
  58052=>"000000011",
  58053=>"100110001",
  58054=>"110110011",
  58055=>"101101101",
  58056=>"101111101",
  58057=>"110001101",
  58058=>"000111111",
  58059=>"110111111",
  58060=>"110111110",
  58061=>"101011011",
  58062=>"001000000",
  58063=>"001111010",
  58064=>"001000011",
  58065=>"001001000",
  58066=>"000101001",
  58067=>"010100111",
  58068=>"101101111",
  58069=>"000110100",
  58070=>"111000000",
  58071=>"010000101",
  58072=>"000000100",
  58073=>"000000001",
  58074=>"100011001",
  58075=>"000110100",
  58076=>"001000001",
  58077=>"101101000",
  58078=>"010000000",
  58079=>"010111101",
  58080=>"000010011",
  58081=>"011111111",
  58082=>"111001101",
  58083=>"000000101",
  58084=>"101000010",
  58085=>"111001011",
  58086=>"101000111",
  58087=>"101000000",
  58088=>"010001100",
  58089=>"101000101",
  58090=>"000110100",
  58091=>"001000000",
  58092=>"000011111",
  58093=>"000000001",
  58094=>"001000100",
  58095=>"000000000",
  58096=>"000000100",
  58097=>"011011000",
  58098=>"000000111",
  58099=>"100000001",
  58100=>"010110010",
  58101=>"000111111",
  58102=>"000000010",
  58103=>"000000100",
  58104=>"111000000",
  58105=>"111111110",
  58106=>"000000001",
  58107=>"000000100",
  58108=>"111111111",
  58109=>"111111111",
  58110=>"001000101",
  58111=>"111111111",
  58112=>"111011111",
  58113=>"010111010",
  58114=>"100000101",
  58115=>"111001101",
  58116=>"101000000",
  58117=>"111101110",
  58118=>"101011101",
  58119=>"011111101",
  58120=>"000101101",
  58121=>"111100110",
  58122=>"000010100",
  58123=>"110001000",
  58124=>"111001000",
  58125=>"110111000",
  58126=>"000000000",
  58127=>"110110110",
  58128=>"111111100",
  58129=>"111111001",
  58130=>"111111000",
  58131=>"011001001",
  58132=>"001000000",
  58133=>"111101101",
  58134=>"001011111",
  58135=>"111110110",
  58136=>"101000000",
  58137=>"111001111",
  58138=>"011110110",
  58139=>"000111111",
  58140=>"101000000",
  58141=>"001111000",
  58142=>"011000101",
  58143=>"110110100",
  58144=>"111001001",
  58145=>"001100111",
  58146=>"110110100",
  58147=>"110110001",
  58148=>"011011011",
  58149=>"000000000",
  58150=>"111101101",
  58151=>"011011000",
  58152=>"111101111",
  58153=>"000000000",
  58154=>"100101000",
  58155=>"000010000",
  58156=>"011111101",
  58157=>"110110000",
  58158=>"111111111",
  58159=>"011101000",
  58160=>"111100000",
  58161=>"111001001",
  58162=>"110000100",
  58163=>"001000000",
  58164=>"101010010",
  58165=>"000101111",
  58166=>"010011010",
  58167=>"010000000",
  58168=>"111001101",
  58169=>"000000000",
  58170=>"000111100",
  58171=>"000011110",
  58172=>"110110111",
  58173=>"101110110",
  58174=>"000000100",
  58175=>"000000101",
  58176=>"011001000",
  58177=>"000010110",
  58178=>"110001101",
  58179=>"100101001",
  58180=>"000110111",
  58181=>"000000100",
  58182=>"000110000",
  58183=>"000110110",
  58184=>"111011111",
  58185=>"000101101",
  58186=>"010000001",
  58187=>"111011010",
  58188=>"000001101",
  58189=>"000101100",
  58190=>"000100100",
  58191=>"000010100",
  58192=>"010000111",
  58193=>"111111010",
  58194=>"000000000",
  58195=>"000011011",
  58196=>"110100111",
  58197=>"110100011",
  58198=>"111110110",
  58199=>"110100000",
  58200=>"110000100",
  58201=>"011001000",
  58202=>"001001001",
  58203=>"001000000",
  58204=>"000010111",
  58205=>"011011010",
  58206=>"111011111",
  58207=>"001001111",
  58208=>"011000000",
  58209=>"010100110",
  58210=>"010001101",
  58211=>"100110000",
  58212=>"100000000",
  58213=>"111101000",
  58214=>"101011110",
  58215=>"000000000",
  58216=>"111101111",
  58217=>"000100010",
  58218=>"111100101",
  58219=>"001010110",
  58220=>"110001000",
  58221=>"000001000",
  58222=>"000000001",
  58223=>"011111111",
  58224=>"001001000",
  58225=>"111100000",
  58226=>"000110111",
  58227=>"100000000",
  58228=>"010111000",
  58229=>"100000000",
  58230=>"111001000",
  58231=>"101101000",
  58232=>"111110110",
  58233=>"011001110",
  58234=>"111100001",
  58235=>"000010101",
  58236=>"001100100",
  58237=>"100110110",
  58238=>"101011110",
  58239=>"010000010",
  58240=>"111101000",
  58241=>"110000000",
  58242=>"000001100",
  58243=>"001110100",
  58244=>"000100111",
  58245=>"111001000",
  58246=>"100000001",
  58247=>"111001001",
  58248=>"100100100",
  58249=>"000000011",
  58250=>"011010000",
  58251=>"110101100",
  58252=>"000001111",
  58253=>"000000100",
  58254=>"111111101",
  58255=>"001101000",
  58256=>"001000000",
  58257=>"000000100",
  58258=>"111010010",
  58259=>"011011000",
  58260=>"111111000",
  58261=>"000000000",
  58262=>"010111000",
  58263=>"110100100",
  58264=>"011100011",
  58265=>"000110110",
  58266=>"111101101",
  58267=>"000000001",
  58268=>"101101101",
  58269=>"111101111",
  58270=>"010101011",
  58271=>"101111111",
  58272=>"001011011",
  58273=>"101111010",
  58274=>"111111010",
  58275=>"111001000",
  58276=>"111001001",
  58277=>"000100100",
  58278=>"000111000",
  58279=>"111100111",
  58280=>"111111111",
  58281=>"110110000",
  58282=>"000111110",
  58283=>"011001111",
  58284=>"111111101",
  58285=>"111101001",
  58286=>"110010011",
  58287=>"110000000",
  58288=>"110101000",
  58289=>"111001111",
  58290=>"101001010",
  58291=>"100000000",
  58292=>"001010000",
  58293=>"111111111",
  58294=>"100111110",
  58295=>"111010111",
  58296=>"110001110",
  58297=>"100111001",
  58298=>"111011000",
  58299=>"111001110",
  58300=>"100000010",
  58301=>"010111111",
  58302=>"100101101",
  58303=>"000010000",
  58304=>"011000000",
  58305=>"010000100",
  58306=>"000000001",
  58307=>"111100100",
  58308=>"111100000",
  58309=>"001110100",
  58310=>"000000011",
  58311=>"111101101",
  58312=>"110111111",
  58313=>"000111100",
  58314=>"101111000",
  58315=>"000010011",
  58316=>"001010001",
  58317=>"110000000",
  58318=>"000110000",
  58319=>"001000000",
  58320=>"110110000",
  58321=>"110011011",
  58322=>"010101100",
  58323=>"000011111",
  58324=>"011001001",
  58325=>"110110110",
  58326=>"010111010",
  58327=>"111010000",
  58328=>"000000000",
  58329=>"100001000",
  58330=>"000110110",
  58331=>"000101101",
  58332=>"011111101",
  58333=>"000000101",
  58334=>"111101000",
  58335=>"111111101",
  58336=>"000110110",
  58337=>"010000101",
  58338=>"110000000",
  58339=>"111111011",
  58340=>"111000000",
  58341=>"000110111",
  58342=>"111001000",
  58343=>"111110110",
  58344=>"111001100",
  58345=>"010011011",
  58346=>"100010010",
  58347=>"101100101",
  58348=>"001000100",
  58349=>"110110010",
  58350=>"111000101",
  58351=>"011001000",
  58352=>"110000000",
  58353=>"011001011",
  58354=>"000111010",
  58355=>"000110100",
  58356=>"111011101",
  58357=>"000110010",
  58358=>"001000000",
  58359=>"011110000",
  58360=>"111001000",
  58361=>"101000010",
  58362=>"000101011",
  58363=>"000011010",
  58364=>"111111111",
  58365=>"000000000",
  58366=>"000000001",
  58367=>"000000000",
  58368=>"001000100",
  58369=>"000000000",
  58370=>"000010010",
  58371=>"000000001",
  58372=>"000111011",
  58373=>"100011111",
  58374=>"010000000",
  58375=>"000111111",
  58376=>"010001101",
  58377=>"000000010",
  58378=>"001011111",
  58379=>"010000000",
  58380=>"110000000",
  58381=>"011111100",
  58382=>"100100111",
  58383=>"111111111",
  58384=>"100111111",
  58385=>"000000000",
  58386=>"000000000",
  58387=>"100000000",
  58388=>"111001011",
  58389=>"000000111",
  58390=>"100000001",
  58391=>"101111111",
  58392=>"101000000",
  58393=>"010000000",
  58394=>"001000000",
  58395=>"000111110",
  58396=>"111101100",
  58397=>"111001111",
  58398=>"101111111",
  58399=>"011111101",
  58400=>"100000011",
  58401=>"000000101",
  58402=>"101111011",
  58403=>"001111111",
  58404=>"011101101",
  58405=>"001001011",
  58406=>"000110111",
  58407=>"110111000",
  58408=>"100110010",
  58409=>"000110110",
  58410=>"100010111",
  58411=>"000000000",
  58412=>"010100100",
  58413=>"111111111",
  58414=>"010000000",
  58415=>"000111001",
  58416=>"111111110",
  58417=>"001101111",
  58418=>"001000000",
  58419=>"111111000",
  58420=>"000011111",
  58421=>"001101111",
  58422=>"100011011",
  58423=>"010010000",
  58424=>"000000000",
  58425=>"010010011",
  58426=>"111001000",
  58427=>"101011100",
  58428=>"010111001",
  58429=>"111111110",
  58430=>"111001000",
  58431=>"001011111",
  58432=>"100000000",
  58433=>"011101111",
  58434=>"111100000",
  58435=>"000111111",
  58436=>"011000000",
  58437=>"011000101",
  58438=>"000011001",
  58439=>"000101000",
  58440=>"110110111",
  58441=>"000000001",
  58442=>"111000000",
  58443=>"000000010",
  58444=>"111010000",
  58445=>"001001001",
  58446=>"100000010",
  58447=>"111111001",
  58448=>"101000000",
  58449=>"111100000",
  58450=>"111000000",
  58451=>"001001000",
  58452=>"111000000",
  58453=>"100110110",
  58454=>"110011001",
  58455=>"101111110",
  58456=>"110010010",
  58457=>"000001111",
  58458=>"001100110",
  58459=>"110110100",
  58460=>"000000000",
  58461=>"110000000",
  58462=>"000111111",
  58463=>"100110101",
  58464=>"111111111",
  58465=>"110111101",
  58466=>"111000000",
  58467=>"111000011",
  58468=>"011100101",
  58469=>"011010000",
  58470=>"011000000",
  58471=>"101110100",
  58472=>"000110100",
  58473=>"111111100",
  58474=>"110111100",
  58475=>"011111111",
  58476=>"101001000",
  58477=>"001111011",
  58478=>"000000000",
  58479=>"100000100",
  58480=>"001001011",
  58481=>"011000010",
  58482=>"001111110",
  58483=>"101000111",
  58484=>"000000000",
  58485=>"000000000",
  58486=>"000110110",
  58487=>"000001111",
  58488=>"010110010",
  58489=>"011101000",
  58490=>"011001001",
  58491=>"001111100",
  58492=>"010000001",
  58493=>"110100000",
  58494=>"010111000",
  58495=>"000000000",
  58496=>"000000000",
  58497=>"000000000",
  58498=>"001000100",
  58499=>"111101111",
  58500=>"111000000",
  58501=>"011000111",
  58502=>"100100110",
  58503=>"000110010",
  58504=>"100100010",
  58505=>"000111111",
  58506=>"100111000",
  58507=>"111001000",
  58508=>"000000000",
  58509=>"000000100",
  58510=>"100000110",
  58511=>"010000000",
  58512=>"111011001",
  58513=>"010010110",
  58514=>"000000111",
  58515=>"011111010",
  58516=>"100111110",
  58517=>"101000100",
  58518=>"000011111",
  58519=>"100001001",
  58520=>"011100110",
  58521=>"000001011",
  58522=>"000110110",
  58523=>"100001000",
  58524=>"000000000",
  58525=>"010000000",
  58526=>"000000001",
  58527=>"101000111",
  58528=>"100101110",
  58529=>"001111000",
  58530=>"001111111",
  58531=>"101101111",
  58532=>"111111110",
  58533=>"101101101",
  58534=>"001101111",
  58535=>"000111111",
  58536=>"111000111",
  58537=>"100001101",
  58538=>"111101100",
  58539=>"000000000",
  58540=>"111111100",
  58541=>"110000000",
  58542=>"010111001",
  58543=>"111000010",
  58544=>"011100100",
  58545=>"111010100",
  58546=>"000000000",
  58547=>"000000100",
  58548=>"111111111",
  58549=>"101111100",
  58550=>"011010000",
  58551=>"011000000",
  58552=>"011111100",
  58553=>"000011010",
  58554=>"000000000",
  58555=>"000111100",
  58556=>"111001100",
  58557=>"100000010",
  58558=>"001100110",
  58559=>"000000000",
  58560=>"111000000",
  58561=>"000100010",
  58562=>"111110000",
  58563=>"110101100",
  58564=>"000000000",
  58565=>"111110001",
  58566=>"010000000",
  58567=>"000010000",
  58568=>"111101000",
  58569=>"000111010",
  58570=>"101110010",
  58571=>"000011011",
  58572=>"000111111",
  58573=>"111000101",
  58574=>"000010010",
  58575=>"111011000",
  58576=>"000000110",
  58577=>"000010110",
  58578=>"000010110",
  58579=>"011101111",
  58580=>"111001100",
  58581=>"010010001",
  58582=>"000011000",
  58583=>"000000101",
  58584=>"000011111",
  58585=>"011000000",
  58586=>"001101110",
  58587=>"111001000",
  58588=>"001000000",
  58589=>"100000101",
  58590=>"101000101",
  58591=>"000000000",
  58592=>"111111000",
  58593=>"111001000",
  58594=>"110100110",
  58595=>"011111111",
  58596=>"111000000",
  58597=>"100110010",
  58598=>"011000011",
  58599=>"111110000",
  58600=>"110101000",
  58601=>"000000011",
  58602=>"100110110",
  58603=>"001001000",
  58604=>"000111111",
  58605=>"110000000",
  58606=>"101000000",
  58607=>"000000000",
  58608=>"110000100",
  58609=>"011011010",
  58610=>"111001001",
  58611=>"100001101",
  58612=>"000100000",
  58613=>"001000101",
  58614=>"101000000",
  58615=>"000000000",
  58616=>"000010010",
  58617=>"100100101",
  58618=>"111100111",
  58619=>"011111101",
  58620=>"100110010",
  58621=>"111111000",
  58622=>"110100101",
  58623=>"011000000",
  58624=>"000001001",
  58625=>"101100011",
  58626=>"000000101",
  58627=>"111101111",
  58628=>"100101011",
  58629=>"110000000",
  58630=>"100001000",
  58631=>"101100000",
  58632=>"000000000",
  58633=>"000000100",
  58634=>"000110000",
  58635=>"010100011",
  58636=>"101000100",
  58637=>"000000000",
  58638=>"101100000",
  58639=>"011010000",
  58640=>"000011001",
  58641=>"110101010",
  58642=>"100000000",
  58643=>"101111101",
  58644=>"000011000",
  58645=>"000000001",
  58646=>"110001101",
  58647=>"010001000",
  58648=>"001111001",
  58649=>"000100100",
  58650=>"000010010",
  58651=>"101101110",
  58652=>"000100000",
  58653=>"000100100",
  58654=>"111011101",
  58655=>"000000000",
  58656=>"100011011",
  58657=>"000010000",
  58658=>"011000010",
  58659=>"111010000",
  58660=>"111111011",
  58661=>"101100000",
  58662=>"000111111",
  58663=>"111111111",
  58664=>"010110110",
  58665=>"000010110",
  58666=>"011000001",
  58667=>"111101000",
  58668=>"001011011",
  58669=>"011101000",
  58670=>"001101100",
  58671=>"000000000",
  58672=>"000001001",
  58673=>"000100110",
  58674=>"000000010",
  58675=>"000000111",
  58676=>"000110111",
  58677=>"110101100",
  58678=>"000010110",
  58679=>"000000000",
  58680=>"011101000",
  58681=>"101001000",
  58682=>"101100110",
  58683=>"101100111",
  58684=>"001001000",
  58685=>"010111101",
  58686=>"001101000",
  58687=>"111000000",
  58688=>"101111011",
  58689=>"010100010",
  58690=>"111111111",
  58691=>"110111111",
  58692=>"011010010",
  58693=>"000100101",
  58694=>"110111010",
  58695=>"010000001",
  58696=>"000000000",
  58697=>"000011011",
  58698=>"000010001",
  58699=>"110010111",
  58700=>"000000000",
  58701=>"100111000",
  58702=>"000101101",
  58703=>"000101000",
  58704=>"010011010",
  58705=>"110111111",
  58706=>"110111010",
  58707=>"001001001",
  58708=>"111101101",
  58709=>"100001110",
  58710=>"111111100",
  58711=>"001001100",
  58712=>"110110000",
  58713=>"101100100",
  58714=>"001001000",
  58715=>"111110100",
  58716=>"010010010",
  58717=>"011001001",
  58718=>"101100111",
  58719=>"001011111",
  58720=>"011011010",
  58721=>"010111110",
  58722=>"101101100",
  58723=>"110110000",
  58724=>"110111110",
  58725=>"010000000",
  58726=>"110110011",
  58727=>"000000000",
  58728=>"010010001",
  58729=>"000100100",
  58730=>"111011110",
  58731=>"000100000",
  58732=>"000010111",
  58733=>"010010010",
  58734=>"000000111",
  58735=>"011000000",
  58736=>"100100101",
  58737=>"111000000",
  58738=>"100110111",
  58739=>"101100111",
  58740=>"111001000",
  58741=>"100000100",
  58742=>"111110101",
  58743=>"011101111",
  58744=>"000000000",
  58745=>"111111100",
  58746=>"011000001",
  58747=>"101000100",
  58748=>"100110111",
  58749=>"000000000",
  58750=>"000001111",
  58751=>"010010010",
  58752=>"101111101",
  58753=>"100101101",
  58754=>"101101111",
  58755=>"111111100",
  58756=>"000001001",
  58757=>"111101111",
  58758=>"001100101",
  58759=>"110000000",
  58760=>"011001111",
  58761=>"010010000",
  58762=>"011111011",
  58763=>"100101111",
  58764=>"100000011",
  58765=>"000110000",
  58766=>"111000000",
  58767=>"000000000",
  58768=>"001011001",
  58769=>"110010000",
  58770=>"000001111",
  58771=>"010000001",
  58772=>"101001000",
  58773=>"100000100",
  58774=>"010110111",
  58775=>"011100110",
  58776=>"010110000",
  58777=>"101100100",
  58778=>"100100101",
  58779=>"100101000",
  58780=>"111111111",
  58781=>"111100001",
  58782=>"111000000",
  58783=>"100111000",
  58784=>"100100111",
  58785=>"100101111",
  58786=>"101100000",
  58787=>"111001000",
  58788=>"101111100",
  58789=>"010011111",
  58790=>"101001011",
  58791=>"000011010",
  58792=>"111111111",
  58793=>"111111010",
  58794=>"000101101",
  58795=>"000101111",
  58796=>"111101111",
  58797=>"111010110",
  58798=>"001111111",
  58799=>"010011010",
  58800=>"101000001",
  58801=>"011011011",
  58802=>"111101011",
  58803=>"101000001",
  58804=>"110110111",
  58805=>"011111000",
  58806=>"001011000",
  58807=>"011100000",
  58808=>"000100000",
  58809=>"110010000",
  58810=>"111000000",
  58811=>"100000001",
  58812=>"000000000",
  58813=>"001111111",
  58814=>"111001001",
  58815=>"111000000",
  58816=>"001001101",
  58817=>"111100001",
  58818=>"100000000",
  58819=>"100110100",
  58820=>"111111011",
  58821=>"100111011",
  58822=>"000101111",
  58823=>"110100100",
  58824=>"000001110",
  58825=>"100100101",
  58826=>"111111010",
  58827=>"111000101",
  58828=>"011011111",
  58829=>"001011111",
  58830=>"000000000",
  58831=>"011011001",
  58832=>"000101111",
  58833=>"111110010",
  58834=>"010010000",
  58835=>"000000010",
  58836=>"100101111",
  58837=>"110110110",
  58838=>"011011000",
  58839=>"101011011",
  58840=>"101101101",
  58841=>"010011000",
  58842=>"101001101",
  58843=>"000111000",
  58844=>"001101011",
  58845=>"001001000",
  58846=>"110111010",
  58847=>"000000100",
  58848=>"000000011",
  58849=>"010010010",
  58850=>"101001101",
  58851=>"111111100",
  58852=>"000000000",
  58853=>"000101111",
  58854=>"011111110",
  58855=>"000111111",
  58856=>"000110110",
  58857=>"000000000",
  58858=>"010011011",
  58859=>"111110010",
  58860=>"110110111",
  58861=>"011011000",
  58862=>"000000000",
  58863=>"000100100",
  58864=>"110101000",
  58865=>"001110110",
  58866=>"011000111",
  58867=>"001001001",
  58868=>"011110100",
  58869=>"111111111",
  58870=>"000000101",
  58871=>"010000100",
  58872=>"101000000",
  58873=>"000001110",
  58874=>"111101000",
  58875=>"111111011",
  58876=>"101111111",
  58877=>"111000000",
  58878=>"011110100",
  58879=>"000001000",
  58880=>"110110100",
  58881=>"000000010",
  58882=>"101000000",
  58883=>"110000010",
  58884=>"000000001",
  58885=>"111101000",
  58886=>"000000110",
  58887=>"110111111",
  58888=>"000000101",
  58889=>"000000111",
  58890=>"011001000",
  58891=>"010000010",
  58892=>"101000000",
  58893=>"001101111",
  58894=>"100100100",
  58895=>"101001010",
  58896=>"111001000",
  58897=>"111000000",
  58898=>"110101001",
  58899=>"000101011",
  58900=>"100000000",
  58901=>"000111111",
  58902=>"000100111",
  58903=>"101000100",
  58904=>"100001000",
  58905=>"001110000",
  58906=>"000000111",
  58907=>"000001101",
  58908=>"000110000",
  58909=>"011101001",
  58910=>"000001001",
  58911=>"000111010",
  58912=>"000100101",
  58913=>"000001111",
  58914=>"000111111",
  58915=>"100111110",
  58916=>"000001011",
  58917=>"000011100",
  58918=>"000010011",
  58919=>"000000000",
  58920=>"100111111",
  58921=>"111111000",
  58922=>"111000111",
  58923=>"010111011",
  58924=>"111111010",
  58925=>"111010010",
  58926=>"110110000",
  58927=>"100101000",
  58928=>"101110000",
  58929=>"000001111",
  58930=>"000000000",
  58931=>"101001111",
  58932=>"101101111",
  58933=>"111111001",
  58934=>"011001000",
  58935=>"000000000",
  58936=>"111110100",
  58937=>"000101000",
  58938=>"111111000",
  58939=>"100101100",
  58940=>"011010001",
  58941=>"011111001",
  58942=>"111000001",
  58943=>"100100010",
  58944=>"000000011",
  58945=>"000101100",
  58946=>"111000101",
  58947=>"100100000",
  58948=>"111000011",
  58949=>"100001000",
  58950=>"000110111",
  58951=>"110111011",
  58952=>"001111111",
  58953=>"011001011",
  58954=>"111101000",
  58955=>"000100001",
  58956=>"000000010",
  58957=>"100100111",
  58958=>"000000110",
  58959=>"111100000",
  58960=>"111110000",
  58961=>"110010000",
  58962=>"001111010",
  58963=>"111100001",
  58964=>"010000101",
  58965=>"000010010",
  58966=>"000101101",
  58967=>"111010000",
  58968=>"001101110",
  58969=>"011011000",
  58970=>"111011010",
  58971=>"000000000",
  58972=>"010000000",
  58973=>"000001001",
  58974=>"010000011",
  58975=>"011001001",
  58976=>"111000101",
  58977=>"001011111",
  58978=>"111000000",
  58979=>"111111001",
  58980=>"011000000",
  58981=>"011100001",
  58982=>"111001111",
  58983=>"010111000",
  58984=>"011010111",
  58985=>"010000000",
  58986=>"000000010",
  58987=>"101000011",
  58988=>"000111110",
  58989=>"111101111",
  58990=>"100101100",
  58991=>"000000001",
  58992=>"100010110",
  58993=>"000000000",
  58994=>"110101001",
  58995=>"010111001",
  58996=>"010011111",
  58997=>"101000000",
  58998=>"001000101",
  58999=>"101001011",
  59000=>"111010000",
  59001=>"010111111",
  59002=>"000000000",
  59003=>"111000111",
  59004=>"110110110",
  59005=>"011001001",
  59006=>"101111111",
  59007=>"111110101",
  59008=>"101101101",
  59009=>"111111100",
  59010=>"000000101",
  59011=>"000000000",
  59012=>"011011010",
  59013=>"111001000",
  59014=>"100100001",
  59015=>"000000000",
  59016=>"011001001",
  59017=>"001101111",
  59018=>"111010010",
  59019=>"111001000",
  59020=>"000000111",
  59021=>"111111111",
  59022=>"010001001",
  59023=>"001001000",
  59024=>"111001111",
  59025=>"000110111",
  59026=>"000100110",
  59027=>"111011101",
  59028=>"100000001",
  59029=>"101001000",
  59030=>"101000000",
  59031=>"000100001",
  59032=>"010001100",
  59033=>"100100010",
  59034=>"101110000",
  59035=>"111010010",
  59036=>"110101111",
  59037=>"111000001",
  59038=>"111111101",
  59039=>"001001001",
  59040=>"000000110",
  59041=>"000101111",
  59042=>"011001111",
  59043=>"000010000",
  59044=>"110110010",
  59045=>"101001100",
  59046=>"001000010",
  59047=>"101001111",
  59048=>"010111100",
  59049=>"101111111",
  59050=>"111100000",
  59051=>"111100000",
  59052=>"110111111",
  59053=>"111101000",
  59054=>"011011110",
  59055=>"101011111",
  59056=>"000011010",
  59057=>"110100111",
  59058=>"011001111",
  59059=>"000010010",
  59060=>"011001010",
  59061=>"111011111",
  59062=>"011111101",
  59063=>"000001111",
  59064=>"110110100",
  59065=>"000000010",
  59066=>"111111010",
  59067=>"011111111",
  59068=>"011111110",
  59069=>"111101111",
  59070=>"001001001",
  59071=>"100010010",
  59072=>"111111101",
  59073=>"000000011",
  59074=>"001001010",
  59075=>"100000101",
  59076=>"101100111",
  59077=>"010001001",
  59078=>"011010000",
  59079=>"110111100",
  59080=>"111100101",
  59081=>"111111010",
  59082=>"111111100",
  59083=>"000000111",
  59084=>"000000000",
  59085=>"011011001",
  59086=>"101111001",
  59087=>"000000000",
  59088=>"101000001",
  59089=>"011100110",
  59090=>"000000000",
  59091=>"100000000",
  59092=>"100000000",
  59093=>"001100101",
  59094=>"111110000",
  59095=>"101011000",
  59096=>"000010111",
  59097=>"000000010",
  59098=>"111001101",
  59099=>"111000111",
  59100=>"000001100",
  59101=>"111111000",
  59102=>"000000000",
  59103=>"000100110",
  59104=>"111010100",
  59105=>"111000000",
  59106=>"100011111",
  59107=>"100000110",
  59108=>"001000001",
  59109=>"111010010",
  59110=>"111101111",
  59111=>"110100101",
  59112=>"010111111",
  59113=>"000101001",
  59114=>"100100001",
  59115=>"110011011",
  59116=>"000000101",
  59117=>"000101111",
  59118=>"000001000",
  59119=>"110001111",
  59120=>"101111111",
  59121=>"100100100",
  59122=>"000000000",
  59123=>"100000110",
  59124=>"001001101",
  59125=>"110000000",
  59126=>"111000000",
  59127=>"011001001",
  59128=>"100100101",
  59129=>"111010111",
  59130=>"011011000",
  59131=>"001100110",
  59132=>"000000000",
  59133=>"000010111",
  59134=>"011000000",
  59135=>"000000101",
  59136=>"001000001",
  59137=>"110111110",
  59138=>"111000111",
  59139=>"110111111",
  59140=>"000100000",
  59141=>"011000110",
  59142=>"101111100",
  59143=>"101001111",
  59144=>"000000000",
  59145=>"111000001",
  59146=>"100110011",
  59147=>"111111000",
  59148=>"101101101",
  59149=>"100111100",
  59150=>"000001110",
  59151=>"111001111",
  59152=>"110000101",
  59153=>"111010111",
  59154=>"101000000",
  59155=>"110111111",
  59156=>"111000110",
  59157=>"100111011",
  59158=>"111101100",
  59159=>"111110111",
  59160=>"000000000",
  59161=>"111111111",
  59162=>"111111111",
  59163=>"000011000",
  59164=>"110100110",
  59165=>"000000000",
  59166=>"111111111",
  59167=>"000000000",
  59168=>"000101101",
  59169=>"101000000",
  59170=>"000000000",
  59171=>"111110100",
  59172=>"000000000",
  59173=>"000001001",
  59174=>"000111111",
  59175=>"101000000",
  59176=>"111110010",
  59177=>"000000000",
  59178=>"111111000",
  59179=>"000010110",
  59180=>"100111110",
  59181=>"111110001",
  59182=>"111101000",
  59183=>"000001010",
  59184=>"111000000",
  59185=>"000000000",
  59186=>"110000111",
  59187=>"111111111",
  59188=>"000000000",
  59189=>"111111000",
  59190=>"010000011",
  59191=>"000000000",
  59192=>"010111111",
  59193=>"000001101",
  59194=>"110000010",
  59195=>"000000100",
  59196=>"111111111",
  59197=>"111000000",
  59198=>"000011000",
  59199=>"001011111",
  59200=>"111111001",
  59201=>"000110010",
  59202=>"111111111",
  59203=>"100110010",
  59204=>"111000000",
  59205=>"100001111",
  59206=>"000111111",
  59207=>"111110010",
  59208=>"100011011",
  59209=>"111111111",
  59210=>"010000011",
  59211=>"000001000",
  59212=>"111000000",
  59213=>"000000000",
  59214=>"000000000",
  59215=>"100101101",
  59216=>"000010000",
  59217=>"111010100",
  59218=>"111100101",
  59219=>"001100110",
  59220=>"111010000",
  59221=>"111111101",
  59222=>"000010100",
  59223=>"101101101",
  59224=>"010001000",
  59225=>"000000011",
  59226=>"000001011",
  59227=>"111111111",
  59228=>"111011111",
  59229=>"000000010",
  59230=>"111111111",
  59231=>"010010111",
  59232=>"111111111",
  59233=>"101101111",
  59234=>"010000010",
  59235=>"000100110",
  59236=>"000000000",
  59237=>"111000011",
  59238=>"011111111",
  59239=>"111001011",
  59240=>"010001011",
  59241=>"111111111",
  59242=>"111111111",
  59243=>"000000111",
  59244=>"101001111",
  59245=>"010010011",
  59246=>"100000000",
  59247=>"010000110",
  59248=>"000000000",
  59249=>"110111111",
  59250=>"100000110",
  59251=>"001001111",
  59252=>"111000010",
  59253=>"000101110",
  59254=>"111111111",
  59255=>"001111001",
  59256=>"111111111",
  59257=>"011001110",
  59258=>"110000010",
  59259=>"000000000",
  59260=>"000000000",
  59261=>"000000000",
  59262=>"000000000",
  59263=>"000000000",
  59264=>"111111010",
  59265=>"111000000",
  59266=>"111111111",
  59267=>"111010000",
  59268=>"111000000",
  59269=>"000010010",
  59270=>"001100100",
  59271=>"100100100",
  59272=>"000000000",
  59273=>"000000000",
  59274=>"111111100",
  59275=>"001001111",
  59276=>"001111111",
  59277=>"000001001",
  59278=>"011111101",
  59279=>"001001001",
  59280=>"000001001",
  59281=>"000000110",
  59282=>"000101111",
  59283=>"000000101",
  59284=>"000000001",
  59285=>"111000111",
  59286=>"111100111",
  59287=>"000000000",
  59288=>"011110110",
  59289=>"110111011",
  59290=>"111110000",
  59291=>"000010010",
  59292=>"100111100",
  59293=>"111110010",
  59294=>"110111111",
  59295=>"000000111",
  59296=>"111001000",
  59297=>"011000001",
  59298=>"111001000",
  59299=>"111011111",
  59300=>"111111010",
  59301=>"000001000",
  59302=>"100111111",
  59303=>"010111111",
  59304=>"111000000",
  59305=>"000000111",
  59306=>"110000000",
  59307=>"010000010",
  59308=>"000011011",
  59309=>"010010000",
  59310=>"000000000",
  59311=>"111111111",
  59312=>"000000111",
  59313=>"000000100",
  59314=>"000000000",
  59315=>"010000010",
  59316=>"010110110",
  59317=>"110000001",
  59318=>"111111110",
  59319=>"000111100",
  59320=>"111111111",
  59321=>"001001000",
  59322=>"101111111",
  59323=>"111000001",
  59324=>"000111110",
  59325=>"111110111",
  59326=>"000110110",
  59327=>"110000000",
  59328=>"111100101",
  59329=>"010110111",
  59330=>"111000111",
  59331=>"000000000",
  59332=>"000001000",
  59333=>"001011001",
  59334=>"001100111",
  59335=>"111110010",
  59336=>"111011001",
  59337=>"000001000",
  59338=>"011001001",
  59339=>"011111111",
  59340=>"000111011",
  59341=>"110001000",
  59342=>"000000010",
  59343=>"011001111",
  59344=>"000000000",
  59345=>"000000100",
  59346=>"111111100",
  59347=>"010100001",
  59348=>"000111100",
  59349=>"000100100",
  59350=>"111101110",
  59351=>"111101111",
  59352=>"101101101",
  59353=>"110011101",
  59354=>"011000000",
  59355=>"111010000",
  59356=>"111011011",
  59357=>"110010011",
  59358=>"010101100",
  59359=>"111111101",
  59360=>"000010111",
  59361=>"111000111",
  59362=>"111001000",
  59363=>"011011010",
  59364=>"000011111",
  59365=>"010111111",
  59366=>"000101110",
  59367=>"000000000",
  59368=>"111110111",
  59369=>"111101110",
  59370=>"011011110",
  59371=>"111111111",
  59372=>"000001111",
  59373=>"111001000",
  59374=>"100000000",
  59375=>"000000111",
  59376=>"101111111",
  59377=>"111111100",
  59378=>"101001000",
  59379=>"001011110",
  59380=>"000100000",
  59381=>"000101110",
  59382=>"101001100",
  59383=>"111111010",
  59384=>"111111101",
  59385=>"000000100",
  59386=>"111010100",
  59387=>"000000000",
  59388=>"110010000",
  59389=>"100111000",
  59390=>"000000000",
  59391=>"000111110",
  59392=>"011001101",
  59393=>"000100110",
  59394=>"101101111",
  59395=>"000000010",
  59396=>"100000011",
  59397=>"000000110",
  59398=>"011111000",
  59399=>"011000100",
  59400=>"010001100",
  59401=>"101100000",
  59402=>"100101001",
  59403=>"110010000",
  59404=>"010111110",
  59405=>"010011000",
  59406=>"101111011",
  59407=>"111000001",
  59408=>"100000101",
  59409=>"000111111",
  59410=>"000000000",
  59411=>"000000000",
  59412=>"101100000",
  59413=>"101000111",
  59414=>"001011100",
  59415=>"101010001",
  59416=>"001101001",
  59417=>"000101111",
  59418=>"111100111",
  59419=>"111101100",
  59420=>"000101000",
  59421=>"000000000",
  59422=>"011010010",
  59423=>"001011000",
  59424=>"010111101",
  59425=>"010010000",
  59426=>"010100000",
  59427=>"000101111",
  59428=>"110110100",
  59429=>"001100110",
  59430=>"000000111",
  59431=>"000111010",
  59432=>"000111111",
  59433=>"011111000",
  59434=>"000010001",
  59435=>"000000101",
  59436=>"111110001",
  59437=>"000101011",
  59438=>"011000111",
  59439=>"011010111",
  59440=>"010000000",
  59441=>"000011001",
  59442=>"111111010",
  59443=>"000000110",
  59444=>"000000000",
  59445=>"100000100",
  59446=>"010100101",
  59447=>"000101111",
  59448=>"111000010",
  59449=>"000000000",
  59450=>"000111000",
  59451=>"000000000",
  59452=>"110110000",
  59453=>"111111101",
  59454=>"000000001",
  59455=>"001001110",
  59456=>"000101000",
  59457=>"101110110",
  59458=>"000111111",
  59459=>"000001000",
  59460=>"001010011",
  59461=>"100000010",
  59462=>"011110100",
  59463=>"110101101",
  59464=>"001111001",
  59465=>"011100000",
  59466=>"000010001",
  59467=>"111101111",
  59468=>"100000000",
  59469=>"011011101",
  59470=>"000100100",
  59471=>"000010111",
  59472=>"101111001",
  59473=>"111101001",
  59474=>"111000010",
  59475=>"011001010",
  59476=>"100101101",
  59477=>"000100011",
  59478=>"011011011",
  59479=>"001001111",
  59480=>"100101000",
  59481=>"001011011",
  59482=>"110000001",
  59483=>"000011001",
  59484=>"000000010",
  59485=>"001001110",
  59486=>"011011010",
  59487=>"000000001",
  59488=>"000100000",
  59489=>"010000000",
  59490=>"111100101",
  59491=>"100100111",
  59492=>"101101001",
  59493=>"010100100",
  59494=>"000000010",
  59495=>"111111000",
  59496=>"000101110",
  59497=>"101111101",
  59498=>"111110110",
  59499=>"010110100",
  59500=>"001000111",
  59501=>"011010010",
  59502=>"011010000",
  59503=>"000000000",
  59504=>"110110000",
  59505=>"000011010",
  59506=>"000000111",
  59507=>"001001000",
  59508=>"101111111",
  59509=>"000100010",
  59510=>"111111110",
  59511=>"110010000",
  59512=>"101000011",
  59513=>"101101111",
  59514=>"000011111",
  59515=>"000011000",
  59516=>"000110110",
  59517=>"110100001",
  59518=>"010010101",
  59519=>"101101101",
  59520=>"010000000",
  59521=>"110000001",
  59522=>"111010000",
  59523=>"001010111",
  59524=>"000000111",
  59525=>"111111000",
  59526=>"100000101",
  59527=>"001001001",
  59528=>"011001000",
  59529=>"110110000",
  59530=>"101000101",
  59531=>"011010000",
  59532=>"000000000",
  59533=>"101000111",
  59534=>"000010010",
  59535=>"000000101",
  59536=>"110110111",
  59537=>"001111101",
  59538=>"001000000",
  59539=>"000000001",
  59540=>"000101101",
  59541=>"001000110",
  59542=>"111110001",
  59543=>"110111100",
  59544=>"010000010",
  59545=>"000010010",
  59546=>"111100000",
  59547=>"001100111",
  59548=>"011010111",
  59549=>"010000000",
  59550=>"110010011",
  59551=>"101000111",
  59552=>"011111000",
  59553=>"111001100",
  59554=>"111110000",
  59555=>"101111111",
  59556=>"010000101",
  59557=>"000100100",
  59558=>"110110000",
  59559=>"000000111",
  59560=>"000000011",
  59561=>"000101101",
  59562=>"000100011",
  59563=>"000000001",
  59564=>"010011000",
  59565=>"000101101",
  59566=>"001000010",
  59567=>"000010111",
  59568=>"000000010",
  59569=>"000110110",
  59570=>"001000000",
  59571=>"100110100",
  59572=>"001011010",
  59573=>"111101111",
  59574=>"111000000",
  59575=>"010011000",
  59576=>"001001000",
  59577=>"000101100",
  59578=>"010010000",
  59579=>"101111111",
  59580=>"000010110",
  59581=>"110100000",
  59582=>"001000011",
  59583=>"000010010",
  59584=>"000101111",
  59585=>"001101011",
  59586=>"101111111",
  59587=>"011111111",
  59588=>"000011010",
  59589=>"010001000",
  59590=>"000000000",
  59591=>"010111100",
  59592=>"111111010",
  59593=>"101000101",
  59594=>"101011010",
  59595=>"111111010",
  59596=>"000000000",
  59597=>"000011110",
  59598=>"111111101",
  59599=>"000110011",
  59600=>"101111111",
  59601=>"100110100",
  59602=>"000010111",
  59603=>"101010000",
  59604=>"010000000",
  59605=>"110111011",
  59606=>"000000111",
  59607=>"110000100",
  59608=>"001000000",
  59609=>"001000111",
  59610=>"100111100",
  59611=>"111101111",
  59612=>"100100000",
  59613=>"000001010",
  59614=>"011101010",
  59615=>"010000000",
  59616=>"101101101",
  59617=>"010101110",
  59618=>"010010010",
  59619=>"010100111",
  59620=>"001101111",
  59621=>"000100111",
  59622=>"111000010",
  59623=>"010100010",
  59624=>"000010000",
  59625=>"111000110",
  59626=>"001000100",
  59627=>"101101101",
  59628=>"101101111",
  59629=>"010010000",
  59630=>"101000000",
  59631=>"000001101",
  59632=>"101000111",
  59633=>"110101100",
  59634=>"000010111",
  59635=>"100110110",
  59636=>"010111010",
  59637=>"111111111",
  59638=>"000010000",
  59639=>"000010011",
  59640=>"000010010",
  59641=>"010010001",
  59642=>"000001000",
  59643=>"100001011",
  59644=>"111011000",
  59645=>"000000111",
  59646=>"011011011",
  59647=>"000000111",
  59648=>"111111011",
  59649=>"000000000",
  59650=>"000000101",
  59651=>"010010000",
  59652=>"111100100",
  59653=>"101000110",
  59654=>"111101101",
  59655=>"000110011",
  59656=>"011001000",
  59657=>"000000001",
  59658=>"001000000",
  59659=>"101101000",
  59660=>"000010000",
  59661=>"001000000",
  59662=>"011111011",
  59663=>"101111010",
  59664=>"000111000",
  59665=>"111000000",
  59666=>"100000000",
  59667=>"000001011",
  59668=>"100000000",
  59669=>"000000100",
  59670=>"111000000",
  59671=>"111111110",
  59672=>"000111110",
  59673=>"111001101",
  59674=>"100000000",
  59675=>"011000000",
  59676=>"000111000",
  59677=>"010000000",
  59678=>"111111010",
  59679=>"111110000",
  59680=>"010101000",
  59681=>"110101010",
  59682=>"111101000",
  59683=>"000010000",
  59684=>"100000000",
  59685=>"111010000",
  59686=>"000010110",
  59687=>"001011100",
  59688=>"000001000",
  59689=>"111001001",
  59690=>"001011001",
  59691=>"111111111",
  59692=>"001111001",
  59693=>"101001111",
  59694=>"111111001",
  59695=>"111001111",
  59696=>"110000000",
  59697=>"010100100",
  59698=>"100110100",
  59699=>"100111010",
  59700=>"001001111",
  59701=>"001011110",
  59702=>"110000001",
  59703=>"000010000",
  59704=>"110101000",
  59705=>"001001000",
  59706=>"100100101",
  59707=>"001001010",
  59708=>"100010100",
  59709=>"010101101",
  59710=>"000000000",
  59711=>"011000000",
  59712=>"001110111",
  59713=>"011010000",
  59714=>"000111111",
  59715=>"001001001",
  59716=>"000000111",
  59717=>"010000100",
  59718=>"001000001",
  59719=>"110010111",
  59720=>"010100100",
  59721=>"010010010",
  59722=>"001101001",
  59723=>"000001111",
  59724=>"001111010",
  59725=>"100100110",
  59726=>"001011011",
  59727=>"100111111",
  59728=>"110010000",
  59729=>"111000010",
  59730=>"000010000",
  59731=>"011001110",
  59732=>"000000111",
  59733=>"100011100",
  59734=>"011011000",
  59735=>"000101100",
  59736=>"001000000",
  59737=>"001101000",
  59738=>"111011000",
  59739=>"011101100",
  59740=>"110111000",
  59741=>"001101000",
  59742=>"000000101",
  59743=>"100100000",
  59744=>"000010110",
  59745=>"110000000",
  59746=>"000010111",
  59747=>"100001011",
  59748=>"100111100",
  59749=>"111110110",
  59750=>"001000110",
  59751=>"000000000",
  59752=>"100111111",
  59753=>"111111111",
  59754=>"000000111",
  59755=>"111101111",
  59756=>"111100000",
  59757=>"111111011",
  59758=>"001000000",
  59759=>"111111000",
  59760=>"100011001",
  59761=>"111111000",
  59762=>"001000110",
  59763=>"110111111",
  59764=>"000111111",
  59765=>"000000100",
  59766=>"000110111",
  59767=>"001000100",
  59768=>"101010010",
  59769=>"000111111",
  59770=>"110000000",
  59771=>"101000001",
  59772=>"000100110",
  59773=>"100100010",
  59774=>"010111111",
  59775=>"111000110",
  59776=>"010111011",
  59777=>"111101000",
  59778=>"111000000",
  59779=>"111110011",
  59780=>"000111111",
  59781=>"000001011",
  59782=>"110011000",
  59783=>"000110000",
  59784=>"101100101",
  59785=>"010110100",
  59786=>"110100100",
  59787=>"101100111",
  59788=>"001000001",
  59789=>"111101111",
  59790=>"111110000",
  59791=>"110001001",
  59792=>"101011000",
  59793=>"010111000",
  59794=>"001001011",
  59795=>"000010010",
  59796=>"000011111",
  59797=>"000111010",
  59798=>"110111011",
  59799=>"111110100",
  59800=>"110111000",
  59801=>"000000010",
  59802=>"110111111",
  59803=>"000000000",
  59804=>"110000000",
  59805=>"000111111",
  59806=>"111110000",
  59807=>"000110111",
  59808=>"000010000",
  59809=>"111111010",
  59810=>"001000101",
  59811=>"101111111",
  59812=>"001011001",
  59813=>"011011011",
  59814=>"100001011",
  59815=>"001110110",
  59816=>"111100101",
  59817=>"001100111",
  59818=>"111100000",
  59819=>"110000000",
  59820=>"111111111",
  59821=>"011111110",
  59822=>"010110011",
  59823=>"010110111",
  59824=>"010000000",
  59825=>"011001111",
  59826=>"011000000",
  59827=>"001001000",
  59828=>"000110110",
  59829=>"000100111",
  59830=>"100001101",
  59831=>"010110100",
  59832=>"001010001",
  59833=>"000110111",
  59834=>"110110101",
  59835=>"101001101",
  59836=>"010111010",
  59837=>"000100111",
  59838=>"111100100",
  59839=>"101001101",
  59840=>"001000101",
  59841=>"000000000",
  59842=>"010000110",
  59843=>"000000100",
  59844=>"010010111",
  59845=>"111111011",
  59846=>"111111000",
  59847=>"000001101",
  59848=>"101111101",
  59849=>"000001111",
  59850=>"110111111",
  59851=>"010000101",
  59852=>"101000010",
  59853=>"001011011",
  59854=>"011001010",
  59855=>"110011111",
  59856=>"000000000",
  59857=>"110011111",
  59858=>"000010001",
  59859=>"111111110",
  59860=>"000100111",
  59861=>"010100110",
  59862=>"000000000",
  59863=>"000000111",
  59864=>"101111001",
  59865=>"000000000",
  59866=>"000110100",
  59867=>"001110000",
  59868=>"011001000",
  59869=>"100100011",
  59870=>"000000000",
  59871=>"001000000",
  59872=>"000000000",
  59873=>"110000000",
  59874=>"010010000",
  59875=>"011111100",
  59876=>"000001111",
  59877=>"011000001",
  59878=>"111000000",
  59879=>"011011101",
  59880=>"000000010",
  59881=>"100101111",
  59882=>"000000011",
  59883=>"111111111",
  59884=>"000001000",
  59885=>"110101111",
  59886=>"000000000",
  59887=>"100100000",
  59888=>"000000010",
  59889=>"011111100",
  59890=>"111100000",
  59891=>"001011011",
  59892=>"110110111",
  59893=>"011101000",
  59894=>"001000011",
  59895=>"010011010",
  59896=>"111000000",
  59897=>"111000000",
  59898=>"111100100",
  59899=>"000111111",
  59900=>"111111111",
  59901=>"111100101",
  59902=>"001001001",
  59903=>"000110111",
  59904=>"100000010",
  59905=>"110000010",
  59906=>"001010000",
  59907=>"000000000",
  59908=>"100000111",
  59909=>"001111000",
  59910=>"011110000",
  59911=>"101101000",
  59912=>"110110101",
  59913=>"000010010",
  59914=>"110111011",
  59915=>"111000000",
  59916=>"000000001",
  59917=>"000000000",
  59918=>"011111001",
  59919=>"111110110",
  59920=>"101111110",
  59921=>"010111110",
  59922=>"000100000",
  59923=>"000010111",
  59924=>"001101011",
  59925=>"000001111",
  59926=>"010011011",
  59927=>"000111111",
  59928=>"011101010",
  59929=>"000000110",
  59930=>"000101111",
  59931=>"000000001",
  59932=>"011110111",
  59933=>"000111001",
  59934=>"011000000",
  59935=>"110111100",
  59936=>"000000101",
  59937=>"000000010",
  59938=>"010010110",
  59939=>"000000001",
  59940=>"010110110",
  59941=>"000001000",
  59942=>"001001111",
  59943=>"001111101",
  59944=>"000111111",
  59945=>"111110000",
  59946=>"000010010",
  59947=>"010000000",
  59948=>"111111001",
  59949=>"101111111",
  59950=>"000101101",
  59951=>"000000110",
  59952=>"100111110",
  59953=>"100000011",
  59954=>"111000010",
  59955=>"010110111",
  59956=>"000001111",
  59957=>"000111111",
  59958=>"000111010",
  59959=>"000000111",
  59960=>"110111001",
  59961=>"000101111",
  59962=>"101111101",
  59963=>"010010110",
  59964=>"110101111",
  59965=>"111111010",
  59966=>"100110000",
  59967=>"110100011",
  59968=>"111111111",
  59969=>"110000001",
  59970=>"001111100",
  59971=>"100000111",
  59972=>"111000000",
  59973=>"111111101",
  59974=>"011010000",
  59975=>"000000000",
  59976=>"001011011",
  59977=>"000000001",
  59978=>"111001000",
  59979=>"100111111",
  59980=>"111110000",
  59981=>"011011111",
  59982=>"111000100",
  59983=>"111001001",
  59984=>"010110010",
  59985=>"010000000",
  59986=>"010111001",
  59987=>"000000101",
  59988=>"001110110",
  59989=>"111000000",
  59990=>"000100000",
  59991=>"110000000",
  59992=>"111001000",
  59993=>"100110000",
  59994=>"111111000",
  59995=>"111110111",
  59996=>"000000000",
  59997=>"100000001",
  59998=>"000000110",
  59999=>"011001110",
  60000=>"010000101",
  60001=>"010000000",
  60002=>"111001000",
  60003=>"111011101",
  60004=>"010101101",
  60005=>"011111100",
  60006=>"000001111",
  60007=>"010101111",
  60008=>"001010010",
  60009=>"011101101",
  60010=>"110111011",
  60011=>"000101000",
  60012=>"001001000",
  60013=>"110011101",
  60014=>"111111000",
  60015=>"110000001",
  60016=>"101000110",
  60017=>"001111001",
  60018=>"001111011",
  60019=>"110000000",
  60020=>"101101111",
  60021=>"101101101",
  60022=>"111110010",
  60023=>"111111111",
  60024=>"000000101",
  60025=>"010000000",
  60026=>"111111000",
  60027=>"000000111",
  60028=>"100101101",
  60029=>"000100101",
  60030=>"011000100",
  60031=>"110000000",
  60032=>"110100110",
  60033=>"010010001",
  60034=>"010100001",
  60035=>"000000101",
  60036=>"101001101",
  60037=>"111111011",
  60038=>"001100100",
  60039=>"100011001",
  60040=>"101001001",
  60041=>"010101110",
  60042=>"010000000",
  60043=>"111000101",
  60044=>"001000111",
  60045=>"010000000",
  60046=>"111000101",
  60047=>"111100100",
  60048=>"100100011",
  60049=>"000111111",
  60050=>"000000010",
  60051=>"101001001",
  60052=>"001000010",
  60053=>"110111000",
  60054=>"111110010",
  60055=>"111111000",
  60056=>"110110000",
  60057=>"010000010",
  60058=>"001000111",
  60059=>"100000100",
  60060=>"111110001",
  60061=>"110000000",
  60062=>"111000111",
  60063=>"011001000",
  60064=>"100111001",
  60065=>"111111000",
  60066=>"110000000",
  60067=>"011011010",
  60068=>"000111010",
  60069=>"001011110",
  60070=>"001111111",
  60071=>"111111000",
  60072=>"010111111",
  60073=>"000000001",
  60074=>"000111110",
  60075=>"001110000",
  60076=>"011111110",
  60077=>"110111000",
  60078=>"010100000",
  60079=>"111000000",
  60080=>"011000001",
  60081=>"110110010",
  60082=>"000001000",
  60083=>"111000000",
  60084=>"011001001",
  60085=>"000111010",
  60086=>"000100100",
  60087=>"000010000",
  60088=>"011011000",
  60089=>"100000010",
  60090=>"000000000",
  60091=>"100001000",
  60092=>"101101111",
  60093=>"111000111",
  60094=>"011111101",
  60095=>"000000101",
  60096=>"000101111",
  60097=>"111111010",
  60098=>"000011101",
  60099=>"001011000",
  60100=>"111001111",
  60101=>"111001000",
  60102=>"111111000",
  60103=>"011000010",
  60104=>"000011111",
  60105=>"001000001",
  60106=>"000001011",
  60107=>"000111111",
  60108=>"000000000",
  60109=>"011010011",
  60110=>"101010000",
  60111=>"001100000",
  60112=>"110010000",
  60113=>"101000110",
  60114=>"001000000",
  60115=>"110100010",
  60116=>"001001101",
  60117=>"001011110",
  60118=>"111101000",
  60119=>"010001000",
  60120=>"000101111",
  60121=>"101001111",
  60122=>"011010111",
  60123=>"101111110",
  60124=>"110110000",
  60125=>"001000000",
  60126=>"101101101",
  60127=>"110101001",
  60128=>"011100100",
  60129=>"011111101",
  60130=>"010000101",
  60131=>"000110111",
  60132=>"000000000",
  60133=>"010000011",
  60134=>"001101111",
  60135=>"100010000",
  60136=>"001111000",
  60137=>"101101010",
  60138=>"111101110",
  60139=>"110111111",
  60140=>"101111101",
  60141=>"101000111",
  60142=>"000000000",
  60143=>"111001101",
  60144=>"001000010",
  60145=>"011000000",
  60146=>"011111101",
  60147=>"100000111",
  60148=>"011000100",
  60149=>"101101000",
  60150=>"111000000",
  60151=>"000100100",
  60152=>"001100110",
  60153=>"001111111",
  60154=>"110110000",
  60155=>"000111101",
  60156=>"000111111",
  60157=>"010000000",
  60158=>"111101100",
  60159=>"010001001",
  60160=>"011011001",
  60161=>"111000000",
  60162=>"101000101",
  60163=>"110000110",
  60164=>"100111111",
  60165=>"010000000",
  60166=>"000000101",
  60167=>"111111000",
  60168=>"110000001",
  60169=>"000000101",
  60170=>"101000010",
  60171=>"110110110",
  60172=>"000000000",
  60173=>"000110110",
  60174=>"100110010",
  60175=>"111001000",
  60176=>"111110100",
  60177=>"111001000",
  60178=>"110111110",
  60179=>"110000000",
  60180=>"100000001",
  60181=>"000000001",
  60182=>"000001111",
  60183=>"111000000",
  60184=>"000001001",
  60185=>"000110000",
  60186=>"000110010",
  60187=>"000010101",
  60188=>"000101110",
  60189=>"000101010",
  60190=>"010011011",
  60191=>"010010011",
  60192=>"000110111",
  60193=>"100110110",
  60194=>"000000000",
  60195=>"101000111",
  60196=>"101100100",
  60197=>"010110100",
  60198=>"010111000",
  60199=>"100110110",
  60200=>"111111000",
  60201=>"001001000",
  60202=>"011000111",
  60203=>"000011010",
  60204=>"001100000",
  60205=>"100110101",
  60206=>"111000001",
  60207=>"111010111",
  60208=>"000000000",
  60209=>"001111011",
  60210=>"110111111",
  60211=>"111001000",
  60212=>"000000100",
  60213=>"000000000",
  60214=>"000000001",
  60215=>"111001101",
  60216=>"001000001",
  60217=>"000000000",
  60218=>"101001101",
  60219=>"000000000",
  60220=>"110110110",
  60221=>"100111111",
  60222=>"000000000",
  60223=>"010110110",
  60224=>"000001001",
  60225=>"111111101",
  60226=>"101000001",
  60227=>"100111011",
  60228=>"101001111",
  60229=>"010110110",
  60230=>"010101110",
  60231=>"000110010",
  60232=>"010111110",
  60233=>"000110010",
  60234=>"111110111",
  60235=>"111111111",
  60236=>"110000111",
  60237=>"101001001",
  60238=>"100101100",
  60239=>"111101000",
  60240=>"101110111",
  60241=>"111111111",
  60242=>"111011111",
  60243=>"011011001",
  60244=>"001000000",
  60245=>"110010110",
  60246=>"011011011",
  60247=>"001111001",
  60248=>"100110110",
  60249=>"001111011",
  60250=>"001011111",
  60251=>"110110111",
  60252=>"101001001",
  60253=>"000000011",
  60254=>"001001001",
  60255=>"110111101",
  60256=>"000000000",
  60257=>"000110010",
  60258=>"101000101",
  60259=>"000100110",
  60260=>"111111110",
  60261=>"101000000",
  60262=>"110110000",
  60263=>"001001101",
  60264=>"000101111",
  60265=>"111111000",
  60266=>"111001111",
  60267=>"110111111",
  60268=>"001111011",
  60269=>"001001001",
  60270=>"000000000",
  60271=>"000000111",
  60272=>"000100100",
  60273=>"011011111",
  60274=>"001001100",
  60275=>"000101111",
  60276=>"001000111",
  60277=>"000000000",
  60278=>"001000111",
  60279=>"000111001",
  60280=>"000000000",
  60281=>"000001011",
  60282=>"111111111",
  60283=>"000000000",
  60284=>"100101110",
  60285=>"010100000",
  60286=>"010110110",
  60287=>"110110110",
  60288=>"010010100",
  60289=>"110110000",
  60290=>"111000101",
  60291=>"000000101",
  60292=>"111110000",
  60293=>"000000101",
  60294=>"000010011",
  60295=>"000100010",
  60296=>"100001001",
  60297=>"000011010",
  60298=>"000100100",
  60299=>"110010000",
  60300=>"001000001",
  60301=>"000001000",
  60302=>"000000101",
  60303=>"000000000",
  60304=>"000000100",
  60305=>"000111000",
  60306=>"111110000",
  60307=>"000100110",
  60308=>"100111110",
  60309=>"111000001",
  60310=>"111001001",
  60311=>"000000010",
  60312=>"010111110",
  60313=>"111011001",
  60314=>"010111110",
  60315=>"000000000",
  60316=>"011101101",
  60317=>"001111011",
  60318=>"000001100",
  60319=>"111001101",
  60320=>"110110010",
  60321=>"010000000",
  60322=>"000001111",
  60323=>"111001000",
  60324=>"001000010",
  60325=>"011001010",
  60326=>"001111010",
  60327=>"100100100",
  60328=>"011111000",
  60329=>"111111010",
  60330=>"010000110",
  60331=>"111000000",
  60332=>"111111101",
  60333=>"000000101",
  60334=>"100101011",
  60335=>"011000001",
  60336=>"001000000",
  60337=>"011010100",
  60338=>"000101110",
  60339=>"010000111",
  60340=>"110101110",
  60341=>"101001001",
  60342=>"000110110",
  60343=>"000111111",
  60344=>"010011011",
  60345=>"001111111",
  60346=>"110111111",
  60347=>"000000110",
  60348=>"000100000",
  60349=>"110110000",
  60350=>"010001000",
  60351=>"000001101",
  60352=>"111000000",
  60353=>"000000111",
  60354=>"111111110",
  60355=>"001100100",
  60356=>"001000000",
  60357=>"110111101",
  60358=>"111101111",
  60359=>"010000001",
  60360=>"000000010",
  60361=>"010000000",
  60362=>"000001101",
  60363=>"101000000",
  60364=>"010010000",
  60365=>"001111110",
  60366=>"001101101",
  60367=>"000111111",
  60368=>"100010000",
  60369=>"000110100",
  60370=>"110111111",
  60371=>"001001000",
  60372=>"110110000",
  60373=>"001000000",
  60374=>"110001000",
  60375=>"000000111",
  60376=>"001001001",
  60377=>"010010000",
  60378=>"000011100",
  60379=>"101001001",
  60380=>"010100010",
  60381=>"001011011",
  60382=>"110111110",
  60383=>"111110101",
  60384=>"111000000",
  60385=>"101011101",
  60386=>"000111110",
  60387=>"001101000",
  60388=>"101000000",
  60389=>"101001001",
  60390=>"101001110",
  60391=>"000010000",
  60392=>"000000100",
  60393=>"000000101",
  60394=>"001000010",
  60395=>"001001111",
  60396=>"000010000",
  60397=>"001000000",
  60398=>"000101000",
  60399=>"010110110",
  60400=>"111000001",
  60401=>"101110010",
  60402=>"010000111",
  60403=>"100100110",
  60404=>"110110011",
  60405=>"000000011",
  60406=>"010110000",
  60407=>"000111111",
  60408=>"000111110",
  60409=>"111101000",
  60410=>"111111111",
  60411=>"000111111",
  60412=>"000100111",
  60413=>"001000010",
  60414=>"001111110",
  60415=>"111100111",
  60416=>"001000100",
  60417=>"101110000",
  60418=>"100000101",
  60419=>"011111000",
  60420=>"011001000",
  60421=>"000101100",
  60422=>"000000000",
  60423=>"001000111",
  60424=>"111110111",
  60425=>"000000111",
  60426=>"111011110",
  60427=>"000101100",
  60428=>"111010010",
  60429=>"111010010",
  60430=>"011011000",
  60431=>"111101111",
  60432=>"110010010",
  60433=>"000101000",
  60434=>"000101110",
  60435=>"100000011",
  60436=>"100000000",
  60437=>"000111111",
  60438=>"111100100",
  60439=>"010111110",
  60440=>"100000000",
  60441=>"110000110",
  60442=>"001000101",
  60443=>"111010110",
  60444=>"000000111",
  60445=>"101111000",
  60446=>"000001010",
  60447=>"111000000",
  60448=>"000000000",
  60449=>"111111010",
  60450=>"001101010",
  60451=>"000000000",
  60452=>"010001001",
  60453=>"100101001",
  60454=>"011110100",
  60455=>"000011101",
  60456=>"100110100",
  60457=>"000010111",
  60458=>"101000001",
  60459=>"000000010",
  60460=>"000101001",
  60461=>"000100000",
  60462=>"010100010",
  60463=>"010001000",
  60464=>"111111000",
  60465=>"001001001",
  60466=>"000111111",
  60467=>"101110110",
  60468=>"100100100",
  60469=>"010110110",
  60470=>"010110001",
  60471=>"101000000",
  60472=>"101000110",
  60473=>"101101111",
  60474=>"101101000",
  60475=>"111011111",
  60476=>"100100011",
  60477=>"011000011",
  60478=>"000000000",
  60479=>"000100100",
  60480=>"111111111",
  60481=>"000101000",
  60482=>"111111010",
  60483=>"100100000",
  60484=>"101111000",
  60485=>"000000000",
  60486=>"111101000",
  60487=>"010100000",
  60488=>"011111111",
  60489=>"111111111",
  60490=>"000101100",
  60491=>"000000001",
  60492=>"000000001",
  60493=>"010101111",
  60494=>"000001100",
  60495=>"101100110",
  60496=>"001111000",
  60497=>"010111110",
  60498=>"111111000",
  60499=>"110000000",
  60500=>"010000100",
  60501=>"000010111",
  60502=>"111001100",
  60503=>"000000111",
  60504=>"111111111",
  60505=>"111100001",
  60506=>"100000000",
  60507=>"111100100",
  60508=>"000000000",
  60509=>"001011010",
  60510=>"011000111",
  60511=>"001001000",
  60512=>"010010000",
  60513=>"010010010",
  60514=>"000000111",
  60515=>"001000000",
  60516=>"110010000",
  60517=>"111100111",
  60518=>"101110110",
  60519=>"111000101",
  60520=>"111111000",
  60521=>"000111111",
  60522=>"101000011",
  60523=>"111111111",
  60524=>"000011110",
  60525=>"111111011",
  60526=>"010000111",
  60527=>"000100000",
  60528=>"001000000",
  60529=>"101101010",
  60530=>"010011100",
  60531=>"111101000",
  60532=>"000111111",
  60533=>"101101111",
  60534=>"101001000",
  60535=>"111011001",
  60536=>"111000000",
  60537=>"001010000",
  60538=>"001000001",
  60539=>"000111111",
  60540=>"111000000",
  60541=>"010100000",
  60542=>"000001111",
  60543=>"010010001",
  60544=>"111111110",
  60545=>"001001111",
  60546=>"000100000",
  60547=>"011010010",
  60548=>"000010010",
  60549=>"111001000",
  60550=>"000110000",
  60551=>"111001011",
  60552=>"000001100",
  60553=>"001111001",
  60554=>"100000000",
  60555=>"011000100",
  60556=>"110010001",
  60557=>"111111101",
  60558=>"011111100",
  60559=>"110100000",
  60560=>"110100100",
  60561=>"001001000",
  60562=>"010001111",
  60563=>"111000000",
  60564=>"001010000",
  60565=>"101000111",
  60566=>"101101101",
  60567=>"011000000",
  60568=>"010000111",
  60569=>"000000111",
  60570=>"000001111",
  60571=>"110111010",
  60572=>"001001111",
  60573=>"000111000",
  60574=>"000001111",
  60575=>"101101101",
  60576=>"111110011",
  60577=>"100101000",
  60578=>"111010000",
  60579=>"001000111",
  60580=>"000111110",
  60581=>"111001001",
  60582=>"100000001",
  60583=>"000111110",
  60584=>"010111111",
  60585=>"111000000",
  60586=>"111101111",
  60587=>"001000000",
  60588=>"111010000",
  60589=>"111010000",
  60590=>"001000000",
  60591=>"011010000",
  60592=>"001100110",
  60593=>"011011110",
  60594=>"100100000",
  60595=>"100000100",
  60596=>"001001011",
  60597=>"000000110",
  60598=>"000110000",
  60599=>"110000111",
  60600=>"011010010",
  60601=>"111000110",
  60602=>"010000000",
  60603=>"000100000",
  60604=>"000000000",
  60605=>"111111000",
  60606=>"111011000",
  60607=>"001101111",
  60608=>"000000111",
  60609=>"001010111",
  60610=>"111111000",
  60611=>"011100000",
  60612=>"011010010",
  60613=>"000010000",
  60614=>"111101011",
  60615=>"000000100",
  60616=>"001000111",
  60617=>"000000000",
  60618=>"111100100",
  60619=>"000101101",
  60620=>"111111101",
  60621=>"111000000",
  60622=>"000000000",
  60623=>"010100000",
  60624=>"111010111",
  60625=>"110110100",
  60626=>"111111010",
  60627=>"111101111",
  60628=>"100000111",
  60629=>"100111000",
  60630=>"000000000",
  60631=>"001111010",
  60632=>"000000101",
  60633=>"110010000",
  60634=>"111111111",
  60635=>"000100010",
  60636=>"101001011",
  60637=>"111111110",
  60638=>"000010001",
  60639=>"001101101",
  60640=>"111010010",
  60641=>"100010110",
  60642=>"111011001",
  60643=>"111111001",
  60644=>"000000101",
  60645=>"000010010",
  60646=>"010010110",
  60647=>"001011111",
  60648=>"000000010",
  60649=>"000000000",
  60650=>"001101111",
  60651=>"111100000",
  60652=>"000010000",
  60653=>"100001001",
  60654=>"000000000",
  60655=>"100000000",
  60656=>"001000000",
  60657=>"001010000",
  60658=>"000001011",
  60659=>"110100000",
  60660=>"101000011",
  60661=>"111111001",
  60662=>"000000010",
  60663=>"000000110",
  60664=>"001000000",
  60665=>"101111110",
  60666=>"111110000",
  60667=>"001010000",
  60668=>"111111111",
  60669=>"001000001",
  60670=>"110001001",
  60671=>"111101000",
  60672=>"100011011",
  60673=>"000100110",
  60674=>"001000001",
  60675=>"000000110",
  60676=>"100110100",
  60677=>"001001001",
  60678=>"111110111",
  60679=>"000110110",
  60680=>"110000000",
  60681=>"011001011",
  60682=>"000100101",
  60683=>"000000001",
  60684=>"000000101",
  60685=>"110110000",
  60686=>"000010100",
  60687=>"111111001",
  60688=>"000100100",
  60689=>"001100110",
  60690=>"011001000",
  60691=>"111100110",
  60692=>"001001101",
  60693=>"001001111",
  60694=>"001011011",
  60695=>"100110110",
  60696=>"011001001",
  60697=>"111111011",
  60698=>"111111110",
  60699=>"000111101",
  60700=>"000111011",
  60701=>"110110100",
  60702=>"001011100",
  60703=>"000010110",
  60704=>"001001001",
  60705=>"000001001",
  60706=>"000000100",
  60707=>"000000100",
  60708=>"001001001",
  60709=>"100100010",
  60710=>"101100110",
  60711=>"110110000",
  60712=>"011010010",
  60713=>"000000000",
  60714=>"000110100",
  60715=>"110000010",
  60716=>"100101110",
  60717=>"011011101",
  60718=>"100001011",
  60719=>"111011100",
  60720=>"110011011",
  60721=>"110111011",
  60722=>"011111001",
  60723=>"011001000",
  60724=>"100110110",
  60725=>"100100100",
  60726=>"000000110",
  60727=>"100110100",
  60728=>"010011001",
  60729=>"000000110",
  60730=>"011001000",
  60731=>"100100101",
  60732=>"000100000",
  60733=>"000111010",
  60734=>"001001000",
  60735=>"100010100",
  60736=>"111001101",
  60737=>"100100110",
  60738=>"001111111",
  60739=>"100110011",
  60740=>"010001010",
  60741=>"100000000",
  60742=>"111111001",
  60743=>"011011010",
  60744=>"110011010",
  60745=>"010011001",
  60746=>"001100111",
  60747=>"111100111",
  60748=>"111001100",
  60749=>"000011011",
  60750=>"000001001",
  60751=>"111010010",
  60752=>"000000010",
  60753=>"110111111",
  60754=>"011011011",
  60755=>"110011001",
  60756=>"001001011",
  60757=>"000111001",
  60758=>"000001100",
  60759=>"011000000",
  60760=>"011111111",
  60761=>"101011011",
  60762=>"000000001",
  60763=>"111111101",
  60764=>"000010010",
  60765=>"110011011",
  60766=>"100110100",
  60767=>"111100000",
  60768=>"110000011",
  60769=>"100000110",
  60770=>"011001101",
  60771=>"001111111",
  60772=>"110010000",
  60773=>"110110000",
  60774=>"000000010",
  60775=>"000110100",
  60776=>"000001111",
  60777=>"011011111",
  60778=>"110000000",
  60779=>"101001111",
  60780=>"011001111",
  60781=>"101100100",
  60782=>"000000000",
  60783=>"000011111",
  60784=>"100011001",
  60785=>"010110110",
  60786=>"010000101",
  60787=>"001000100",
  60788=>"111111010",
  60789=>"011001100",
  60790=>"011000111",
  60791=>"110000011",
  60792=>"011111001",
  60793=>"001111110",
  60794=>"111111011",
  60795=>"110011011",
  60796=>"000100110",
  60797=>"100000000",
  60798=>"111110010",
  60799=>"001000001",
  60800=>"100000111",
  60801=>"011001000",
  60802=>"001001000",
  60803=>"100000000",
  60804=>"001110100",
  60805=>"101001101",
  60806=>"100101111",
  60807=>"000000001",
  60808=>"000000000",
  60809=>"100110010",
  60810=>"111011001",
  60811=>"110001001",
  60812=>"000100110",
  60813=>"001001011",
  60814=>"011111000",
  60815=>"000000000",
  60816=>"111011001",
  60817=>"000100100",
  60818=>"110110011",
  60819=>"000110010",
  60820=>"010100010",
  60821=>"001001100",
  60822=>"000100100",
  60823=>"110100100",
  60824=>"110010000",
  60825=>"011011001",
  60826=>"001011110",
  60827=>"011011000",
  60828=>"100110111",
  60829=>"111001111",
  60830=>"110110010",
  60831=>"000100100",
  60832=>"011011001",
  60833=>"001101111",
  60834=>"100011011",
  60835=>"000011010",
  60836=>"011011111",
  60837=>"000000000",
  60838=>"101001100",
  60839=>"100100100",
  60840=>"101001110",
  60841=>"011001011",
  60842=>"011001001",
  60843=>"001000100",
  60844=>"000001000",
  60845=>"110010011",
  60846=>"000100100",
  60847=>"000011111",
  60848=>"000000010",
  60849=>"111110000",
  60850=>"110011011",
  60851=>"000001000",
  60852=>"110111101",
  60853=>"010101000",
  60854=>"000101011",
  60855=>"110010010",
  60856=>"110101111",
  60857=>"100100000",
  60858=>"110010111",
  60859=>"011011011",
  60860=>"001110010",
  60861=>"011101001",
  60862=>"010000011",
  60863=>"000100111",
  60864=>"011001001",
  60865=>"000000010",
  60866=>"001101110",
  60867=>"110011011",
  60868=>"100010000",
  60869=>"010011011",
  60870=>"110111111",
  60871=>"011101111",
  60872=>"110010011",
  60873=>"000100110",
  60874=>"011001000",
  60875=>"000100001",
  60876=>"100110010",
  60877=>"010000100",
  60878=>"000100000",
  60879=>"111101000",
  60880=>"000100000",
  60881=>"100010100",
  60882=>"001100011",
  60883=>"111111000",
  60884=>"100101001",
  60885=>"001000001",
  60886=>"000010001",
  60887=>"100101111",
  60888=>"100110110",
  60889=>"110100100",
  60890=>"000001001",
  60891=>"011001101",
  60892=>"000010000",
  60893=>"001101011",
  60894=>"000101111",
  60895=>"100011000",
  60896=>"000100000",
  60897=>"001001000",
  60898=>"100110110",
  60899=>"111001001",
  60900=>"001000011",
  60901=>"111011011",
  60902=>"100110110",
  60903=>"110111011",
  60904=>"111111100",
  60905=>"100110101",
  60906=>"101110010",
  60907=>"011001001",
  60908=>"100100100",
  60909=>"100110110",
  60910=>"000000001",
  60911=>"100010010",
  60912=>"100110110",
  60913=>"111011011",
  60914=>"000111000",
  60915=>"100010000",
  60916=>"101101001",
  60917=>"011000001",
  60918=>"101000000",
  60919=>"010110010",
  60920=>"000100110",
  60921=>"000110110",
  60922=>"111001111",
  60923=>"110111001",
  60924=>"001111011",
  60925=>"000001010",
  60926=>"111001001",
  60927=>"100110010",
  60928=>"100000110",
  60929=>"000000001",
  60930=>"011000001",
  60931=>"111111111",
  60932=>"101101001",
  60933=>"100001000",
  60934=>"000111111",
  60935=>"111001110",
  60936=>"000000000",
  60937=>"000000000",
  60938=>"100100100",
  60939=>"000000111",
  60940=>"000000111",
  60941=>"111010111",
  60942=>"100000100",
  60943=>"100000000",
  60944=>"001001001",
  60945=>"000000000",
  60946=>"000000000",
  60947=>"000000000",
  60948=>"001000011",
  60949=>"111001111",
  60950=>"101001001",
  60951=>"000000100",
  60952=>"001000000",
  60953=>"111111010",
  60954=>"100001000",
  60955=>"000001000",
  60956=>"110101001",
  60957=>"111101100",
  60958=>"000001000",
  60959=>"110010010",
  60960=>"001001000",
  60961=>"111101111",
  60962=>"110011111",
  60963=>"000001010",
  60964=>"111111111",
  60965=>"000000011",
  60966=>"001100001",
  60967=>"000001111",
  60968=>"111101000",
  60969=>"110100000",
  60970=>"000000010",
  60971=>"011010001",
  60972=>"101000100",
  60973=>"000000111",
  60974=>"101101100",
  60975=>"111011001",
  60976=>"000000000",
  60977=>"001000000",
  60978=>"000111110",
  60979=>"111110110",
  60980=>"000100100",
  60981=>"110101111",
  60982=>"000000100",
  60983=>"000111111",
  60984=>"000000011",
  60985=>"100100111",
  60986=>"101100111",
  60987=>"000100010",
  60988=>"001001111",
  60989=>"110010010",
  60990=>"000001101",
  60991=>"000100110",
  60992=>"111100001",
  60993=>"000000101",
  60994=>"111101101",
  60995=>"000000000",
  60996=>"111011111",
  60997=>"111100001",
  60998=>"000110100",
  60999=>"011100010",
  61000=>"001001111",
  61001=>"000000000",
  61002=>"001000110",
  61003=>"111111010",
  61004=>"000000000",
  61005=>"001001001",
  61006=>"100101100",
  61007=>"111111010",
  61008=>"010110000",
  61009=>"110000000",
  61010=>"010001101",
  61011=>"001000010",
  61012=>"110100000",
  61013=>"001010011",
  61014=>"111111110",
  61015=>"000010110",
  61016=>"000000000",
  61017=>"001000000",
  61018=>"001001001",
  61019=>"101100100",
  61020=>"000000000",
  61021=>"000000000",
  61022=>"111111111",
  61023=>"000000000",
  61024=>"000010000",
  61025=>"110010011",
  61026=>"000001000",
  61027=>"001000000",
  61028=>"000000011",
  61029=>"101111100",
  61030=>"000011111",
  61031=>"111110100",
  61032=>"001101111",
  61033=>"100001111",
  61034=>"000000000",
  61035=>"100001111",
  61036=>"110110101",
  61037=>"111100000",
  61038=>"001000001",
  61039=>"101000000",
  61040=>"001001100",
  61041=>"000000001",
  61042=>"000000000",
  61043=>"111000000",
  61044=>"000000010",
  61045=>"100000100",
  61046=>"011001000",
  61047=>"001111111",
  61048=>"001000000",
  61049=>"111000000",
  61050=>"111111111",
  61051=>"000010011",
  61052=>"011001001",
  61053=>"000001010",
  61054=>"000001101",
  61055=>"001001000",
  61056=>"101000000",
  61057=>"000000000",
  61058=>"000000000",
  61059=>"111110010",
  61060=>"111001000",
  61061=>"111011000",
  61062=>"000000000",
  61063=>"100100101",
  61064=>"000001100",
  61065=>"101000001",
  61066=>"101111111",
  61067=>"000000000",
  61068=>"111111000",
  61069=>"000000000",
  61070=>"001101101",
  61071=>"001001001",
  61072=>"100100100",
  61073=>"000000000",
  61074=>"000000111",
  61075=>"001001111",
  61076=>"111000000",
  61077=>"000000000",
  61078=>"111001111",
  61079=>"001100101",
  61080=>"111001000",
  61081=>"001101011",
  61082=>"000000000",
  61083=>"111111011",
  61084=>"100111111",
  61085=>"101101111",
  61086=>"010110111",
  61087=>"000000001",
  61088=>"111111111",
  61089=>"111101001",
  61090=>"000000010",
  61091=>"001111011",
  61092=>"000000011",
  61093=>"011011111",
  61094=>"011000000",
  61095=>"110000010",
  61096=>"000000101",
  61097=>"001001001",
  61098=>"101101000",
  61099=>"000001000",
  61100=>"111001000",
  61101=>"001111001",
  61102=>"100100100",
  61103=>"111111111",
  61104=>"111111111",
  61105=>"100110111",
  61106=>"001010101",
  61107=>"000000100",
  61108=>"100000010",
  61109=>"100111110",
  61110=>"111110001",
  61111=>"100111111",
  61112=>"100101111",
  61113=>"000000010",
  61114=>"101111011",
  61115=>"000000010",
  61116=>"111111111",
  61117=>"111110110",
  61118=>"100110011",
  61119=>"000001000",
  61120=>"000000100",
  61121=>"000101111",
  61122=>"000000111",
  61123=>"111111110",
  61124=>"000000011",
  61125=>"100000011",
  61126=>"000000001",
  61127=>"000000000",
  61128=>"010010001",
  61129=>"101101101",
  61130=>"000001110",
  61131=>"000111110",
  61132=>"000101101",
  61133=>"110100000",
  61134=>"111111111",
  61135=>"001110010",
  61136=>"110000110",
  61137=>"011111011",
  61138=>"111101111",
  61139=>"101000010",
  61140=>"000000001",
  61141=>"011111110",
  61142=>"000001111",
  61143=>"000010010",
  61144=>"000000111",
  61145=>"110100110",
  61146=>"111111111",
  61147=>"111110000",
  61148=>"000001000",
  61149=>"111111111",
  61150=>"110110000",
  61151=>"011110111",
  61152=>"100000000",
  61153=>"111111101",
  61154=>"111111111",
  61155=>"011010011",
  61156=>"000100111",
  61157=>"011111111",
  61158=>"000000000",
  61159=>"001011001",
  61160=>"111000011",
  61161=>"000000000",
  61162=>"001001001",
  61163=>"000101000",
  61164=>"111101111",
  61165=>"111110011",
  61166=>"010000000",
  61167=>"000000111",
  61168=>"000000010",
  61169=>"001001101",
  61170=>"000000111",
  61171=>"000000000",
  61172=>"000110101",
  61173=>"111011111",
  61174=>"000000010",
  61175=>"111000011",
  61176=>"000000101",
  61177=>"000010110",
  61178=>"111110010",
  61179=>"000000111",
  61180=>"101101101",
  61181=>"100111001",
  61182=>"101000000",
  61183=>"111101010",
  61184=>"001010110",
  61185=>"000111111",
  61186=>"001100111",
  61187=>"000111111",
  61188=>"011001000",
  61189=>"000000000",
  61190=>"101111111",
  61191=>"111010000",
  61192=>"110001111",
  61193=>"100000111",
  61194=>"100111110",
  61195=>"110000000",
  61196=>"111110000",
  61197=>"110010000",
  61198=>"110110011",
  61199=>"110000000",
  61200=>"011001000",
  61201=>"111000000",
  61202=>"001101111",
  61203=>"000001101",
  61204=>"110111111",
  61205=>"000000111",
  61206=>"000100111",
  61207=>"111010111",
  61208=>"111111111",
  61209=>"110011000",
  61210=>"110110111",
  61211=>"110000011",
  61212=>"111111000",
  61213=>"100111111",
  61214=>"000101101",
  61215=>"011111111",
  61216=>"000000010",
  61217=>"000000001",
  61218=>"000001000",
  61219=>"101111000",
  61220=>"011000001",
  61221=>"000000010",
  61222=>"000001111",
  61223=>"111000000",
  61224=>"101111111",
  61225=>"110010110",
  61226=>"000010000",
  61227=>"000101111",
  61228=>"111000111",
  61229=>"101110111",
  61230=>"111001001",
  61231=>"011010001",
  61232=>"000010000",
  61233=>"011011001",
  61234=>"000111101",
  61235=>"111111101",
  61236=>"101110110",
  61237=>"101110011",
  61238=>"000001111",
  61239=>"110101011",
  61240=>"011100011",
  61241=>"010000000",
  61242=>"000111011",
  61243=>"010011011",
  61244=>"110000000",
  61245=>"111110000",
  61246=>"000001011",
  61247=>"100100000",
  61248=>"100100101",
  61249=>"010110000",
  61250=>"000101010",
  61251=>"000000000",
  61252=>"010000000",
  61253=>"111110000",
  61254=>"000000000",
  61255=>"101101101",
  61256=>"101111001",
  61257=>"011111111",
  61258=>"000000000",
  61259=>"111111010",
  61260=>"111100100",
  61261=>"100001000",
  61262=>"110100000",
  61263=>"101111111",
  61264=>"001000111",
  61265=>"111110000",
  61266=>"101000000",
  61267=>"001001001",
  61268=>"000011000",
  61269=>"000111111",
  61270=>"110110010",
  61271=>"111001000",
  61272=>"110001001",
  61273=>"001011101",
  61274=>"111111111",
  61275=>"100000000",
  61276=>"000100111",
  61277=>"001000011",
  61278=>"111111110",
  61279=>"000000110",
  61280=>"100111111",
  61281=>"001011111",
  61282=>"100000000",
  61283=>"001100100",
  61284=>"001001000",
  61285=>"111101100",
  61286=>"110111111",
  61287=>"010001011",
  61288=>"000111111",
  61289=>"001001000",
  61290=>"111000100",
  61291=>"101100000",
  61292=>"110100111",
  61293=>"001000010",
  61294=>"000100111",
  61295=>"001111111",
  61296=>"001000001",
  61297=>"000110000",
  61298=>"000100010",
  61299=>"101011000",
  61300=>"010000000",
  61301=>"000000000",
  61302=>"110110000",
  61303=>"100010010",
  61304=>"000110011",
  61305=>"110100000",
  61306=>"001000000",
  61307=>"011010000",
  61308=>"100000000",
  61309=>"100000010",
  61310=>"000000111",
  61311=>"111111110",
  61312=>"000000000",
  61313=>"101101000",
  61314=>"100000100",
  61315=>"000111111",
  61316=>"110000100",
  61317=>"111010110",
  61318=>"100000110",
  61319=>"011000000",
  61320=>"110110100",
  61321=>"010001011",
  61322=>"111011011",
  61323=>"010000001",
  61324=>"001001110",
  61325=>"100000100",
  61326=>"000000000",
  61327=>"000010010",
  61328=>"111101000",
  61329=>"111000000",
  61330=>"001001011",
  61331=>"000110011",
  61332=>"110000000",
  61333=>"101001001",
  61334=>"101101010",
  61335=>"011010100",
  61336=>"000000000",
  61337=>"000001001",
  61338=>"000100111",
  61339=>"101000000",
  61340=>"101011111",
  61341=>"010000000",
  61342=>"000011000",
  61343=>"111110100",
  61344=>"001011011",
  61345=>"000000111",
  61346=>"011010111",
  61347=>"001001000",
  61348=>"000001111",
  61349=>"110000100",
  61350=>"001111010",
  61351=>"000101111",
  61352=>"100100001",
  61353=>"110110100",
  61354=>"101101111",
  61355=>"010000100",
  61356=>"110111110",
  61357=>"111000000",
  61358=>"000010111",
  61359=>"101100000",
  61360=>"000000000",
  61361=>"000000000",
  61362=>"111000010",
  61363=>"110000101",
  61364=>"001011111",
  61365=>"101111111",
  61366=>"000000001",
  61367=>"110011010",
  61368=>"011100111",
  61369=>"010111000",
  61370=>"010000111",
  61371=>"111011111",
  61372=>"001000010",
  61373=>"111000100",
  61374=>"000000000",
  61375=>"000011111",
  61376=>"101101111",
  61377=>"000000010",
  61378=>"100000000",
  61379=>"001011000",
  61380=>"011011111",
  61381=>"000100010",
  61382=>"011011000",
  61383=>"000101110",
  61384=>"010000000",
  61385=>"100100000",
  61386=>"001110111",
  61387=>"110000000",
  61388=>"011111000",
  61389=>"001010110",
  61390=>"000000000",
  61391=>"000100111",
  61392=>"000110000",
  61393=>"000110010",
  61394=>"010011001",
  61395=>"111000110",
  61396=>"111000000",
  61397=>"000111011",
  61398=>"110110111",
  61399=>"001101110",
  61400=>"111011000",
  61401=>"000100100",
  61402=>"110101111",
  61403=>"101111011",
  61404=>"001100110",
  61405=>"011010111",
  61406=>"000100000",
  61407=>"001000000",
  61408=>"011101010",
  61409=>"101001011",
  61410=>"111110100",
  61411=>"011111111",
  61412=>"111001000",
  61413=>"111000000",
  61414=>"111100000",
  61415=>"100000010",
  61416=>"101000000",
  61417=>"001000101",
  61418=>"101111111",
  61419=>"000101110",
  61420=>"111110010",
  61421=>"011111001",
  61422=>"111000000",
  61423=>"111100000",
  61424=>"101111011",
  61425=>"011011111",
  61426=>"111000110",
  61427=>"110100000",
  61428=>"101000011",
  61429=>"101010011",
  61430=>"111000000",
  61431=>"100000000",
  61432=>"000000000",
  61433=>"110110111",
  61434=>"101000000",
  61435=>"101001000",
  61436=>"000000010",
  61437=>"010000000",
  61438=>"001000011",
  61439=>"010000000",
  61440=>"111011111",
  61441=>"111110000",
  61442=>"101000000",
  61443=>"000110110",
  61444=>"100110110",
  61445=>"000100111",
  61446=>"110111000",
  61447=>"111011111",
  61448=>"100110011",
  61449=>"000000100",
  61450=>"101000000",
  61451=>"000000000",
  61452=>"100001001",
  61453=>"111110000",
  61454=>"011000011",
  61455=>"001000000",
  61456=>"110111100",
  61457=>"001000000",
  61458=>"100001000",
  61459=>"001111110",
  61460=>"111101101",
  61461=>"110110110",
  61462=>"010000000",
  61463=>"001011111",
  61464=>"101001000",
  61465=>"000000000",
  61466=>"000000011",
  61467=>"001111111",
  61468=>"000000101",
  61469=>"011001000",
  61470=>"111111111",
  61471=>"011000000",
  61472=>"000000000",
  61473=>"110101000",
  61474=>"000000101",
  61475=>"000000000",
  61476=>"100111101",
  61477=>"110111111",
  61478=>"110010000",
  61479=>"111111111",
  61480=>"111001111",
  61481=>"111111111",
  61482=>"101111111",
  61483=>"001000000",
  61484=>"110100100",
  61485=>"000110010",
  61486=>"110110101",
  61487=>"000101000",
  61488=>"111111110",
  61489=>"110100000",
  61490=>"000010010",
  61491=>"000110111",
  61492=>"000000000",
  61493=>"001001001",
  61494=>"000000001",
  61495=>"110111110",
  61496=>"000111111",
  61497=>"110110010",
  61498=>"000101111",
  61499=>"000000000",
  61500=>"100001000",
  61501=>"111111011",
  61502=>"001000100",
  61503=>"110111001",
  61504=>"110011001",
  61505=>"001001101",
  61506=>"111111100",
  61507=>"110110001",
  61508=>"001111100",
  61509=>"001101000",
  61510=>"000111010",
  61511=>"000111110",
  61512=>"110111011",
  61513=>"010000001",
  61514=>"111001000",
  61515=>"111111110",
  61516=>"111111111",
  61517=>"100011011",
  61518=>"010011101",
  61519=>"001001101",
  61520=>"001100111",
  61521=>"111111111",
  61522=>"111111111",
  61523=>"111101101",
  61524=>"001001010",
  61525=>"001111110",
  61526=>"001011111",
  61527=>"001000001",
  61528=>"100100100",
  61529=>"000100110",
  61530=>"000101001",
  61531=>"011011111",
  61532=>"111111110",
  61533=>"001001001",
  61534=>"000110010",
  61535=>"110110100",
  61536=>"000000001",
  61537=>"010110111",
  61538=>"000000000",
  61539=>"000011001",
  61540=>"110111111",
  61541=>"010100100",
  61542=>"101001001",
  61543=>"111111000",
  61544=>"110010010",
  61545=>"001000000",
  61546=>"111111111",
  61547=>"110001101",
  61548=>"111000001",
  61549=>"001001000",
  61550=>"010111110",
  61551=>"100101111",
  61552=>"011111011",
  61553=>"010101111",
  61554=>"000100010",
  61555=>"101001001",
  61556=>"111110110",
  61557=>"001000001",
  61558=>"110111101",
  61559=>"100001111",
  61560=>"000000000",
  61561=>"111001000",
  61562=>"001011010",
  61563=>"110111100",
  61564=>"110100100",
  61565=>"110100100",
  61566=>"000101000",
  61567=>"101110000",
  61568=>"000001001",
  61569=>"111111111",
  61570=>"111010010",
  61571=>"111111111",
  61572=>"000111110",
  61573=>"000111110",
  61574=>"010000101",
  61575=>"001001001",
  61576=>"110110111",
  61577=>"111000010",
  61578=>"101101100",
  61579=>"001101000",
  61580=>"000000000",
  61581=>"111101000",
  61582=>"000110010",
  61583=>"000001001",
  61584=>"000001010",
  61585=>"000100111",
  61586=>"011010011",
  61587=>"110101001",
  61588=>"111010010",
  61589=>"000000001",
  61590=>"000000000",
  61591=>"110011110",
  61592=>"000000000",
  61593=>"100001101",
  61594=>"010111110",
  61595=>"000000000",
  61596=>"001111111",
  61597=>"000001000",
  61598=>"111111111",
  61599=>"101001001",
  61600=>"100000100",
  61601=>"010001010",
  61602=>"111111100",
  61603=>"010011000",
  61604=>"111111111",
  61605=>"001001011",
  61606=>"100110100",
  61607=>"111011100",
  61608=>"001100110",
  61609=>"111111101",
  61610=>"001001001",
  61611=>"001000000",
  61612=>"000111111",
  61613=>"111110110",
  61614=>"100101111",
  61615=>"100101111",
  61616=>"111111100",
  61617=>"011011001",
  61618=>"111011011",
  61619=>"110100100",
  61620=>"111101100",
  61621=>"000000000",
  61622=>"000000000",
  61623=>"000000000",
  61624=>"001000000",
  61625=>"101100100",
  61626=>"010010000",
  61627=>"110000011",
  61628=>"000001000",
  61629=>"001010011",
  61630=>"001111000",
  61631=>"111011001",
  61632=>"000110010",
  61633=>"000000000",
  61634=>"010110111",
  61635=>"111011001",
  61636=>"001000111",
  61637=>"001100110",
  61638=>"111110001",
  61639=>"100110111",
  61640=>"110010111",
  61641=>"110110111",
  61642=>"000000000",
  61643=>"000010000",
  61644=>"111010000",
  61645=>"011001001",
  61646=>"000000000",
  61647=>"111000000",
  61648=>"110111111",
  61649=>"110101011",
  61650=>"000000111",
  61651=>"011101111",
  61652=>"000000111",
  61653=>"100001000",
  61654=>"101110111",
  61655=>"111101111",
  61656=>"000000000",
  61657=>"000000010",
  61658=>"010000010",
  61659=>"001001101",
  61660=>"001100110",
  61661=>"001001000",
  61662=>"110100110",
  61663=>"110111100",
  61664=>"111110001",
  61665=>"000100000",
  61666=>"000000001",
  61667=>"101001000",
  61668=>"000000000",
  61669=>"000001101",
  61670=>"000100110",
  61671=>"111011101",
  61672=>"111001101",
  61673=>"000001001",
  61674=>"001000000",
  61675=>"001000001",
  61676=>"000000000",
  61677=>"000111001",
  61678=>"111000000",
  61679=>"111000001",
  61680=>"000000000",
  61681=>"000011110",
  61682=>"111111110",
  61683=>"011011011",
  61684=>"101100100",
  61685=>"001000010",
  61686=>"011000001",
  61687=>"000111010",
  61688=>"100111111",
  61689=>"011111101",
  61690=>"101111010",
  61691=>"001001000",
  61692=>"110110110",
  61693=>"001000000",
  61694=>"111100111",
  61695=>"111000001",
  61696=>"011001011",
  61697=>"110111111",
  61698=>"000001111",
  61699=>"000000000",
  61700=>"001000011",
  61701=>"000111101",
  61702=>"111000000",
  61703=>"111111101",
  61704=>"010010000",
  61705=>"000000000",
  61706=>"001000110",
  61707=>"000011000",
  61708=>"000100111",
  61709=>"000000001",
  61710=>"100011001",
  61711=>"001000000",
  61712=>"111111111",
  61713=>"000000110",
  61714=>"000001000",
  61715=>"101111110",
  61716=>"011000000",
  61717=>"000000111",
  61718=>"101011111",
  61719=>"100111111",
  61720=>"000010000",
  61721=>"000001000",
  61722=>"000101111",
  61723=>"000000101",
  61724=>"001000000",
  61725=>"100101111",
  61726=>"000000000",
  61727=>"000101000",
  61728=>"010101101",
  61729=>"011111111",
  61730=>"100101100",
  61731=>"000000111",
  61732=>"011001011",
  61733=>"101111000",
  61734=>"000101111",
  61735=>"001000010",
  61736=>"100111111",
  61737=>"000111111",
  61738=>"111000000",
  61739=>"110110110",
  61740=>"111011000",
  61741=>"110010000",
  61742=>"010110111",
  61743=>"000000000",
  61744=>"100111000",
  61745=>"001000000",
  61746=>"010000100",
  61747=>"000111000",
  61748=>"000111111",
  61749=>"111111111",
  61750=>"001111100",
  61751=>"110010000",
  61752=>"010000000",
  61753=>"000100110",
  61754=>"100100100",
  61755=>"000000000",
  61756=>"111110010",
  61757=>"110110110",
  61758=>"000000011",
  61759=>"111110000",
  61760=>"110011111",
  61761=>"111111001",
  61762=>"010010010",
  61763=>"011000000",
  61764=>"100110110",
  61765=>"000000010",
  61766=>"001001000",
  61767=>"110100001",
  61768=>"100010001",
  61769=>"111000000",
  61770=>"000000010",
  61771=>"000010111",
  61772=>"000001000",
  61773=>"111000000",
  61774=>"111000000",
  61775=>"001000010",
  61776=>"111101010",
  61777=>"111010010",
  61778=>"100111111",
  61779=>"001001000",
  61780=>"001111000",
  61781=>"001010110",
  61782=>"010100111",
  61783=>"101101101",
  61784=>"000011011",
  61785=>"100110111",
  61786=>"111110101",
  61787=>"100100110",
  61788=>"110000000",
  61789=>"001011011",
  61790=>"111110000",
  61791=>"100001010",
  61792=>"010000000",
  61793=>"000000000",
  61794=>"001101111",
  61795=>"010010110",
  61796=>"101000000",
  61797=>"001001010",
  61798=>"110111000",
  61799=>"101111011",
  61800=>"110110010",
  61801=>"010000000",
  61802=>"110111110",
  61803=>"111010111",
  61804=>"111111111",
  61805=>"111101011",
  61806=>"101000000",
  61807=>"000010001",
  61808=>"111000001",
  61809=>"000000111",
  61810=>"001110011",
  61811=>"001001001",
  61812=>"000000000",
  61813=>"000101001",
  61814=>"101001110",
  61815=>"000000010",
  61816=>"000001111",
  61817=>"010000010",
  61818=>"110011101",
  61819=>"111000000",
  61820=>"011111110",
  61821=>"100000100",
  61822=>"000000111",
  61823=>"000000010",
  61824=>"001001000",
  61825=>"101001001",
  61826=>"010010000",
  61827=>"111000010",
  61828=>"100110010",
  61829=>"111000000",
  61830=>"111111001",
  61831=>"111000100",
  61832=>"110110001",
  61833=>"000111111",
  61834=>"000001101",
  61835=>"011000101",
  61836=>"000000110",
  61837=>"111110000",
  61838=>"111010000",
  61839=>"000000000",
  61840=>"101111011",
  61841=>"110010011",
  61842=>"000110111",
  61843=>"010001000",
  61844=>"010111110",
  61845=>"000000111",
  61846=>"111000000",
  61847=>"011011001",
  61848=>"010011000",
  61849=>"010110000",
  61850=>"000010111",
  61851=>"111000000",
  61852=>"011010111",
  61853=>"010010000",
  61854=>"000001000",
  61855=>"101101111",
  61856=>"011001001",
  61857=>"000111111",
  61858=>"110000000",
  61859=>"100101101",
  61860=>"011001000",
  61861=>"101000000",
  61862=>"110000001",
  61863=>"111000000",
  61864=>"000000101",
  61865=>"110110000",
  61866=>"001101111",
  61867=>"000000000",
  61868=>"110000000",
  61869=>"100111100",
  61870=>"110110011",
  61871=>"110001000",
  61872=>"010001000",
  61873=>"110000000",
  61874=>"101001101",
  61875=>"001000110",
  61876=>"111011000",
  61877=>"000000110",
  61878=>"000000000",
  61879=>"000011100",
  61880=>"010101010",
  61881=>"111011000",
  61882=>"111010000",
  61883=>"110000100",
  61884=>"110001001",
  61885=>"101111111",
  61886=>"110000000",
  61887=>"000000000",
  61888=>"000101111",
  61889=>"100111111",
  61890=>"011111000",
  61891=>"001011111",
  61892=>"100000000",
  61893=>"100101100",
  61894=>"111111010",
  61895=>"001111111",
  61896=>"001000100",
  61897=>"110111101",
  61898=>"000101111",
  61899=>"111011000",
  61900=>"010010000",
  61901=>"111100110",
  61902=>"000001111",
  61903=>"101000000",
  61904=>"000101111",
  61905=>"110110110",
  61906=>"000000110",
  61907=>"011000000",
  61908=>"001011011",
  61909=>"110110110",
  61910=>"000010111",
  61911=>"010110111",
  61912=>"000001110",
  61913=>"110111000",
  61914=>"100100110",
  61915=>"000000111",
  61916=>"000100011",
  61917=>"010000000",
  61918=>"000000010",
  61919=>"000000000",
  61920=>"000101111",
  61921=>"000100000",
  61922=>"000001001",
  61923=>"011011001",
  61924=>"000111111",
  61925=>"010111010",
  61926=>"000000101",
  61927=>"010000100",
  61928=>"111011101",
  61929=>"010111111",
  61930=>"000100011",
  61931=>"000100111",
  61932=>"000000101",
  61933=>"000111111",
  61934=>"101000010",
  61935=>"101100100",
  61936=>"000000000",
  61937=>"011011011",
  61938=>"000001001",
  61939=>"011011000",
  61940=>"111010000",
  61941=>"000111111",
  61942=>"000110111",
  61943=>"100000000",
  61944=>"111111010",
  61945=>"000101000",
  61946=>"100110111",
  61947=>"011111101",
  61948=>"000000111",
  61949=>"111010000",
  61950=>"011011100",
  61951=>"110101000",
  61952=>"011000100",
  61953=>"011000001",
  61954=>"001001111",
  61955=>"000010010",
  61956=>"111111000",
  61957=>"110110000",
  61958=>"010000001",
  61959=>"111111110",
  61960=>"100110000",
  61961=>"101001100",
  61962=>"100000001",
  61963=>"111000000",
  61964=>"000001110",
  61965=>"110110000",
  61966=>"011001101",
  61967=>"000000000",
  61968=>"110110000",
  61969=>"000001101",
  61970=>"000111111",
  61971=>"110110000",
  61972=>"000001100",
  61973=>"111111111",
  61974=>"011111111",
  61975=>"011111111",
  61976=>"100110110",
  61977=>"111111111",
  61978=>"101000111",
  61979=>"000101111",
  61980=>"100100001",
  61981=>"110101000",
  61982=>"100001001",
  61983=>"000111111",
  61984=>"001001001",
  61985=>"111110001",
  61986=>"000000000",
  61987=>"100110110",
  61988=>"000001000",
  61989=>"110100000",
  61990=>"001000110",
  61991=>"000110000",
  61992=>"011111010",
  61993=>"101110111",
  61994=>"000001111",
  61995=>"000000000",
  61996=>"010011000",
  61997=>"000010011",
  61998=>"111000000",
  61999=>"000110111",
  62000=>"000111110",
  62001=>"111111010",
  62002=>"001001000",
  62003=>"001111111",
  62004=>"011001111",
  62005=>"111101000",
  62006=>"110100001",
  62007=>"001001001",
  62008=>"001000010",
  62009=>"001001111",
  62010=>"011111110",
  62011=>"011111011",
  62012=>"000110100",
  62013=>"010111010",
  62014=>"000000011",
  62015=>"000010000",
  62016=>"111111101",
  62017=>"111111111",
  62018=>"110000001",
  62019=>"110111001",
  62020=>"010000010",
  62021=>"100100000",
  62022=>"110111111",
  62023=>"111111001",
  62024=>"001110000",
  62025=>"110001110",
  62026=>"111001111",
  62027=>"101001101",
  62028=>"101000000",
  62029=>"111111100",
  62030=>"100110100",
  62031=>"111011001",
  62032=>"110110000",
  62033=>"101001110",
  62034=>"001000000",
  62035=>"010010000",
  62036=>"000000110",
  62037=>"101110011",
  62038=>"011011010",
  62039=>"111001111",
  62040=>"100100111",
  62041=>"001011111",
  62042=>"110100100",
  62043=>"011101000",
  62044=>"000001111",
  62045=>"000000000",
  62046=>"111110000",
  62047=>"110110101",
  62048=>"000010000",
  62049=>"000010111",
  62050=>"000000011",
  62051=>"011000011",
  62052=>"000000000",
  62053=>"011111000",
  62054=>"000101000",
  62055=>"000101000",
  62056=>"110111110",
  62057=>"111000000",
  62058=>"110110000",
  62059=>"111011001",
  62060=>"100110111",
  62061=>"001001101",
  62062=>"000001100",
  62063=>"001111110",
  62064=>"101001100",
  62065=>"111001001",
  62066=>"001111100",
  62067=>"000001111",
  62068=>"010000000",
  62069=>"000001001",
  62070=>"110000001",
  62071=>"000110000",
  62072=>"000010110",
  62073=>"010000000",
  62074=>"001000000",
  62075=>"110110001",
  62076=>"100000110",
  62077=>"110111000",
  62078=>"010100111",
  62079=>"101110101",
  62080=>"111001000",
  62081=>"110000001",
  62082=>"101000000",
  62083=>"000011010",
  62084=>"110110101",
  62085=>"001001111",
  62086=>"011011000",
  62087=>"001001011",
  62088=>"101001011",
  62089=>"010110000",
  62090=>"001001111",
  62091=>"111110111",
  62092=>"000000000",
  62093=>"001001001",
  62094=>"000000111",
  62095=>"001001001",
  62096=>"111111000",
  62097=>"000100100",
  62098=>"001000000",
  62099=>"010111111",
  62100=>"001111100",
  62101=>"111001101",
  62102=>"101101111",
  62103=>"011010000",
  62104=>"001111111",
  62105=>"001110110",
  62106=>"111101101",
  62107=>"010000000",
  62108=>"001001001",
  62109=>"000000000",
  62110=>"001111110",
  62111=>"001000111",
  62112=>"101011111",
  62113=>"110110111",
  62114=>"000000000",
  62115=>"000011101",
  62116=>"000111001",
  62117=>"001000100",
  62118=>"000000000",
  62119=>"111000000",
  62120=>"001001001",
  62121=>"100000001",
  62122=>"111111111",
  62123=>"001000001",
  62124=>"001111101",
  62125=>"001000110",
  62126=>"110100011",
  62127=>"000000001",
  62128=>"010111101",
  62129=>"101011000",
  62130=>"010010010",
  62131=>"000000000",
  62132=>"000110000",
  62133=>"010010010",
  62134=>"010111010",
  62135=>"110000101",
  62136=>"010011011",
  62137=>"000100101",
  62138=>"011001001",
  62139=>"110010110",
  62140=>"000001000",
  62141=>"010010000",
  62142=>"010110000",
  62143=>"000000100",
  62144=>"100000001",
  62145=>"000001111",
  62146=>"110101001",
  62147=>"111010000",
  62148=>"000001011",
  62149=>"101000101",
  62150=>"110000000",
  62151=>"110000000",
  62152=>"110110110",
  62153=>"111011001",
  62154=>"110110110",
  62155=>"000111110",
  62156=>"000111110",
  62157=>"011000001",
  62158=>"001000010",
  62159=>"110111110",
  62160=>"110010000",
  62161=>"110101110",
  62162=>"101111111",
  62163=>"101101101",
  62164=>"000000001",
  62165=>"000000010",
  62166=>"101000101",
  62167=>"010001111",
  62168=>"001101110",
  62169=>"000000000",
  62170=>"011110100",
  62171=>"101101111",
  62172=>"101101110",
  62173=>"011110111",
  62174=>"000001001",
  62175=>"101001111",
  62176=>"111111010",
  62177=>"001000111",
  62178=>"110111000",
  62179=>"011111000",
  62180=>"000000001",
  62181=>"110010000",
  62182=>"111000000",
  62183=>"000001111",
  62184=>"001000000",
  62185=>"000000000",
  62186=>"001001000",
  62187=>"111111111",
  62188=>"000000000",
  62189=>"011100001",
  62190=>"000000010",
  62191=>"111010010",
  62192=>"111101110",
  62193=>"011001011",
  62194=>"000100101",
  62195=>"110110110",
  62196=>"110000100",
  62197=>"001000000",
  62198=>"101000101",
  62199=>"000011000",
  62200=>"000111010",
  62201=>"110110000",
  62202=>"101001011",
  62203=>"001011010",
  62204=>"100101111",
  62205=>"111111110",
  62206=>"100100000",
  62207=>"001000111",
  62208=>"000000000",
  62209=>"100000001",
  62210=>"001000101",
  62211=>"101001011",
  62212=>"000111000",
  62213=>"100101001",
  62214=>"000111111",
  62215=>"110111111",
  62216=>"010011110",
  62217=>"111001111",
  62218=>"011011010",
  62219=>"111111111",
  62220=>"100000000",
  62221=>"111111101",
  62222=>"100110100",
  62223=>"011011111",
  62224=>"011101110",
  62225=>"011001000",
  62226=>"000000000",
  62227=>"000011010",
  62228=>"101111000",
  62229=>"001000001",
  62230=>"001000000",
  62231=>"111111001",
  62232=>"000000100",
  62233=>"111000011",
  62234=>"010000101",
  62235=>"000111101",
  62236=>"001000101",
  62237=>"000000010",
  62238=>"000000000",
  62239=>"111111111",
  62240=>"111100010",
  62241=>"111111111",
  62242=>"000000111",
  62243=>"000001000",
  62244=>"001111011",
  62245=>"011000001",
  62246=>"001101001",
  62247=>"000010110",
  62248=>"000001011",
  62249=>"100101111",
  62250=>"000000000",
  62251=>"101101101",
  62252=>"110001011",
  62253=>"001010000",
  62254=>"001000000",
  62255=>"110110100",
  62256=>"000111100",
  62257=>"001000011",
  62258=>"000111111",
  62259=>"011001101",
  62260=>"000111000",
  62261=>"101001000",
  62262=>"110110100",
  62263=>"000000100",
  62264=>"111111111",
  62265=>"000000000",
  62266=>"000000001",
  62267=>"000000110",
  62268=>"001000111",
  62269=>"111110011",
  62270=>"000001101",
  62271=>"100100100",
  62272=>"101001111",
  62273=>"000000000",
  62274=>"111111010",
  62275=>"010000001",
  62276=>"000000011",
  62277=>"000000000",
  62278=>"000011100",
  62279=>"101111111",
  62280=>"000010000",
  62281=>"000110111",
  62282=>"100000001",
  62283=>"011111010",
  62284=>"111111110",
  62285=>"001101100",
  62286=>"001111110",
  62287=>"000000010",
  62288=>"000000001",
  62289=>"011110111",
  62290=>"101101000",
  62291=>"110011011",
  62292=>"100100101",
  62293=>"001001000",
  62294=>"000010010",
  62295=>"101001101",
  62296=>"111001000",
  62297=>"010111011",
  62298=>"010000000",
  62299=>"111110000",
  62300=>"000000100",
  62301=>"000000010",
  62302=>"110010000",
  62303=>"000000000",
  62304=>"000010000",
  62305=>"001000101",
  62306=>"000000011",
  62307=>"011000010",
  62308=>"111111111",
  62309=>"010011110",
  62310=>"011111111",
  62311=>"001000111",
  62312=>"011111101",
  62313=>"111111111",
  62314=>"111000000",
  62315=>"000000001",
  62316=>"001100110",
  62317=>"111111101",
  62318=>"111000001",
  62319=>"010111111",
  62320=>"110011110",
  62321=>"111111011",
  62322=>"011011111",
  62323=>"000000000",
  62324=>"111010000",
  62325=>"000000111",
  62326=>"011110000",
  62327=>"000000111",
  62328=>"101000000",
  62329=>"011111100",
  62330=>"111111111",
  62331=>"001110110",
  62332=>"011001011",
  62333=>"001001000",
  62334=>"010101111",
  62335=>"000000010",
  62336=>"000000001",
  62337=>"101100111",
  62338=>"000000000",
  62339=>"000000010",
  62340=>"011001001",
  62341=>"111101011",
  62342=>"100000100",
  62343=>"111111111",
  62344=>"000010010",
  62345=>"010111000",
  62346=>"011111000",
  62347=>"001000101",
  62348=>"111100000",
  62349=>"000000000",
  62350=>"111000000",
  62351=>"000000111",
  62352=>"111011011",
  62353=>"000000000",
  62354=>"111111000",
  62355=>"000000011",
  62356=>"111111101",
  62357=>"101001001",
  62358=>"111111100",
  62359=>"110100001",
  62360=>"000000001",
  62361=>"000011001",
  62362=>"101000101",
  62363=>"100111101",
  62364=>"100110100",
  62365=>"010000010",
  62366=>"101111111",
  62367=>"100000111",
  62368=>"000000000",
  62369=>"111101000",
  62370=>"101111111",
  62371=>"000010000",
  62372=>"001111101",
  62373=>"010111111",
  62374=>"000000010",
  62375=>"101101111",
  62376=>"101001001",
  62377=>"111101001",
  62378=>"111100101",
  62379=>"101000000",
  62380=>"110010000",
  62381=>"000011001",
  62382=>"011111111",
  62383=>"010100111",
  62384=>"001000101",
  62385=>"100100111",
  62386=>"101111001",
  62387=>"001011111",
  62388=>"110010110",
  62389=>"010000000",
  62390=>"000000000",
  62391=>"111000011",
  62392=>"000000011",
  62393=>"111111111",
  62394=>"000100111",
  62395=>"010011111",
  62396=>"100000000",
  62397=>"101011000",
  62398=>"001010010",
  62399=>"000101100",
  62400=>"000000000",
  62401=>"001000000",
  62402=>"111111010",
  62403=>"000100000",
  62404=>"000111001",
  62405=>"111111111",
  62406=>"110011111",
  62407=>"111111111",
  62408=>"000000010",
  62409=>"101101000",
  62410=>"000011000",
  62411=>"100010000",
  62412=>"000111100",
  62413=>"100100110",
  62414=>"111101111",
  62415=>"010000100",
  62416=>"111011100",
  62417=>"000010100",
  62418=>"111111111",
  62419=>"111111010",
  62420=>"111001101",
  62421=>"001001000",
  62422=>"101100000",
  62423=>"110111101",
  62424=>"000001001",
  62425=>"000101010",
  62426=>"001011011",
  62427=>"101101001",
  62428=>"100000110",
  62429=>"110011101",
  62430=>"110101010",
  62431=>"000101110",
  62432=>"000000000",
  62433=>"111110000",
  62434=>"110010000",
  62435=>"000011011",
  62436=>"000000000",
  62437=>"000010111",
  62438=>"101111100",
  62439=>"100010011",
  62440=>"110001100",
  62441=>"111110100",
  62442=>"100100000",
  62443=>"000000001",
  62444=>"001000111",
  62445=>"101101001",
  62446=>"111011011",
  62447=>"000000001",
  62448=>"011001001",
  62449=>"111111111",
  62450=>"000000101",
  62451=>"011111010",
  62452=>"000000111",
  62453=>"010010010",
  62454=>"000000111",
  62455=>"000000000",
  62456=>"100000101",
  62457=>"111111000",
  62458=>"111101000",
  62459=>"111111111",
  62460=>"011111011",
  62461=>"000010000",
  62462=>"000000000",
  62463=>"000000000",
  62464=>"010100110",
  62465=>"010111111",
  62466=>"101000100",
  62467=>"010000000",
  62468=>"111011011",
  62469=>"011000000",
  62470=>"111111011",
  62471=>"000111011",
  62472=>"000000100",
  62473=>"000101001",
  62474=>"111101101",
  62475=>"111100000",
  62476=>"100111111",
  62477=>"111111000",
  62478=>"111101100",
  62479=>"000010000",
  62480=>"010000000",
  62481=>"101000100",
  62482=>"000101000",
  62483=>"110100000",
  62484=>"000011111",
  62485=>"000100110",
  62486=>"000101101",
  62487=>"101101101",
  62488=>"111000100",
  62489=>"110010000",
  62490=>"010100000",
  62491=>"111000000",
  62492=>"111101001",
  62493=>"000100111",
  62494=>"110000000",
  62495=>"000110111",
  62496=>"011101000",
  62497=>"111111011",
  62498=>"000100111",
  62499=>"000110000",
  62500=>"011000001",
  62501=>"011001010",
  62502=>"000000001",
  62503=>"111011000",
  62504=>"111111001",
  62505=>"100111010",
  62506=>"000001000",
  62507=>"110000000",
  62508=>"111110100",
  62509=>"101010101",
  62510=>"000000000",
  62511=>"101111101",
  62512=>"000001111",
  62513=>"111100000",
  62514=>"000111111",
  62515=>"011000111",
  62516=>"111001000",
  62517=>"111111101",
  62518=>"110000000",
  62519=>"000110111",
  62520=>"100010001",
  62521=>"000000000",
  62522=>"011100101",
  62523=>"000100001",
  62524=>"110000000",
  62525=>"000111111",
  62526=>"100000000",
  62527=>"111111111",
  62528=>"100101100",
  62529=>"110000011",
  62530=>"010010010",
  62531=>"011100000",
  62532=>"000000000",
  62533=>"000011100",
  62534=>"111000000",
  62535=>"001000101",
  62536=>"000101111",
  62537=>"011000000",
  62538=>"001000111",
  62539=>"000000000",
  62540=>"111000000",
  62541=>"000001100",
  62542=>"110111100",
  62543=>"111110101",
  62544=>"101101000",
  62545=>"111100000",
  62546=>"010101100",
  62547=>"010011001",
  62548=>"101101100",
  62549=>"001110111",
  62550=>"001001000",
  62551=>"111000000",
  62552=>"111111000",
  62553=>"111101100",
  62554=>"111111101",
  62555=>"001011011",
  62556=>"000000010",
  62557=>"000001001",
  62558=>"000111111",
  62559=>"000000000",
  62560=>"011111110",
  62561=>"001111110",
  62562=>"111100000",
  62563=>"100101111",
  62564=>"100001010",
  62565=>"010000000",
  62566=>"111000000",
  62567=>"000000011",
  62568=>"111100110",
  62569=>"000000000",
  62570=>"101000010",
  62571=>"000111101",
  62572=>"000000111",
  62573=>"101000000",
  62574=>"000000000",
  62575=>"001000011",
  62576=>"000000011",
  62577=>"001000001",
  62578=>"011000000",
  62579=>"000000000",
  62580=>"011011001",
  62581=>"000000000",
  62582=>"111111101",
  62583=>"000010011",
  62584=>"111101000",
  62585=>"110010111",
  62586=>"000100000",
  62587=>"001100111",
  62588=>"111100000",
  62589=>"000010000",
  62590=>"000011011",
  62591=>"101101100",
  62592=>"100000000",
  62593=>"000111010",
  62594=>"000000011",
  62595=>"000001010",
  62596=>"111100000",
  62597=>"000100010",
  62598=>"010001011",
  62599=>"000001001",
  62600=>"111111110",
  62601=>"011000000",
  62602=>"000000011",
  62603=>"000010000",
  62604=>"000010010",
  62605=>"000000110",
  62606=>"100010111",
  62607=>"110000000",
  62608=>"100001001",
  62609=>"110110111",
  62610=>"101101100",
  62611=>"100101000",
  62612=>"100110100",
  62613=>"111000000",
  62614=>"110000000",
  62615=>"000000011",
  62616=>"000000000",
  62617=>"000100011",
  62618=>"111100000",
  62619=>"011000000",
  62620=>"011000111",
  62621=>"111100000",
  62622=>"001111111",
  62623=>"000001111",
  62624=>"001001011",
  62625=>"101000011",
  62626=>"000011111",
  62627=>"000100111",
  62628=>"011011000",
  62629=>"010111111",
  62630=>"001010011",
  62631=>"010101001",
  62632=>"111000100",
  62633=>"000010011",
  62634=>"111111100",
  62635=>"111000000",
  62636=>"000010011",
  62637=>"111100000",
  62638=>"110000001",
  62639=>"000111111",
  62640=>"000000100",
  62641=>"000100011",
  62642=>"111100100",
  62643=>"000100000",
  62644=>"010011011",
  62645=>"111011111",
  62646=>"000111010",
  62647=>"111001000",
  62648=>"011011000",
  62649=>"000100011",
  62650=>"111000101",
  62651=>"111111111",
  62652=>"011011010",
  62653=>"111010000",
  62654=>"000011110",
  62655=>"000010011",
  62656=>"101100100",
  62657=>"101100100",
  62658=>"111101111",
  62659=>"000100000",
  62660=>"000000000",
  62661=>"111100101",
  62662=>"000000011",
  62663=>"111100100",
  62664=>"111111000",
  62665=>"100011000",
  62666=>"110111001",
  62667=>"000011010",
  62668=>"011000110",
  62669=>"110111001",
  62670=>"111101101",
  62671=>"011111111",
  62672=>"011000100",
  62673=>"010000100",
  62674=>"010000000",
  62675=>"001010111",
  62676=>"101100101",
  62677=>"000100111",
  62678=>"111100000",
  62679=>"001000000",
  62680=>"000111011",
  62681=>"000100111",
  62682=>"100111111",
  62683=>"100100000",
  62684=>"110011001",
  62685=>"111011101",
  62686=>"000111111",
  62687=>"011000000",
  62688=>"111111000",
  62689=>"000000100",
  62690=>"101000111",
  62691=>"011001011",
  62692=>"001000000",
  62693=>"000110010",
  62694=>"101101000",
  62695=>"000110100",
  62696=>"000000000",
  62697=>"011000000",
  62698=>"111110101",
  62699=>"011011000",
  62700=>"000111000",
  62701=>"111000000",
  62702=>"000001001",
  62703=>"010101101",
  62704=>"011111101",
  62705=>"101001011",
  62706=>"011011000",
  62707=>"001111101",
  62708=>"010001001",
  62709=>"011101000",
  62710=>"010000100",
  62711=>"001001000",
  62712=>"111101000",
  62713=>"000101100",
  62714=>"000011000",
  62715=>"000111001",
  62716=>"011000000",
  62717=>"101000001",
  62718=>"000110111",
  62719=>"111100011",
  62720=>"001001001",
  62721=>"101111111",
  62722=>"100101111",
  62723=>"001111111",
  62724=>"111110011",
  62725=>"000000001",
  62726=>"100100110",
  62727=>"111111101",
  62728=>"000000110",
  62729=>"000000000",
  62730=>"111011000",
  62731=>"101101000",
  62732=>"101011110",
  62733=>"000000000",
  62734=>"110100100",
  62735=>"111110000",
  62736=>"101000111",
  62737=>"111011111",
  62738=>"001110111",
  62739=>"111011000",
  62740=>"000111110",
  62741=>"101111111",
  62742=>"001001111",
  62743=>"010111101",
  62744=>"000000000",
  62745=>"101001111",
  62746=>"000000000",
  62747=>"000000100",
  62748=>"101101000",
  62749=>"011011111",
  62750=>"111000000",
  62751=>"000001111",
  62752=>"110000101",
  62753=>"000000001",
  62754=>"000111001",
  62755=>"000000111",
  62756=>"000000000",
  62757=>"110011001",
  62758=>"110011010",
  62759=>"000001101",
  62760=>"101111000",
  62761=>"010111000",
  62762=>"111101101",
  62763=>"000000011",
  62764=>"111111010",
  62765=>"001111111",
  62766=>"000000011",
  62767=>"110100111",
  62768=>"111001000",
  62769=>"000111110",
  62770=>"000111101",
  62771=>"000000000",
  62772=>"111111101",
  62773=>"101000000",
  62774=>"110110110",
  62775=>"010000001",
  62776=>"000111111",
  62777=>"000001000",
  62778=>"101111111",
  62779=>"000111001",
  62780=>"111001001",
  62781=>"000011000",
  62782=>"000000111",
  62783=>"010111001",
  62784=>"000000000",
  62785=>"111111110",
  62786=>"110111000",
  62787=>"010001001",
  62788=>"000000000",
  62789=>"000001000",
  62790=>"111111000",
  62791=>"101000110",
  62792=>"111011001",
  62793=>"001000001",
  62794=>"000101011",
  62795=>"110000000",
  62796=>"010110111",
  62797=>"001000010",
  62798=>"111111110",
  62799=>"101110111",
  62800=>"111110111",
  62801=>"011111100",
  62802=>"111000111",
  62803=>"000100111",
  62804=>"000000010",
  62805=>"100111110",
  62806=>"011111100",
  62807=>"000000000",
  62808=>"000000111",
  62809=>"100110111",
  62810=>"111000000",
  62811=>"111000000",
  62812=>"001000000",
  62813=>"001000111",
  62814=>"011010010",
  62815=>"010100100",
  62816=>"111111000",
  62817=>"100001000",
  62818=>"000000011",
  62819=>"011110110",
  62820=>"011010001",
  62821=>"000101101",
  62822=>"000000111",
  62823=>"000010110",
  62824=>"000101000",
  62825=>"011000101",
  62826=>"111110000",
  62827=>"000000000",
  62828=>"001000100",
  62829=>"110000111",
  62830=>"110000000",
  62831=>"111001000",
  62832=>"011011001",
  62833=>"001100101",
  62834=>"111011001",
  62835=>"001000100",
  62836=>"011111110",
  62837=>"000111111",
  62838=>"111111000",
  62839=>"011000000",
  62840=>"101001110",
  62841=>"000000111",
  62842=>"000000000",
  62843=>"000111111",
  62844=>"000010011",
  62845=>"100000000",
  62846=>"010001111",
  62847=>"000000011",
  62848=>"000000000",
  62849=>"011011000",
  62850=>"010010111",
  62851=>"010001110",
  62852=>"001100111",
  62853=>"000000000",
  62854=>"001110000",
  62855=>"110000000",
  62856=>"111101000",
  62857=>"000000011",
  62858=>"000000111",
  62859=>"000001111",
  62860=>"000000001",
  62861=>"010111101",
  62862=>"111111111",
  62863=>"000000011",
  62864=>"100100110",
  62865=>"000001000",
  62866=>"010111001",
  62867=>"000001000",
  62868=>"000001001",
  62869=>"111001101",
  62870=>"111010000",
  62871=>"011011010",
  62872=>"111101000",
  62873=>"000111000",
  62874=>"111011010",
  62875=>"000111100",
  62876=>"011111000",
  62877=>"000000000",
  62878=>"110101100",
  62879=>"000010110",
  62880=>"101111000",
  62881=>"100110111",
  62882=>"011000000",
  62883=>"001001101",
  62884=>"001011011",
  62885=>"001000001",
  62886=>"111111101",
  62887=>"010010001",
  62888=>"000111111",
  62889=>"111111111",
  62890=>"101000111",
  62891=>"000000110",
  62892=>"111010000",
  62893=>"001101111",
  62894=>"000000111",
  62895=>"000000001",
  62896=>"111101101",
  62897=>"011001000",
  62898=>"010100111",
  62899=>"100010011",
  62900=>"111100110",
  62901=>"111001101",
  62902=>"011000001",
  62903=>"001000111",
  62904=>"110100100",
  62905=>"011100100",
  62906=>"111111110",
  62907=>"001101001",
  62908=>"111000011",
  62909=>"010011000",
  62910=>"100100100",
  62911=>"001000001",
  62912=>"000000110",
  62913=>"100000000",
  62914=>"010111100",
  62915=>"001001000",
  62916=>"000000111",
  62917=>"110001111",
  62918=>"100101111",
  62919=>"010111111",
  62920=>"111111000",
  62921=>"000000100",
  62922=>"111011111",
  62923=>"111111001",
  62924=>"010100101",
  62925=>"011010100",
  62926=>"111000110",
  62927=>"000111110",
  62928=>"000010000",
  62929=>"111110010",
  62930=>"101101101",
  62931=>"111101100",
  62932=>"111001111",
  62933=>"100110000",
  62934=>"000101111",
  62935=>"110111000",
  62936=>"001111001",
  62937=>"101000111",
  62938=>"101100000",
  62939=>"000000101",
  62940=>"001110111",
  62941=>"000010111",
  62942=>"001001111",
  62943=>"001011111",
  62944=>"000000000",
  62945=>"001000010",
  62946=>"101111111",
  62947=>"111011000",
  62948=>"001101001",
  62949=>"001000001",
  62950=>"111110000",
  62951=>"000010110",
  62952=>"011110100",
  62953=>"000111011",
  62954=>"111111000",
  62955=>"111000000",
  62956=>"000000000",
  62957=>"000000111",
  62958=>"000010000",
  62959=>"111100010",
  62960=>"111111000",
  62961=>"010001011",
  62962=>"110101111",
  62963=>"111111111",
  62964=>"101101111",
  62965=>"000000100",
  62966=>"000000101",
  62967=>"000110100",
  62968=>"111101001",
  62969=>"111111101",
  62970=>"100000000",
  62971=>"110101111",
  62972=>"110110000",
  62973=>"111000000",
  62974=>"001111100",
  62975=>"110111000",
  62976=>"110110110",
  62977=>"101101010",
  62978=>"000000000",
  62979=>"111010100",
  62980=>"111100001",
  62981=>"111111000",
  62982=>"011111011",
  62983=>"010001100",
  62984=>"111111100",
  62985=>"001000000",
  62986=>"000001111",
  62987=>"101101000",
  62988=>"100100101",
  62989=>"000000010",
  62990=>"011010110",
  62991=>"111101000",
  62992=>"011111000",
  62993=>"000011011",
  62994=>"101101110",
  62995=>"010000100",
  62996=>"111111111",
  62997=>"101001001",
  62998=>"011111011",
  62999=>"110000010",
  63000=>"111000101",
  63001=>"001000101",
  63002=>"100000011",
  63003=>"101011010",
  63004=>"000110000",
  63005=>"111110000",
  63006=>"100000101",
  63007=>"100000100",
  63008=>"011011000",
  63009=>"111100000",
  63010=>"111000101",
  63011=>"011111111",
  63012=>"000001101",
  63013=>"100101010",
  63014=>"111100100",
  63015=>"000000111",
  63016=>"111111000",
  63017=>"100100111",
  63018=>"101101010",
  63019=>"110000000",
  63020=>"001111111",
  63021=>"010111111",
  63022=>"011001100",
  63023=>"000010010",
  63024=>"100111101",
  63025=>"111111011",
  63026=>"000000111",
  63027=>"111011111",
  63028=>"011000000",
  63029=>"100111011",
  63030=>"010000000",
  63031=>"000000100",
  63032=>"001000000",
  63033=>"100101101",
  63034=>"111110100",
  63035=>"101100110",
  63036=>"100001101",
  63037=>"100111010",
  63038=>"001000000",
  63039=>"100110111",
  63040=>"011000000",
  63041=>"010000111",
  63042=>"000111101",
  63043=>"011011110",
  63044=>"100100100",
  63045=>"100111000",
  63046=>"010010000",
  63047=>"010101011",
  63048=>"111101001",
  63049=>"011010000",
  63050=>"111100000",
  63051=>"000100000",
  63052=>"100100000",
  63053=>"000100100",
  63054=>"011011110",
  63055=>"010101111",
  63056=>"000100001",
  63057=>"010011010",
  63058=>"011101010",
  63059=>"011100101",
  63060=>"111100000",
  63061=>"100111100",
  63062=>"010000100",
  63063=>"111111011",
  63064=>"111101111",
  63065=>"111111111",
  63066=>"011011111",
  63067=>"010000101",
  63068=>"000010000",
  63069=>"101101001",
  63070=>"100100111",
  63071=>"110110001",
  63072=>"000011110",
  63073=>"000000000",
  63074=>"111000101",
  63075=>"111110100",
  63076=>"000010000",
  63077=>"011011101",
  63078=>"110110001",
  63079=>"011011000",
  63080=>"001011110",
  63081=>"100100000",
  63082=>"000000011",
  63083=>"111111111",
  63084=>"111100110",
  63085=>"000011111",
  63086=>"001000000",
  63087=>"100000000",
  63088=>"111110000",
  63089=>"100000111",
  63090=>"011010110",
  63091=>"000011101",
  63092=>"000000110",
  63093=>"000000000",
  63094=>"100000000",
  63095=>"000101111",
  63096=>"000100111",
  63097=>"001100101",
  63098=>"101001000",
  63099=>"100010111",
  63100=>"010110001",
  63101=>"010010000",
  63102=>"010010010",
  63103=>"111011010",
  63104=>"000010111",
  63105=>"010000000",
  63106=>"011010000",
  63107=>"111011101",
  63108=>"010000001",
  63109=>"110000111",
  63110=>"011001011",
  63111=>"100000001",
  63112=>"001011000",
  63113=>"000000000",
  63114=>"011011011",
  63115=>"111101111",
  63116=>"000011000",
  63117=>"100100001",
  63118=>"111111110",
  63119=>"110100000",
  63120=>"110011001",
  63121=>"110110111",
  63122=>"111001010",
  63123=>"111011000",
  63124=>"111101011",
  63125=>"101111000",
  63126=>"000101000",
  63127=>"101100000",
  63128=>"001101001",
  63129=>"100000111",
  63130=>"001111111",
  63131=>"000000000",
  63132=>"000000100",
  63133=>"100000000",
  63134=>"000000110",
  63135=>"111111000",
  63136=>"110011001",
  63137=>"111011100",
  63138=>"111101111",
  63139=>"000000111",
  63140=>"000000111",
  63141=>"011011110",
  63142=>"111001001",
  63143=>"000100000",
  63144=>"100111111",
  63145=>"000101100",
  63146=>"111111111",
  63147=>"111111010",
  63148=>"001000000",
  63149=>"000000000",
  63150=>"110110010",
  63151=>"000000000",
  63152=>"000000000",
  63153=>"001100110",
  63154=>"000000000",
  63155=>"000110100",
  63156=>"111111111",
  63157=>"000011111",
  63158=>"000011000",
  63159=>"101100111",
  63160=>"100110101",
  63161=>"011101100",
  63162=>"010101100",
  63163=>"001111111",
  63164=>"111011011",
  63165=>"111111011",
  63166=>"010011001",
  63167=>"100010011",
  63168=>"000000000",
  63169=>"111110010",
  63170=>"111000011",
  63171=>"111100011",
  63172=>"000000111",
  63173=>"111111101",
  63174=>"000000000",
  63175=>"000000110",
  63176=>"100111000",
  63177=>"000001100",
  63178=>"000000010",
  63179=>"111101000",
  63180=>"000011011",
  63181=>"010011111",
  63182=>"011011011",
  63183=>"000000010",
  63184=>"010010000",
  63185=>"010011011",
  63186=>"111111000",
  63187=>"111100000",
  63188=>"000000100",
  63189=>"001011101",
  63190=>"011111111",
  63191=>"010000000",
  63192=>"000000100",
  63193=>"000000000",
  63194=>"000001000",
  63195=>"101000101",
  63196=>"011010000",
  63197=>"000000101",
  63198=>"000000000",
  63199=>"000010000",
  63200=>"000000000",
  63201=>"100100111",
  63202=>"101101001",
  63203=>"110111100",
  63204=>"000111000",
  63205=>"111111111",
  63206=>"100000000",
  63207=>"011111101",
  63208=>"100111101",
  63209=>"100000000",
  63210=>"100110010",
  63211=>"011011111",
  63212=>"011111111",
  63213=>"100000101",
  63214=>"000000000",
  63215=>"000000100",
  63216=>"000010000",
  63217=>"111111011",
  63218=>"000000000",
  63219=>"011011011",
  63220=>"000111000",
  63221=>"111111000",
  63222=>"000100000",
  63223=>"000000001",
  63224=>"000000000",
  63225=>"110000000",
  63226=>"010111111",
  63227=>"011011000",
  63228=>"000101000",
  63229=>"111010100",
  63230=>"000001111",
  63231=>"000100100",
  63232=>"100110011",
  63233=>"011000010",
  63234=>"100101111",
  63235=>"111010010",
  63236=>"001001101",
  63237=>"110000001",
  63238=>"001011101",
  63239=>"000011111",
  63240=>"100110010",
  63241=>"001001000",
  63242=>"100100000",
  63243=>"100100100",
  63244=>"100100110",
  63245=>"111110000",
  63246=>"001101101",
  63247=>"000010010",
  63248=>"110111001",
  63249=>"001111001",
  63250=>"100000000",
  63251=>"000000011",
  63252=>"011001010",
  63253=>"111110110",
  63254=>"001010000",
  63255=>"000111110",
  63256=>"011000000",
  63257=>"001001001",
  63258=>"000011000",
  63259=>"001011111",
  63260=>"100101101",
  63261=>"011010000",
  63262=>"100000101",
  63263=>"100110110",
  63264=>"111000111",
  63265=>"110110100",
  63266=>"000010100",
  63267=>"000100100",
  63268=>"011111111",
  63269=>"111110010",
  63270=>"011000001",
  63271=>"000111011",
  63272=>"001011010",
  63273=>"010000111",
  63274=>"000010110",
  63275=>"101100000",
  63276=>"111100010",
  63277=>"011000000",
  63278=>"001100111",
  63279=>"100010000",
  63280=>"011000001",
  63281=>"101100100",
  63282=>"000011011",
  63283=>"001011011",
  63284=>"110100000",
  63285=>"011010000",
  63286=>"000010110",
  63287=>"000011111",
  63288=>"110100100",
  63289=>"011011111",
  63290=>"001001100",
  63291=>"011111111",
  63292=>"100000001",
  63293=>"010110100",
  63294=>"100100000",
  63295=>"011110010",
  63296=>"100100111",
  63297=>"111100011",
  63298=>"101111111",
  63299=>"100100111",
  63300=>"111100000",
  63301=>"000000111",
  63302=>"000001011",
  63303=>"011111111",
  63304=>"100110110",
  63305=>"000010000",
  63306=>"110100111",
  63307=>"100100110",
  63308=>"100100110",
  63309=>"111111101",
  63310=>"100110110",
  63311=>"111111011",
  63312=>"100000111",
  63313=>"110100000",
  63314=>"011011111",
  63315=>"001000000",
  63316=>"011101110",
  63317=>"110000110",
  63318=>"100001101",
  63319=>"001001101",
  63320=>"111000000",
  63321=>"001000000",
  63322=>"000000110",
  63323=>"001111111",
  63324=>"000000001",
  63325=>"000000000",
  63326=>"111111111",
  63327=>"000000101",
  63328=>"000000000",
  63329=>"111000000",
  63330=>"100100110",
  63331=>"111111111",
  63332=>"110010010",
  63333=>"011101100",
  63334=>"011010011",
  63335=>"011000011",
  63336=>"001100111",
  63337=>"001011011",
  63338=>"000011011",
  63339=>"100100000",
  63340=>"000000111",
  63341=>"011011000",
  63342=>"000001001",
  63343=>"000011011",
  63344=>"011011100",
  63345=>"001111101",
  63346=>"100110001",
  63347=>"011111000",
  63348=>"001011010",
  63349=>"100100000",
  63350=>"100011101",
  63351=>"110100111",
  63352=>"100100110",
  63353=>"000011111",
  63354=>"001111110",
  63355=>"011110110",
  63356=>"100001001",
  63357=>"110100100",
  63358=>"100100100",
  63359=>"100100100",
  63360=>"100100010",
  63361=>"110100110",
  63362=>"000001011",
  63363=>"001010000",
  63364=>"000111011",
  63365=>"010000000",
  63366=>"101001011",
  63367=>"100100100",
  63368=>"011101011",
  63369=>"011011010",
  63370=>"001001000",
  63371=>"000001111",
  63372=>"100111000",
  63373=>"101111000",
  63374=>"011100100",
  63375=>"001011000",
  63376=>"001011000",
  63377=>"110110000",
  63378=>"100110000",
  63379=>"110110001",
  63380=>"010010000",
  63381=>"100100111",
  63382=>"000001000",
  63383=>"111110110",
  63384=>"000100100",
  63385=>"110110100",
  63386=>"110100100",
  63387=>"000101111",
  63388=>"011111101",
  63389=>"100110111",
  63390=>"000000110",
  63391=>"100000000",
  63392=>"001000100",
  63393=>"111101011",
  63394=>"100000110",
  63395=>"100000001",
  63396=>"000000111",
  63397=>"111001011",
  63398=>"010010000",
  63399=>"000000011",
  63400=>"001011011",
  63401=>"000000000",
  63402=>"110110111",
  63403=>"100100100",
  63404=>"110100000",
  63405=>"110100001",
  63406=>"110000111",
  63407=>"000001000",
  63408=>"100000011",
  63409=>"000001001",
  63410=>"110100100",
  63411=>"100100001",
  63412=>"001010000",
  63413=>"011101100",
  63414=>"000001001",
  63415=>"010111001",
  63416=>"110110110",
  63417=>"101111000",
  63418=>"111111000",
  63419=>"100100110",
  63420=>"011011001",
  63421=>"100100110",
  63422=>"001001111",
  63423=>"001011001",
  63424=>"111110111",
  63425=>"000001001",
  63426=>"001111011",
  63427=>"101111010",
  63428=>"011011100",
  63429=>"100110111",
  63430=>"111011000",
  63431=>"110100010",
  63432=>"000001001",
  63433=>"100110110",
  63434=>"011011001",
  63435=>"001111101",
  63436=>"011011010",
  63437=>"010110110",
  63438=>"100110111",
  63439=>"100110110",
  63440=>"001111111",
  63441=>"110110000",
  63442=>"000001001",
  63443=>"011000000",
  63444=>"110100111",
  63445=>"000000010",
  63446=>"100101111",
  63447=>"000000001",
  63448=>"000110111",
  63449=>"000010000",
  63450=>"111110100",
  63451=>"001011001",
  63452=>"100100111",
  63453=>"111011000",
  63454=>"010011011",
  63455=>"110111001",
  63456=>"100110110",
  63457=>"101000111",
  63458=>"000000110",
  63459=>"111101011",
  63460=>"011011000",
  63461=>"100000011",
  63462=>"011011011",
  63463=>"001001111",
  63464=>"001000111",
  63465=>"011000010",
  63466=>"000001001",
  63467=>"000001001",
  63468=>"110110111",
  63469=>"011010000",
  63470=>"100000000",
  63471=>"100001000",
  63472=>"001111111",
  63473=>"000001110",
  63474=>"000011111",
  63475=>"111100000",
  63476=>"011000010",
  63477=>"000011010",
  63478=>"001100001",
  63479=>"011100101",
  63480=>"100100110",
  63481=>"010000011",
  63482=>"111111101",
  63483=>"011011010",
  63484=>"011000000",
  63485=>"000000001",
  63486=>"011111111",
  63487=>"111101101",
  63488=>"100110110",
  63489=>"000010000",
  63490=>"011000000",
  63491=>"001100100",
  63492=>"000000001",
  63493=>"000010001",
  63494=>"111001110",
  63495=>"000000000",
  63496=>"000000000",
  63497=>"000100111",
  63498=>"100111111",
  63499=>"000010111",
  63500=>"011111011",
  63501=>"101000111",
  63502=>"011110110",
  63503=>"101010000",
  63504=>"000011111",
  63505=>"111110110",
  63506=>"111011011",
  63507=>"000000001",
  63508=>"001100111",
  63509=>"000011000",
  63510=>"111111001",
  63511=>"101101101",
  63512=>"000000101",
  63513=>"000000001",
  63514=>"000111111",
  63515=>"111100100",
  63516=>"111010101",
  63517=>"000111111",
  63518=>"000010011",
  63519=>"100111111",
  63520=>"111101101",
  63521=>"000111010",
  63522=>"111100111",
  63523=>"000111101",
  63524=>"001001010",
  63525=>"000011010",
  63526=>"000000000",
  63527=>"000000000",
  63528=>"010101110",
  63529=>"111101010",
  63530=>"111110111",
  63531=>"111111111",
  63532=>"001111111",
  63533=>"000111001",
  63534=>"011111000",
  63535=>"111111101",
  63536=>"000100100",
  63537=>"000111000",
  63538=>"111101101",
  63539=>"111111011",
  63540=>"010000110",
  63541=>"000000000",
  63542=>"010110110",
  63543=>"000010110",
  63544=>"000110111",
  63545=>"101000100",
  63546=>"000000000",
  63547=>"111111111",
  63548=>"101111111",
  63549=>"111111111",
  63550=>"101000111",
  63551=>"001100111",
  63552=>"000111010",
  63553=>"000111010",
  63554=>"111010110",
  63555=>"110111110",
  63556=>"000100111",
  63557=>"000111111",
  63558=>"101000100",
  63559=>"001111000",
  63560=>"001011111",
  63561=>"000000010",
  63562=>"001011000",
  63563=>"010010111",
  63564=>"111111100",
  63565=>"100001011",
  63566=>"001100110",
  63567=>"000111010",
  63568=>"111111100",
  63569=>"010111100",
  63570=>"000000001",
  63571=>"000010011",
  63572=>"000000000",
  63573=>"011111110",
  63574=>"000110100",
  63575=>"010101000",
  63576=>"010000011",
  63577=>"111000010",
  63578=>"110011111",
  63579=>"101110111",
  63580=>"001100100",
  63581=>"100100100",
  63582=>"000000000",
  63583=>"011001011",
  63584=>"111111111",
  63585=>"110110110",
  63586=>"000111011",
  63587=>"111101001",
  63588=>"000000110",
  63589=>"111100000",
  63590=>"000000000",
  63591=>"100101110",
  63592=>"000100100",
  63593=>"111001011",
  63594=>"010100000",
  63595=>"000010100",
  63596=>"101000000",
  63597=>"100000110",
  63598=>"000000000",
  63599=>"000110011",
  63600=>"011011111",
  63601=>"010000000",
  63602=>"000011111",
  63603=>"100111111",
  63604=>"101110110",
  63605=>"010010110",
  63606=>"100000111",
  63607=>"000000011",
  63608=>"011000110",
  63609=>"100000000",
  63610=>"010110111",
  63611=>"000100111",
  63612=>"010001000",
  63613=>"001011010",
  63614=>"000111010",
  63615=>"110100110",
  63616=>"001111111",
  63617=>"010010010",
  63618=>"000000000",
  63619=>"000111011",
  63620=>"001111111",
  63621=>"111111101",
  63622=>"100110111",
  63623=>"111110000",
  63624=>"101110101",
  63625=>"111001001",
  63626=>"000000000",
  63627=>"011110000",
  63628=>"001101100",
  63629=>"000000000",
  63630=>"000000101",
  63631=>"001000001",
  63632=>"011011011",
  63633=>"010110010",
  63634=>"101000111",
  63635=>"010001001",
  63636=>"000100100",
  63637=>"111100000",
  63638=>"011010010",
  63639=>"110111111",
  63640=>"111101111",
  63641=>"010000010",
  63642=>"011011010",
  63643=>"010011010",
  63644=>"110100000",
  63645=>"100010011",
  63646=>"111101101",
  63647=>"111010001",
  63648=>"111011001",
  63649=>"110110000",
  63650=>"011111011",
  63651=>"011000000",
  63652=>"100000000",
  63653=>"011011111",
  63654=>"001011011",
  63655=>"101000110",
  63656=>"011011111",
  63657=>"111101100",
  63658=>"000000010",
  63659=>"101110101",
  63660=>"011110011",
  63661=>"000101101",
  63662=>"101010000",
  63663=>"110111011",
  63664=>"011011000",
  63665=>"111001100",
  63666=>"000100111",
  63667=>"111011011",
  63668=>"000011110",
  63669=>"000101010",
  63670=>"010011100",
  63671=>"000100110",
  63672=>"100100000",
  63673=>"001001001",
  63674=>"000000000",
  63675=>"000101111",
  63676=>"101111111",
  63677=>"100010110",
  63678=>"110100110",
  63679=>"100101000",
  63680=>"111001000",
  63681=>"000111010",
  63682=>"001100000",
  63683=>"111001101",
  63684=>"101101101",
  63685=>"010001111",
  63686=>"111100000",
  63687=>"100111011",
  63688=>"000000000",
  63689=>"111010111",
  63690=>"101001001",
  63691=>"000000000",
  63692=>"000000010",
  63693=>"100000000",
  63694=>"000110110",
  63695=>"000111011",
  63696=>"101100111",
  63697=>"111111111",
  63698=>"101001000",
  63699=>"101001111",
  63700=>"010010010",
  63701=>"001001000",
  63702=>"111111011",
  63703=>"000110111",
  63704=>"000000100",
  63705=>"000001001",
  63706=>"111111001",
  63707=>"111000101",
  63708=>"110111110",
  63709=>"111111100",
  63710=>"000000000",
  63711=>"100110111",
  63712=>"000001001",
  63713=>"000100010",
  63714=>"000000000",
  63715=>"000011000",
  63716=>"011000101",
  63717=>"101100000",
  63718=>"110000001",
  63719=>"000000010",
  63720=>"011111100",
  63721=>"001000000",
  63722=>"001000111",
  63723=>"000100000",
  63724=>"011000000",
  63725=>"000001001",
  63726=>"110111101",
  63727=>"000000000",
  63728=>"010010000",
  63729=>"011100110",
  63730=>"011010111",
  63731=>"000000111",
  63732=>"001011011",
  63733=>"011011000",
  63734=>"111011011",
  63735=>"101010010",
  63736=>"000000000",
  63737=>"111111111",
  63738=>"101100111",
  63739=>"100010100",
  63740=>"101000101",
  63741=>"101101110",
  63742=>"100100100",
  63743=>"111111111",
  63744=>"011001000",
  63745=>"110110110",
  63746=>"001100011",
  63747=>"100010110",
  63748=>"001011111",
  63749=>"100010010",
  63750=>"111011001",
  63751=>"010111001",
  63752=>"000000010",
  63753=>"100110100",
  63754=>"111100001",
  63755=>"010001111",
  63756=>"111110110",
  63757=>"111000000",
  63758=>"101011101",
  63759=>"011101111",
  63760=>"110010010",
  63761=>"100110000",
  63762=>"001001001",
  63763=>"000110110",
  63764=>"001111101",
  63765=>"100111110",
  63766=>"111001011",
  63767=>"001111001",
  63768=>"101001001",
  63769=>"101101001",
  63770=>"111111110",
  63771=>"110110110",
  63772=>"001001001",
  63773=>"111000011",
  63774=>"110100110",
  63775=>"001000001",
  63776=>"001100100",
  63777=>"101001101",
  63778=>"011011000",
  63779=>"100110110",
  63780=>"001011011",
  63781=>"001001011",
  63782=>"110110110",
  63783=>"110110100",
  63784=>"001011001",
  63785=>"000000000",
  63786=>"110110100",
  63787=>"110011110",
  63788=>"101111111",
  63789=>"001110111",
  63790=>"110000010",
  63791=>"001001011",
  63792=>"111001101",
  63793=>"001101001",
  63794=>"110101111",
  63795=>"110010100",
  63796=>"100010100",
  63797=>"010110000",
  63798=>"100110110",
  63799=>"110110100",
  63800=>"110100000",
  63801=>"100000001",
  63802=>"001001001",
  63803=>"110010100",
  63804=>"100111100",
  63805=>"001001011",
  63806=>"100010010",
  63807=>"010000000",
  63808=>"110101111",
  63809=>"111110110",
  63810=>"111111001",
  63811=>"111110100",
  63812=>"001001011",
  63813=>"010000000",
  63814=>"001111111",
  63815=>"111000000",
  63816=>"111011110",
  63817=>"000111110",
  63818=>"100010000",
  63819=>"000000100",
  63820=>"110110110",
  63821=>"011001001",
  63822=>"001001000",
  63823=>"011001111",
  63824=>"011010001",
  63825=>"000001000",
  63826=>"110111111",
  63827=>"111001001",
  63828=>"000000011",
  63829=>"110110110",
  63830=>"011001001",
  63831=>"100000000",
  63832=>"100000010",
  63833=>"001011111",
  63834=>"000100101",
  63835=>"101000100",
  63836=>"110110110",
  63837=>"001001011",
  63838=>"110110110",
  63839=>"110110111",
  63840=>"110110110",
  63841=>"100110110",
  63842=>"101110111",
  63843=>"001001111",
  63844=>"001000000",
  63845=>"101010100",
  63846=>"100001000",
  63847=>"110000000",
  63848=>"110110100",
  63849=>"010100101",
  63850=>"110110111",
  63851=>"010110111",
  63852=>"011011110",
  63853=>"001101001",
  63854=>"000000110",
  63855=>"011011110",
  63856=>"011101011",
  63857=>"110110111",
  63858=>"110100100",
  63859=>"001011011",
  63860=>"110110110",
  63861=>"001100000",
  63862=>"100100111",
  63863=>"110110110",
  63864=>"110110010",
  63865=>"001001111",
  63866=>"001001100",
  63867=>"001001001",
  63868=>"010010010",
  63869=>"100000000",
  63870=>"110000001",
  63871=>"110000001",
  63872=>"010000000",
  63873=>"000000110",
  63874=>"110110110",
  63875=>"000010110",
  63876=>"111000100",
  63877=>"001101011",
  63878=>"001011010",
  63879=>"000100001",
  63880=>"001011011",
  63881=>"010110110",
  63882=>"011111001",
  63883=>"000110111",
  63884=>"011011001",
  63885=>"100100111",
  63886=>"111101101",
  63887=>"010000110",
  63888=>"101001001",
  63889=>"001101111",
  63890=>"011010111",
  63891=>"110101110",
  63892=>"000101010",
  63893=>"100110110",
  63894=>"001111101",
  63895=>"001011111",
  63896=>"001011100",
  63897=>"111000111",
  63898=>"101001101",
  63899=>"010000010",
  63900=>"000111100",
  63901=>"110110100",
  63902=>"110110110",
  63903=>"001000000",
  63904=>"001001001",
  63905=>"001001010",
  63906=>"011010001",
  63907=>"101111111",
  63908=>"110000111",
  63909=>"000001000",
  63910=>"010001011",
  63911=>"101101011",
  63912=>"110010010",
  63913=>"000110110",
  63914=>"001001000",
  63915=>"000010010",
  63916=>"011001000",
  63917=>"011011110",
  63918=>"000010010",
  63919=>"000000000",
  63920=>"011111000",
  63921=>"111110010",
  63922=>"001001001",
  63923=>"000000000",
  63924=>"001110000",
  63925=>"111111111",
  63926=>"111111000",
  63927=>"001011111",
  63928=>"011001001",
  63929=>"111001111",
  63930=>"111101001",
  63931=>"110111000",
  63932=>"000000000",
  63933=>"001011011",
  63934=>"011111111",
  63935=>"110000001",
  63936=>"001011011",
  63937=>"110110110",
  63938=>"010111111",
  63939=>"011011000",
  63940=>"001001001",
  63941=>"000000111",
  63942=>"101111111",
  63943=>"101101101",
  63944=>"010001001",
  63945=>"011001000",
  63946=>"110101100",
  63947=>"110010110",
  63948=>"001011011",
  63949=>"111111111",
  63950=>"110110100",
  63951=>"111110000",
  63952=>"001001001",
  63953=>"010001000",
  63954=>"110011011",
  63955=>"001001001",
  63956=>"101100111",
  63957=>"100110101",
  63958=>"100101110",
  63959=>"110110110",
  63960=>"000001011",
  63961=>"010010110",
  63962=>"001001000",
  63963=>"001111001",
  63964=>"111111000",
  63965=>"111011001",
  63966=>"011001001",
  63967=>"110110110",
  63968=>"000010010",
  63969=>"000000100",
  63970=>"110000000",
  63971=>"001101001",
  63972=>"011110110",
  63973=>"110011011",
  63974=>"011000000",
  63975=>"111101110",
  63976=>"111000110",
  63977=>"111010010",
  63978=>"101101001",
  63979=>"001001001",
  63980=>"000110110",
  63981=>"010111111",
  63982=>"001001011",
  63983=>"001000100",
  63984=>"010100111",
  63985=>"111011001",
  63986=>"110010100",
  63987=>"111111000",
  63988=>"000001111",
  63989=>"100100111",
  63990=>"000100110",
  63991=>"010110000",
  63992=>"100110111",
  63993=>"100101110",
  63994=>"101101001",
  63995=>"111011101",
  63996=>"011011011",
  63997=>"001001001",
  63998=>"001001101",
  63999=>"001011000",
  64000=>"001001101",
  64001=>"100111111",
  64002=>"000000100",
  64003=>"000000110",
  64004=>"001001000",
  64005=>"000100000",
  64006=>"000000111",
  64007=>"011000000",
  64008=>"010100111",
  64009=>"111111100",
  64010=>"000000000",
  64011=>"000100111",
  64012=>"100000111",
  64013=>"000101111",
  64014=>"000000011",
  64015=>"100111111",
  64016=>"111110000",
  64017=>"101000000",
  64018=>"111101111",
  64019=>"111001000",
  64020=>"011111111",
  64021=>"100000000",
  64022=>"011011001",
  64023=>"000111111",
  64024=>"000000011",
  64025=>"001101001",
  64026=>"000000010",
  64027=>"011011000",
  64028=>"000000010",
  64029=>"000100000",
  64030=>"100100111",
  64031=>"111010000",
  64032=>"000000101",
  64033=>"110101111",
  64034=>"111111001",
  64035=>"010000000",
  64036=>"011011011",
  64037=>"000001001",
  64038=>"011111000",
  64039=>"010011101",
  64040=>"111111000",
  64041=>"111111101",
  64042=>"100110100",
  64043=>"011000000",
  64044=>"110100110",
  64045=>"100111111",
  64046=>"101101101",
  64047=>"100100000",
  64048=>"000100111",
  64049=>"011010100",
  64050=>"100110111",
  64051=>"111000000",
  64052=>"000000000",
  64053=>"111101000",
  64054=>"011011011",
  64055=>"101111111",
  64056=>"001000100",
  64057=>"000000101",
  64058=>"100001011",
  64059=>"010111000",
  64060=>"110011111",
  64061=>"110111110",
  64062=>"000100111",
  64063=>"110111010",
  64064=>"011000101",
  64065=>"100001010",
  64066=>"110000101",
  64067=>"010010100",
  64068=>"111100000",
  64069=>"100100110",
  64070=>"000100101",
  64071=>"011001011",
  64072=>"001010101",
  64073=>"000000101",
  64074=>"000000000",
  64075=>"100100110",
  64076=>"100000000",
  64077=>"110100100",
  64078=>"111011000",
  64079=>"101101111",
  64080=>"100000001",
  64081=>"010001000",
  64082=>"000101110",
  64083=>"001000000",
  64084=>"000000000",
  64085=>"110011011",
  64086=>"101110011",
  64087=>"000000010",
  64088=>"111111110",
  64089=>"110000111",
  64090=>"011111100",
  64091=>"111110000",
  64092=>"000000011",
  64093=>"000000111",
  64094=>"011011000",
  64095=>"011010001",
  64096=>"111111011",
  64097=>"110101101",
  64098=>"000000111",
  64099=>"110101100",
  64100=>"100000011",
  64101=>"111101000",
  64102=>"000000011",
  64103=>"011000000",
  64104=>"111111111",
  64105=>"111000100",
  64106=>"111000000",
  64107=>"000000001",
  64108=>"111011111",
  64109=>"000000011",
  64110=>"111111001",
  64111=>"001001111",
  64112=>"101111000",
  64113=>"100111111",
  64114=>"000010110",
  64115=>"011000000",
  64116=>"000000111",
  64117=>"100000000",
  64118=>"001000100",
  64119=>"001000001",
  64120=>"000100000",
  64121=>"011000110",
  64122=>"111111111",
  64123=>"101100000",
  64124=>"111110011",
  64125=>"100100000",
  64126=>"010010001",
  64127=>"000000100",
  64128=>"111111000",
  64129=>"100001110",
  64130=>"111000011",
  64131=>"111001100",
  64132=>"101100000",
  64133=>"101101110",
  64134=>"100000000",
  64135=>"010100000",
  64136=>"100100110",
  64137=>"000000000",
  64138=>"000000000",
  64139=>"111000011",
  64140=>"000110000",
  64141=>"000000000",
  64142=>"100000111",
  64143=>"000000000",
  64144=>"110011011",
  64145=>"111111111",
  64146=>"000110010",
  64147=>"101100101",
  64148=>"100100100",
  64149=>"000100000",
  64150=>"000111111",
  64151=>"001001010",
  64152=>"000001111",
  64153=>"000000111",
  64154=>"101100111",
  64155=>"000100111",
  64156=>"111100101",
  64157=>"111100001",
  64158=>"000111011",
  64159=>"011010011",
  64160=>"100111111",
  64161=>"000010110",
  64162=>"111001000",
  64163=>"000000101",
  64164=>"100101110",
  64165=>"011001100",
  64166=>"110110000",
  64167=>"110100000",
  64168=>"100101111",
  64169=>"100011010",
  64170=>"111011010",
  64171=>"010110110",
  64172=>"111100010",
  64173=>"000000101",
  64174=>"011001001",
  64175=>"011000011",
  64176=>"000100011",
  64177=>"110000001",
  64178=>"000000010",
  64179=>"110010111",
  64180=>"001000101",
  64181=>"000000111",
  64182=>"111110100",
  64183=>"100100001",
  64184=>"011100001",
  64185=>"001111110",
  64186=>"001111001",
  64187=>"100000000",
  64188=>"000000000",
  64189=>"111111111",
  64190=>"111101001",
  64191=>"010011100",
  64192=>"100000101",
  64193=>"100000111",
  64194=>"000010011",
  64195=>"000000011",
  64196=>"000101111",
  64197=>"101101111",
  64198=>"110100110",
  64199=>"011000000",
  64200=>"111111111",
  64201=>"011011010",
  64202=>"101111111",
  64203=>"100101111",
  64204=>"001100110",
  64205=>"111111000",
  64206=>"101010011",
  64207=>"011111111",
  64208=>"010000000",
  64209=>"110000100",
  64210=>"111101101",
  64211=>"111111011",
  64212=>"011000000",
  64213=>"101100110",
  64214=>"000000111",
  64215=>"000101111",
  64216=>"011010000",
  64217=>"101100110",
  64218=>"111101111",
  64219=>"000000100",
  64220=>"111011100",
  64221=>"111000010",
  64222=>"110100011",
  64223=>"000000000",
  64224=>"000010010",
  64225=>"000100101",
  64226=>"010010000",
  64227=>"000010110",
  64228=>"100000000",
  64229=>"111011100",
  64230=>"001000000",
  64231=>"001100101",
  64232=>"111100000",
  64233=>"001001001",
  64234=>"100100000",
  64235=>"100000101",
  64236=>"111111000",
  64237=>"111111000",
  64238=>"100000000",
  64239=>"101011111",
  64240=>"111111000",
  64241=>"110101111",
  64242=>"101000000",
  64243=>"110000100",
  64244=>"000100100",
  64245=>"010000001",
  64246=>"000000000",
  64247=>"011001111",
  64248=>"000011111",
  64249=>"111100110",
  64250=>"100000010",
  64251=>"000101101",
  64252=>"110110111",
  64253=>"101000000",
  64254=>"000000001",
  64255=>"000000000",
  64256=>"100101101",
  64257=>"111000010",
  64258=>"010010000",
  64259=>"100000000",
  64260=>"111111110",
  64261=>"111101101",
  64262=>"101111110",
  64263=>"110100000",
  64264=>"111110111",
  64265=>"000000100",
  64266=>"100100011",
  64267=>"000000000",
  64268=>"111000100",
  64269=>"000001101",
  64270=>"000100011",
  64271=>"111101111",
  64272=>"000110111",
  64273=>"000000011",
  64274=>"000000011",
  64275=>"111000100",
  64276=>"000010000",
  64277=>"111110111",
  64278=>"111111011",
  64279=>"101111011",
  64280=>"101000011",
  64281=>"000000001",
  64282=>"111000011",
  64283=>"000000000",
  64284=>"101100000",
  64285=>"111111111",
  64286=>"000001110",
  64287=>"000000001",
  64288=>"111011000",
  64289=>"000000000",
  64290=>"110000101",
  64291=>"101000111",
  64292=>"000110010",
  64293=>"001001000",
  64294=>"110010010",
  64295=>"000000000",
  64296=>"111111010",
  64297=>"000000011",
  64298=>"000000101",
  64299=>"110001000",
  64300=>"010010001",
  64301=>"111000111",
  64302=>"110000101",
  64303=>"000000000",
  64304=>"111011000",
  64305=>"011101111",
  64306=>"011011011",
  64307=>"000110100",
  64308=>"100101111",
  64309=>"101101111",
  64310=>"010011011",
  64311=>"000100001",
  64312=>"110101100",
  64313=>"000000001",
  64314=>"011000000",
  64315=>"010000000",
  64316=>"001000001",
  64317=>"111111111",
  64318=>"101000001",
  64319=>"111101101",
  64320=>"110100010",
  64321=>"111000010",
  64322=>"000100100",
  64323=>"100001101",
  64324=>"101100100",
  64325=>"000000001",
  64326=>"101101111",
  64327=>"111001101",
  64328=>"001110010",
  64329=>"100000000",
  64330=>"101100000",
  64331=>"101010010",
  64332=>"010000000",
  64333=>"100100111",
  64334=>"101011111",
  64335=>"000100000",
  64336=>"100101101",
  64337=>"111111000",
  64338=>"100000000",
  64339=>"110001000",
  64340=>"111111000",
  64341=>"100111111",
  64342=>"000011011",
  64343=>"000000100",
  64344=>"001000101",
  64345=>"000000001",
  64346=>"011101011",
  64347=>"010011111",
  64348=>"011000100",
  64349=>"010110100",
  64350=>"000111010",
  64351=>"101000110",
  64352=>"111100101",
  64353=>"000000000",
  64354=>"100000100",
  64355=>"011011001",
  64356=>"001001001",
  64357=>"000010111",
  64358=>"000000000",
  64359=>"100111011",
  64360=>"000000101",
  64361=>"100111010",
  64362=>"111010010",
  64363=>"000000000",
  64364=>"000000000",
  64365=>"000111011",
  64366=>"000000000",
  64367=>"000000111",
  64368=>"100100110",
  64369=>"000000010",
  64370=>"110010110",
  64371=>"000001010",
  64372=>"111110000",
  64373=>"000101101",
  64374=>"111000101",
  64375=>"000000000",
  64376=>"111111000",
  64377=>"100101010",
  64378=>"000110111",
  64379=>"111101111",
  64380=>"001111110",
  64381=>"011011001",
  64382=>"011011111",
  64383=>"101000101",
  64384=>"000000101",
  64385=>"000000000",
  64386=>"000000110",
  64387=>"000000100",
  64388=>"000101000",
  64389=>"110011000",
  64390=>"100100010",
  64391=>"000000000",
  64392=>"000000000",
  64393=>"000000100",
  64394=>"100111010",
  64395=>"001101010",
  64396=>"000111101",
  64397=>"111100101",
  64398=>"111101000",
  64399=>"000000101",
  64400=>"101000000",
  64401=>"111111111",
  64402=>"011011101",
  64403=>"111111100",
  64404=>"000100000",
  64405=>"101101110",
  64406=>"101000000",
  64407=>"011111101",
  64408=>"111101101",
  64409=>"111011011",
  64410=>"111010000",
  64411=>"010000000",
  64412=>"101000000",
  64413=>"000100000",
  64414=>"111111110",
  64415=>"101100101",
  64416=>"110111011",
  64417=>"011011111",
  64418=>"111000001",
  64419=>"000000000",
  64420=>"000010111",
  64421=>"011100001",
  64422=>"010010000",
  64423=>"011100000",
  64424=>"000101110",
  64425=>"111001100",
  64426=>"111000100",
  64427=>"101000100",
  64428=>"000001001",
  64429=>"111000000",
  64430=>"011111111",
  64431=>"000000101",
  64432=>"111000101",
  64433=>"000000100",
  64434=>"011101101",
  64435=>"000100110",
  64436=>"011001000",
  64437=>"111100111",
  64438=>"000000100",
  64439=>"000011100",
  64440=>"000100100",
  64441=>"001001011",
  64442=>"011111111",
  64443=>"011011000",
  64444=>"100111000",
  64445=>"000000000",
  64446=>"111100111",
  64447=>"000111111",
  64448=>"000100100",
  64449=>"000000000",
  64450=>"000111011",
  64451=>"010000100",
  64452=>"000000001",
  64453=>"011000010",
  64454=>"000000000",
  64455=>"111000000",
  64456=>"111101111",
  64457=>"000000000",
  64458=>"000101111",
  64459=>"100000000",
  64460=>"111111011",
  64461=>"110100001",
  64462=>"100000000",
  64463=>"000111011",
  64464=>"000010010",
  64465=>"100001000",
  64466=>"000000000",
  64467=>"001111011",
  64468=>"000000000",
  64469=>"101101001",
  64470=>"111000000",
  64471=>"011111011",
  64472=>"111011111",
  64473=>"000010111",
  64474=>"011110111",
  64475=>"111110000",
  64476=>"111111110",
  64477=>"001111100",
  64478=>"000000100",
  64479=>"000110110",
  64480=>"010000010",
  64481=>"000000011",
  64482=>"111111111",
  64483=>"001101110",
  64484=>"001011010",
  64485=>"000100101",
  64486=>"000000100",
  64487=>"100110100",
  64488=>"011011000",
  64489=>"111111100",
  64490=>"001011111",
  64491=>"101000100",
  64492=>"001000110",
  64493=>"000100000",
  64494=>"111111001",
  64495=>"111000001",
  64496=>"000000010",
  64497=>"110100001",
  64498=>"100101100",
  64499=>"110110101",
  64500=>"001111011",
  64501=>"110011110",
  64502=>"000000001",
  64503=>"000111111",
  64504=>"000100010",
  64505=>"011010110",
  64506=>"111000111",
  64507=>"000110011",
  64508=>"111011011",
  64509=>"100010111",
  64510=>"111010000",
  64511=>"100000100",
  64512=>"100101000",
  64513=>"000000100",
  64514=>"111000001",
  64515=>"011000000",
  64516=>"010111011",
  64517=>"000000111",
  64518=>"111111000",
  64519=>"110111111",
  64520=>"100110110",
  64521=>"010000001",
  64522=>"100000001",
  64523=>"100100101",
  64524=>"000110010",
  64525=>"000010111",
  64526=>"000001100",
  64527=>"111111000",
  64528=>"010000000",
  64529=>"010000000",
  64530=>"110111000",
  64531=>"000000111",
  64532=>"111000111",
  64533=>"111000000",
  64534=>"111101100",
  64535=>"110111011",
  64536=>"010111010",
  64537=>"001000000",
  64538=>"111000000",
  64539=>"000000010",
  64540=>"010000010",
  64541=>"001101000",
  64542=>"000000000",
  64543=>"001001000",
  64544=>"111111001",
  64545=>"101010010",
  64546=>"000101101",
  64547=>"001111001",
  64548=>"010011001",
  64549=>"111000111",
  64550=>"111101000",
  64551=>"011011000",
  64552=>"111100000",
  64553=>"010000001",
  64554=>"101101000",
  64555=>"000000000",
  64556=>"010111101",
  64557=>"111000111",
  64558=>"100111001",
  64559=>"000110110",
  64560=>"111000110",
  64561=>"100111011",
  64562=>"101101000",
  64563=>"000000100",
  64564=>"001001000",
  64565=>"001101101",
  64566=>"000100000",
  64567=>"010000001",
  64568=>"110110100",
  64569=>"001001000",
  64570=>"000101101",
  64571=>"000010100",
  64572=>"001110111",
  64573=>"010111111",
  64574=>"101001101",
  64575=>"111011111",
  64576=>"000101111",
  64577=>"010111101",
  64578=>"010010001",
  64579=>"010111001",
  64580=>"111101000",
  64581=>"101000001",
  64582=>"010110111",
  64583=>"000111101",
  64584=>"011001101",
  64585=>"101010010",
  64586=>"000001011",
  64587=>"111001000",
  64588=>"111101001",
  64589=>"011011011",
  64590=>"110111110",
  64591=>"101111010",
  64592=>"111100000",
  64593=>"110111111",
  64594=>"111101001",
  64595=>"000001000",
  64596=>"000000000",
  64597=>"011000000",
  64598=>"100100000",
  64599=>"010000000",
  64600=>"111011000",
  64601=>"000110001",
  64602=>"111111000",
  64603=>"110110111",
  64604=>"110111001",
  64605=>"100110100",
  64606=>"010011110",
  64607=>"000000001",
  64608=>"101100000",
  64609=>"110100000",
  64610=>"000010010",
  64611=>"111111001",
  64612=>"000000000",
  64613=>"000001101",
  64614=>"000000111",
  64615=>"001001100",
  64616=>"110000010",
  64617=>"000111111",
  64618=>"111111101",
  64619=>"010111001",
  64620=>"111111001",
  64621=>"011100110",
  64622=>"000000011",
  64623=>"110000110",
  64624=>"011110110",
  64625=>"010111111",
  64626=>"010000000",
  64627=>"000000001",
  64628=>"000001110",
  64629=>"111001101",
  64630=>"101000010",
  64631=>"101111001",
  64632=>"010111110",
  64633=>"101110101",
  64634=>"101101000",
  64635=>"000000111",
  64636=>"001000100",
  64637=>"010000001",
  64638=>"011110100",
  64639=>"111000000",
  64640=>"000011011",
  64641=>"011111000",
  64642=>"010110110",
  64643=>"000111111",
  64644=>"001010111",
  64645=>"011011101",
  64646=>"110111111",
  64647=>"111000000",
  64648=>"100011011",
  64649=>"111000111",
  64650=>"111100100",
  64651=>"010000111",
  64652=>"000000001",
  64653=>"111111101",
  64654=>"011000001",
  64655=>"100001000",
  64656=>"001111110",
  64657=>"000011111",
  64658=>"000000101",
  64659=>"101100000",
  64660=>"111000110",
  64661=>"000110001",
  64662=>"111111111",
  64663=>"100111100",
  64664=>"101100001",
  64665=>"000101000",
  64666=>"000000011",
  64667=>"000010010",
  64668=>"011101000",
  64669=>"110110110",
  64670=>"011001000",
  64671=>"111101001",
  64672=>"011101111",
  64673=>"111101011",
  64674=>"000111101",
  64675=>"111100000",
  64676=>"000000001",
  64677=>"010000011",
  64678=>"111011001",
  64679=>"000000000",
  64680=>"000000000",
  64681=>"111000000",
  64682=>"000010110",
  64683=>"111001001",
  64684=>"110101110",
  64685=>"111101100",
  64686=>"101011001",
  64687=>"111000000",
  64688=>"100111111",
  64689=>"110110000",
  64690=>"110100000",
  64691=>"000000100",
  64692=>"101111110",
  64693=>"001001011",
  64694=>"111101100",
  64695=>"001011010",
  64696=>"100011011",
  64697=>"111000001",
  64698=>"000111110",
  64699=>"011010010",
  64700=>"001001011",
  64701=>"111111111",
  64702=>"000000011",
  64703=>"000110111",
  64704=>"111100100",
  64705=>"000000000",
  64706=>"110011010",
  64707=>"001011011",
  64708=>"111000101",
  64709=>"111001010",
  64710=>"000111111",
  64711=>"000010010",
  64712=>"100110000",
  64713=>"000000000",
  64714=>"010101000",
  64715=>"111101101",
  64716=>"011111111",
  64717=>"100001001",
  64718=>"111111110",
  64719=>"111001010",
  64720=>"000000111",
  64721=>"011001001",
  64722=>"111000010",
  64723=>"111111100",
  64724=>"000010111",
  64725=>"010011011",
  64726=>"000000000",
  64727=>"111111111",
  64728=>"000000101",
  64729=>"111100111",
  64730=>"000100101",
  64731=>"110000111",
  64732=>"100101001",
  64733=>"111101010",
  64734=>"111101100",
  64735=>"001000000",
  64736=>"111110111",
  64737=>"001111010",
  64738=>"001000000",
  64739=>"111000000",
  64740=>"010000000",
  64741=>"000000101",
  64742=>"100000000",
  64743=>"111111100",
  64744=>"000111111",
  64745=>"111111101",
  64746=>"011100100",
  64747=>"001000000",
  64748=>"101111000",
  64749=>"111100001",
  64750=>"110000101",
  64751=>"000000000",
  64752=>"111101100",
  64753=>"100100100",
  64754=>"101001000",
  64755=>"000010110",
  64756=>"001101000",
  64757=>"010111101",
  64758=>"111000000",
  64759=>"000000010",
  64760=>"111111000",
  64761=>"010110111",
  64762=>"100000000",
  64763=>"111101111",
  64764=>"111111000",
  64765=>"000010000",
  64766=>"101111110",
  64767=>"110000000",
  64768=>"001000000",
  64769=>"000000111",
  64770=>"000100100",
  64771=>"000011001",
  64772=>"011000100",
  64773=>"111000000",
  64774=>"000000011",
  64775=>"100110110",
  64776=>"000000001",
  64777=>"000011001",
  64778=>"011111010",
  64779=>"000011000",
  64780=>"000100101",
  64781=>"000000010",
  64782=>"001011001",
  64783=>"110111010",
  64784=>"010011011",
  64785=>"010011011",
  64786=>"000100111",
  64787=>"011100111",
  64788=>"000100000",
  64789=>"100100101",
  64790=>"111001010",
  64791=>"001000011",
  64792=>"011000011",
  64793=>"100100111",
  64794=>"010000110",
  64795=>"011011000",
  64796=>"000000001",
  64797=>"101101100",
  64798=>"011000000",
  64799=>"000100100",
  64800=>"000000000",
  64801=>"010000111",
  64802=>"101010011",
  64803=>"111101010",
  64804=>"010100000",
  64805=>"011001001",
  64806=>"100100110",
  64807=>"000111010",
  64808=>"010100101",
  64809=>"011111011",
  64810=>"100010000",
  64811=>"111110111",
  64812=>"011011011",
  64813=>"111100000",
  64814=>"101101100",
  64815=>"110100000",
  64816=>"010000011",
  64817=>"111111111",
  64818=>"100100010",
  64819=>"000111111",
  64820=>"011111000",
  64821=>"011111101",
  64822=>"110000001",
  64823=>"000100000",
  64824=>"000001000",
  64825=>"000000110",
  64826=>"100100111",
  64827=>"000010110",
  64828=>"110111000",
  64829=>"100100110",
  64830=>"000000000",
  64831=>"001001101",
  64832=>"111111011",
  64833=>"011001000",
  64834=>"100001010",
  64835=>"001011000",
  64836=>"000000000",
  64837=>"001000000",
  64838=>"000100011",
  64839=>"011111001",
  64840=>"100101101",
  64841=>"010001111",
  64842=>"101100000",
  64843=>"000000111",
  64844=>"010011010",
  64845=>"110011111",
  64846=>"100110110",
  64847=>"010010011",
  64848=>"100100100",
  64849=>"010000011",
  64850=>"111011101",
  64851=>"001000000",
  64852=>"000010000",
  64853=>"110100001",
  64854=>"010001000",
  64855=>"000010000",
  64856=>"000101001",
  64857=>"110010010",
  64858=>"010110000",
  64859=>"110110110",
  64860=>"101100101",
  64861=>"000000000",
  64862=>"011011010",
  64863=>"110011000",
  64864=>"101001001",
  64865=>"010101111",
  64866=>"101001101",
  64867=>"001011000",
  64868=>"000000000",
  64869=>"000001000",
  64870=>"000100010",
  64871=>"100101101",
  64872=>"000011010",
  64873=>"000100100",
  64874=>"111011010",
  64875=>"011011101",
  64876=>"000101000",
  64877=>"111111000",
  64878=>"100100111",
  64879=>"011011111",
  64880=>"110001001",
  64881=>"000010011",
  64882=>"001100110",
  64883=>"101000000",
  64884=>"000000011",
  64885=>"100100010",
  64886=>"000111111",
  64887=>"111000000",
  64888=>"011000100",
  64889=>"111000000",
  64890=>"000001011",
  64891=>"111100101",
  64892=>"000110010",
  64893=>"110000000",
  64894=>"100100111",
  64895=>"100001100",
  64896=>"011010000",
  64897=>"011011000",
  64898=>"000000111",
  64899=>"111101100",
  64900=>"100000100",
  64901=>"100111100",
  64902=>"011110100",
  64903=>"000001100",
  64904=>"110000100",
  64905=>"000111111",
  64906=>"000000000",
  64907=>"011000110",
  64908=>"100100000",
  64909=>"101100101",
  64910=>"111011010",
  64911=>"100001001",
  64912=>"011001101",
  64913=>"000010011",
  64914=>"000000000",
  64915=>"100000011",
  64916=>"100111011",
  64917=>"000000000",
  64918=>"111011011",
  64919=>"101001000",
  64920=>"011011000",
  64921=>"110101111",
  64922=>"100000010",
  64923=>"011010000",
  64924=>"100100000",
  64925=>"011011010",
  64926=>"000111110",
  64927=>"100101100",
  64928=>"001001110",
  64929=>"010011010",
  64930=>"100100000",
  64931=>"000000010",
  64932=>"010100111",
  64933=>"000000000",
  64934=>"010011101",
  64935=>"000000000",
  64936=>"011010111",
  64937=>"011111011",
  64938=>"110100101",
  64939=>"000000000",
  64940=>"111111000",
  64941=>"100000000",
  64942=>"100101001",
  64943=>"000000000",
  64944=>"100100010",
  64945=>"000110110",
  64946=>"000100000",
  64947=>"000100000",
  64948=>"111110100",
  64949=>"101111111",
  64950=>"111100100",
  64951=>"001011001",
  64952=>"101101100",
  64953=>"101111111",
  64954=>"011001000",
  64955=>"011000000",
  64956=>"000101100",
  64957=>"111111111",
  64958=>"110110010",
  64959=>"100111111",
  64960=>"000100111",
  64961=>"000000000",
  64962=>"000000101",
  64963=>"100100100",
  64964=>"000000010",
  64965=>"010010000",
  64966=>"011000001",
  64967=>"000001111",
  64968=>"101101011",
  64969=>"111000000",
  64970=>"000000100",
  64971=>"101011010",
  64972=>"100001111",
  64973=>"000001011",
  64974=>"000110000",
  64975=>"100011111",
  64976=>"000110111",
  64977=>"110110100",
  64978=>"000110011",
  64979=>"010111010",
  64980=>"000100111",
  64981=>"100101100",
  64982=>"000111011",
  64983=>"000001011",
  64984=>"100101111",
  64985=>"111100100",
  64986=>"010100000",
  64987=>"100100110",
  64988=>"111011011",
  64989=>"011111100",
  64990=>"111111111",
  64991=>"010011001",
  64992=>"000000100",
  64993=>"000000011",
  64994=>"111100111",
  64995=>"000101001",
  64996=>"000100000",
  64997=>"000001111",
  64998=>"000000011",
  64999=>"001000100",
  65000=>"100100000",
  65001=>"100100111",
  65002=>"111111110",
  65003=>"001100111",
  65004=>"001000000",
  65005=>"000010111",
  65006=>"000100000",
  65007=>"101111100",
  65008=>"011010011",
  65009=>"111011101",
  65010=>"000010111",
  65011=>"101011101",
  65012=>"110110000",
  65013=>"111111111",
  65014=>"100110000",
  65015=>"011011101",
  65016=>"000000101",
  65017=>"000101011",
  65018=>"110100100",
  65019=>"011111111",
  65020=>"111011000",
  65021=>"011111000",
  65022=>"111110000",
  65023=>"111010000",
  65024=>"011100100",
  65025=>"011000010",
  65026=>"100101101",
  65027=>"000000000",
  65028=>"111011000",
  65029=>"000001110",
  65030=>"100100111",
  65031=>"000000010",
  65032=>"000000010",
  65033=>"000000110",
  65034=>"110110010",
  65035=>"111000101",
  65036=>"111111000",
  65037=>"111101100",
  65038=>"010000000",
  65039=>"001101111",
  65040=>"110000010",
  65041=>"111111000",
  65042=>"101001101",
  65043=>"110011001",
  65044=>"101000101",
  65045=>"100000000",
  65046=>"011111110",
  65047=>"111010000",
  65048=>"111110000",
  65049=>"110110011",
  65050=>"000011011",
  65051=>"011000000",
  65052=>"011011001",
  65053=>"111110110",
  65054=>"001000011",
  65055=>"000110101",
  65056=>"101101111",
  65057=>"010110111",
  65058=>"011100111",
  65059=>"111000000",
  65060=>"001001011",
  65061=>"110110100",
  65062=>"000010010",
  65063=>"111111010",
  65064=>"000111111",
  65065=>"000001011",
  65066=>"010011111",
  65067=>"000000000",
  65068=>"011011011",
  65069=>"111111001",
  65070=>"011000000",
  65071=>"111111111",
  65072=>"111111001",
  65073=>"011111111",
  65074=>"000000010",
  65075=>"010010010",
  65076=>"010100111",
  65077=>"000000000",
  65078=>"011000100",
  65079=>"010011111",
  65080=>"001011010",
  65081=>"010111111",
  65082=>"000000100",
  65083=>"001000010",
  65084=>"110101000",
  65085=>"110111111",
  65086=>"010000011",
  65087=>"001111111",
  65088=>"000000111",
  65089=>"111111000",
  65090=>"101101111",
  65091=>"110001101",
  65092=>"001101001",
  65093=>"000111111",
  65094=>"110000010",
  65095=>"100101100",
  65096=>"000000000",
  65097=>"111101111",
  65098=>"010000011",
  65099=>"000010111",
  65100=>"000010010",
  65101=>"011001000",
  65102=>"100110111",
  65103=>"111111111",
  65104=>"100100111",
  65105=>"110111000",
  65106=>"000000000",
  65107=>"001011000",
  65108=>"010000111",
  65109=>"110111000",
  65110=>"100110110",
  65111=>"111100100",
  65112=>"000000000",
  65113=>"010011100",
  65114=>"000010110",
  65115=>"100100111",
  65116=>"011101111",
  65117=>"001001001",
  65118=>"000010010",
  65119=>"010100101",
  65120=>"111100111",
  65121=>"111111001",
  65122=>"111000000",
  65123=>"000100110",
  65124=>"100001010",
  65125=>"000111101",
  65126=>"000100000",
  65127=>"000000000",
  65128=>"101111011",
  65129=>"000000010",
  65130=>"110000111",
  65131=>"100010110",
  65132=>"000010000",
  65133=>"101111111",
  65134=>"010000001",
  65135=>"111111010",
  65136=>"001001011",
  65137=>"000000000",
  65138=>"111000011",
  65139=>"101110111",
  65140=>"000100001",
  65141=>"000010000",
  65142=>"000001000",
  65143=>"001000110",
  65144=>"101000000",
  65145=>"000000000",
  65146=>"111111111",
  65147=>"111101000",
  65148=>"001001110",
  65149=>"100001010",
  65150=>"111101111",
  65151=>"000101111",
  65152=>"011000101",
  65153=>"001010000",
  65154=>"010000000",
  65155=>"010010110",
  65156=>"000000010",
  65157=>"111101001",
  65158=>"111111001",
  65159=>"001001001",
  65160=>"100110011",
  65161=>"000000000",
  65162=>"000110110",
  65163=>"100101111",
  65164=>"000000000",
  65165=>"000000000",
  65166=>"000000001",
  65167=>"000000011",
  65168=>"100111011",
  65169=>"110010001",
  65170=>"001000001",
  65171=>"010111011",
  65172=>"011010000",
  65173=>"010110111",
  65174=>"011111000",
  65175=>"000000100",
  65176=>"000000000",
  65177=>"000000000",
  65178=>"110111111",
  65179=>"111000000",
  65180=>"000010011",
  65181=>"000000010",
  65182=>"000100010",
  65183=>"101001000",
  65184=>"001101101",
  65185=>"110000100",
  65186=>"111101101",
  65187=>"111111111",
  65188=>"110011010",
  65189=>"100111111",
  65190=>"111110011",
  65191=>"000011011",
  65192=>"110010000",
  65193=>"000000010",
  65194=>"000101111",
  65195=>"110111111",
  65196=>"010110000",
  65197=>"000100111",
  65198=>"110110110",
  65199=>"001000111",
  65200=>"111111011",
  65201=>"000110110",
  65202=>"111100101",
  65203=>"100110010",
  65204=>"111111110",
  65205=>"110010000",
  65206=>"111011000",
  65207=>"011001001",
  65208=>"001000000",
  65209=>"010010110",
  65210=>"010000000",
  65211=>"010001001",
  65212=>"101000000",
  65213=>"000000000",
  65214=>"001111011",
  65215=>"000000000",
  65216=>"101000111",
  65217=>"000011111",
  65218=>"010010010",
  65219=>"011111110",
  65220=>"000010101",
  65221=>"110110010",
  65222=>"011011000",
  65223=>"000000000",
  65224=>"111111111",
  65225=>"010010001",
  65226=>"100111010",
  65227=>"111111101",
  65228=>"111100111",
  65229=>"111000000",
  65230=>"000101101",
  65231=>"100010110",
  65232=>"100110100",
  65233=>"100100111",
  65234=>"000110001",
  65235=>"010001111",
  65236=>"111000111",
  65237=>"000110110",
  65238=>"011111001",
  65239=>"111111001",
  65240=>"111111000",
  65241=>"111111001",
  65242=>"110111111",
  65243=>"000000010",
  65244=>"001101000",
  65245=>"001010000",
  65246=>"101010000",
  65247=>"000000010",
  65248=>"111111000",
  65249=>"010100110",
  65250=>"111000001",
  65251=>"111111010",
  65252=>"110000011",
  65253=>"000000000",
  65254=>"101011000",
  65255=>"001001011",
  65256=>"111000001",
  65257=>"000000011",
  65258=>"000011011",
  65259=>"111101101",
  65260=>"010111101",
  65261=>"011010111",
  65262=>"100000000",
  65263=>"111001000",
  65264=>"110111001",
  65265=>"011011110",
  65266=>"111000110",
  65267=>"101011011",
  65268=>"111011001",
  65269=>"000000111",
  65270=>"101101111",
  65271=>"111111101",
  65272=>"111011000",
  65273=>"000101001",
  65274=>"010001111",
  65275=>"101110110",
  65276=>"111111111",
  65277=>"111110011",
  65278=>"000000011",
  65279=>"000010010",
  65280=>"011010011",
  65281=>"000000110",
  65282=>"100110101",
  65283=>"000101111",
  65284=>"000000000",
  65285=>"000001010",
  65286=>"111000111",
  65287=>"011111111",
  65288=>"100101111",
  65289=>"000000101",
  65290=>"110011011",
  65291=>"100000001",
  65292=>"000010000",
  65293=>"000100111",
  65294=>"001111111",
  65295=>"110000110",
  65296=>"000000000",
  65297=>"000000000",
  65298=>"111111111",
  65299=>"001001010",
  65300=>"011111000",
  65301=>"001000000",
  65302=>"010001110",
  65303=>"010010111",
  65304=>"000001101",
  65305=>"111111111",
  65306=>"000100100",
  65307=>"111111111",
  65308=>"100111111",
  65309=>"101101111",
  65310=>"111111110",
  65311=>"000000000",
  65312=>"000000000",
  65313=>"010001001",
  65314=>"000000101",
  65315=>"000100001",
  65316=>"110011011",
  65317=>"000010110",
  65318=>"000000000",
  65319=>"010111111",
  65320=>"000000111",
  65321=>"111111111",
  65322=>"111110111",
  65323=>"000000000",
  65324=>"011011011",
  65325=>"000001111",
  65326=>"001100000",
  65327=>"011110001",
  65328=>"100011000",
  65329=>"110011011",
  65330=>"000000101",
  65331=>"111001000",
  65332=>"101000000",
  65333=>"110010010",
  65334=>"100000010",
  65335=>"111111110",
  65336=>"111111011",
  65337=>"011011111",
  65338=>"111100111",
  65339=>"000000000",
  65340=>"111101011",
  65341=>"011111111",
  65342=>"000000100",
  65343=>"000111100",
  65344=>"000000000",
  65345=>"011111111",
  65346=>"111111111",
  65347=>"111101010",
  65348=>"111110010",
  65349=>"000000000",
  65350=>"101000000",
  65351=>"010000000",
  65352=>"111001111",
  65353=>"010010000",
  65354=>"010111111",
  65355=>"000001000",
  65356=>"011011000",
  65357=>"000100011",
  65358=>"111111011",
  65359=>"101101101",
  65360=>"001000000",
  65361=>"011111111",
  65362=>"010111111",
  65363=>"111101011",
  65364=>"011011011",
  65365=>"110001000",
  65366=>"110000100",
  65367=>"000111111",
  65368=>"100000010",
  65369=>"111110110",
  65370=>"110000000",
  65371=>"001110111",
  65372=>"111111000",
  65373=>"010001011",
  65374=>"000000000",
  65375=>"011111101",
  65376=>"111101011",
  65377=>"110001101",
  65378=>"000100000",
  65379=>"110100010",
  65380=>"100100110",
  65381=>"111111111",
  65382=>"111001000",
  65383=>"111101111",
  65384=>"111111110",
  65385=>"000000000",
  65386=>"110111111",
  65387=>"011010010",
  65388=>"110111001",
  65389=>"101100000",
  65390=>"000000000",
  65391=>"111011000",
  65392=>"111111011",
  65393=>"011000100",
  65394=>"000000010",
  65395=>"111101111",
  65396=>"010000000",
  65397=>"101100000",
  65398=>"111111111",
  65399=>"000111010",
  65400=>"000000000",
  65401=>"111111000",
  65402=>"000101101",
  65403=>"000000010",
  65404=>"100100001",
  65405=>"111111000",
  65406=>"000000000",
  65407=>"111111010",
  65408=>"111111000",
  65409=>"010111000",
  65410=>"000001111",
  65411=>"000000001",
  65412=>"101011111",
  65413=>"110011111",
  65414=>"110110111",
  65415=>"111011001",
  65416=>"001111011",
  65417=>"101000000",
  65418=>"110100110",
  65419=>"111111000",
  65420=>"000000000",
  65421=>"000000000",
  65422=>"011010000",
  65423=>"111000100",
  65424=>"001011111",
  65425=>"001011000",
  65426=>"101000000",
  65427=>"111000010",
  65428=>"010100100",
  65429=>"010111111",
  65430=>"111111010",
  65431=>"101001110",
  65432=>"000000001",
  65433=>"111100101",
  65434=>"101100100",
  65435=>"000000000",
  65436=>"111000100",
  65437=>"111111111",
  65438=>"111111111",
  65439=>"000010011",
  65440=>"011010001",
  65441=>"110100100",
  65442=>"111111011",
  65443=>"111101111",
  65444=>"110010001",
  65445=>"110110110",
  65446=>"000000111",
  65447=>"100000000",
  65448=>"000000011",
  65449=>"000000111",
  65450=>"111111100",
  65451=>"000100100",
  65452=>"111001011",
  65453=>"111111111",
  65454=>"001011011",
  65455=>"111001111",
  65456=>"000000000",
  65457=>"111111001",
  65458=>"111100110",
  65459=>"110011001",
  65460=>"000001001",
  65461=>"101101110",
  65462=>"000001001",
  65463=>"000100000",
  65464=>"110110101",
  65465=>"110110101",
  65466=>"110000000",
  65467=>"111010011",
  65468=>"111000000",
  65469=>"000011000",
  65470=>"000010100",
  65471=>"101000000",
  65472=>"000000000",
  65473=>"000000000",
  65474=>"011011111",
  65475=>"110100010",
  65476=>"000001100",
  65477=>"011001001",
  65478=>"000011010",
  65479=>"000100110",
  65480=>"101111000",
  65481=>"011111010",
  65482=>"010010001",
  65483=>"000011010",
  65484=>"000010000",
  65485=>"001101100",
  65486=>"111100001",
  65487=>"110100100",
  65488=>"111101111",
  65489=>"100100011",
  65490=>"010010111",
  65491=>"010010001",
  65492=>"100100111",
  65493=>"100110000",
  65494=>"010111001",
  65495=>"000101111",
  65496=>"000000010",
  65497=>"111011101",
  65498=>"100110010",
  65499=>"100000000",
  65500=>"000100001",
  65501=>"000000010",
  65502=>"011111010",
  65503=>"000001000",
  65504=>"010010100",
  65505=>"111100100",
  65506=>"001010110",
  65507=>"100110010",
  65508=>"000000100",
  65509=>"100000000",
  65510=>"000010010",
  65511=>"011011111",
  65512=>"010011111",
  65513=>"100000011",
  65514=>"001110110",
  65515=>"000100100",
  65516=>"011111111",
  65517=>"010000001",
  65518=>"001101001",
  65519=>"101100000",
  65520=>"100111010",
  65521=>"100110000",
  65522=>"111111111",
  65523=>"000010010",
  65524=>"110101111",
  65525=>"000000000",
  65526=>"111000000",
  65527=>"111111111",
  65528=>"000000100",
  65529=>"111111111",
  65530=>"010010000",
  65531=>"010111010",
  65532=>"100000100",
  65533=>"000000000",
  65534=>"110000110",
  65535=>"001111111");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;