LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L7_2_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(7) - 1 DOWNTO 0));
END L7_2_WROM;

ARCHITECTURE RTL OF L7_2_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"111111100",
  1=>"001001111",
  2=>"111111111",
  3=>"111101001",
  4=>"111111111",
  5=>"101111111",
  6=>"111111111",
  7=>"101101111",
  8=>"001000000",
  9=>"001111111",
  10=>"101000000",
  11=>"111111111",
  12=>"000000000",
  13=>"000111111",
  14=>"111111111",
  15=>"010011011",
  16=>"111100000",
  17=>"001000000",
  18=>"111111111",
  19=>"000111111",
  20=>"111111001",
  21=>"111111111",
  22=>"100000111",
  23=>"000000000",
  24=>"100111111",
  25=>"000000010",
  26=>"010000000",
  27=>"011111110",
  28=>"111101000",
  29=>"111111101",
  30=>"000000000",
  31=>"000000000",
  32=>"000000000",
  33=>"000000001",
  34=>"110110111",
  35=>"100100100",
  36=>"111000000",
  37=>"001001000",
  38=>"000001111",
  39=>"001000000",
  40=>"100000000",
  41=>"111111110",
  42=>"000001000",
  43=>"111111111",
  44=>"000000111",
  45=>"011111110",
  46=>"001000000",
  47=>"101001000",
  48=>"111001111",
  49=>"000000000",
  50=>"010000000",
  51=>"000001111",
  52=>"001001000",
  53=>"110000000",
  54=>"111001000",
  55=>"000000000",
  56=>"111011001",
  57=>"101111000",
  58=>"111111111",
  59=>"001111111",
  60=>"000000000",
  61=>"000000000",
  62=>"100110111",
  63=>"111011000",
  64=>"000000000",
  65=>"001111001",
  66=>"000000000",
  67=>"000000000",
  68=>"000000000",
  69=>"111111010",
  70=>"000000000",
  71=>"111111111",
  72=>"000001000",
  73=>"000000000",
  74=>"111111111",
  75=>"110111001",
  76=>"110100100",
  77=>"000000000",
  78=>"111011011",
  79=>"000000000",
  80=>"000011111",
  81=>"111111111",
  82=>"111110000",
  83=>"100111111",
  84=>"111111111",
  85=>"010111000",
  86=>"000101101",
  87=>"111100100",
  88=>"110111111",
  89=>"111101101",
  90=>"000000000",
  91=>"100110111",
  92=>"000000000",
  93=>"000101101",
  94=>"000001111",
  95=>"100000000",
  96=>"001100101",
  97=>"000000000",
  98=>"000000000",
  99=>"000000000",
  100=>"011111111",
  101=>"111111000",
  102=>"111111111",
  103=>"111100111",
  104=>"000000001",
  105=>"111111011",
  106=>"000001111",
  107=>"101101111",
  108=>"001101111",
  109=>"111100101",
  110=>"111111111",
  111=>"000000000",
  112=>"000001000",
  113=>"111000111",
  114=>"000011111",
  115=>"010110111",
  116=>"111110000",
  117=>"100100100",
  118=>"000000000",
  119=>"011011100",
  120=>"000000000",
  121=>"000111000",
  122=>"000100000",
  123=>"000000000",
  124=>"101111111",
  125=>"100111000",
  126=>"111000001",
  127=>"000000000",
  128=>"000000111",
  129=>"000000111",
  130=>"000000111",
  131=>"001011000",
  132=>"011111000",
  133=>"111111101",
  134=>"001001000",
  135=>"000000001",
  136=>"001000000",
  137=>"000111000",
  138=>"000000000",
  139=>"000100110",
  140=>"111111111",
  141=>"011001000",
  142=>"100011000",
  143=>"111000000",
  144=>"111111011",
  145=>"011111111",
  146=>"000000000",
  147=>"110000000",
  148=>"000000000",
  149=>"000010111",
  150=>"001111111",
  151=>"111101100",
  152=>"101001000",
  153=>"000101001",
  154=>"111111000",
  155=>"111011000",
  156=>"111111101",
  157=>"001000000",
  158=>"110110111",
  159=>"000000011",
  160=>"000010000",
  161=>"000000111",
  162=>"000011111",
  163=>"111111111",
  164=>"011000000",
  165=>"000011111",
  166=>"111000000",
  167=>"111101111",
  168=>"000001000",
  169=>"111011111",
  170=>"111100110",
  171=>"000000000",
  172=>"000000000",
  173=>"100100000",
  174=>"111111111",
  175=>"011001001",
  176=>"000000111",
  177=>"000000000",
  178=>"110111111",
  179=>"111110111",
  180=>"001000000",
  181=>"000000111",
  182=>"000000000",
  183=>"111111111",
  184=>"111111010",
  185=>"111111111",
  186=>"000000000",
  187=>"111000101",
  188=>"000000000",
  189=>"111011001",
  190=>"000000000",
  191=>"110111011",
  192=>"111111110",
  193=>"000000000",
  194=>"111101111",
  195=>"000000000",
  196=>"111111111",
  197=>"000000000",
  198=>"000101101",
  199=>"111111111",
  200=>"111000100",
  201=>"100111111",
  202=>"000000000",
  203=>"000000000",
  204=>"000001111",
  205=>"001101111",
  206=>"011011000",
  207=>"111111111",
  208=>"000111111",
  209=>"111000111",
  210=>"111111111",
  211=>"000000000",
  212=>"011011111",
  213=>"110110110",
  214=>"111100100",
  215=>"000111111",
  216=>"000000000",
  217=>"111111111",
  218=>"111111000",
  219=>"000100110",
  220=>"000000000",
  221=>"000000111",
  222=>"111011111",
  223=>"111111111",
  224=>"111111111",
  225=>"111111111",
  226=>"111111111",
  227=>"000000000",
  228=>"111111100",
  229=>"000111011",
  230=>"001000000",
  231=>"110111111",
  232=>"001101000",
  233=>"000000000",
  234=>"111001001",
  235=>"001000000",
  236=>"111011000",
  237=>"111111111",
  238=>"111111001",
  239=>"111111001",
  240=>"001111111",
  241=>"001000000",
  242=>"111111111",
  243=>"111000100",
  244=>"111111111",
  245=>"100000000",
  246=>"000111011",
  247=>"111111111",
  248=>"111001001",
  249=>"001000000",
  250=>"000000000",
  251=>"111111111",
  252=>"000100100",
  253=>"110110110",
  254=>"000110111",
  255=>"111111111",
  256=>"000000000",
  257=>"011011011",
  258=>"111111111",
  259=>"000000000",
  260=>"000000000",
  261=>"000010011",
  262=>"011111111",
  263=>"000000000",
  264=>"000000001",
  265=>"000000000",
  266=>"111111101",
  267=>"111111111",
  268=>"101100100",
  269=>"111111100",
  270=>"111111111",
  271=>"011111011",
  272=>"111111111",
  273=>"011000000",
  274=>"000000000",
  275=>"111000110",
  276=>"100100000",
  277=>"000000000",
  278=>"100100100",
  279=>"111111111",
  280=>"110111111",
  281=>"101000000",
  282=>"000001001",
  283=>"001000111",
  284=>"111001100",
  285=>"111000000",
  286=>"111111000",
  287=>"000000111",
  288=>"110100111",
  289=>"111111111",
  290=>"000000000",
  291=>"111111111",
  292=>"111111100",
  293=>"101100100",
  294=>"111111111",
  295=>"010000000",
  296=>"000000000",
  297=>"111111100",
  298=>"111111111",
  299=>"101000101",
  300=>"000001000",
  301=>"000110101",
  302=>"101111111",
  303=>"111111000",
  304=>"000110110",
  305=>"111000000",
  306=>"000000000",
  307=>"111111111",
  308=>"001000011",
  309=>"011111111",
  310=>"000000000",
  311=>"100000000",
  312=>"000000000",
  313=>"111111111",
  314=>"111001000",
  315=>"111001000",
  316=>"001001111",
  317=>"111111011",
  318=>"000100000",
  319=>"000111111",
  320=>"000000000",
  321=>"111111010",
  322=>"111111101",
  323=>"000000000",
  324=>"000001001",
  325=>"000000000",
  326=>"000000110",
  327=>"111111111",
  328=>"000000000",
  329=>"000000111",
  330=>"001111111",
  331=>"000000000",
  332=>"101000000",
  333=>"000000000",
  334=>"000001111",
  335=>"000000000",
  336=>"000000000",
  337=>"000000000",
  338=>"000000000",
  339=>"110110000",
  340=>"111111110",
  341=>"011001011",
  342=>"000011111",
  343=>"111011111",
  344=>"001111111",
  345=>"111100000",
  346=>"000000000",
  347=>"000100100",
  348=>"111100000",
  349=>"111101000",
  350=>"101101101",
  351=>"111101111",
  352=>"000000000",
  353=>"000000000",
  354=>"000000000",
  355=>"001001000",
  356=>"100100111",
  357=>"111111111",
  358=>"111111111",
  359=>"100000000",
  360=>"100000000",
  361=>"111111000",
  362=>"001000000",
  363=>"000000000",
  364=>"111111111",
  365=>"000000000",
  366=>"000000000",
  367=>"000000000",
  368=>"000000111",
  369=>"000000000",
  370=>"000000000",
  371=>"011011111",
  372=>"111111001",
  373=>"111101000",
  374=>"011111000",
  375=>"001101101",
  376=>"100100110",
  377=>"000000000",
  378=>"110110111",
  379=>"000000000",
  380=>"011011000",
  381=>"111100000",
  382=>"111111001",
  383=>"001001111",
  384=>"010010000",
  385=>"110111101",
  386=>"111111010",
  387=>"111111111",
  388=>"000000100",
  389=>"111111011",
  390=>"000000000",
  391=>"000000000",
  392=>"111111111",
  393=>"111111100",
  394=>"100101001",
  395=>"000000110",
  396=>"101111111",
  397=>"111111111",
  398=>"000100100",
  399=>"111111111",
  400=>"000000000",
  401=>"111101000",
  402=>"111111111",
  403=>"110110111",
  404=>"100101111",
  405=>"000000000",
  406=>"111111111",
  407=>"111111111",
  408=>"100111000",
  409=>"000110110",
  410=>"110111110",
  411=>"100111111",
  412=>"000000000",
  413=>"011000000",
  414=>"111111111",
  415=>"001000000",
  416=>"000011111",
  417=>"001001001",
  418=>"001000000",
  419=>"011110110",
  420=>"100111111",
  421=>"000111111",
  422=>"000000000",
  423=>"111111111",
  424=>"000000100",
  425=>"000000100",
  426=>"111111111",
  427=>"111100111",
  428=>"000000000",
  429=>"000000000",
  430=>"000000111",
  431=>"000000000",
  432=>"000000000",
  433=>"000000000",
  434=>"100000000",
  435=>"000000000",
  436=>"000100111",
  437=>"001000101",
  438=>"001111111",
  439=>"000010000",
  440=>"111111000",
  441=>"000000000",
  442=>"011000000",
  443=>"111111111",
  444=>"001111101",
  445=>"111110000",
  446=>"000000111",
  447=>"100111111",
  448=>"000100000",
  449=>"001111111",
  450=>"000000000",
  451=>"001000000",
  452=>"100110111",
  453=>"100100000",
  454=>"000000000",
  455=>"111111111",
  456=>"000000100",
  457=>"000000000",
  458=>"000001001",
  459=>"111111111",
  460=>"011011011",
  461=>"110100100",
  462=>"000000000",
  463=>"111111111",
  464=>"011000000",
  465=>"000000000",
  466=>"000000000",
  467=>"100101000",
  468=>"101001010",
  469=>"000111111",
  470=>"011001000",
  471=>"000000000",
  472=>"111111111",
  473=>"111110110",
  474=>"110111000",
  475=>"000000111",
  476=>"011000000",
  477=>"111000000",
  478=>"000000000",
  479=>"010110000",
  480=>"111000000",
  481=>"111100100",
  482=>"000010011",
  483=>"001111111",
  484=>"000000001",
  485=>"000111111",
  486=>"000010011",
  487=>"000000001",
  488=>"111111011",
  489=>"100000001",
  490=>"000000000",
  491=>"001001111",
  492=>"100101111",
  493=>"111111111",
  494=>"111111111",
  495=>"011011111",
  496=>"111111111",
  497=>"000000001",
  498=>"101111101",
  499=>"011000000",
  500=>"000100111",
  501=>"000000000",
  502=>"111111111",
  503=>"001001000",
  504=>"000000000",
  505=>"001001001",
  506=>"000100110",
  507=>"100110000",
  508=>"000111111",
  509=>"000000000",
  510=>"100110000",
  511=>"000000000",
  512=>"001111111",
  513=>"000000011",
  514=>"111111111",
  515=>"000000001",
  516=>"011111111",
  517=>"100000000",
  518=>"000000000",
  519=>"000000000",
  520=>"111111111",
  521=>"111111111",
  522=>"000001001",
  523=>"111111101",
  524=>"000000000",
  525=>"110111110",
  526=>"011001001",
  527=>"000000111",
  528=>"000100111",
  529=>"001000111",
  530=>"000100101",
  531=>"111101111",
  532=>"111001000",
  533=>"111100111",
  534=>"001000000",
  535=>"111111110",
  536=>"110110000",
  537=>"000000000",
  538=>"100100000",
  539=>"111111111",
  540=>"000000000",
  541=>"100111111",
  542=>"111100000",
  543=>"001100000",
  544=>"111111010",
  545=>"100001111",
  546=>"100000100",
  547=>"111111111",
  548=>"110111110",
  549=>"111111111",
  550=>"111100000",
  551=>"000000000",
  552=>"000001011",
  553=>"000000000",
  554=>"000000000",
  555=>"000000000",
  556=>"111000111",
  557=>"000000000",
  558=>"111111011",
  559=>"101100000",
  560=>"000000001",
  561=>"010001101",
  562=>"010011001",
  563=>"000100000",
  564=>"000000000",
  565=>"110111010",
  566=>"011111111",
  567=>"000000000",
  568=>"111111000",
  569=>"111111111",
  570=>"111111111",
  571=>"000000000",
  572=>"001000000",
  573=>"111111111",
  574=>"111111111",
  575=>"111000001",
  576=>"000010000",
  577=>"000000111",
  578=>"110111111",
  579=>"100100110",
  580=>"110111111",
  581=>"000000110",
  582=>"111111111",
  583=>"100000000",
  584=>"001100100",
  585=>"000000111",
  586=>"000000000",
  587=>"000000000",
  588=>"111111111",
  589=>"000000001",
  590=>"000000011",
  591=>"110101111",
  592=>"011011011",
  593=>"000000111",
  594=>"000000000",
  595=>"111111111",
  596=>"000000000",
  597=>"011000000",
  598=>"111111111",
  599=>"001000000",
  600=>"000000000",
  601=>"001000000",
  602=>"111111111",
  603=>"000111111",
  604=>"000000000",
  605=>"000000111",
  606=>"000000110",
  607=>"110111010",
  608=>"000000000",
  609=>"000000000",
  610=>"000001111",
  611=>"101111111",
  612=>"101001000",
  613=>"001111111",
  614=>"111110111",
  615=>"111111111",
  616=>"111111111",
  617=>"111111111",
  618=>"111111111",
  619=>"111111111",
  620=>"111111110",
  621=>"100100111",
  622=>"111111111",
  623=>"000000111",
  624=>"111000000",
  625=>"000000000",
  626=>"011010011",
  627=>"111011011",
  628=>"011001000",
  629=>"000000000",
  630=>"011000000",
  631=>"000000000",
  632=>"000000000",
  633=>"110000101",
  634=>"000000111",
  635=>"001001001",
  636=>"000001001",
  637=>"111111010",
  638=>"011011111",
  639=>"110100000",
  640=>"111001001",
  641=>"111111000",
  642=>"111110100",
  643=>"011111111",
  644=>"100110111",
  645=>"000101000",
  646=>"111111111",
  647=>"011000000",
  648=>"110111111",
  649=>"000000000",
  650=>"000000001",
  651=>"111000111",
  652=>"011000010",
  653=>"110000000",
  654=>"101001000",
  655=>"000000000",
  656=>"111111111",
  657=>"011011001",
  658=>"000100100",
  659=>"000000000",
  660=>"000110111",
  661=>"000100100",
  662=>"111111111",
  663=>"111111100",
  664=>"000000010",
  665=>"000000000",
  666=>"000000111",
  667=>"111111000",
  668=>"101111111",
  669=>"110110000",
  670=>"101100110",
  671=>"111001001",
  672=>"111111111",
  673=>"000000000",
  674=>"000000000",
  675=>"000000000",
  676=>"000000100",
  677=>"000100111",
  678=>"000000001",
  679=>"000100110",
  680=>"111111110",
  681=>"000000000",
  682=>"000000000",
  683=>"101000100",
  684=>"001100111",
  685=>"111111001",
  686=>"100111111",
  687=>"111111100",
  688=>"000110111",
  689=>"110111111",
  690=>"111011111",
  691=>"000001001",
  692=>"101100100",
  693=>"111111100",
  694=>"000000000",
  695=>"111111000",
  696=>"110100110",
  697=>"111100101",
  698=>"000100111",
  699=>"000000111",
  700=>"000000000",
  701=>"100000010",
  702=>"000000000",
  703=>"111111001",
  704=>"010011000",
  705=>"000111111",
  706=>"011011011",
  707=>"111000000",
  708=>"111101010",
  709=>"000000000",
  710=>"000000000",
  711=>"000000000",
  712=>"111000000",
  713=>"111011000",
  714=>"001000110",
  715=>"110011111",
  716=>"000000000",
  717=>"001000000",
  718=>"000000000",
  719=>"000000100",
  720=>"111111111",
  721=>"001001111",
  722=>"000000111",
  723=>"111111011",
  724=>"000000000",
  725=>"111000100",
  726=>"000001000",
  727=>"111111111",
  728=>"000000000",
  729=>"110111111",
  730=>"000000000",
  731=>"111111111",
  732=>"111111111",
  733=>"111001000",
  734=>"000000111",
  735=>"100000000",
  736=>"000000000",
  737=>"000000000",
  738=>"111111100",
  739=>"000000000",
  740=>"011011011",
  741=>"000000000",
  742=>"000000000",
  743=>"011011100",
  744=>"111111111",
  745=>"111111111",
  746=>"000000000",
  747=>"000000000",
  748=>"000000000",
  749=>"000000111",
  750=>"000110111",
  751=>"000000000",
  752=>"110110010",
  753=>"111011000",
  754=>"111111111",
  755=>"010100100",
  756=>"111101100",
  757=>"011111111",
  758=>"000000000",
  759=>"000100000",
  760=>"000000000",
  761=>"111101101",
  762=>"111111111",
  763=>"000000000",
  764=>"001001001",
  765=>"100100011",
  766=>"000000000",
  767=>"000000000",
  768=>"000000000",
  769=>"000000000",
  770=>"000000111",
  771=>"010000000",
  772=>"000000000",
  773=>"000000000",
  774=>"111000000",
  775=>"000000000",
  776=>"110110010",
  777=>"111000000",
  778=>"111111111",
  779=>"110111100",
  780=>"111000000",
  781=>"110100000",
  782=>"000000111",
  783=>"000000110",
  784=>"111011000",
  785=>"001000001",
  786=>"011000000",
  787=>"111110001",
  788=>"111111111",
  789=>"011111111",
  790=>"111111111",
  791=>"100111111",
  792=>"110111111",
  793=>"111000000",
  794=>"001000000",
  795=>"111111111",
  796=>"000000000",
  797=>"110110000",
  798=>"000000000",
  799=>"111111001",
  800=>"111111111",
  801=>"111111111",
  802=>"111111000",
  803=>"101111111",
  804=>"111111111",
  805=>"000000000",
  806=>"110110111",
  807=>"111111111",
  808=>"111111111",
  809=>"000000001",
  810=>"100111011",
  811=>"111111111",
  812=>"111111110",
  813=>"000001101",
  814=>"111101111",
  815=>"000000000",
  816=>"001011110",
  817=>"111111111",
  818=>"111011001",
  819=>"000001100",
  820=>"111111111",
  821=>"110111111",
  822=>"000000100",
  823=>"110000101",
  824=>"000000000",
  825=>"111111111",
  826=>"111001000",
  827=>"000000000",
  828=>"111101000",
  829=>"000000000",
  830=>"101000000",
  831=>"111111111",
  832=>"000000000",
  833=>"111110100",
  834=>"000000011",
  835=>"000000000",
  836=>"000000011",
  837=>"000001111",
  838=>"011011011",
  839=>"001001101",
  840=>"000000000",
  841=>"000000000",
  842=>"000011111",
  843=>"100100100",
  844=>"101111001",
  845=>"000000111",
  846=>"111111111",
  847=>"110000110",
  848=>"100010011",
  849=>"111111111",
  850=>"000010110",
  851=>"111111101",
  852=>"000111111",
  853=>"111111111",
  854=>"000001111",
  855=>"111111111",
  856=>"000000000",
  857=>"111000000",
  858=>"110010110",
  859=>"111111111",
  860=>"010000000",
  861=>"111000000",
  862=>"000011011",
  863=>"000000000",
  864=>"000000000",
  865=>"111001101",
  866=>"011011001",
  867=>"111111000",
  868=>"111111000",
  869=>"000000000",
  870=>"000000111",
  871=>"111111111",
  872=>"001001100",
  873=>"011000100",
  874=>"111111111",
  875=>"000000011",
  876=>"000100110",
  877=>"000000100",
  878=>"111000000",
  879=>"111000111",
  880=>"111001111",
  881=>"000000000",
  882=>"111000000",
  883=>"001000001",
  884=>"111111111",
  885=>"111111111",
  886=>"010111111",
  887=>"000000000",
  888=>"101000000",
  889=>"011101100",
  890=>"001001001",
  891=>"001111110",
  892=>"111111000",
  893=>"001000101",
  894=>"101111111",
  895=>"100000111",
  896=>"100000011",
  897=>"001000000",
  898=>"100110110",
  899=>"111000000",
  900=>"000000101",
  901=>"111111111",
  902=>"101111011",
  903=>"000111111",
  904=>"000000000",
  905=>"000000000",
  906=>"001000010",
  907=>"100100100",
  908=>"111111111",
  909=>"001001000",
  910=>"011111111",
  911=>"011010000",
  912=>"001000001",
  913=>"111111111",
  914=>"111000111",
  915=>"110100100",
  916=>"111111111",
  917=>"000000000",
  918=>"000110111",
  919=>"111111011",
  920=>"111101110",
  921=>"000000000",
  922=>"111111110",
  923=>"000000000",
  924=>"101000000",
  925=>"011000001",
  926=>"011111111",
  927=>"000110111",
  928=>"111000100",
  929=>"001011111",
  930=>"000111111",
  931=>"000000000",
  932=>"000111110",
  933=>"000000000",
  934=>"111111111",
  935=>"000000111",
  936=>"100000000",
  937=>"100100000",
  938=>"001000000",
  939=>"000000000",
  940=>"111111001",
  941=>"010000010",
  942=>"000000000",
  943=>"111111110",
  944=>"111111111",
  945=>"111111111",
  946=>"000000000",
  947=>"111111001",
  948=>"001000000",
  949=>"000001000",
  950=>"110111111",
  951=>"111111111",
  952=>"111111111",
  953=>"111111111",
  954=>"000100111",
  955=>"111110100",
  956=>"111111111",
  957=>"100101101",
  958=>"111111111",
  959=>"101000100",
  960=>"000000000",
  961=>"111111111",
  962=>"111111111",
  963=>"110110111",
  964=>"001001111",
  965=>"100100100",
  966=>"000000000",
  967=>"000000000",
  968=>"000000000",
  969=>"111111001",
  970=>"000000000",
  971=>"111111111",
  972=>"000000111",
  973=>"111111000",
  974=>"000000100",
  975=>"000000000",
  976=>"001011111",
  977=>"001000110",
  978=>"001001000",
  979=>"000000000",
  980=>"111001100",
  981=>"111000111",
  982=>"111101000",
  983=>"001011101",
  984=>"000000000",
  985=>"111111011",
  986=>"111100111",
  987=>"000011111",
  988=>"000000000",
  989=>"100000000",
  990=>"111111111",
  991=>"000110110",
  992=>"000000111",
  993=>"111111111",
  994=>"011000111",
  995=>"010111111",
  996=>"001011111",
  997=>"100000000",
  998=>"000000000",
  999=>"000000000",
  1000=>"000001001",
  1001=>"000000010",
  1002=>"010111111",
  1003=>"000000000",
  1004=>"100001101",
  1005=>"110111100",
  1006=>"111111111",
  1007=>"101111111",
  1008=>"000111110",
  1009=>"100110000",
  1010=>"000111111",
  1011=>"110100100",
  1012=>"000000000",
  1013=>"111111111",
  1014=>"110100100",
  1015=>"110100100",
  1016=>"111111111",
  1017=>"100100000",
  1018=>"000100000",
  1019=>"111111111",
  1020=>"000000000",
  1021=>"000011011",
  1022=>"111111111",
  1023=>"110110110",
  1024=>"000111111",
  1025=>"000000000",
  1026=>"101101111",
  1027=>"011011011",
  1028=>"000100100",
  1029=>"110110111",
  1030=>"111111010",
  1031=>"111111111",
  1032=>"111111111",
  1033=>"111111111",
  1034=>"110010000",
  1035=>"111111111",
  1036=>"110000100",
  1037=>"000000000",
  1038=>"001010111",
  1039=>"011011011",
  1040=>"111111110",
  1041=>"000010000",
  1042=>"111111111",
  1043=>"111111111",
  1044=>"111111111",
  1045=>"111111111",
  1046=>"000001001",
  1047=>"111111111",
  1048=>"100100100",
  1049=>"111011001",
  1050=>"111111111",
  1051=>"110000000",
  1052=>"000111111",
  1053=>"110000110",
  1054=>"111110000",
  1055=>"000000000",
  1056=>"101101111",
  1057=>"110110000",
  1058=>"000000000",
  1059=>"000110111",
  1060=>"001000000",
  1061=>"111011000",
  1062=>"000000000",
  1063=>"000000000",
  1064=>"011111111",
  1065=>"001001000",
  1066=>"000000000",
  1067=>"000000000",
  1068=>"101111111",
  1069=>"000000000",
  1070=>"110111000",
  1071=>"000100000",
  1072=>"111111111",
  1073=>"001111111",
  1074=>"000000100",
  1075=>"000110111",
  1076=>"000000000",
  1077=>"000000001",
  1078=>"111011000",
  1079=>"000000000",
  1080=>"100000000",
  1081=>"001000110",
  1082=>"000110110",
  1083=>"111111111",
  1084=>"000000000",
  1085=>"000000111",
  1086=>"111111111",
  1087=>"000000000",
  1088=>"011011111",
  1089=>"011101111",
  1090=>"000111111",
  1091=>"111111111",
  1092=>"111110110",
  1093=>"000000000",
  1094=>"111111111",
  1095=>"100111111",
  1096=>"111111111",
  1097=>"111111111",
  1098=>"000011111",
  1099=>"000001111",
  1100=>"100111000",
  1101=>"000000000",
  1102=>"100000000",
  1103=>"111111111",
  1104=>"111000000",
  1105=>"000000111",
  1106=>"111111110",
  1107=>"000000000",
  1108=>"111000000",
  1109=>"000000110",
  1110=>"101101111",
  1111=>"111001000",
  1112=>"000000000",
  1113=>"100100000",
  1114=>"111111000",
  1115=>"111101001",
  1116=>"000011011",
  1117=>"110111011",
  1118=>"000001100",
  1119=>"001001011",
  1120=>"111111010",
  1121=>"000001111",
  1122=>"010110000",
  1123=>"000000000",
  1124=>"000100111",
  1125=>"000100100",
  1126=>"000100000",
  1127=>"000100110",
  1128=>"111111111",
  1129=>"000000000",
  1130=>"000000111",
  1131=>"101111111",
  1132=>"000101110",
  1133=>"111111110",
  1134=>"000000000",
  1135=>"000011010",
  1136=>"000011110",
  1137=>"111111111",
  1138=>"011000000",
  1139=>"111111111",
  1140=>"111000000",
  1141=>"001000110",
  1142=>"000001001",
  1143=>"000000111",
  1144=>"000001101",
  1145=>"000001111",
  1146=>"000100101",
  1147=>"111111111",
  1148=>"100111111",
  1149=>"110110110",
  1150=>"110111111",
  1151=>"010000000",
  1152=>"000000000",
  1153=>"011001100",
  1154=>"001000110",
  1155=>"000000001",
  1156=>"000000000",
  1157=>"000000100",
  1158=>"110110000",
  1159=>"000111111",
  1160=>"000000000",
  1161=>"100011011",
  1162=>"000111111",
  1163=>"000000000",
  1164=>"111111111",
  1165=>"111111111",
  1166=>"111111111",
  1167=>"110110110",
  1168=>"111111111",
  1169=>"000000000",
  1170=>"000010011",
  1171=>"000000001",
  1172=>"111111011",
  1173=>"000010010",
  1174=>"000000000",
  1175=>"100000000",
  1176=>"111111100",
  1177=>"111111001",
  1178=>"111010000",
  1179=>"011111111",
  1180=>"000010111",
  1181=>"011001001",
  1182=>"111111111",
  1183=>"001000000",
  1184=>"111111001",
  1185=>"110111111",
  1186=>"000000111",
  1187=>"000000000",
  1188=>"000010111",
  1189=>"000010111",
  1190=>"101000101",
  1191=>"010000000",
  1192=>"000000000",
  1193=>"000001111",
  1194=>"000011011",
  1195=>"110111000",
  1196=>"010000110",
  1197=>"000000000",
  1198=>"111011011",
  1199=>"000000111",
  1200=>"000000000",
  1201=>"110110010",
  1202=>"111111111",
  1203=>"000100000",
  1204=>"100111011",
  1205=>"111111111",
  1206=>"000000000",
  1207=>"000000000",
  1208=>"000000100",
  1209=>"111111111",
  1210=>"000111101",
  1211=>"111111100",
  1212=>"000000000",
  1213=>"000000000",
  1214=>"000010000",
  1215=>"000000000",
  1216=>"000000000",
  1217=>"010000000",
  1218=>"111111111",
  1219=>"000000000",
  1220=>"000000000",
  1221=>"111111111",
  1222=>"000000110",
  1223=>"111111111",
  1224=>"000110000",
  1225=>"000100100",
  1226=>"000000000",
  1227=>"111111111",
  1228=>"111111111",
  1229=>"111111111",
  1230=>"000001111",
  1231=>"000000000",
  1232=>"000011011",
  1233=>"111111010",
  1234=>"000111111",
  1235=>"000000000",
  1236=>"000000100",
  1237=>"011011100",
  1238=>"111111011",
  1239=>"001111111",
  1240=>"100100000",
  1241=>"000111111",
  1242=>"111111110",
  1243=>"000000000",
  1244=>"010111111",
  1245=>"110111111",
  1246=>"000000000",
  1247=>"000000100",
  1248=>"011011111",
  1249=>"000111011",
  1250=>"100000111",
  1251=>"000100000",
  1252=>"000000000",
  1253=>"111111000",
  1254=>"001001001",
  1255=>"111111101",
  1256=>"000100100",
  1257=>"000000111",
  1258=>"100111111",
  1259=>"011001001",
  1260=>"100000100",
  1261=>"111111110",
  1262=>"101101000",
  1263=>"111111111",
  1264=>"001000000",
  1265=>"011000000",
  1266=>"000000000",
  1267=>"000000100",
  1268=>"111111111",
  1269=>"000100110",
  1270=>"001000011",
  1271=>"000000000",
  1272=>"000000000",
  1273=>"000000000",
  1274=>"001011111",
  1275=>"101111110",
  1276=>"100100000",
  1277=>"111011111",
  1278=>"011111111",
  1279=>"000100111",
  1280=>"011111111",
  1281=>"000100101",
  1282=>"111111111",
  1283=>"111101111",
  1284=>"000000100",
  1285=>"000000000",
  1286=>"000000000",
  1287=>"011001111",
  1288=>"110110000",
  1289=>"001000111",
  1290=>"111111111",
  1291=>"000000000",
  1292=>"111111000",
  1293=>"111110110",
  1294=>"111111110",
  1295=>"111101000",
  1296=>"011001000",
  1297=>"000000010",
  1298=>"111111111",
  1299=>"000000001",
  1300=>"111111111",
  1301=>"111001001",
  1302=>"110110110",
  1303=>"111110111",
  1304=>"010010111",
  1305=>"000110000",
  1306=>"111111111",
  1307=>"000000111",
  1308=>"100000111",
  1309=>"000000000",
  1310=>"010111111",
  1311=>"111111111",
  1312=>"000111111",
  1313=>"110001101",
  1314=>"000000000",
  1315=>"011000000",
  1316=>"100000100",
  1317=>"000000001",
  1318=>"000001001",
  1319=>"010000101",
  1320=>"001101100",
  1321=>"111111010",
  1322=>"111111111",
  1323=>"111111111",
  1324=>"000000000",
  1325=>"100111111",
  1326=>"111101000",
  1327=>"111111111",
  1328=>"111111111",
  1329=>"001001111",
  1330=>"000000000",
  1331=>"111111100",
  1332=>"111001001",
  1333=>"111111111",
  1334=>"000000000",
  1335=>"111111111",
  1336=>"000000000",
  1337=>"000000100",
  1338=>"000000000",
  1339=>"001001001",
  1340=>"000000000",
  1341=>"100100110",
  1342=>"000000000",
  1343=>"000000000",
  1344=>"000100111",
  1345=>"111110110",
  1346=>"111111110",
  1347=>"111111011",
  1348=>"000111000",
  1349=>"000001001",
  1350=>"000000011",
  1351=>"101100111",
  1352=>"000000000",
  1353=>"000000001",
  1354=>"000000000",
  1355=>"111111011",
  1356=>"011111111",
  1357=>"000000000",
  1358=>"111111111",
  1359=>"111001000",
  1360=>"111011110",
  1361=>"111101000",
  1362=>"011011000",
  1363=>"000000000",
  1364=>"111111111",
  1365=>"111110111",
  1366=>"000000000",
  1367=>"111111111",
  1368=>"111111100",
  1369=>"110111111",
  1370=>"111111111",
  1371=>"000101111",
  1372=>"111100100",
  1373=>"000000110",
  1374=>"000111101",
  1375=>"000000110",
  1376=>"000000011",
  1377=>"111111111",
  1378=>"100000000",
  1379=>"000000000",
  1380=>"000000000",
  1381=>"001000000",
  1382=>"000111111",
  1383=>"110000000",
  1384=>"111111111",
  1385=>"000001001",
  1386=>"011011011",
  1387=>"011111110",
  1388=>"100000000",
  1389=>"010110100",
  1390=>"111111000",
  1391=>"111111111",
  1392=>"000101111",
  1393=>"111001001",
  1394=>"001001001",
  1395=>"000111111",
  1396=>"000000000",
  1397=>"010111110",
  1398=>"010111101",
  1399=>"111111000",
  1400=>"110111111",
  1401=>"101111010",
  1402=>"111111111",
  1403=>"011111011",
  1404=>"110110110",
  1405=>"111111111",
  1406=>"000000000",
  1407=>"000000101",
  1408=>"010010000",
  1409=>"001111111",
  1410=>"000000000",
  1411=>"000000000",
  1412=>"000000000",
  1413=>"111111111",
  1414=>"111111111",
  1415=>"111111111",
  1416=>"111111111",
  1417=>"100010000",
  1418=>"000000000",
  1419=>"100111111",
  1420=>"111111111",
  1421=>"001000110",
  1422=>"110100111",
  1423=>"000000000",
  1424=>"001101001",
  1425=>"111111110",
  1426=>"000001000",
  1427=>"000000000",
  1428=>"000000000",
  1429=>"001001001",
  1430=>"011111111",
  1431=>"110110111",
  1432=>"000100000",
  1433=>"101100000",
  1434=>"000100110",
  1435=>"111111111",
  1436=>"000000000",
  1437=>"111111111",
  1438=>"111011111",
  1439=>"111111111",
  1440=>"000000000",
  1441=>"111101100",
  1442=>"101000101",
  1443=>"111001000",
  1444=>"000001000",
  1445=>"111111000",
  1446=>"001001100",
  1447=>"111001001",
  1448=>"111111000",
  1449=>"000000111",
  1450=>"000000000",
  1451=>"000100111",
  1452=>"000000010",
  1453=>"110000000",
  1454=>"000000111",
  1455=>"000000000",
  1456=>"000000000",
  1457=>"000000000",
  1458=>"000100111",
  1459=>"011000000",
  1460=>"001000000",
  1461=>"000000101",
  1462=>"000101101",
  1463=>"000100000",
  1464=>"000111110",
  1465=>"110111111",
  1466=>"000101100",
  1467=>"111111111",
  1468=>"000100111",
  1469=>"111111111",
  1470=>"000000000",
  1471=>"111110100",
  1472=>"000000000",
  1473=>"000111111",
  1474=>"000000000",
  1475=>"000000000",
  1476=>"000100100",
  1477=>"001011011",
  1478=>"001001111",
  1479=>"100000000",
  1480=>"111101111",
  1481=>"001001011",
  1482=>"001000101",
  1483=>"110111111",
  1484=>"000111111",
  1485=>"000000000",
  1486=>"000000000",
  1487=>"000011111",
  1488=>"101100000",
  1489=>"111100100",
  1490=>"111111111",
  1491=>"001001001",
  1492=>"110110110",
  1493=>"000000001",
  1494=>"100111111",
  1495=>"011000001",
  1496=>"000111111",
  1497=>"111111011",
  1498=>"000000000",
  1499=>"000000000",
  1500=>"111111111",
  1501=>"111111111",
  1502=>"000000000",
  1503=>"000000000",
  1504=>"111110111",
  1505=>"111111111",
  1506=>"011111111",
  1507=>"101001000",
  1508=>"011111111",
  1509=>"101111001",
  1510=>"110110000",
  1511=>"000000000",
  1512=>"100111111",
  1513=>"000000000",
  1514=>"000011000",
  1515=>"000000000",
  1516=>"000000000",
  1517=>"011101101",
  1518=>"111111111",
  1519=>"111111111",
  1520=>"001011001",
  1521=>"000000000",
  1522=>"110111111",
  1523=>"000101100",
  1524=>"000011111",
  1525=>"000000000",
  1526=>"000000001",
  1527=>"011011010",
  1528=>"000000000",
  1529=>"001011011",
  1530=>"110110111",
  1531=>"001000001",
  1532=>"111101111",
  1533=>"010111110",
  1534=>"011010111",
  1535=>"000000111",
  1536=>"000000000",
  1537=>"001000000",
  1538=>"000101100",
  1539=>"001000011",
  1540=>"000000011",
  1541=>"111111111",
  1542=>"111001000",
  1543=>"000000101",
  1544=>"000000000",
  1545=>"110111111",
  1546=>"011000000",
  1547=>"111111001",
  1548=>"110111111",
  1549=>"101010010",
  1550=>"000011101",
  1551=>"001011111",
  1552=>"111111000",
  1553=>"000100010",
  1554=>"000000000",
  1555=>"000000111",
  1556=>"111000000",
  1557=>"000000000",
  1558=>"000000111",
  1559=>"100100110",
  1560=>"100100110",
  1561=>"111111000",
  1562=>"000000000",
  1563=>"111011111",
  1564=>"000000000",
  1565=>"011010000",
  1566=>"110100110",
  1567=>"000000001",
  1568=>"000000000",
  1569=>"000000001",
  1570=>"000000001",
  1571=>"000000011",
  1572=>"111111011",
  1573=>"000000111",
  1574=>"111000000",
  1575=>"101101100",
  1576=>"111111001",
  1577=>"000000111",
  1578=>"000000000",
  1579=>"111111111",
  1580=>"110000100",
  1581=>"001001000",
  1582=>"000111111",
  1583=>"111000000",
  1584=>"100110110",
  1585=>"000000111",
  1586=>"000111110",
  1587=>"000011011",
  1588=>"111111000",
  1589=>"111100101",
  1590=>"000000000",
  1591=>"000011111",
  1592=>"000001000",
  1593=>"000000000",
  1594=>"111111111",
  1595=>"111110110",
  1596=>"000000111",
  1597=>"000000000",
  1598=>"111011001",
  1599=>"100100111",
  1600=>"000110110",
  1601=>"111111111",
  1602=>"111111111",
  1603=>"000000000",
  1604=>"000000000",
  1605=>"111000000",
  1606=>"110100111",
  1607=>"000000000",
  1608=>"011000000",
  1609=>"100000111",
  1610=>"000111110",
  1611=>"000000000",
  1612=>"000000100",
  1613=>"000000000",
  1614=>"100100000",
  1615=>"100000000",
  1616=>"000000000",
  1617=>"001001001",
  1618=>"111100000",
  1619=>"111100000",
  1620=>"000000001",
  1621=>"111110111",
  1622=>"001110100",
  1623=>"111111111",
  1624=>"011000101",
  1625=>"101100111",
  1626=>"111000000",
  1627=>"011001001",
  1628=>"000000000",
  1629=>"110110110",
  1630=>"111111000",
  1631=>"100100100",
  1632=>"111111111",
  1633=>"000000011",
  1634=>"111111100",
  1635=>"000000110",
  1636=>"101101111",
  1637=>"000110111",
  1638=>"111110110",
  1639=>"110111010",
  1640=>"111111111",
  1641=>"111111000",
  1642=>"000000001",
  1643=>"111111000",
  1644=>"111111000",
  1645=>"111011000",
  1646=>"000000000",
  1647=>"100000000",
  1648=>"010000111",
  1649=>"100111111",
  1650=>"111111111",
  1651=>"010111011",
  1652=>"000010000",
  1653=>"011011000",
  1654=>"111011111",
  1655=>"000000000",
  1656=>"110100111",
  1657=>"000000000",
  1658=>"101101000",
  1659=>"110111000",
  1660=>"110111100",
  1661=>"000000000",
  1662=>"000000000",
  1663=>"010111110",
  1664=>"000000000",
  1665=>"111000110",
  1666=>"000000000",
  1667=>"011010001",
  1668=>"111011011",
  1669=>"000000111",
  1670=>"111111110",
  1671=>"111111000",
  1672=>"111000000",
  1673=>"110000110",
  1674=>"011001001",
  1675=>"100111111",
  1676=>"001000001",
  1677=>"000010000",
  1678=>"111110000",
  1679=>"111010010",
  1680=>"000000000",
  1681=>"000000010",
  1682=>"000111111",
  1683=>"000111111",
  1684=>"110010011",
  1685=>"110111000",
  1686=>"111111100",
  1687=>"111000000",
  1688=>"111001001",
  1689=>"111110000",
  1690=>"111111111",
  1691=>"111000000",
  1692=>"011000000",
  1693=>"000000000",
  1694=>"000000000",
  1695=>"000000000",
  1696=>"110110101",
  1697=>"000110000",
  1698=>"010010000",
  1699=>"111111000",
  1700=>"000000000",
  1701=>"111111110",
  1702=>"000100110",
  1703=>"011011001",
  1704=>"000000000",
  1705=>"000000000",
  1706=>"000000000",
  1707=>"000000011",
  1708=>"111000000",
  1709=>"010110110",
  1710=>"000000000",
  1711=>"000000001",
  1712=>"000001000",
  1713=>"001011110",
  1714=>"110111000",
  1715=>"000000000",
  1716=>"100000100",
  1717=>"000111111",
  1718=>"000111111",
  1719=>"000101111",
  1720=>"011001001",
  1721=>"000000000",
  1722=>"000000000",
  1723=>"110000000",
  1724=>"000001111",
  1725=>"001001000",
  1726=>"000000000",
  1727=>"111111000",
  1728=>"011111111",
  1729=>"100110111",
  1730=>"011101101",
  1731=>"111000000",
  1732=>"111110000",
  1733=>"000000000",
  1734=>"100000000",
  1735=>"110110111",
  1736=>"111111110",
  1737=>"011011000",
  1738=>"000000000",
  1739=>"111001111",
  1740=>"111111101",
  1741=>"000111111",
  1742=>"111000110",
  1743=>"011000000",
  1744=>"101001000",
  1745=>"000001011",
  1746=>"111111111",
  1747=>"111111111",
  1748=>"111010000",
  1749=>"000000111",
  1750=>"000000000",
  1751=>"111010000",
  1752=>"010000000",
  1753=>"000100111",
  1754=>"000000101",
  1755=>"101111110",
  1756=>"000000000",
  1757=>"010010001",
  1758=>"000000000",
  1759=>"000000000",
  1760=>"001001111",
  1761=>"000111110",
  1762=>"111111111",
  1763=>"111111000",
  1764=>"001101111",
  1765=>"110000000",
  1766=>"111111111",
  1767=>"111001000",
  1768=>"000000000",
  1769=>"101111011",
  1770=>"000000101",
  1771=>"100000000",
  1772=>"011000000",
  1773=>"000000110",
  1774=>"000010001",
  1775=>"001111111",
  1776=>"100000000",
  1777=>"100101011",
  1778=>"111111000",
  1779=>"000100111",
  1780=>"011111100",
  1781=>"010110010",
  1782=>"011001011",
  1783=>"011011110",
  1784=>"010000000",
  1785=>"110111111",
  1786=>"111110100",
  1787=>"000000000",
  1788=>"010001100",
  1789=>"110111111",
  1790=>"101111001",
  1791=>"011010011",
  1792=>"000000011",
  1793=>"011011001",
  1794=>"000111111",
  1795=>"000110101",
  1796=>"000000000",
  1797=>"110111000",
  1798=>"111101000",
  1799=>"111100000",
  1800=>"000000000",
  1801=>"000000000",
  1802=>"001010000",
  1803=>"000000111",
  1804=>"111101111",
  1805=>"000000010",
  1806=>"111001111",
  1807=>"110001111",
  1808=>"000110000",
  1809=>"111111111",
  1810=>"111111111",
  1811=>"000000110",
  1812=>"111111000",
  1813=>"111000111",
  1814=>"111100000",
  1815=>"111111111",
  1816=>"100111111",
  1817=>"111111000",
  1818=>"111110111",
  1819=>"000000000",
  1820=>"001001000",
  1821=>"111000111",
  1822=>"000000111",
  1823=>"111111111",
  1824=>"111111100",
  1825=>"001010111",
  1826=>"000011111",
  1827=>"111111000",
  1828=>"111110010",
  1829=>"111101101",
  1830=>"000000001",
  1831=>"111111101",
  1832=>"000011011",
  1833=>"000000000",
  1834=>"101101111",
  1835=>"111100000",
  1836=>"111111000",
  1837=>"001111011",
  1838=>"000001111",
  1839=>"000000000",
  1840=>"100100110",
  1841=>"000100110",
  1842=>"000000001",
  1843=>"110110011",
  1844=>"111101111",
  1845=>"001011000",
  1846=>"100111111",
  1847=>"000000111",
  1848=>"110000000",
  1849=>"011101111",
  1850=>"000001000",
  1851=>"001000110",
  1852=>"000000110",
  1853=>"111111000",
  1854=>"100111111",
  1855=>"000000000",
  1856=>"000111111",
  1857=>"111111111",
  1858=>"111111000",
  1859=>"000110111",
  1860=>"000000111",
  1861=>"000000100",
  1862=>"000000110",
  1863=>"111111000",
  1864=>"000000110",
  1865=>"111111111",
  1866=>"111111111",
  1867=>"001001110",
  1868=>"101000000",
  1869=>"111011000",
  1870=>"110111111",
  1871=>"100100001",
  1872=>"110110000",
  1873=>"000000011",
  1874=>"000000111",
  1875=>"100000000",
  1876=>"001001001",
  1877=>"011001001",
  1878=>"111111000",
  1879=>"111111000",
  1880=>"111111000",
  1881=>"101101101",
  1882=>"000000001",
  1883=>"000000000",
  1884=>"011111001",
  1885=>"111000000",
  1886=>"001111111",
  1887=>"110110100",
  1888=>"000001101",
  1889=>"000000000",
  1890=>"111001111",
  1891=>"111101111",
  1892=>"111111000",
  1893=>"111111111",
  1894=>"000000000",
  1895=>"000110111",
  1896=>"001111011",
  1897=>"000000011",
  1898=>"000011011",
  1899=>"000101101",
  1900=>"011100100",
  1901=>"000000000",
  1902=>"100111111",
  1903=>"011000111",
  1904=>"011000000",
  1905=>"101000000",
  1906=>"111000000",
  1907=>"011001010",
  1908=>"111111001",
  1909=>"001001001",
  1910=>"110000000",
  1911=>"000000000",
  1912=>"000000000",
  1913=>"111011000",
  1914=>"000010000",
  1915=>"100111110",
  1916=>"111011001",
  1917=>"111010111",
  1918=>"111111111",
  1919=>"111001000",
  1920=>"000100110",
  1921=>"111010000",
  1922=>"111001000",
  1923=>"111100110",
  1924=>"111111111",
  1925=>"000000000",
  1926=>"111111000",
  1927=>"100111111",
  1928=>"100000100",
  1929=>"000111111",
  1930=>"000000000",
  1931=>"111111111",
  1932=>"101110111",
  1933=>"011010000",
  1934=>"001011001",
  1935=>"000000000",
  1936=>"000000000",
  1937=>"000000000",
  1938=>"111010010",
  1939=>"000110111",
  1940=>"000111001",
  1941=>"000111000",
  1942=>"011011001",
  1943=>"000100110",
  1944=>"111111111",
  1945=>"000110110",
  1946=>"000000010",
  1947=>"000110000",
  1948=>"000000000",
  1949=>"111111111",
  1950=>"000000000",
  1951=>"000111111",
  1952=>"111000000",
  1953=>"100110110",
  1954=>"111111111",
  1955=>"111111000",
  1956=>"111111110",
  1957=>"111111111",
  1958=>"111111111",
  1959=>"000000110",
  1960=>"000000000",
  1961=>"101111100",
  1962=>"111111101",
  1963=>"000100100",
  1964=>"000000011",
  1965=>"101100100",
  1966=>"000000000",
  1967=>"000000000",
  1968=>"110111000",
  1969=>"111011011",
  1970=>"000000000",
  1971=>"000100110",
  1972=>"111110111",
  1973=>"000000111",
  1974=>"000000001",
  1975=>"110111111",
  1976=>"000000011",
  1977=>"000000100",
  1978=>"111000000",
  1979=>"111111011",
  1980=>"011111111",
  1981=>"001000111",
  1982=>"011111111",
  1983=>"001000001",
  1984=>"000000111",
  1985=>"011000000",
  1986=>"000010111",
  1987=>"010000000",
  1988=>"000100100",
  1989=>"100000001",
  1990=>"111110010",
  1991=>"011101000",
  1992=>"000000000",
  1993=>"011000100",
  1994=>"000000110",
  1995=>"111111011",
  1996=>"111111000",
  1997=>"110111010",
  1998=>"100010110",
  1999=>"101111100",
  2000=>"111000000",
  2001=>"111111011",
  2002=>"011111011",
  2003=>"011111110",
  2004=>"000000110",
  2005=>"000101111",
  2006=>"000000000",
  2007=>"000000000",
  2008=>"000000101",
  2009=>"000000000",
  2010=>"000010000",
  2011=>"000111111",
  2012=>"000001011",
  2013=>"000000000",
  2014=>"111000000",
  2015=>"011011011",
  2016=>"000011000",
  2017=>"000100000",
  2018=>"110100111",
  2019=>"100011111",
  2020=>"111110000",
  2021=>"111110110",
  2022=>"111110100",
  2023=>"100110110",
  2024=>"000110111",
  2025=>"000110110",
  2026=>"011011011",
  2027=>"000000011",
  2028=>"001000111",
  2029=>"000011011",
  2030=>"000000101",
  2031=>"000000000",
  2032=>"000011001",
  2033=>"111111111",
  2034=>"011011011",
  2035=>"101100111",
  2036=>"000000000",
  2037=>"111111111",
  2038=>"000001111",
  2039=>"011111111",
  2040=>"000001110",
  2041=>"101101001",
  2042=>"000000000",
  2043=>"111111111",
  2044=>"000011011",
  2045=>"111110110",
  2046=>"101111110",
  2047=>"000001111",
  2048=>"001000000",
  2049=>"110000000",
  2050=>"111111111",
  2051=>"110111111",
  2052=>"111111111",
  2053=>"000010011",
  2054=>"111101000",
  2055=>"000000111",
  2056=>"000000011",
  2057=>"111111001",
  2058=>"000111111",
  2059=>"111111111",
  2060=>"111111111",
  2061=>"101111101",
  2062=>"000100111",
  2063=>"000000000",
  2064=>"110000000",
  2065=>"000101111",
  2066=>"000000101",
  2067=>"100110110",
  2068=>"000000111",
  2069=>"111001000",
  2070=>"111111111",
  2071=>"001000000",
  2072=>"111111001",
  2073=>"111111000",
  2074=>"111111110",
  2075=>"011000111",
  2076=>"000101111",
  2077=>"101101000",
  2078=>"011000011",
  2079=>"000111010",
  2080=>"111111111",
  2081=>"000111111",
  2082=>"000000110",
  2083=>"111000001",
  2084=>"000001000",
  2085=>"111111111",
  2086=>"011000001",
  2087=>"111000000",
  2088=>"011100111",
  2089=>"111000000",
  2090=>"001001111",
  2091=>"000100110",
  2092=>"010110111",
  2093=>"111001000",
  2094=>"000111111",
  2095=>"000000111",
  2096=>"000000111",
  2097=>"110111000",
  2098=>"101111011",
  2099=>"111111111",
  2100=>"011001001",
  2101=>"111111011",
  2102=>"000011111",
  2103=>"000010110",
  2104=>"000001000",
  2105=>"100000101",
  2106=>"101101100",
  2107=>"111011010",
  2108=>"000000000",
  2109=>"001001001",
  2110=>"011111111",
  2111=>"111001000",
  2112=>"000111111",
  2113=>"001111111",
  2114=>"100100111",
  2115=>"000110111",
  2116=>"100111110",
  2117=>"000000000",
  2118=>"000000000",
  2119=>"111111000",
  2120=>"111111111",
  2121=>"100100101",
  2122=>"000000000",
  2123=>"001000000",
  2124=>"000111111",
  2125=>"101000000",
  2126=>"111000000",
  2127=>"001101101",
  2128=>"000100111",
  2129=>"001111111",
  2130=>"110110100",
  2131=>"111111000",
  2132=>"111000000",
  2133=>"000100100",
  2134=>"111000000",
  2135=>"111010000",
  2136=>"000000001",
  2137=>"111111101",
  2138=>"110010010",
  2139=>"111100000",
  2140=>"111111111",
  2141=>"010000000",
  2142=>"000110110",
  2143=>"000111110",
  2144=>"101011111",
  2145=>"011011100",
  2146=>"110111111",
  2147=>"111000110",
  2148=>"001101111",
  2149=>"100000111",
  2150=>"111111110",
  2151=>"000000101",
  2152=>"110111001",
  2153=>"110111111",
  2154=>"000000000",
  2155=>"000000010",
  2156=>"101000111",
  2157=>"111110111",
  2158=>"000000000",
  2159=>"000010111",
  2160=>"011100111",
  2161=>"111110111",
  2162=>"111000000",
  2163=>"110111000",
  2164=>"111111010",
  2165=>"110100000",
  2166=>"111111000",
  2167=>"000000111",
  2168=>"000000111",
  2169=>"111010111",
  2170=>"100000000",
  2171=>"000000000",
  2172=>"000111111",
  2173=>"111111100",
  2174=>"110111111",
  2175=>"011010000",
  2176=>"111111000",
  2177=>"001010111",
  2178=>"111001011",
  2179=>"001010010",
  2180=>"111000000",
  2181=>"111000000",
  2182=>"000011110",
  2183=>"000111111",
  2184=>"111111111",
  2185=>"111000100",
  2186=>"111111000",
  2187=>"000000001",
  2188=>"011111111",
  2189=>"000111110",
  2190=>"111111111",
  2191=>"000000000",
  2192=>"111000000",
  2193=>"001000000",
  2194=>"000111111",
  2195=>"000000111",
  2196=>"111000001",
  2197=>"001100100",
  2198=>"000001000",
  2199=>"111101000",
  2200=>"111000110",
  2201=>"000001011",
  2202=>"110010000",
  2203=>"000011011",
  2204=>"111110110",
  2205=>"100000001",
  2206=>"000100000",
  2207=>"000010111",
  2208=>"000000000",
  2209=>"111100111",
  2210=>"000000000",
  2211=>"000001000",
  2212=>"110011011",
  2213=>"111111111",
  2214=>"110111111",
  2215=>"111111000",
  2216=>"000000100",
  2217=>"000111111",
  2218=>"000000000",
  2219=>"100111010",
  2220=>"010111111",
  2221=>"010111010",
  2222=>"111111101",
  2223=>"100111111",
  2224=>"000000111",
  2225=>"111111011",
  2226=>"111111111",
  2227=>"111111111",
  2228=>"111011000",
  2229=>"100000000",
  2230=>"000111000",
  2231=>"101000111",
  2232=>"000101111",
  2233=>"000000111",
  2234=>"110100100",
  2235=>"110000100",
  2236=>"110110111",
  2237=>"011111111",
  2238=>"000110110",
  2239=>"001011011",
  2240=>"111000000",
  2241=>"110111111",
  2242=>"000111011",
  2243=>"000010010",
  2244=>"001000111",
  2245=>"000111111",
  2246=>"001000000",
  2247=>"011011101",
  2248=>"000000111",
  2249=>"000000111",
  2250=>"110000110",
  2251=>"101000000",
  2252=>"100111111",
  2253=>"000000111",
  2254=>"000000111",
  2255=>"110000000",
  2256=>"001001000",
  2257=>"001000000",
  2258=>"100100111",
  2259=>"000000111",
  2260=>"111111001",
  2261=>"110110111",
  2262=>"001000111",
  2263=>"000000111",
  2264=>"000000000",
  2265=>"011111111",
  2266=>"000000000",
  2267=>"000000000",
  2268=>"111010110",
  2269=>"000000000",
  2270=>"000111111",
  2271=>"010010000",
  2272=>"101111111",
  2273=>"000111101",
  2274=>"000111110",
  2275=>"110101000",
  2276=>"111111100",
  2277=>"011000001",
  2278=>"000000000",
  2279=>"111111000",
  2280=>"000111111",
  2281=>"111111010",
  2282=>"111111111",
  2283=>"001111111",
  2284=>"110101001",
  2285=>"011111011",
  2286=>"111111111",
  2287=>"111111111",
  2288=>"000000000",
  2289=>"000000001",
  2290=>"111110111",
  2291=>"111100100",
  2292=>"100010110",
  2293=>"100111111",
  2294=>"000100100",
  2295=>"000000001",
  2296=>"111000111",
  2297=>"111011111",
  2298=>"000000110",
  2299=>"110111110",
  2300=>"111000001",
  2301=>"100111111",
  2302=>"110110000",
  2303=>"000101100",
  2304=>"111111111",
  2305=>"110000000",
  2306=>"100111111",
  2307=>"111100100",
  2308=>"011111111",
  2309=>"000000000",
  2310=>"000111111",
  2311=>"010000000",
  2312=>"110111000",
  2313=>"111000110",
  2314=>"011111111",
  2315=>"111111001",
  2316=>"111000111",
  2317=>"000011111",
  2318=>"111111111",
  2319=>"111100110",
  2320=>"101000000",
  2321=>"100110111",
  2322=>"111000000",
  2323=>"111000110",
  2324=>"000110100",
  2325=>"000101111",
  2326=>"101100000",
  2327=>"111111111",
  2328=>"111000000",
  2329=>"110000100",
  2330=>"000111110",
  2331=>"000000111",
  2332=>"000100010",
  2333=>"110111011",
  2334=>"000100111",
  2335=>"111111111",
  2336=>"000001111",
  2337=>"000100000",
  2338=>"000111100",
  2339=>"100100111",
  2340=>"000000000",
  2341=>"111111111",
  2342=>"011111011",
  2343=>"010111110",
  2344=>"111000000",
  2345=>"111111000",
  2346=>"000000110",
  2347=>"001000111",
  2348=>"111010000",
  2349=>"111011111",
  2350=>"111001001",
  2351=>"000000111",
  2352=>"000000000",
  2353=>"011000000",
  2354=>"110010111",
  2355=>"100000111",
  2356=>"111111000",
  2357=>"111110000",
  2358=>"011001001",
  2359=>"000110111",
  2360=>"100100000",
  2361=>"111111101",
  2362=>"111000000",
  2363=>"000111111",
  2364=>"100101111",
  2365=>"001000010",
  2366=>"000000000",
  2367=>"111111110",
  2368=>"111010000",
  2369=>"111011011",
  2370=>"111111111",
  2371=>"111000000",
  2372=>"010000000",
  2373=>"000000000",
  2374=>"000000000",
  2375=>"111110001",
  2376=>"000000110",
  2377=>"000111111",
  2378=>"000111111",
  2379=>"000000111",
  2380=>"000000111",
  2381=>"011111000",
  2382=>"000000000",
  2383=>"000000001",
  2384=>"100111100",
  2385=>"010000100",
  2386=>"010111110",
  2387=>"110110111",
  2388=>"000000110",
  2389=>"001011011",
  2390=>"000000100",
  2391=>"111111000",
  2392=>"000000111",
  2393=>"111111000",
  2394=>"111110111",
  2395=>"111111111",
  2396=>"111101001",
  2397=>"111111111",
  2398=>"110111111",
  2399=>"011011000",
  2400=>"000001111",
  2401=>"111001000",
  2402=>"100000100",
  2403=>"000000000",
  2404=>"001001001",
  2405=>"111110000",
  2406=>"000100111",
  2407=>"101000111",
  2408=>"000000111",
  2409=>"101000111",
  2410=>"000000000",
  2411=>"111111110",
  2412=>"000001101",
  2413=>"000000000",
  2414=>"000000000",
  2415=>"111101000",
  2416=>"000011110",
  2417=>"000000000",
  2418=>"000000111",
  2419=>"111111100",
  2420=>"111111110",
  2421=>"110000111",
  2422=>"100000000",
  2423=>"011000000",
  2424=>"000101001",
  2425=>"100111001",
  2426=>"100000000",
  2427=>"111111110",
  2428=>"111001111",
  2429=>"011001000",
  2430=>"000111111",
  2431=>"000100111",
  2432=>"000011011",
  2433=>"100000000",
  2434=>"000000111",
  2435=>"111001000",
  2436=>"000111111",
  2437=>"000111111",
  2438=>"000111110",
  2439=>"000000110",
  2440=>"111000000",
  2441=>"011111101",
  2442=>"111111111",
  2443=>"000000000",
  2444=>"111111001",
  2445=>"011011011",
  2446=>"111100111",
  2447=>"000000010",
  2448=>"001011000",
  2449=>"000110110",
  2450=>"000000111",
  2451=>"111110100",
  2452=>"000001111",
  2453=>"101110000",
  2454=>"111110111",
  2455=>"110100001",
  2456=>"000000111",
  2457=>"100000111",
  2458=>"001000111",
  2459=>"110111111",
  2460=>"000000000",
  2461=>"000000000",
  2462=>"111111000",
  2463=>"000000000",
  2464=>"100000000",
  2465=>"111111100",
  2466=>"111001000",
  2467=>"001000000",
  2468=>"110000111",
  2469=>"111111000",
  2470=>"011011000",
  2471=>"001000000",
  2472=>"101000000",
  2473=>"011000000",
  2474=>"100110110",
  2475=>"111100000",
  2476=>"000111111",
  2477=>"000001000",
  2478=>"000111111",
  2479=>"011111000",
  2480=>"111111111",
  2481=>"011110111",
  2482=>"000000000",
  2483=>"011000000",
  2484=>"001111111",
  2485=>"111111111",
  2486=>"110000111",
  2487=>"101110000",
  2488=>"000000111",
  2489=>"010000111",
  2490=>"111111111",
  2491=>"110110000",
  2492=>"000000111",
  2493=>"011001111",
  2494=>"111000000",
  2495=>"100110000",
  2496=>"000011011",
  2497=>"000111111",
  2498=>"000111111",
  2499=>"110111000",
  2500=>"111000000",
  2501=>"010000000",
  2502=>"001000000",
  2503=>"111000000",
  2504=>"100000100",
  2505=>"000000111",
  2506=>"111111000",
  2507=>"111111111",
  2508=>"000111110",
  2509=>"000111111",
  2510=>"011111000",
  2511=>"001000000",
  2512=>"000111111",
  2513=>"001111000",
  2514=>"001111111",
  2515=>"101000101",
  2516=>"100111100",
  2517=>"000000000",
  2518=>"100000000",
  2519=>"111001011",
  2520=>"000100000",
  2521=>"101111111",
  2522=>"111111000",
  2523=>"111000000",
  2524=>"110111100",
  2525=>"001000101",
  2526=>"111111011",
  2527=>"111111000",
  2528=>"011011111",
  2529=>"111000000",
  2530=>"111101101",
  2531=>"101111111",
  2532=>"111110110",
  2533=>"111100000",
  2534=>"111111111",
  2535=>"000000111",
  2536=>"000110111",
  2537=>"000000000",
  2538=>"000000011",
  2539=>"000001001",
  2540=>"000110111",
  2541=>"011111010",
  2542=>"111111101",
  2543=>"111111111",
  2544=>"111000000",
  2545=>"000000000",
  2546=>"111000000",
  2547=>"000001101",
  2548=>"000000100",
  2549=>"000000000",
  2550=>"111111111",
  2551=>"000000111",
  2552=>"000111100",
  2553=>"010111111",
  2554=>"110111111",
  2555=>"000000000",
  2556=>"111111000",
  2557=>"000110100",
  2558=>"111111100",
  2559=>"111000000",
  2560=>"000010100",
  2561=>"111111110",
  2562=>"101101101",
  2563=>"110110110",
  2564=>"000000110",
  2565=>"000000000",
  2566=>"111111011",
  2567=>"101001101",
  2568=>"010110111",
  2569=>"000000111",
  2570=>"111111111",
  2571=>"111111001",
  2572=>"110110110",
  2573=>"000000000",
  2574=>"000101111",
  2575=>"010010111",
  2576=>"100000100",
  2577=>"111010110",
  2578=>"111000000",
  2579=>"100100100",
  2580=>"101100100",
  2581=>"111000111",
  2582=>"011001001",
  2583=>"101011011",
  2584=>"000100110",
  2585=>"100000000",
  2586=>"000000100",
  2587=>"110100000",
  2588=>"100000000",
  2589=>"111111111",
  2590=>"111111011",
  2591=>"110000000",
  2592=>"111111111",
  2593=>"110100010",
  2594=>"110111111",
  2595=>"000001001",
  2596=>"000001001",
  2597=>"001000000",
  2598=>"100000101",
  2599=>"000100010",
  2600=>"111111111",
  2601=>"111011001",
  2602=>"000000000",
  2603=>"110010010",
  2604=>"111111110",
  2605=>"111111100",
  2606=>"101001001",
  2607=>"111111111",
  2608=>"001001001",
  2609=>"111111011",
  2610=>"111101001",
  2611=>"000100100",
  2612=>"111111111",
  2613=>"111000000",
  2614=>"110110000",
  2615=>"010000110",
  2616=>"101000000",
  2617=>"100000001",
  2618=>"010110111",
  2619=>"000100101",
  2620=>"111111010",
  2621=>"010000001",
  2622=>"011000000",
  2623=>"100111111",
  2624=>"000000001",
  2625=>"001000000",
  2626=>"001001111",
  2627=>"000111111",
  2628=>"110110110",
  2629=>"001001011",
  2630=>"000000110",
  2631=>"101101101",
  2632=>"000001101",
  2633=>"001001011",
  2634=>"111111111",
  2635=>"101101101",
  2636=>"000111110",
  2637=>"000000000",
  2638=>"111110110",
  2639=>"101001001",
  2640=>"101101101",
  2641=>"001000000",
  2642=>"000000000",
  2643=>"100110110",
  2644=>"010010010",
  2645=>"100000001",
  2646=>"100100100",
  2647=>"001001011",
  2648=>"110110010",
  2649=>"101000111",
  2650=>"111011010",
  2651=>"011011011",
  2652=>"101000000",
  2653=>"000000000",
  2654=>"000000010",
  2655=>"111011111",
  2656=>"000010010",
  2657=>"000000000",
  2658=>"011000000",
  2659=>"111111111",
  2660=>"000000010",
  2661=>"000111111",
  2662=>"011001110",
  2663=>"111100000",
  2664=>"000111111",
  2665=>"101111111",
  2666=>"000000100",
  2667=>"111111110",
  2668=>"000000000",
  2669=>"111111111",
  2670=>"111011111",
  2671=>"010010110",
  2672=>"110000000",
  2673=>"001001111",
  2674=>"111011111",
  2675=>"011000010",
  2676=>"000001011",
  2677=>"110110110",
  2678=>"000000000",
  2679=>"111100000",
  2680=>"111101101",
  2681=>"111111001",
  2682=>"011001000",
  2683=>"000000000",
  2684=>"110001000",
  2685=>"111111010",
  2686=>"001000000",
  2687=>"001001000",
  2688=>"000000001",
  2689=>"000000000",
  2690=>"000000000",
  2691=>"011011011",
  2692=>"111100000",
  2693=>"111010110",
  2694=>"101111111",
  2695=>"111000000",
  2696=>"010000000",
  2697=>"101101101",
  2698=>"110110010",
  2699=>"111111011",
  2700=>"100100101",
  2701=>"000000000",
  2702=>"000100110",
  2703=>"111000000",
  2704=>"101000100",
  2705=>"111101101",
  2706=>"110111000",
  2707=>"000000011",
  2708=>"111111111",
  2709=>"111000000",
  2710=>"000000000",
  2711=>"000101101",
  2712=>"000001100",
  2713=>"111001001",
  2714=>"111110010",
  2715=>"000000000",
  2716=>"000000100",
  2717=>"100100001",
  2718=>"111010111",
  2719=>"010010111",
  2720=>"111111111",
  2721=>"000000000",
  2722=>"110111010",
  2723=>"111111111",
  2724=>"110000001",
  2725=>"011111100",
  2726=>"001001000",
  2727=>"110110110",
  2728=>"000010000",
  2729=>"101100101",
  2730=>"000000000",
  2731=>"100001111",
  2732=>"000011000",
  2733=>"100110111",
  2734=>"000000000",
  2735=>"101101101",
  2736=>"100100110",
  2737=>"001111001",
  2738=>"011111011",
  2739=>"100000000",
  2740=>"111111000",
  2741=>"000000000",
  2742=>"010010011",
  2743=>"100011111",
  2744=>"101111101",
  2745=>"110111111",
  2746=>"111101101",
  2747=>"010010110",
  2748=>"000000000",
  2749=>"010110010",
  2750=>"111111110",
  2751=>"001000000",
  2752=>"010111010",
  2753=>"001000000",
  2754=>"111000000",
  2755=>"001000001",
  2756=>"111111111",
  2757=>"001001000",
  2758=>"010010011",
  2759=>"101001001",
  2760=>"000000001",
  2761=>"101101000",
  2762=>"000001111",
  2763=>"111111111",
  2764=>"110111110",
  2765=>"001001110",
  2766=>"001000000",
  2767=>"000001000",
  2768=>"000000100",
  2769=>"100100111",
  2770=>"000000000",
  2771=>"000000000",
  2772=>"100110010",
  2773=>"000001001",
  2774=>"111111001",
  2775=>"011011011",
  2776=>"111111001",
  2777=>"000110110",
  2778=>"110111111",
  2779=>"100101001",
  2780=>"000000100",
  2781=>"111001100",
  2782=>"000000000",
  2783=>"001000100",
  2784=>"000000000",
  2785=>"000000010",
  2786=>"111111111",
  2787=>"000000000",
  2788=>"010110010",
  2789=>"000100001",
  2790=>"000000010",
  2791=>"001001001",
  2792=>"000000000",
  2793=>"111111010",
  2794=>"111110010",
  2795=>"101100100",
  2796=>"101101111",
  2797=>"111111101",
  2798=>"000100111",
  2799=>"111100000",
  2800=>"100000100",
  2801=>"011100100",
  2802=>"111111010",
  2803=>"111001000",
  2804=>"000000001",
  2805=>"001000110",
  2806=>"010110111",
  2807=>"000000101",
  2808=>"111111111",
  2809=>"100111111",
  2810=>"000000000",
  2811=>"100100100",
  2812=>"001000000",
  2813=>"000000000",
  2814=>"000111111",
  2815=>"000000000",
  2816=>"001001001",
  2817=>"011001000",
  2818=>"000111111",
  2819=>"010111011",
  2820=>"111111010",
  2821=>"000000000",
  2822=>"000000101",
  2823=>"010010000",
  2824=>"110110110",
  2825=>"010011111",
  2826=>"111111110",
  2827=>"110010010",
  2828=>"000000001",
  2829=>"001000010",
  2830=>"000001001",
  2831=>"001001100",
  2832=>"001111111",
  2833=>"000000000",
  2834=>"001000000",
  2835=>"111110111",
  2836=>"010011011",
  2837=>"111111111",
  2838=>"000000000",
  2839=>"010000000",
  2840=>"100100100",
  2841=>"101000000",
  2842=>"000010000",
  2843=>"000000100",
  2844=>"110100100",
  2845=>"000010000",
  2846=>"010000000",
  2847=>"111001100",
  2848=>"100100011",
  2849=>"000111111",
  2850=>"000110110",
  2851=>"001111110",
  2852=>"110110110",
  2853=>"000010111",
  2854=>"001000011",
  2855=>"000111110",
  2856=>"000001000",
  2857=>"101001000",
  2858=>"010010010",
  2859=>"000000010",
  2860=>"000000000",
  2861=>"010110100",
  2862=>"000000111",
  2863=>"000001001",
  2864=>"000000000",
  2865=>"000010011",
  2866=>"111001101",
  2867=>"111000000",
  2868=>"010111110",
  2869=>"111110000",
  2870=>"111111101",
  2871=>"010110111",
  2872=>"000000000",
  2873=>"101001111",
  2874=>"101101101",
  2875=>"010110010",
  2876=>"110010011",
  2877=>"001011000",
  2878=>"000000000",
  2879=>"000000000",
  2880=>"000000000",
  2881=>"000000000",
  2882=>"000000000",
  2883=>"000000000",
  2884=>"010110111",
  2885=>"111111111",
  2886=>"000000000",
  2887=>"111110010",
  2888=>"111111111",
  2889=>"111111111",
  2890=>"111100100",
  2891=>"001101101",
  2892=>"000000001",
  2893=>"001000001",
  2894=>"111111001",
  2895=>"110100100",
  2896=>"011011011",
  2897=>"001001001",
  2898=>"000101111",
  2899=>"101000001",
  2900=>"000000001",
  2901=>"011111000",
  2902=>"111111111",
  2903=>"001001000",
  2904=>"110111111",
  2905=>"000000101",
  2906=>"110110111",
  2907=>"100101100",
  2908=>"000110111",
  2909=>"000000100",
  2910=>"111011011",
  2911=>"111111100",
  2912=>"001111111",
  2913=>"111100100",
  2914=>"111111110",
  2915=>"000000101",
  2916=>"110110110",
  2917=>"010010011",
  2918=>"001000000",
  2919=>"010110111",
  2920=>"000100000",
  2921=>"011010010",
  2922=>"001000101",
  2923=>"100101111",
  2924=>"011010110",
  2925=>"110101101",
  2926=>"000010010",
  2927=>"000100101",
  2928=>"101001000",
  2929=>"000000000",
  2930=>"111111011",
  2931=>"011011011",
  2932=>"111000000",
  2933=>"001111111",
  2934=>"000000000",
  2935=>"010000000",
  2936=>"101100101",
  2937=>"111001101",
  2938=>"101001001",
  2939=>"001101101",
  2940=>"101100111",
  2941=>"111111000",
  2942=>"010010111",
  2943=>"001100001",
  2944=>"110110110",
  2945=>"101001001",
  2946=>"000000000",
  2947=>"000000000",
  2948=>"011101111",
  2949=>"100101100",
  2950=>"111000000",
  2951=>"111111101",
  2952=>"110110110",
  2953=>"111111011",
  2954=>"001001000",
  2955=>"111111111",
  2956=>"000111111",
  2957=>"011111010",
  2958=>"001111111",
  2959=>"000000000",
  2960=>"100100100",
  2961=>"000000000",
  2962=>"100111110",
  2963=>"000000000",
  2964=>"110000100",
  2965=>"000010000",
  2966=>"011001001",
  2967=>"110100100",
  2968=>"101101101",
  2969=>"000000100",
  2970=>"010110010",
  2971=>"010010010",
  2972=>"010011011",
  2973=>"111101111",
  2974=>"101101111",
  2975=>"111111111",
  2976=>"001000000",
  2977=>"101110100",
  2978=>"010110010",
  2979=>"111111111",
  2980=>"011111010",
  2981=>"101101111",
  2982=>"100000111",
  2983=>"100111111",
  2984=>"100000000",
  2985=>"001001000",
  2986=>"110110010",
  2987=>"000000000",
  2988=>"111001001",
  2989=>"000000110",
  2990=>"100010011",
  2991=>"001000000",
  2992=>"000000100",
  2993=>"111111011",
  2994=>"000000101",
  2995=>"000000000",
  2996=>"000000101",
  2997=>"000000000",
  2998=>"110000100",
  2999=>"111101101",
  3000=>"111111110",
  3001=>"111101101",
  3002=>"100000001",
  3003=>"010011111",
  3004=>"000010000",
  3005=>"001001001",
  3006=>"000101111",
  3007=>"000000000",
  3008=>"001011001",
  3009=>"001001001",
  3010=>"011111111",
  3011=>"001000000",
  3012=>"110111010",
  3013=>"000001001",
  3014=>"000000000",
  3015=>"000101111",
  3016=>"000001001",
  3017=>"000110101",
  3018=>"000000101",
  3019=>"111011111",
  3020=>"010010000",
  3021=>"101111000",
  3022=>"001001101",
  3023=>"111111111",
  3024=>"100100000",
  3025=>"100100100",
  3026=>"001001011",
  3027=>"000000101",
  3028=>"000000011",
  3029=>"000010110",
  3030=>"111111110",
  3031=>"011011011",
  3032=>"000101111",
  3033=>"100101001",
  3034=>"000001011",
  3035=>"001000110",
  3036=>"000000011",
  3037=>"000000000",
  3038=>"011011111",
  3039=>"011001001",
  3040=>"000000111",
  3041=>"111111111",
  3042=>"001001001",
  3043=>"000000100",
  3044=>"110111101",
  3045=>"111001111",
  3046=>"000000000",
  3047=>"000100000",
  3048=>"111111111",
  3049=>"010000010",
  3050=>"110000000",
  3051=>"011111111",
  3052=>"000000111",
  3053=>"010100101",
  3054=>"111111111",
  3055=>"101000000",
  3056=>"001000000",
  3057=>"000000000",
  3058=>"000000000",
  3059=>"001111011",
  3060=>"111111111",
  3061=>"011111010",
  3062=>"000000001",
  3063=>"101101101",
  3064=>"011011111",
  3065=>"000101101",
  3066=>"111000001",
  3067=>"000000000",
  3068=>"111000010",
  3069=>"000000000",
  3070=>"100111111",
  3071=>"000101111",
  3072=>"000000000",
  3073=>"000100111",
  3074=>"111000000",
  3075=>"111111111",
  3076=>"111001111",
  3077=>"111101111",
  3078=>"111101001",
  3079=>"100000111",
  3080=>"000000111",
  3081=>"111111111",
  3082=>"000000000",
  3083=>"110100100",
  3084=>"000000000",
  3085=>"001001100",
  3086=>"100110111",
  3087=>"001001001",
  3088=>"000000000",
  3089=>"000111111",
  3090=>"000000000",
  3091=>"111111111",
  3092=>"000000000",
  3093=>"000000000",
  3094=>"011111100",
  3095=>"111011001",
  3096=>"100001111",
  3097=>"111001000",
  3098=>"111111111",
  3099=>"000100100",
  3100=>"111111111",
  3101=>"110000001",
  3102=>"101100000",
  3103=>"000110000",
  3104=>"000000000",
  3105=>"111110110",
  3106=>"000000111",
  3107=>"111111111",
  3108=>"000000000",
  3109=>"110000000",
  3110=>"001001111",
  3111=>"000000000",
  3112=>"100100000",
  3113=>"000000000",
  3114=>"010100110",
  3115=>"111111111",
  3116=>"111011111",
  3117=>"111111111",
  3118=>"110100000",
  3119=>"111001000",
  3120=>"100100000",
  3121=>"010111010",
  3122=>"001111100",
  3123=>"000000101",
  3124=>"000110110",
  3125=>"000000000",
  3126=>"000000101",
  3127=>"111111000",
  3128=>"111000000",
  3129=>"011111111",
  3130=>"111111111",
  3131=>"000000000",
  3132=>"000111111",
  3133=>"001001000",
  3134=>"000000111",
  3135=>"111111011",
  3136=>"101001100",
  3137=>"000010111",
  3138=>"111000011",
  3139=>"111100111",
  3140=>"000010011",
  3141=>"001011011",
  3142=>"000000111",
  3143=>"111111111",
  3144=>"111111111",
  3145=>"000000111",
  3146=>"000000100",
  3147=>"000000000",
  3148=>"001000000",
  3149=>"000000111",
  3150=>"000000000",
  3151=>"000111011",
  3152=>"000000001",
  3153=>"111000000",
  3154=>"000000111",
  3155=>"000000001",
  3156=>"110110110",
  3157=>"000000110",
  3158=>"001000110",
  3159=>"110111111",
  3160=>"011111111",
  3161=>"000000101",
  3162=>"000000000",
  3163=>"100100100",
  3164=>"001011111",
  3165=>"001111011",
  3166=>"000000111",
  3167=>"000000000",
  3168=>"000000111",
  3169=>"010000000",
  3170=>"000000000",
  3171=>"111111111",
  3172=>"011000100",
  3173=>"111111111",
  3174=>"111111111",
  3175=>"110110000",
  3176=>"000000010",
  3177=>"111110111",
  3178=>"111111011",
  3179=>"100110011",
  3180=>"001001011",
  3181=>"000000000",
  3182=>"000000000",
  3183=>"100111111",
  3184=>"110100100",
  3185=>"000011111",
  3186=>"000000111",
  3187=>"111101111",
  3188=>"111111111",
  3189=>"111011000",
  3190=>"000000000",
  3191=>"111111111",
  3192=>"000000001",
  3193=>"111111111",
  3194=>"000000000",
  3195=>"111000001",
  3196=>"100000100",
  3197=>"000000000",
  3198=>"000110000",
  3199=>"000000111",
  3200=>"111111000",
  3201=>"000010111",
  3202=>"111000000",
  3203=>"000000000",
  3204=>"001000111",
  3205=>"111000001",
  3206=>"001001110",
  3207=>"000000001",
  3208=>"111111001",
  3209=>"000000000",
  3210=>"000000000",
  3211=>"111001001",
  3212=>"111111111",
  3213=>"111111010",
  3214=>"000000111",
  3215=>"111011111",
  3216=>"000000000",
  3217=>"000000100",
  3218=>"000000000",
  3219=>"000000000",
  3220=>"111111111",
  3221=>"111111111",
  3222=>"111011011",
  3223=>"000000000",
  3224=>"000001101",
  3225=>"111110111",
  3226=>"111111111",
  3227=>"000000000",
  3228=>"111110111",
  3229=>"100000000",
  3230=>"111011001",
  3231=>"001000100",
  3232=>"000000000",
  3233=>"111001001",
  3234=>"000000000",
  3235=>"000100111",
  3236=>"000000000",
  3237=>"111110111",
  3238=>"111111111",
  3239=>"000000001",
  3240=>"000000100",
  3241=>"101101101",
  3242=>"100000110",
  3243=>"111111111",
  3244=>"011111111",
  3245=>"110110111",
  3246=>"111111111",
  3247=>"101000000",
  3248=>"000000000",
  3249=>"111000000",
  3250=>"011111111",
  3251=>"111111100",
  3252=>"000000011",
  3253=>"000000000",
  3254=>"000111000",
  3255=>"111110010",
  3256=>"001111111",
  3257=>"111011111",
  3258=>"000000000",
  3259=>"001000000",
  3260=>"000000000",
  3261=>"000000000",
  3262=>"000000000",
  3263=>"000000000",
  3264=>"000000001",
  3265=>"001001111",
  3266=>"000000000",
  3267=>"100111111",
  3268=>"001000000",
  3269=>"000000000",
  3270=>"000000000",
  3271=>"000000000",
  3272=>"000000000",
  3273=>"111111101",
  3274=>"100100101",
  3275=>"000000000",
  3276=>"001101101",
  3277=>"000000010",
  3278=>"111111111",
  3279=>"011000000",
  3280=>"000000000",
  3281=>"000000000",
  3282=>"001111111",
  3283=>"000000100",
  3284=>"000000000",
  3285=>"111111001",
  3286=>"000000000",
  3287=>"111101111",
  3288=>"000000100",
  3289=>"111111110",
  3290=>"111000000",
  3291=>"000000000",
  3292=>"000000001",
  3293=>"000000101",
  3294=>"011111111",
  3295=>"110111111",
  3296=>"000000000",
  3297=>"000111111",
  3298=>"000010010",
  3299=>"111011111",
  3300=>"111111111",
  3301=>"011000000",
  3302=>"111111110",
  3303=>"111111100",
  3304=>"000000000",
  3305=>"011111011",
  3306=>"111111111",
  3307=>"111000000",
  3308=>"111111111",
  3309=>"000000000",
  3310=>"111100000",
  3311=>"001000111",
  3312=>"100101111",
  3313=>"111111111",
  3314=>"000111111",
  3315=>"000000001",
  3316=>"111111111",
  3317=>"000000001",
  3318=>"111111010",
  3319=>"001111111",
  3320=>"000000000",
  3321=>"110100000",
  3322=>"001000000",
  3323=>"000000000",
  3324=>"111110000",
  3325=>"111011001",
  3326=>"001000000",
  3327=>"111111000",
  3328=>"001000000",
  3329=>"000100111",
  3330=>"110000000",
  3331=>"100001001",
  3332=>"000100111",
  3333=>"000010110",
  3334=>"111000000",
  3335=>"110110111",
  3336=>"111011000",
  3337=>"010000000",
  3338=>"000000100",
  3339=>"001110100",
  3340=>"101000001",
  3341=>"111110100",
  3342=>"111111111",
  3343=>"111110110",
  3344=>"000000000",
  3345=>"111111111",
  3346=>"110010000",
  3347=>"000000000",
  3348=>"111111000",
  3349=>"111000000",
  3350=>"111001111",
  3351=>"111111000",
  3352=>"111111100",
  3353=>"000000000",
  3354=>"111111001",
  3355=>"111111000",
  3356=>"110100000",
  3357=>"000000000",
  3358=>"111111000",
  3359=>"111111111",
  3360=>"111110010",
  3361=>"001000000",
  3362=>"111111111",
  3363=>"111001000",
  3364=>"111000100",
  3365=>"001111111",
  3366=>"111111110",
  3367=>"011001111",
  3368=>"000000001",
  3369=>"011111100",
  3370=>"000000000",
  3371=>"000000111",
  3372=>"010010000",
  3373=>"111101000",
  3374=>"111111111",
  3375=>"000000001",
  3376=>"010001111",
  3377=>"111111111",
  3378=>"000000000",
  3379=>"000000000",
  3380=>"111111111",
  3381=>"000111111",
  3382=>"000000000",
  3383=>"101001111",
  3384=>"000000000",
  3385=>"000000000",
  3386=>"111110010",
  3387=>"001111111",
  3388=>"000000100",
  3389=>"111111011",
  3390=>"000000100",
  3391=>"111110111",
  3392=>"001000100",
  3393=>"111111000",
  3394=>"111101111",
  3395=>"000000000",
  3396=>"000000000",
  3397=>"000000000",
  3398=>"111111011",
  3399=>"000000001",
  3400=>"111111111",
  3401=>"001011111",
  3402=>"111000000",
  3403=>"000000000",
  3404=>"000001000",
  3405=>"000000100",
  3406=>"001000100",
  3407=>"110111111",
  3408=>"001000000",
  3409=>"000100110",
  3410=>"001001011",
  3411=>"000000111",
  3412=>"111000000",
  3413=>"011011011",
  3414=>"111111111",
  3415=>"111101101",
  3416=>"101111111",
  3417=>"110110111",
  3418=>"101001101",
  3419=>"111111111",
  3420=>"000111111",
  3421=>"111111111",
  3422=>"000000000",
  3423=>"111111011",
  3424=>"110111110",
  3425=>"101101110",
  3426=>"011011011",
  3427=>"111000000",
  3428=>"000000110",
  3429=>"000000000",
  3430=>"000000000",
  3431=>"001001111",
  3432=>"101000001",
  3433=>"000000000",
  3434=>"100000000",
  3435=>"111001001",
  3436=>"110001001",
  3437=>"001111101",
  3438=>"110000000",
  3439=>"111010110",
  3440=>"000000111",
  3441=>"000011111",
  3442=>"000000000",
  3443=>"000000000",
  3444=>"111111100",
  3445=>"111111111",
  3446=>"010000000",
  3447=>"011111111",
  3448=>"111000001",
  3449=>"110110001",
  3450=>"000111110",
  3451=>"000000001",
  3452=>"111111000",
  3453=>"111111110",
  3454=>"101000000",
  3455=>"111001001",
  3456=>"111011000",
  3457=>"000000111",
  3458=>"110110010",
  3459=>"000001111",
  3460=>"000000111",
  3461=>"010010000",
  3462=>"000000000",
  3463=>"111111111",
  3464=>"000001111",
  3465=>"111111111",
  3466=>"101100101",
  3467=>"000000000",
  3468=>"101001111",
  3469=>"101100000",
  3470=>"111110000",
  3471=>"010011111",
  3472=>"000100111",
  3473=>"000010000",
  3474=>"000000000",
  3475=>"010000000",
  3476=>"111111000",
  3477=>"000010010",
  3478=>"111001001",
  3479=>"111111001",
  3480=>"111000000",
  3481=>"011111101",
  3482=>"110000000",
  3483=>"000000100",
  3484=>"111111001",
  3485=>"000000000",
  3486=>"110111100",
  3487=>"000000111",
  3488=>"111111010",
  3489=>"000000011",
  3490=>"111111111",
  3491=>"001010010",
  3492=>"011111111",
  3493=>"111111111",
  3494=>"000000111",
  3495=>"000110111",
  3496=>"100100101",
  3497=>"000111111",
  3498=>"111110111",
  3499=>"001000000",
  3500=>"000000110",
  3501=>"111001000",
  3502=>"000000111",
  3503=>"111111111",
  3504=>"011011111",
  3505=>"000000000",
  3506=>"111010000",
  3507=>"111111111",
  3508=>"011011000",
  3509=>"000000000",
  3510=>"111111111",
  3511=>"001001111",
  3512=>"111111111",
  3513=>"011011111",
  3514=>"111111001",
  3515=>"111111001",
  3516=>"000000000",
  3517=>"000000000",
  3518=>"000000000",
  3519=>"000000000",
  3520=>"111111000",
  3521=>"111000110",
  3522=>"000000111",
  3523=>"000000100",
  3524=>"111000111",
  3525=>"011011111",
  3526=>"001001111",
  3527=>"110000000",
  3528=>"000000000",
  3529=>"000000110",
  3530=>"000000000",
  3531=>"000000000",
  3532=>"111000000",
  3533=>"000000101",
  3534=>"000111101",
  3535=>"000010110",
  3536=>"001000110",
  3537=>"001111000",
  3538=>"111100110",
  3539=>"000000000",
  3540=>"001000100",
  3541=>"111111110",
  3542=>"111000111",
  3543=>"000000010",
  3544=>"000000100",
  3545=>"100110000",
  3546=>"000000111",
  3547=>"000000000",
  3548=>"110100111",
  3549=>"111111111",
  3550=>"001000111",
  3551=>"000110111",
  3552=>"011111111",
  3553=>"011101101",
  3554=>"000011011",
  3555=>"111111001",
  3556=>"000000000",
  3557=>"000000000",
  3558=>"111011000",
  3559=>"001000000",
  3560=>"000000111",
  3561=>"111111111",
  3562=>"100000011",
  3563=>"111111111",
  3564=>"000000000",
  3565=>"111111101",
  3566=>"000001001",
  3567=>"000001001",
  3568=>"000000000",
  3569=>"000000000",
  3570=>"111111000",
  3571=>"000000111",
  3572=>"000111100",
  3573=>"000000000",
  3574=>"000000000",
  3575=>"000011111",
  3576=>"010011001",
  3577=>"001000000",
  3578=>"000110111",
  3579=>"110010111",
  3580=>"111111100",
  3581=>"000000001",
  3582=>"011111100",
  3583=>"100000000",
  3584=>"000100000",
  3585=>"000000000",
  3586=>"000000100",
  3587=>"000000010",
  3588=>"000000000",
  3589=>"011011001",
  3590=>"000000011",
  3591=>"111111111",
  3592=>"000010111",
  3593=>"111110111",
  3594=>"000111111",
  3595=>"000001000",
  3596=>"000100100",
  3597=>"110111111",
  3598=>"111111011",
  3599=>"000000000",
  3600=>"111111111",
  3601=>"110011011",
  3602=>"111011000",
  3603=>"011000111",
  3604=>"000010000",
  3605=>"101101111",
  3606=>"000000000",
  3607=>"100000000",
  3608=>"000001111",
  3609=>"111000100",
  3610=>"100101001",
  3611=>"111001101",
  3612=>"001000111",
  3613=>"100000000",
  3614=>"010000000",
  3615=>"111111111",
  3616=>"111011000",
  3617=>"111011000",
  3618=>"100000010",
  3619=>"110110100",
  3620=>"000000000",
  3621=>"001000000",
  3622=>"010011111",
  3623=>"111111111",
  3624=>"110000100",
  3625=>"000000000",
  3626=>"000111111",
  3627=>"000100000",
  3628=>"111010000",
  3629=>"111111111",
  3630=>"110100000",
  3631=>"001001000",
  3632=>"111110110",
  3633=>"111111001",
  3634=>"001011010",
  3635=>"111111110",
  3636=>"000010000",
  3637=>"000001000",
  3638=>"000110111",
  3639=>"100110110",
  3640=>"000100000",
  3641=>"100000000",
  3642=>"000000001",
  3643=>"001101111",
  3644=>"001111111",
  3645=>"011111111",
  3646=>"000000000",
  3647=>"000000000",
  3648=>"000000000",
  3649=>"000000111",
  3650=>"001111111",
  3651=>"001111111",
  3652=>"000100100",
  3653=>"100100000",
  3654=>"111110100",
  3655=>"000000000",
  3656=>"110110100",
  3657=>"000000111",
  3658=>"000000110",
  3659=>"000100000",
  3660=>"011011011",
  3661=>"000000111",
  3662=>"111110110",
  3663=>"111111111",
  3664=>"000000000",
  3665=>"000000000",
  3666=>"000011001",
  3667=>"100100100",
  3668=>"000110110",
  3669=>"000000111",
  3670=>"011111000",
  3671=>"001000000",
  3672=>"111111111",
  3673=>"111000000",
  3674=>"000000000",
  3675=>"001000000",
  3676=>"011011100",
  3677=>"111001000",
  3678=>"011000000",
  3679=>"000000110",
  3680=>"000100100",
  3681=>"111101001",
  3682=>"011110110",
  3683=>"000000100",
  3684=>"000000000",
  3685=>"000100111",
  3686=>"000001111",
  3687=>"000111000",
  3688=>"111100100",
  3689=>"000101111",
  3690=>"111111000",
  3691=>"000000000",
  3692=>"110111011",
  3693=>"000100111",
  3694=>"111111111",
  3695=>"100000000",
  3696=>"111111111",
  3697=>"101100000",
  3698=>"111111111",
  3699=>"111111100",
  3700=>"001011011",
  3701=>"000101101",
  3702=>"000000000",
  3703=>"000100100",
  3704=>"110000000",
  3705=>"000001111",
  3706=>"111011010",
  3707=>"001000000",
  3708=>"000001000",
  3709=>"011001000",
  3710=>"000111000",
  3711=>"000001000",
  3712=>"000010110",
  3713=>"011111111",
  3714=>"100110111",
  3715=>"000011000",
  3716=>"011111111",
  3717=>"000000100",
  3718=>"000011011",
  3719=>"111111111",
  3720=>"010111111",
  3721=>"000000000",
  3722=>"011111111",
  3723=>"110111111",
  3724=>"000000000",
  3725=>"000000000",
  3726=>"011000000",
  3727=>"011011011",
  3728=>"000000111",
  3729=>"000000000",
  3730=>"000110000",
  3731=>"110000000",
  3732=>"111111111",
  3733=>"111111111",
  3734=>"111111100",
  3735=>"001000000",
  3736=>"000011111",
  3737=>"111111001",
  3738=>"111111111",
  3739=>"111111100",
  3740=>"111111111",
  3741=>"000000000",
  3742=>"011001001",
  3743=>"000001111",
  3744=>"100100100",
  3745=>"110100100",
  3746=>"000000111",
  3747=>"000000111",
  3748=>"110000000",
  3749=>"111101011",
  3750=>"111111111",
  3751=>"100100000",
  3752=>"111111111",
  3753=>"111111100",
  3754=>"000100011",
  3755=>"111111111",
  3756=>"111111111",
  3757=>"110110110",
  3758=>"111111100",
  3759=>"110100100",
  3760=>"000111001",
  3761=>"000010011",
  3762=>"011111111",
  3763=>"111111111",
  3764=>"111111111",
  3765=>"111110000",
  3766=>"000000000",
  3767=>"100100001",
  3768=>"000000000",
  3769=>"111111111",
  3770=>"111111111",
  3771=>"111111111",
  3772=>"111111000",
  3773=>"011011111",
  3774=>"111111111",
  3775=>"111011000",
  3776=>"111110100",
  3777=>"110111101",
  3778=>"111111111",
  3779=>"000000000",
  3780=>"111111100",
  3781=>"000000000",
  3782=>"111111101",
  3783=>"010001000",
  3784=>"110001000",
  3785=>"001000110",
  3786=>"010110010",
  3787=>"011001111",
  3788=>"001100101",
  3789=>"111111001",
  3790=>"000001011",
  3791=>"001000110",
  3792=>"010011001",
  3793=>"111111111",
  3794=>"000011011",
  3795=>"111111111",
  3796=>"001001111",
  3797=>"011001011",
  3798=>"111111111",
  3799=>"111000100",
  3800=>"001001000",
  3801=>"100100111",
  3802=>"000000000",
  3803=>"000011111",
  3804=>"111111000",
  3805=>"001100000",
  3806=>"001001011",
  3807=>"011000001",
  3808=>"000000000",
  3809=>"111100000",
  3810=>"110111111",
  3811=>"000110110",
  3812=>"001111111",
  3813=>"100100110",
  3814=>"000000000",
  3815=>"011111000",
  3816=>"111111111",
  3817=>"000001101",
  3818=>"001000100",
  3819=>"000000101",
  3820=>"010000000",
  3821=>"000000000",
  3822=>"111111111",
  3823=>"111000001",
  3824=>"111110101",
  3825=>"111110000",
  3826=>"000011111",
  3827=>"000000000",
  3828=>"111111000",
  3829=>"000000110",
  3830=>"011011000",
  3831=>"000000000",
  3832=>"110000000",
  3833=>"111001000",
  3834=>"000110111",
  3835=>"000010010",
  3836=>"101100000",
  3837=>"111101111",
  3838=>"001111101",
  3839=>"000100100",
  3840=>"000000000",
  3841=>"011010000",
  3842=>"000011011",
  3843=>"111111111",
  3844=>"110111111",
  3845=>"010111111",
  3846=>"000000000",
  3847=>"011111111",
  3848=>"000111110",
  3849=>"000000000",
  3850=>"110100000",
  3851=>"011011111",
  3852=>"001001010",
  3853=>"111111111",
  3854=>"110101000",
  3855=>"011110000",
  3856=>"000000000",
  3857=>"000111111",
  3858=>"111111111",
  3859=>"000010000",
  3860=>"010111111",
  3861=>"110001111",
  3862=>"010000000",
  3863=>"000000000",
  3864=>"111101101",
  3865=>"000111000",
  3866=>"100000111",
  3867=>"101001001",
  3868=>"110010011",
  3869=>"000000000",
  3870=>"001111111",
  3871=>"011111000",
  3872=>"000110011",
  3873=>"000000000",
  3874=>"000000001",
  3875=>"000000000",
  3876=>"110010111",
  3877=>"111111111",
  3878=>"000111000",
  3879=>"111101110",
  3880=>"000000100",
  3881=>"111000000",
  3882=>"000100110",
  3883=>"011110111",
  3884=>"111111000",
  3885=>"011000000",
  3886=>"000000111",
  3887=>"000000000",
  3888=>"011001000",
  3889=>"111111111",
  3890=>"101000001",
  3891=>"000000000",
  3892=>"110100000",
  3893=>"111010000",
  3894=>"110111011",
  3895=>"000000100",
  3896=>"110111111",
  3897=>"011001111",
  3898=>"111111111",
  3899=>"000110110",
  3900=>"000000000",
  3901=>"000001001",
  3902=>"111111111",
  3903=>"111000000",
  3904=>"010000000",
  3905=>"000011011",
  3906=>"110111110",
  3907=>"111010000",
  3908=>"000000110",
  3909=>"111111111",
  3910=>"111111000",
  3911=>"011000111",
  3912=>"110110010",
  3913=>"111111111",
  3914=>"111111111",
  3915=>"100000111",
  3916=>"001111111",
  3917=>"111111001",
  3918=>"011111111",
  3919=>"000011001",
  3920=>"000110110",
  3921=>"111111111",
  3922=>"110000000",
  3923=>"000000001",
  3924=>"101001000",
  3925=>"111111001",
  3926=>"111111110",
  3927=>"110100101",
  3928=>"111011111",
  3929=>"111000000",
  3930=>"111111111",
  3931=>"001001111",
  3932=>"111101101",
  3933=>"000000100",
  3934=>"111101100",
  3935=>"000000000",
  3936=>"111111111",
  3937=>"000000000",
  3938=>"100000011",
  3939=>"000010111",
  3940=>"110110100",
  3941=>"000100000",
  3942=>"011011000",
  3943=>"111111111",
  3944=>"101111111",
  3945=>"000000000",
  3946=>"111111000",
  3947=>"110110100",
  3948=>"000000000",
  3949=>"000000000",
  3950=>"111101111",
  3951=>"010000000",
  3952=>"001001000",
  3953=>"111111000",
  3954=>"111111111",
  3955=>"011000000",
  3956=>"101101111",
  3957=>"110100100",
  3958=>"100111111",
  3959=>"000011010",
  3960=>"111111000",
  3961=>"111001111",
  3962=>"111111111",
  3963=>"011110110",
  3964=>"111111111",
  3965=>"111111111",
  3966=>"111111111",
  3967=>"111111111",
  3968=>"100100100",
  3969=>"101101111",
  3970=>"000000000",
  3971=>"000000000",
  3972=>"111110101",
  3973=>"111111111",
  3974=>"001100100",
  3975=>"111111111",
  3976=>"100101101",
  3977=>"110011011",
  3978=>"111001001",
  3979=>"110111111",
  3980=>"111111111",
  3981=>"000110110",
  3982=>"110110110",
  3983=>"111111111",
  3984=>"000001001",
  3985=>"110000000",
  3986=>"110110100",
  3987=>"000000000",
  3988=>"000000000",
  3989=>"000011000",
  3990=>"111111111",
  3991=>"000000010",
  3992=>"011111111",
  3993=>"111111111",
  3994=>"000001111",
  3995=>"100110000",
  3996=>"011111010",
  3997=>"101111111",
  3998=>"000001000",
  3999=>"110110111",
  4000=>"110110000",
  4001=>"111111111",
  4002=>"010001111",
  4003=>"000000011",
  4004=>"100100111",
  4005=>"000000000",
  4006=>"001001111",
  4007=>"111101111",
  4008=>"111111011",
  4009=>"110110100",
  4010=>"000000000",
  4011=>"000000000",
  4012=>"000000000",
  4013=>"100000100",
  4014=>"000000110",
  4015=>"111111111",
  4016=>"011000101",
  4017=>"000000000",
  4018=>"001011011",
  4019=>"000111111",
  4020=>"000000111",
  4021=>"110110111",
  4022=>"000000011",
  4023=>"111111111",
  4024=>"000000000",
  4025=>"000000000",
  4026=>"111001111",
  4027=>"110110111",
  4028=>"100111110",
  4029=>"111111111",
  4030=>"011110110",
  4031=>"001001001",
  4032=>"101101000",
  4033=>"001001011",
  4034=>"000011111",
  4035=>"000000000",
  4036=>"000000111",
  4037=>"111011011",
  4038=>"100101111",
  4039=>"000010000",
  4040=>"000000000",
  4041=>"011011111",
  4042=>"000101111",
  4043=>"000000000",
  4044=>"111111111",
  4045=>"000000000",
  4046=>"000101101",
  4047=>"110001001",
  4048=>"000000011",
  4049=>"111111111",
  4050=>"100111111",
  4051=>"000000000",
  4052=>"000000000",
  4053=>"111100111",
  4054=>"111011011",
  4055=>"000111111",
  4056=>"000001001",
  4057=>"011011111",
  4058=>"111111111",
  4059=>"111111111",
  4060=>"110110000",
  4061=>"000000000",
  4062=>"010011111",
  4063=>"000000000",
  4064=>"101110100",
  4065=>"111111111",
  4066=>"101110101",
  4067=>"010000000",
  4068=>"000000000",
  4069=>"000011110",
  4070=>"100101111",
  4071=>"000000000",
  4072=>"011100100",
  4073=>"000000000",
  4074=>"000011011",
  4075=>"000000001",
  4076=>"000000000",
  4077=>"001111111",
  4078=>"001011000",
  4079=>"000100111",
  4080=>"111111111",
  4081=>"111000000",
  4082=>"011111111",
  4083=>"000000000",
  4084=>"011011111",
  4085=>"000100111",
  4086=>"111111111",
  4087=>"111100110",
  4088=>"111111101",
  4089=>"000111111",
  4090=>"111110000",
  4091=>"000101101",
  4092=>"000000000",
  4093=>"111111110",
  4094=>"000001111",
  4095=>"011111111",
  4096=>"000000000",
  4097=>"000000000",
  4098=>"000000000",
  4099=>"011111111",
  4100=>"111111111",
  4101=>"111001011",
  4102=>"111000000",
  4103=>"111101111",
  4104=>"000000011",
  4105=>"111011111",
  4106=>"111111111",
  4107=>"000000111",
  4108=>"000000000",
  4109=>"111101111",
  4110=>"111011011",
  4111=>"111111110",
  4112=>"111111111",
  4113=>"111110110",
  4114=>"101000100",
  4115=>"010100110",
  4116=>"000000000",
  4117=>"110011011",
  4118=>"111111001",
  4119=>"011011001",
  4120=>"010000100",
  4121=>"110110100",
  4122=>"000001010",
  4123=>"100001001",
  4124=>"111111111",
  4125=>"111111011",
  4126=>"110110100",
  4127=>"111111111",
  4128=>"000000000",
  4129=>"111111111",
  4130=>"110000000",
  4131=>"111111111",
  4132=>"011111111",
  4133=>"100000000",
  4134=>"001001101",
  4135=>"000110110",
  4136=>"111000000",
  4137=>"000111111",
  4138=>"111111111",
  4139=>"111111111",
  4140=>"111110111",
  4141=>"111111010",
  4142=>"000000011",
  4143=>"111111000",
  4144=>"001111111",
  4145=>"111011111",
  4146=>"001000001",
  4147=>"011011001",
  4148=>"101001101",
  4149=>"011011011",
  4150=>"111110111",
  4151=>"101111111",
  4152=>"000000000",
  4153=>"000000100",
  4154=>"111111111",
  4155=>"001001001",
  4156=>"000001111",
  4157=>"111001111",
  4158=>"111111010",
  4159=>"000000000",
  4160=>"111101111",
  4161=>"100111100",
  4162=>"111111111",
  4163=>"000000111",
  4164=>"111000000",
  4165=>"001001011",
  4166=>"110110000",
  4167=>"111111111",
  4168=>"111101101",
  4169=>"111100000",
  4170=>"110111110",
  4171=>"000001111",
  4172=>"111111111",
  4173=>"111000000",
  4174=>"000001000",
  4175=>"110110110",
  4176=>"000000000",
  4177=>"000000000",
  4178=>"000000000",
  4179=>"111000011",
  4180=>"011000000",
  4181=>"000110111",
  4182=>"110000000",
  4183=>"011011000",
  4184=>"010011001",
  4185=>"000000000",
  4186=>"111110100",
  4187=>"000110000",
  4188=>"000000000",
  4189=>"000000000",
  4190=>"010000000",
  4191=>"000111111",
  4192=>"000111111",
  4193=>"111111111",
  4194=>"111111111",
  4195=>"100000000",
  4196=>"000000110",
  4197=>"101111111",
  4198=>"000010011",
  4199=>"111111000",
  4200=>"000000000",
  4201=>"000000000",
  4202=>"110101111",
  4203=>"000000010",
  4204=>"111001100",
  4205=>"100001000",
  4206=>"111111111",
  4207=>"100000000",
  4208=>"000000100",
  4209=>"100100111",
  4210=>"111100110",
  4211=>"111110111",
  4212=>"111000000",
  4213=>"100000110",
  4214=>"111111000",
  4215=>"001000011",
  4216=>"000001011",
  4217=>"000100100",
  4218=>"000000000",
  4219=>"000000001",
  4220=>"011011001",
  4221=>"000000000",
  4222=>"110101000",
  4223=>"111111111",
  4224=>"000000000",
  4225=>"111111111",
  4226=>"101100011",
  4227=>"000100100",
  4228=>"000001000",
  4229=>"111111110",
  4230=>"000000001",
  4231=>"111111011",
  4232=>"111111111",
  4233=>"000000000",
  4234=>"000000000",
  4235=>"111111111",
  4236=>"111111111",
  4237=>"000000000",
  4238=>"011001000",
  4239=>"000000000",
  4240=>"101111000",
  4241=>"000100100",
  4242=>"111111111",
  4243=>"110110100",
  4244=>"001101000",
  4245=>"111001011",
  4246=>"000000000",
  4247=>"000000000",
  4248=>"000010000",
  4249=>"000000000",
  4250=>"111110111",
  4251=>"111111111",
  4252=>"010011001",
  4253=>"001001100",
  4254=>"000110110",
  4255=>"111111011",
  4256=>"111000100",
  4257=>"111011011",
  4258=>"110001000",
  4259=>"001000000",
  4260=>"001000100",
  4261=>"100101011",
  4262=>"000000101",
  4263=>"110110111",
  4264=>"000000000",
  4265=>"101111111",
  4266=>"000000000",
  4267=>"000000001",
  4268=>"111111111",
  4269=>"111111011",
  4270=>"000000001",
  4271=>"101100000",
  4272=>"000010000",
  4273=>"001000000",
  4274=>"111111111",
  4275=>"000000000",
  4276=>"011011101",
  4277=>"011011111",
  4278=>"111111111",
  4279=>"000000111",
  4280=>"111011011",
  4281=>"000011011",
  4282=>"100110000",
  4283=>"100100010",
  4284=>"000000000",
  4285=>"000110000",
  4286=>"000000000",
  4287=>"111111111",
  4288=>"100000000",
  4289=>"111000000",
  4290=>"111011111",
  4291=>"001000001",
  4292=>"000000000",
  4293=>"000000000",
  4294=>"000111111",
  4295=>"110100111",
  4296=>"000000001",
  4297=>"011010000",
  4298=>"000000000",
  4299=>"111100100",
  4300=>"111011000",
  4301=>"111111000",
  4302=>"011011111",
  4303=>"110110110",
  4304=>"011011111",
  4305=>"110000000",
  4306=>"000000000",
  4307=>"000000100",
  4308=>"001000000",
  4309=>"000001001",
  4310=>"000000000",
  4311=>"000000110",
  4312=>"111111111",
  4313=>"100111111",
  4314=>"000000000",
  4315=>"000000000",
  4316=>"000000000",
  4317=>"111111111",
  4318=>"111011011",
  4319=>"000010000",
  4320=>"000000000",
  4321=>"000010000",
  4322=>"000110000",
  4323=>"011010000",
  4324=>"111101100",
  4325=>"001001001",
  4326=>"111111111",
  4327=>"111011011",
  4328=>"001011011",
  4329=>"101101001",
  4330=>"111010011",
  4331=>"000000000",
  4332=>"011011011",
  4333=>"111111111",
  4334=>"000000111",
  4335=>"111111010",
  4336=>"000000111",
  4337=>"100000000",
  4338=>"100000000",
  4339=>"111111001",
  4340=>"000000000",
  4341=>"100000000",
  4342=>"011001001",
  4343=>"000000001",
  4344=>"000000000",
  4345=>"111110000",
  4346=>"111001000",
  4347=>"011111001",
  4348=>"101000000",
  4349=>"110111111",
  4350=>"110001000",
  4351=>"111101111",
  4352=>"010010011",
  4353=>"000001000",
  4354=>"110100100",
  4355=>"000000111",
  4356=>"000000000",
  4357=>"001001101",
  4358=>"000011111",
  4359=>"111111111",
  4360=>"001000100",
  4361=>"000000000",
  4362=>"111110000",
  4363=>"111111000",
  4364=>"000000000",
  4365=>"111000000",
  4366=>"010011100",
  4367=>"111111111",
  4368=>"110000000",
  4369=>"111011000",
  4370=>"111111111",
  4371=>"011000000",
  4372=>"111111111",
  4373=>"000000000",
  4374=>"000000000",
  4375=>"011111010",
  4376=>"111101111",
  4377=>"000110000",
  4378=>"101100000",
  4379=>"101001001",
  4380=>"000000000",
  4381=>"000000001",
  4382=>"000000000",
  4383=>"001000001",
  4384=>"110111111",
  4385=>"011010010",
  4386=>"000000001",
  4387=>"100000000",
  4388=>"100000100",
  4389=>"100000000",
  4390=>"001001000",
  4391=>"101011001",
  4392=>"100111111",
  4393=>"111111110",
  4394=>"111111111",
  4395=>"011111111",
  4396=>"001011110",
  4397=>"111001000",
  4398=>"000000000",
  4399=>"000000011",
  4400=>"111000000",
  4401=>"111111111",
  4402=>"111100000",
  4403=>"001001001",
  4404=>"000000000",
  4405=>"000000111",
  4406=>"100000001",
  4407=>"110111111",
  4408=>"000000000",
  4409=>"001011011",
  4410=>"111001000",
  4411=>"000000000",
  4412=>"100000111",
  4413=>"000000010",
  4414=>"001000000",
  4415=>"111111110",
  4416=>"000000111",
  4417=>"001000000",
  4418=>"000001000",
  4419=>"111111111",
  4420=>"111111111",
  4421=>"000000000",
  4422=>"011011000",
  4423=>"001101100",
  4424=>"000111111",
  4425=>"100000000",
  4426=>"000000000",
  4427=>"110100100",
  4428=>"010000001",
  4429=>"100101000",
  4430=>"110110010",
  4431=>"001000000",
  4432=>"111001001",
  4433=>"100111111",
  4434=>"000000001",
  4435=>"011000000",
  4436=>"000000000",
  4437=>"001001011",
  4438=>"001111011",
  4439=>"111110111",
  4440=>"111111111",
  4441=>"111111111",
  4442=>"111111111",
  4443=>"010010110",
  4444=>"011011101",
  4445=>"000000000",
  4446=>"000000000",
  4447=>"111110000",
  4448=>"000100111",
  4449=>"111111111",
  4450=>"001011011",
  4451=>"000000000",
  4452=>"111111111",
  4453=>"000000111",
  4454=>"111111011",
  4455=>"111011011",
  4456=>"000000111",
  4457=>"111111000",
  4458=>"000000000",
  4459=>"011000000",
  4460=>"110111001",
  4461=>"001000000",
  4462=>"111111111",
  4463=>"000000001",
  4464=>"111111111",
  4465=>"000000001",
  4466=>"101111111",
  4467=>"011001000",
  4468=>"111111100",
  4469=>"111001000",
  4470=>"011111011",
  4471=>"111111111",
  4472=>"010111111",
  4473=>"000000000",
  4474=>"111111111",
  4475=>"000000000",
  4476=>"110111100",
  4477=>"111111110",
  4478=>"100111111",
  4479=>"000000000",
  4480=>"000000000",
  4481=>"111111110",
  4482=>"000000111",
  4483=>"110111111",
  4484=>"010000000",
  4485=>"111111010",
  4486=>"100001000",
  4487=>"000001001",
  4488=>"100100111",
  4489=>"110111111",
  4490=>"111011010",
  4491=>"100001001",
  4492=>"101101001",
  4493=>"110110110",
  4494=>"000000000",
  4495=>"111111111",
  4496=>"000000000",
  4497=>"000000000",
  4498=>"000010011",
  4499=>"000000011",
  4500=>"001011111",
  4501=>"010000011",
  4502=>"011110110",
  4503=>"000000001",
  4504=>"110110111",
  4505=>"110110110",
  4506=>"111111111",
  4507=>"111111111",
  4508=>"111111110",
  4509=>"111111111",
  4510=>"100101000",
  4511=>"011111010",
  4512=>"000000000",
  4513=>"010110110",
  4514=>"111000001",
  4515=>"010111011",
  4516=>"000010000",
  4517=>"000000000",
  4518=>"000000000",
  4519=>"000000000",
  4520=>"111111001",
  4521=>"000000000",
  4522=>"000110010",
  4523=>"000101101",
  4524=>"000111100",
  4525=>"111111111",
  4526=>"000111111",
  4527=>"010011001",
  4528=>"101101000",
  4529=>"000000111",
  4530=>"111000000",
  4531=>"111110110",
  4532=>"011000000",
  4533=>"000000001",
  4534=>"011000000",
  4535=>"000000000",
  4536=>"001001001",
  4537=>"001111111",
  4538=>"001000000",
  4539=>"101101111",
  4540=>"000111111",
  4541=>"000000000",
  4542=>"011000000",
  4543=>"010010010",
  4544=>"000000001",
  4545=>"000000000",
  4546=>"000000011",
  4547=>"111111111",
  4548=>"010000000",
  4549=>"001011111",
  4550=>"000001010",
  4551=>"000000000",
  4552=>"011011011",
  4553=>"000000110",
  4554=>"100111100",
  4555=>"000000001",
  4556=>"111111111",
  4557=>"010000000",
  4558=>"110010111",
  4559=>"111100110",
  4560=>"011100101",
  4561=>"101101001",
  4562=>"000000000",
  4563=>"100100000",
  4564=>"111111111",
  4565=>"111100100",
  4566=>"011111011",
  4567=>"111001001",
  4568=>"000000000",
  4569=>"111100000",
  4570=>"110010010",
  4571=>"100100100",
  4572=>"110001011",
  4573=>"100001100",
  4574=>"000000000",
  4575=>"000000111",
  4576=>"000000000",
  4577=>"011000000",
  4578=>"110110110",
  4579=>"000011101",
  4580=>"000000110",
  4581=>"001001001",
  4582=>"000100001",
  4583=>"000000000",
  4584=>"001001000",
  4585=>"011011111",
  4586=>"000000000",
  4587=>"111111111",
  4588=>"011001001",
  4589=>"111010010",
  4590=>"000000000",
  4591=>"000000000",
  4592=>"111111011",
  4593=>"111111001",
  4594=>"010000000",
  4595=>"011101101",
  4596=>"110110111",
  4597=>"000100111",
  4598=>"000000000",
  4599=>"110111100",
  4600=>"111111111",
  4601=>"001100110",
  4602=>"111000100",
  4603=>"000001000",
  4604=>"000000000",
  4605=>"000000100",
  4606=>"000000100",
  4607=>"000000000",
  4608=>"000000000",
  4609=>"000000000",
  4610=>"101111111",
  4611=>"001111111",
  4612=>"000000000",
  4613=>"010010000",
  4614=>"000100000",
  4615=>"111111111",
  4616=>"111111010",
  4617=>"000000111",
  4618=>"000111100",
  4619=>"000000100",
  4620=>"000000010",
  4621=>"011011111",
  4622=>"011001000",
  4623=>"000000000",
  4624=>"000000000",
  4625=>"000101111",
  4626=>"000000000",
  4627=>"100110111",
  4628=>"110111000",
  4629=>"000000000",
  4630=>"000000000",
  4631=>"111111100",
  4632=>"111111011",
  4633=>"000000000",
  4634=>"111000000",
  4635=>"011001000",
  4636=>"001111111",
  4637=>"111100111",
  4638=>"111111111",
  4639=>"111101101",
  4640=>"000000000",
  4641=>"111111111",
  4642=>"111111110",
  4643=>"111001001",
  4644=>"111111111",
  4645=>"000000000",
  4646=>"111100000",
  4647=>"000000000",
  4648=>"111011001",
  4649=>"111111111",
  4650=>"111000000",
  4651=>"000110100",
  4652=>"000111111",
  4653=>"001111111",
  4654=>"011011011",
  4655=>"111111111",
  4656=>"011111111",
  4657=>"000000000",
  4658=>"101101100",
  4659=>"110111111",
  4660=>"000000010",
  4661=>"000000010",
  4662=>"111111001",
  4663=>"000000111",
  4664=>"111111000",
  4665=>"000011000",
  4666=>"000000000",
  4667=>"000000110",
  4668=>"000000000",
  4669=>"000000111",
  4670=>"000000000",
  4671=>"111000000",
  4672=>"000010000",
  4673=>"000000100",
  4674=>"001011111",
  4675=>"110111010",
  4676=>"000001110",
  4677=>"100100000",
  4678=>"111111111",
  4679=>"111111111",
  4680=>"011000100",
  4681=>"111001111",
  4682=>"000010011",
  4683=>"000000000",
  4684=>"111111000",
  4685=>"110110110",
  4686=>"100100100",
  4687=>"000001000",
  4688=>"000000101",
  4689=>"000000000",
  4690=>"111111000",
  4691=>"000000000",
  4692=>"000111111",
  4693=>"000000100",
  4694=>"111111100",
  4695=>"000000000",
  4696=>"111100000",
  4697=>"111101111",
  4698=>"111111110",
  4699=>"011111000",
  4700=>"001000000",
  4701=>"111111111",
  4702=>"111111111",
  4703=>"000000000",
  4704=>"000000000",
  4705=>"111111111",
  4706=>"010000000",
  4707=>"001110111",
  4708=>"001111011",
  4709=>"000000101",
  4710=>"111111111",
  4711=>"000000000",
  4712=>"000000000",
  4713=>"111101111",
  4714=>"111111111",
  4715=>"000000100",
  4716=>"000000000",
  4717=>"000000000",
  4718=>"111111100",
  4719=>"000100101",
  4720=>"000010111",
  4721=>"000000000",
  4722=>"011011111",
  4723=>"111110100",
  4724=>"000000010",
  4725=>"111110111",
  4726=>"111111000",
  4727=>"000011101",
  4728=>"000000010",
  4729=>"110010000",
  4730=>"011011000",
  4731=>"111111111",
  4732=>"111111011",
  4733=>"000011111",
  4734=>"001000000",
  4735=>"000001000",
  4736=>"111111111",
  4737=>"011111000",
  4738=>"001000000",
  4739=>"000000000",
  4740=>"111110100",
  4741=>"111000000",
  4742=>"110000000",
  4743=>"011111111",
  4744=>"111111111",
  4745=>"000000000",
  4746=>"000000000",
  4747=>"000000000",
  4748=>"111101011",
  4749=>"111111111",
  4750=>"100000001",
  4751=>"000000000",
  4752=>"111111111",
  4753=>"000000000",
  4754=>"000000000",
  4755=>"111111110",
  4756=>"000100100",
  4757=>"011001111",
  4758=>"111111111",
  4759=>"111111010",
  4760=>"111111110",
  4761=>"000000111",
  4762=>"000000000",
  4763=>"000011111",
  4764=>"110110111",
  4765=>"000000000",
  4766=>"111111111",
  4767=>"000000000",
  4768=>"000000000",
  4769=>"111111111",
  4770=>"000000000",
  4771=>"111111111",
  4772=>"000100110",
  4773=>"100100000",
  4774=>"111111111",
  4775=>"111110111",
  4776=>"101000000",
  4777=>"111111111",
  4778=>"000000000",
  4779=>"001001101",
  4780=>"111101000",
  4781=>"001111111",
  4782=>"111111111",
  4783=>"110100111",
  4784=>"000000000",
  4785=>"000000000",
  4786=>"101101101",
  4787=>"111111110",
  4788=>"000000000",
  4789=>"000101001",
  4790=>"000000000",
  4791=>"100100000",
  4792=>"011000000",
  4793=>"000000000",
  4794=>"000000000",
  4795=>"001000000",
  4796=>"111101111",
  4797=>"100000000",
  4798=>"000100100",
  4799=>"000000000",
  4800=>"100100111",
  4801=>"111111111",
  4802=>"000110110",
  4803=>"111111000",
  4804=>"100100000",
  4805=>"111111101",
  4806=>"111111111",
  4807=>"010011000",
  4808=>"000000000",
  4809=>"110000000",
  4810=>"110010010",
  4811=>"000000000",
  4812=>"111111111",
  4813=>"000000111",
  4814=>"111111111",
  4815=>"011111111",
  4816=>"000000000",
  4817=>"111000000",
  4818=>"111111111",
  4819=>"000010111",
  4820=>"001000000",
  4821=>"111101001",
  4822=>"000000000",
  4823=>"100000000",
  4824=>"011111000",
  4825=>"111111000",
  4826=>"000000000",
  4827=>"000100111",
  4828=>"000101111",
  4829=>"111111111",
  4830=>"000000000",
  4831=>"110110111",
  4832=>"111111111",
  4833=>"000000000",
  4834=>"101000000",
  4835=>"111111100",
  4836=>"111010111",
  4837=>"100000000",
  4838=>"000000000",
  4839=>"111111100",
  4840=>"000000000",
  4841=>"000000011",
  4842=>"111111111",
  4843=>"111111011",
  4844=>"000110110",
  4845=>"000011011",
  4846=>"111111110",
  4847=>"001000100",
  4848=>"110100100",
  4849=>"111111111",
  4850=>"111111111",
  4851=>"000000001",
  4852=>"000000000",
  4853=>"100000000",
  4854=>"001000011",
  4855=>"000000000",
  4856=>"000111111",
  4857=>"100000000",
  4858=>"000000010",
  4859=>"010010000",
  4860=>"011011011",
  4861=>"111110110",
  4862=>"100000100",
  4863=>"000000000",
  4864=>"000111000",
  4865=>"101111111",
  4866=>"111111010",
  4867=>"000001101",
  4868=>"110100111",
  4869=>"111110110",
  4870=>"111111111",
  4871=>"111111111",
  4872=>"000000000",
  4873=>"101000111",
  4874=>"111100001",
  4875=>"000000000",
  4876=>"001001111",
  4877=>"000001101",
  4878=>"110110111",
  4879=>"111111111",
  4880=>"100111111",
  4881=>"011111111",
  4882=>"110010110",
  4883=>"000111101",
  4884=>"000000000",
  4885=>"100101111",
  4886=>"010010000",
  4887=>"010000000",
  4888=>"000100111",
  4889=>"000111111",
  4890=>"110011101",
  4891=>"110100000",
  4892=>"110110111",
  4893=>"000000010",
  4894=>"111111111",
  4895=>"010010110",
  4896=>"000011000",
  4897=>"111100000",
  4898=>"100111011",
  4899=>"011110010",
  4900=>"011011111",
  4901=>"010000111",
  4902=>"000000000",
  4903=>"000000000",
  4904=>"011110111",
  4905=>"000000000",
  4906=>"111100000",
  4907=>"000000000",
  4908=>"110000000",
  4909=>"111111011",
  4910=>"001000000",
  4911=>"000000000",
  4912=>"101100100",
  4913=>"000000111",
  4914=>"000000001",
  4915=>"111111111",
  4916=>"101000100",
  4917=>"000000000",
  4918=>"000000000",
  4919=>"100100000",
  4920=>"000000000",
  4921=>"010010111",
  4922=>"000000000",
  4923=>"100111111",
  4924=>"111111111",
  4925=>"111100111",
  4926=>"011011111",
  4927=>"000000000",
  4928=>"111100000",
  4929=>"111111111",
  4930=>"111100000",
  4931=>"000000000",
  4932=>"000000100",
  4933=>"000000111",
  4934=>"000010111",
  4935=>"000001000",
  4936=>"111111000",
  4937=>"011111111",
  4938=>"110000000",
  4939=>"111111000",
  4940=>"011010011",
  4941=>"111000000",
  4942=>"111111100",
  4943=>"101000000",
  4944=>"100000000",
  4945=>"001000000",
  4946=>"111110111",
  4947=>"000000101",
  4948=>"000000000",
  4949=>"011011011",
  4950=>"000000000",
  4951=>"111111100",
  4952=>"111111000",
  4953=>"000000000",
  4954=>"111010000",
  4955=>"111111111",
  4956=>"101101101",
  4957=>"010110011",
  4958=>"000000001",
  4959=>"000000110",
  4960=>"111111111",
  4961=>"111111111",
  4962=>"111100101",
  4963=>"111111111",
  4964=>"000000000",
  4965=>"000000001",
  4966=>"111111111",
  4967=>"111111000",
  4968=>"110111001",
  4969=>"100100000",
  4970=>"011111111",
  4971=>"000001011",
  4972=>"000000000",
  4973=>"111111111",
  4974=>"000000000",
  4975=>"111110111",
  4976=>"111111111",
  4977=>"111111111",
  4978=>"001101000",
  4979=>"001000000",
  4980=>"100000000",
  4981=>"111111111",
  4982=>"001000101",
  4983=>"100000000",
  4984=>"111111111",
  4985=>"001101101",
  4986=>"111101111",
  4987=>"011000000",
  4988=>"111110000",
  4989=>"111111111",
  4990=>"001011111",
  4991=>"111111111",
  4992=>"111001001",
  4993=>"100101001",
  4994=>"011011011",
  4995=>"111111011",
  4996=>"000000000",
  4997=>"000000000",
  4998=>"110011111",
  4999=>"111111111",
  5000=>"000001111",
  5001=>"111110000",
  5002=>"110000000",
  5003=>"100100110",
  5004=>"111111111",
  5005=>"000010000",
  5006=>"111111111",
  5007=>"111111000",
  5008=>"000000011",
  5009=>"001001111",
  5010=>"011101000",
  5011=>"111111111",
  5012=>"000100111",
  5013=>"000000000",
  5014=>"111111111",
  5015=>"000000000",
  5016=>"000000000",
  5017=>"111001111",
  5018=>"111111111",
  5019=>"011001001",
  5020=>"110110111",
  5021=>"111111111",
  5022=>"000000001",
  5023=>"000000100",
  5024=>"000000000",
  5025=>"000000110",
  5026=>"000101000",
  5027=>"111111101",
  5028=>"100100100",
  5029=>"010010010",
  5030=>"000000101",
  5031=>"110000000",
  5032=>"100000111",
  5033=>"000000000",
  5034=>"111111111",
  5035=>"111111111",
  5036=>"111000000",
  5037=>"111100111",
  5038=>"111111111",
  5039=>"000000100",
  5040=>"000100000",
  5041=>"110110111",
  5042=>"000000000",
  5043=>"000000000",
  5044=>"000000110",
  5045=>"111111111",
  5046=>"111111111",
  5047=>"111101000",
  5048=>"111111111",
  5049=>"101111111",
  5050=>"110010000",
  5051=>"101001111",
  5052=>"111111111",
  5053=>"110110100",
  5054=>"000000000",
  5055=>"001001001",
  5056=>"110110000",
  5057=>"111111010",
  5058=>"111111111",
  5059=>"111111000",
  5060=>"111111111",
  5061=>"001001101",
  5062=>"011111010",
  5063=>"000000111",
  5064=>"001000000",
  5065=>"100111110",
  5066=>"100100111",
  5067=>"111111111",
  5068=>"000000000",
  5069=>"100111111",
  5070=>"111111000",
  5071=>"111111111",
  5072=>"111101111",
  5073=>"100100100",
  5074=>"000000000",
  5075=>"111011000",
  5076=>"000000000",
  5077=>"111111100",
  5078=>"000000000",
  5079=>"011011111",
  5080=>"111110110",
  5081=>"100000111",
  5082=>"000000111",
  5083=>"111110010",
  5084=>"000011001",
  5085=>"110000000",
  5086=>"000000100",
  5087=>"001001001",
  5088=>"000000000",
  5089=>"000000001",
  5090=>"000000110",
  5091=>"010000111",
  5092=>"111111111",
  5093=>"000000110",
  5094=>"010010110",
  5095=>"000000000",
  5096=>"001001001",
  5097=>"000000000",
  5098=>"111111111",
  5099=>"111111101",
  5100=>"111111111",
  5101=>"000000000",
  5102=>"000000111",
  5103=>"110111111",
  5104=>"000000001",
  5105=>"111111111",
  5106=>"001011000",
  5107=>"000110000",
  5108=>"000000000",
  5109=>"111111111",
  5110=>"111111000",
  5111=>"111011000",
  5112=>"110110000",
  5113=>"111101101",
  5114=>"100110100",
  5115=>"011001100",
  5116=>"111111000",
  5117=>"010101011",
  5118=>"000000101",
  5119=>"000000000",
  5120=>"100011011",
  5121=>"111000000",
  5122=>"111111111",
  5123=>"000101001",
  5124=>"111111001",
  5125=>"111111111",
  5126=>"000010111",
  5127=>"111111111",
  5128=>"000000000",
  5129=>"111011011",
  5130=>"010110110",
  5131=>"011110110",
  5132=>"000010110",
  5133=>"000000100",
  5134=>"100100110",
  5135=>"111111111",
  5136=>"100000011",
  5137=>"101011111",
  5138=>"111011000",
  5139=>"111111111",
  5140=>"000001100",
  5141=>"011001000",
  5142=>"000000000",
  5143=>"011111011",
  5144=>"110110000",
  5145=>"110100101",
  5146=>"000000000",
  5147=>"110011100",
  5148=>"000000001",
  5149=>"111110100",
  5150=>"110000000",
  5151=>"000111111",
  5152=>"001111111",
  5153=>"100100000",
  5154=>"000000000",
  5155=>"111111001",
  5156=>"000010000",
  5157=>"000000000",
  5158=>"111100111",
  5159=>"000000000",
  5160=>"000010011",
  5161=>"000000010",
  5162=>"000000000",
  5163=>"111111100",
  5164=>"000000000",
  5165=>"000000110",
  5166=>"000000000",
  5167=>"111110111",
  5168=>"111111111",
  5169=>"111111111",
  5170=>"001001111",
  5171=>"111111111",
  5172=>"000000000",
  5173=>"110110111",
  5174=>"110100100",
  5175=>"010000111",
  5176=>"000001111",
  5177=>"111000011",
  5178=>"111111111",
  5179=>"011011111",
  5180=>"111001011",
  5181=>"111111111",
  5182=>"111101111",
  5183=>"000000000",
  5184=>"000111111",
  5185=>"110000010",
  5186=>"000110110",
  5187=>"110101001",
  5188=>"111011100",
  5189=>"100100101",
  5190=>"110111011",
  5191=>"000000001",
  5192=>"000000010",
  5193=>"111111111",
  5194=>"111111011",
  5195=>"111111111",
  5196=>"001011111",
  5197=>"110111111",
  5198=>"111111111",
  5199=>"001001001",
  5200=>"111110111",
  5201=>"111101001",
  5202=>"111111111",
  5203=>"111111111",
  5204=>"111111111",
  5205=>"100111111",
  5206=>"001000000",
  5207=>"111100100",
  5208=>"111111111",
  5209=>"000000100",
  5210=>"100111111",
  5211=>"000101001",
  5212=>"000000001",
  5213=>"111011001",
  5214=>"000001001",
  5215=>"100000111",
  5216=>"111111111",
  5217=>"111111000",
  5218=>"111110111",
  5219=>"111110111",
  5220=>"000000100",
  5221=>"011001001",
  5222=>"100000000",
  5223=>"110111101",
  5224=>"000000000",
  5225=>"010000000",
  5226=>"011000000",
  5227=>"000111111",
  5228=>"111011001",
  5229=>"111111000",
  5230=>"111111111",
  5231=>"110111111",
  5232=>"111111111",
  5233=>"100000000",
  5234=>"000000000",
  5235=>"110110000",
  5236=>"111110000",
  5237=>"000000000",
  5238=>"111000010",
  5239=>"000000000",
  5240=>"000000000",
  5241=>"110000000",
  5242=>"000010000",
  5243=>"111111100",
  5244=>"110100100",
  5245=>"111111110",
  5246=>"000010011",
  5247=>"111110100",
  5248=>"111111111",
  5249=>"111110111",
  5250=>"000000000",
  5251=>"111111111",
  5252=>"001000000",
  5253=>"111111111",
  5254=>"011011111",
  5255=>"011011111",
  5256=>"000001111",
  5257=>"000000000",
  5258=>"011010000",
  5259=>"000011011",
  5260=>"111111011",
  5261=>"000000000",
  5262=>"010000000",
  5263=>"111100110",
  5264=>"010110000",
  5265=>"001000000",
  5266=>"111111111",
  5267=>"100110111",
  5268=>"101000000",
  5269=>"000110111",
  5270=>"111111001",
  5271=>"111101000",
  5272=>"111110110",
  5273=>"011000000",
  5274=>"001000000",
  5275=>"111000111",
  5276=>"010000100",
  5277=>"010000000",
  5278=>"010000000",
  5279=>"111111111",
  5280=>"000100110",
  5281=>"011111111",
  5282=>"111111111",
  5283=>"111001101",
  5284=>"111111110",
  5285=>"011011111",
  5286=>"111110000",
  5287=>"101111101",
  5288=>"000000101",
  5289=>"001000110",
  5290=>"000111110",
  5291=>"111111110",
  5292=>"100111111",
  5293=>"110100100",
  5294=>"000010011",
  5295=>"111111111",
  5296=>"000000000",
  5297=>"100100001",
  5298=>"000000000",
  5299=>"011111111",
  5300=>"111111111",
  5301=>"111111111",
  5302=>"000100111",
  5303=>"000100000",
  5304=>"111111111",
  5305=>"111111111",
  5306=>"000000010",
  5307=>"000000001",
  5308=>"000111011",
  5309=>"111100111",
  5310=>"000000000",
  5311=>"011001001",
  5312=>"111111111",
  5313=>"111000000",
  5314=>"111011101",
  5315=>"000000000",
  5316=>"110110110",
  5317=>"000000000",
  5318=>"001000010",
  5319=>"111111111",
  5320=>"000000001",
  5321=>"000000000",
  5322=>"111111100",
  5323=>"111111111",
  5324=>"111011001",
  5325=>"001001000",
  5326=>"111111101",
  5327=>"000000000",
  5328=>"111111111",
  5329=>"100100111",
  5330=>"011110111",
  5331=>"111111111",
  5332=>"001000001",
  5333=>"000000000",
  5334=>"000000011",
  5335=>"110111111",
  5336=>"111111111",
  5337=>"011011111",
  5338=>"000000000",
  5339=>"011000000",
  5340=>"000000100",
  5341=>"100000000",
  5342=>"000000000",
  5343=>"010110100",
  5344=>"000000000",
  5345=>"000000111",
  5346=>"000000010",
  5347=>"110100110",
  5348=>"001111100",
  5349=>"011011111",
  5350=>"000000000",
  5351=>"111110100",
  5352=>"111111111",
  5353=>"000000000",
  5354=>"010000000",
  5355=>"000000001",
  5356=>"010000000",
  5357=>"100100000",
  5358=>"011111111",
  5359=>"000000000",
  5360=>"111011111",
  5361=>"010011111",
  5362=>"000000000",
  5363=>"000011000",
  5364=>"001011000",
  5365=>"010000110",
  5366=>"001011011",
  5367=>"000000000",
  5368=>"000000000",
  5369=>"001000000",
  5370=>"111111111",
  5371=>"111011111",
  5372=>"011010100",
  5373=>"001011110",
  5374=>"001100000",
  5375=>"110000000",
  5376=>"111110100",
  5377=>"100100111",
  5378=>"000111111",
  5379=>"110110101",
  5380=>"011011000",
  5381=>"000000000",
  5382=>"001001011",
  5383=>"110000111",
  5384=>"111110001",
  5385=>"000000111",
  5386=>"011001101",
  5387=>"000000000",
  5388=>"011011001",
  5389=>"011110000",
  5390=>"000000000",
  5391=>"000000111",
  5392=>"000000111",
  5393=>"011111111",
  5394=>"111111010",
  5395=>"011110110",
  5396=>"111111111",
  5397=>"000011000",
  5398=>"100100100",
  5399=>"110100111",
  5400=>"000000001",
  5401=>"000000000",
  5402=>"111111010",
  5403=>"000100111",
  5404=>"111111111",
  5405=>"110111011",
  5406=>"111111111",
  5407=>"101001001",
  5408=>"100000011",
  5409=>"111111111",
  5410=>"000000111",
  5411=>"000010111",
  5412=>"000000000",
  5413=>"101111110",
  5414=>"101001000",
  5415=>"111001000",
  5416=>"000000000",
  5417=>"111101100",
  5418=>"011111110",
  5419=>"101111111",
  5420=>"111000111",
  5421=>"100000000",
  5422=>"111111111",
  5423=>"101000111",
  5424=>"111111111",
  5425=>"110111110",
  5426=>"111111111",
  5427=>"111110000",
  5428=>"100000000",
  5429=>"011000100",
  5430=>"111111100",
  5431=>"001000110",
  5432=>"000000111",
  5433=>"111111111",
  5434=>"000000000",
  5435=>"101110111",
  5436=>"110110100",
  5437=>"110110000",
  5438=>"000111001",
  5439=>"111111111",
  5440=>"110011000",
  5441=>"111111111",
  5442=>"010000000",
  5443=>"111000000",
  5444=>"111111111",
  5445=>"111011001",
  5446=>"110111000",
  5447=>"000000000",
  5448=>"111111111",
  5449=>"000110111",
  5450=>"000000000",
  5451=>"010111101",
  5452=>"000000110",
  5453=>"111111011",
  5454=>"001000100",
  5455=>"000000001",
  5456=>"000000100",
  5457=>"001001000",
  5458=>"101111101",
  5459=>"000111000",
  5460=>"111111111",
  5461=>"011000011",
  5462=>"111111001",
  5463=>"000000000",
  5464=>"000000000",
  5465=>"001011011",
  5466=>"100110110",
  5467=>"011000001",
  5468=>"111111011",
  5469=>"111111111",
  5470=>"000000000",
  5471=>"100000000",
  5472=>"011111011",
  5473=>"000011000",
  5474=>"111001001",
  5475=>"111111111",
  5476=>"110000000",
  5477=>"100110000",
  5478=>"000100101",
  5479=>"011110110",
  5480=>"110110101",
  5481=>"111111111",
  5482=>"111111111",
  5483=>"000000000",
  5484=>"010011001",
  5485=>"000000000",
  5486=>"000010111",
  5487=>"111101111",
  5488=>"000000100",
  5489=>"111111111",
  5490=>"011011000",
  5491=>"011001000",
  5492=>"000000000",
  5493=>"011000100",
  5494=>"000000101",
  5495=>"110101101",
  5496=>"000000000",
  5497=>"111111111",
  5498=>"111111010",
  5499=>"011111111",
  5500=>"000011011",
  5501=>"010000000",
  5502=>"111111111",
  5503=>"000000111",
  5504=>"111110100",
  5505=>"011001111",
  5506=>"111111111",
  5507=>"000000000",
  5508=>"010000111",
  5509=>"111111111",
  5510=>"000010011",
  5511=>"101101101",
  5512=>"010000000",
  5513=>"010000000",
  5514=>"111011001",
  5515=>"110111111",
  5516=>"111000100",
  5517=>"111101001",
  5518=>"000000000",
  5519=>"010010011",
  5520=>"000010010",
  5521=>"000001001",
  5522=>"111111111",
  5523=>"011111111",
  5524=>"011001000",
  5525=>"000001001",
  5526=>"111110100",
  5527=>"110110111",
  5528=>"100001111",
  5529=>"000000011",
  5530=>"101011111",
  5531=>"000100111",
  5532=>"000000011",
  5533=>"000001111",
  5534=>"000000000",
  5535=>"111111111",
  5536=>"000111111",
  5537=>"111001100",
  5538=>"111000001",
  5539=>"000001111",
  5540=>"111111000",
  5541=>"101101111",
  5542=>"111111111",
  5543=>"110110110",
  5544=>"001001001",
  5545=>"111110110",
  5546=>"111111110",
  5547=>"000000001",
  5548=>"111111111",
  5549=>"000001001",
  5550=>"000000000",
  5551=>"000001111",
  5552=>"111011011",
  5553=>"010000000",
  5554=>"000000000",
  5555=>"011010110",
  5556=>"111111111",
  5557=>"111001000",
  5558=>"000111000",
  5559=>"111111111",
  5560=>"001110111",
  5561=>"011011010",
  5562=>"010110110",
  5563=>"111111111",
  5564=>"000000011",
  5565=>"000000000",
  5566=>"101011011",
  5567=>"100100101",
  5568=>"000000000",
  5569=>"000000000",
  5570=>"111111111",
  5571=>"111011010",
  5572=>"001000111",
  5573=>"000000000",
  5574=>"010000000",
  5575=>"101101111",
  5576=>"011110101",
  5577=>"000000101",
  5578=>"010000011",
  5579=>"111111111",
  5580=>"111111000",
  5581=>"000100101",
  5582=>"011110111",
  5583=>"000000000",
  5584=>"000000000",
  5585=>"011011101",
  5586=>"111111111",
  5587=>"111111111",
  5588=>"100100100",
  5589=>"111001111",
  5590=>"111100110",
  5591=>"001001011",
  5592=>"110101100",
  5593=>"000111111",
  5594=>"000000000",
  5595=>"000000100",
  5596=>"010010111",
  5597=>"000001001",
  5598=>"011111111",
  5599=>"000100101",
  5600=>"000000000",
  5601=>"000000000",
  5602=>"000000111",
  5603=>"000000001",
  5604=>"000000000",
  5605=>"111111011",
  5606=>"111110100",
  5607=>"000100100",
  5608=>"011011000",
  5609=>"111111111",
  5610=>"110000001",
  5611=>"110111111",
  5612=>"100000000",
  5613=>"111101111",
  5614=>"101000000",
  5615=>"111000000",
  5616=>"000000000",
  5617=>"000001101",
  5618=>"001001000",
  5619=>"000101111",
  5620=>"011000111",
  5621=>"000000010",
  5622=>"000000000",
  5623=>"111111010",
  5624=>"111111111",
  5625=>"010010011",
  5626=>"011011000",
  5627=>"111111111",
  5628=>"111111111",
  5629=>"111011111",
  5630=>"101110111",
  5631=>"000000000",
  5632=>"111111110",
  5633=>"000000000",
  5634=>"000000000",
  5635=>"010011111",
  5636=>"111111001",
  5637=>"100000111",
  5638=>"000000000",
  5639=>"111111110",
  5640=>"100101000",
  5641=>"111111111",
  5642=>"000101111",
  5643=>"011011111",
  5644=>"001001111",
  5645=>"000100111",
  5646=>"101111111",
  5647=>"111111000",
  5648=>"000000000",
  5649=>"001011011",
  5650=>"100100000",
  5651=>"111110000",
  5652=>"000000000",
  5653=>"000011000",
  5654=>"000000000",
  5655=>"011011011",
  5656=>"001001000",
  5657=>"000000000",
  5658=>"111111111",
  5659=>"110111100",
  5660=>"111111101",
  5661=>"111111000",
  5662=>"101101111",
  5663=>"000100000",
  5664=>"011000000",
  5665=>"111111110",
  5666=>"110111111",
  5667=>"000000000",
  5668=>"110111111",
  5669=>"110110000",
  5670=>"000110111",
  5671=>"000000111",
  5672=>"011011001",
  5673=>"111000000",
  5674=>"111001111",
  5675=>"111000000",
  5676=>"010000000",
  5677=>"100110111",
  5678=>"100100110",
  5679=>"000000000",
  5680=>"111111111",
  5681=>"001000011",
  5682=>"111111111",
  5683=>"111111000",
  5684=>"000000000",
  5685=>"100100111",
  5686=>"111111001",
  5687=>"000000000",
  5688=>"111111111",
  5689=>"111101100",
  5690=>"000000000",
  5691=>"001000000",
  5692=>"111111111",
  5693=>"101110110",
  5694=>"111111001",
  5695=>"000000000",
  5696=>"001001000",
  5697=>"001001001",
  5698=>"000010111",
  5699=>"111000000",
  5700=>"111111011",
  5701=>"111111111",
  5702=>"000000000",
  5703=>"000000000",
  5704=>"111111011",
  5705=>"000000000",
  5706=>"111111111",
  5707=>"000000000",
  5708=>"111111111",
  5709=>"011111111",
  5710=>"000000000",
  5711=>"111011111",
  5712=>"111111000",
  5713=>"000100111",
  5714=>"000001111",
  5715=>"000001111",
  5716=>"000000000",
  5717=>"101111011",
  5718=>"001001000",
  5719=>"000000000",
  5720=>"011000001",
  5721=>"100110000",
  5722=>"000000000",
  5723=>"111001001",
  5724=>"000001001",
  5725=>"110101111",
  5726=>"111111111",
  5727=>"000111111",
  5728=>"100000000",
  5729=>"111000100",
  5730=>"000011111",
  5731=>"111111010",
  5732=>"001001010",
  5733=>"111111111",
  5734=>"111111111",
  5735=>"000001011",
  5736=>"000000000",
  5737=>"100000010",
  5738=>"111001111",
  5739=>"011111111",
  5740=>"111111111",
  5741=>"001000101",
  5742=>"000000101",
  5743=>"000001111",
  5744=>"100110101",
  5745=>"110111110",
  5746=>"000001011",
  5747=>"111000011",
  5748=>"000100000",
  5749=>"000000111",
  5750=>"111111111",
  5751=>"000000110",
  5752=>"000010000",
  5753=>"000000100",
  5754=>"000000111",
  5755=>"000000000",
  5756=>"101101100",
  5757=>"111111111",
  5758=>"000000111",
  5759=>"110111111",
  5760=>"000000000",
  5761=>"011111011",
  5762=>"110111101",
  5763=>"111111111",
  5764=>"111110000",
  5765=>"111100110",
  5766=>"000000000",
  5767=>"000011000",
  5768=>"111000000",
  5769=>"111111111",
  5770=>"000001111",
  5771=>"101001000",
  5772=>"111110110",
  5773=>"110000111",
  5774=>"110110000",
  5775=>"000000000",
  5776=>"100001101",
  5777=>"001000001",
  5778=>"000000111",
  5779=>"111111001",
  5780=>"001000000",
  5781=>"011111000",
  5782=>"000000000",
  5783=>"111111000",
  5784=>"001000001",
  5785=>"000000000",
  5786=>"000010001",
  5787=>"111010000",
  5788=>"000000000",
  5789=>"111111000",
  5790=>"110000000",
  5791=>"111111111",
  5792=>"000000001",
  5793=>"000000000",
  5794=>"011111111",
  5795=>"000000000",
  5796=>"001000111",
  5797=>"101111111",
  5798=>"101111010",
  5799=>"111111111",
  5800=>"000000100",
  5801=>"100111111",
  5802=>"001000000",
  5803=>"000000000",
  5804=>"001110111",
  5805=>"100100000",
  5806=>"000111111",
  5807=>"111111000",
  5808=>"111111000",
  5809=>"001111111",
  5810=>"011111111",
  5811=>"011000000",
  5812=>"100100001",
  5813=>"110110110",
  5814=>"000000000",
  5815=>"001101000",
  5816=>"000000000",
  5817=>"000000000",
  5818=>"000000101",
  5819=>"111111000",
  5820=>"111111111",
  5821=>"000000000",
  5822=>"111110111",
  5823=>"000000111",
  5824=>"100100100",
  5825=>"011111111",
  5826=>"111111111",
  5827=>"101111100",
  5828=>"000000000",
  5829=>"111000000",
  5830=>"000000111",
  5831=>"111111011",
  5832=>"000000000",
  5833=>"111111111",
  5834=>"000010110",
  5835=>"000000111",
  5836=>"100100110",
  5837=>"000000000",
  5838=>"000110110",
  5839=>"011011000",
  5840=>"100000000",
  5841=>"001010010",
  5842=>"000000010",
  5843=>"000000000",
  5844=>"000000100",
  5845=>"111111011",
  5846=>"111111100",
  5847=>"111110000",
  5848=>"000000111",
  5849=>"111111100",
  5850=>"110101111",
  5851=>"000111111",
  5852=>"100100111",
  5853=>"111111000",
  5854=>"110111000",
  5855=>"010000110",
  5856=>"000000000",
  5857=>"111011011",
  5858=>"111001001",
  5859=>"100111111",
  5860=>"000000000",
  5861=>"100011001",
  5862=>"000000000",
  5863=>"111111111",
  5864=>"000000000",
  5865=>"111111001",
  5866=>"000111111",
  5867=>"000000111",
  5868=>"000110110",
  5869=>"111111111",
  5870=>"111111100",
  5871=>"000000000",
  5872=>"000000000",
  5873=>"001000111",
  5874=>"111111111",
  5875=>"000000001",
  5876=>"111111011",
  5877=>"000111111",
  5878=>"110001001",
  5879=>"000000001",
  5880=>"000111111",
  5881=>"000000000",
  5882=>"101111011",
  5883=>"000000000",
  5884=>"100110110",
  5885=>"111111001",
  5886=>"111101111",
  5887=>"000000000",
  5888=>"001000001",
  5889=>"111001001",
  5890=>"000000000",
  5891=>"101000000",
  5892=>"000000000",
  5893=>"000000100",
  5894=>"111111100",
  5895=>"111110000",
  5896=>"001011111",
  5897=>"000000000",
  5898=>"111111100",
  5899=>"111111010",
  5900=>"000000000",
  5901=>"100000111",
  5902=>"000110110",
  5903=>"100110110",
  5904=>"010010000",
  5905=>"001100000",
  5906=>"011111111",
  5907=>"011001001",
  5908=>"110110000",
  5909=>"000000111",
  5910=>"110100000",
  5911=>"000000111",
  5912=>"000000111",
  5913=>"110000000",
  5914=>"111111001",
  5915=>"111111110",
  5916=>"111111111",
  5917=>"110000000",
  5918=>"000011101",
  5919=>"000000000",
  5920=>"100100000",
  5921=>"001000000",
  5922=>"100100111",
  5923=>"000010000",
  5924=>"111000000",
  5925=>"000000000",
  5926=>"111100100",
  5927=>"111010000",
  5928=>"111111111",
  5929=>"000111000",
  5930=>"000000110",
  5931=>"011010010",
  5932=>"000011111",
  5933=>"110000000",
  5934=>"000010000",
  5935=>"101001001",
  5936=>"101001001",
  5937=>"011111001",
  5938=>"111111011",
  5939=>"011001011",
  5940=>"111111000",
  5941=>"110110010",
  5942=>"000000101",
  5943=>"000000000",
  5944=>"000000100",
  5945=>"001000111",
  5946=>"010010000",
  5947=>"100111111",
  5948=>"011001000",
  5949=>"111111101",
  5950=>"010111111",
  5951=>"000000000",
  5952=>"111111100",
  5953=>"111111110",
  5954=>"000111111",
  5955=>"000000000",
  5956=>"101110000",
  5957=>"000000001",
  5958=>"000000111",
  5959=>"000000111",
  5960=>"000111011",
  5961=>"000000000",
  5962=>"111111010",
  5963=>"100110100",
  5964=>"000000000",
  5965=>"111111011",
  5966=>"000000000",
  5967=>"000000110",
  5968=>"100101111",
  5969=>"000000000",
  5970=>"110010111",
  5971=>"111001000",
  5972=>"001001111",
  5973=>"011011011",
  5974=>"111111110",
  5975=>"101111111",
  5976=>"000101000",
  5977=>"000000000",
  5978=>"110100000",
  5979=>"001111011",
  5980=>"000000000",
  5981=>"000000000",
  5982=>"111110110",
  5983=>"111101111",
  5984=>"100000001",
  5985=>"000011110",
  5986=>"110100000",
  5987=>"000000000",
  5988=>"101100000",
  5989=>"100000000",
  5990=>"000000011",
  5991=>"111111000",
  5992=>"111111111",
  5993=>"011111001",
  5994=>"110110000",
  5995=>"000010001",
  5996=>"111111011",
  5997=>"000000000",
  5998=>"000000000",
  5999=>"000000000",
  6000=>"000000111",
  6001=>"111110111",
  6002=>"000100000",
  6003=>"000000110",
  6004=>"000000011",
  6005=>"111111101",
  6006=>"001001000",
  6007=>"001011011",
  6008=>"001001111",
  6009=>"000000000",
  6010=>"111111011",
  6011=>"110111100",
  6012=>"111111111",
  6013=>"011010010",
  6014=>"111110000",
  6015=>"111111111",
  6016=>"000100100",
  6017=>"000000011",
  6018=>"111111111",
  6019=>"000000000",
  6020=>"000111111",
  6021=>"000000000",
  6022=>"000111111",
  6023=>"001000000",
  6024=>"111111111",
  6025=>"000001001",
  6026=>"001001000",
  6027=>"111000000",
  6028=>"111011111",
  6029=>"100100111",
  6030=>"000000000",
  6031=>"001011001",
  6032=>"000111111",
  6033=>"100000000",
  6034=>"111001011",
  6035=>"100000000",
  6036=>"100101111",
  6037=>"000000000",
  6038=>"111111111",
  6039=>"111011111",
  6040=>"000111011",
  6041=>"000110001",
  6042=>"111111011",
  6043=>"111010111",
  6044=>"000000001",
  6045=>"111111000",
  6046=>"000000000",
  6047=>"000000110",
  6048=>"001001111",
  6049=>"111111000",
  6050=>"100000000",
  6051=>"001000000",
  6052=>"000000000",
  6053=>"011111000",
  6054=>"000000000",
  6055=>"100111000",
  6056=>"000000000",
  6057=>"111111111",
  6058=>"000110111",
  6059=>"000000000",
  6060=>"000000001",
  6061=>"000000000",
  6062=>"000000000",
  6063=>"111111111",
  6064=>"101000000",
  6065=>"000111011",
  6066=>"000111000",
  6067=>"000111101",
  6068=>"000111111",
  6069=>"111111000",
  6070=>"111111101",
  6071=>"111111111",
  6072=>"000000000",
  6073=>"011011111",
  6074=>"111111111",
  6075=>"000000111",
  6076=>"111001001",
  6077=>"111111011",
  6078=>"000000101",
  6079=>"111111101",
  6080=>"000000001",
  6081=>"000000000",
  6082=>"000000101",
  6083=>"111100000",
  6084=>"111010000",
  6085=>"111101000",
  6086=>"000000001",
  6087=>"000000000",
  6088=>"001000111",
  6089=>"000000110",
  6090=>"101000101",
  6091=>"110111011",
  6092=>"111000000",
  6093=>"111111001",
  6094=>"000000000",
  6095=>"111111111",
  6096=>"110000110",
  6097=>"111111111",
  6098=>"010111011",
  6099=>"011000000",
  6100=>"101000000",
  6101=>"000111010",
  6102=>"000000000",
  6103=>"000111110",
  6104=>"111111100",
  6105=>"000011001",
  6106=>"011000011",
  6107=>"000000000",
  6108=>"000000000",
  6109=>"111110000",
  6110=>"111111001",
  6111=>"001000001",
  6112=>"001000100",
  6113=>"111011001",
  6114=>"000111111",
  6115=>"111101001",
  6116=>"100111100",
  6117=>"000001000",
  6118=>"110111111",
  6119=>"000000111",
  6120=>"000000000",
  6121=>"001111111",
  6122=>"111011000",
  6123=>"000000000",
  6124=>"100000000",
  6125=>"000000000",
  6126=>"000111011",
  6127=>"111110110",
  6128=>"001000000",
  6129=>"100000000",
  6130=>"000000100",
  6131=>"001111111",
  6132=>"000000111",
  6133=>"000000000",
  6134=>"100101111",
  6135=>"100111110",
  6136=>"000000000",
  6137=>"000000000",
  6138=>"000000000",
  6139=>"100000000",
  6140=>"111000111",
  6141=>"111111100",
  6142=>"000111111",
  6143=>"000000000",
  6144=>"111111011",
  6145=>"011010000",
  6146=>"111111111",
  6147=>"101000000",
  6148=>"000001111",
  6149=>"100000000",
  6150=>"000111000",
  6151=>"000000111",
  6152=>"000000000",
  6153=>"111111111",
  6154=>"111000000",
  6155=>"110010110",
  6156=>"001001011",
  6157=>"111111111",
  6158=>"111011011",
  6159=>"111111111",
  6160=>"000000000",
  6161=>"011111000",
  6162=>"000111111",
  6163=>"101000000",
  6164=>"000000001",
  6165=>"000000000",
  6166=>"110100000",
  6167=>"000001000",
  6168=>"010100100",
  6169=>"111111001",
  6170=>"000001000",
  6171=>"000000000",
  6172=>"000000001",
  6173=>"000111100",
  6174=>"000011111",
  6175=>"100100111",
  6176=>"100000000",
  6177=>"000001111",
  6178=>"111111111",
  6179=>"111000111",
  6180=>"000000000",
  6181=>"000111111",
  6182=>"111111011",
  6183=>"110111111",
  6184=>"000000100",
  6185=>"000111111",
  6186=>"000000000",
  6187=>"101111111",
  6188=>"111111110",
  6189=>"111111111",
  6190=>"000000000",
  6191=>"111111110",
  6192=>"000000000",
  6193=>"000111111",
  6194=>"000010010",
  6195=>"000001011",
  6196=>"110110000",
  6197=>"000010011",
  6198=>"000000100",
  6199=>"001000000",
  6200=>"111111010",
  6201=>"110111011",
  6202=>"000000111",
  6203=>"000000000",
  6204=>"000000000",
  6205=>"111110100",
  6206=>"111100110",
  6207=>"111000000",
  6208=>"000001000",
  6209=>"001000110",
  6210=>"001001000",
  6211=>"100100100",
  6212=>"100000000",
  6213=>"011011111",
  6214=>"011000000",
  6215=>"111111111",
  6216=>"110110110",
  6217=>"000000111",
  6218=>"001000101",
  6219=>"111100100",
  6220=>"110100110",
  6221=>"000101111",
  6222=>"001000000",
  6223=>"110010000",
  6224=>"000000000",
  6225=>"101111111",
  6226=>"000000000",
  6227=>"000000000",
  6228=>"111101111",
  6229=>"001000000",
  6230=>"011001111",
  6231=>"111111000",
  6232=>"110111111",
  6233=>"111101111",
  6234=>"111111111",
  6235=>"111111011",
  6236=>"000000000",
  6237=>"010000100",
  6238=>"000100010",
  6239=>"100100000",
  6240=>"000111111",
  6241=>"110111000",
  6242=>"000000000",
  6243=>"000000000",
  6244=>"011110001",
  6245=>"000000000",
  6246=>"111110100",
  6247=>"111100100",
  6248=>"000000000",
  6249=>"111111000",
  6250=>"111111110",
  6251=>"111111111",
  6252=>"001011111",
  6253=>"000111111",
  6254=>"001000000",
  6255=>"000000000",
  6256=>"111111011",
  6257=>"000110110",
  6258=>"001001000",
  6259=>"101100000",
  6260=>"100111111",
  6261=>"000000000",
  6262=>"001000000",
  6263=>"000000110",
  6264=>"000111000",
  6265=>"001111111",
  6266=>"101001000",
  6267=>"000111111",
  6268=>"111101001",
  6269=>"111100100",
  6270=>"001001011",
  6271=>"111001110",
  6272=>"111111111",
  6273=>"111100111",
  6274=>"111111111",
  6275=>"000000110",
  6276=>"011001000",
  6277=>"001000111",
  6278=>"110000001",
  6279=>"111111000",
  6280=>"010110111",
  6281=>"000000000",
  6282=>"000000001",
  6283=>"110111111",
  6284=>"110111111",
  6285=>"110000000",
  6286=>"110111000",
  6287=>"000101111",
  6288=>"111111111",
  6289=>"111111111",
  6290=>"000000000",
  6291=>"111000010",
  6292=>"000111111",
  6293=>"011011000",
  6294=>"111111011",
  6295=>"111111000",
  6296=>"000000010",
  6297=>"111101110",
  6298=>"100101011",
  6299=>"000111111",
  6300=>"000000110",
  6301=>"000000000",
  6302=>"001111110",
  6303=>"111111111",
  6304=>"000000110",
  6305=>"111111001",
  6306=>"111010000",
  6307=>"110000000",
  6308=>"100110000",
  6309=>"100110000",
  6310=>"000000000",
  6311=>"111110110",
  6312=>"000000000",
  6313=>"000000000",
  6314=>"101001000",
  6315=>"001111111",
  6316=>"100111100",
  6317=>"111110100",
  6318=>"000000000",
  6319=>"111111000",
  6320=>"111100111",
  6321=>"010111110",
  6322=>"111111111",
  6323=>"111000000",
  6324=>"000000000",
  6325=>"000000000",
  6326=>"110000000",
  6327=>"110110000",
  6328=>"111111111",
  6329=>"111111101",
  6330=>"110000010",
  6331=>"110010110",
  6332=>"000000000",
  6333=>"111111110",
  6334=>"111111101",
  6335=>"000000000",
  6336=>"111011001",
  6337=>"000110000",
  6338=>"000000000",
  6339=>"101111111",
  6340=>"110110000",
  6341=>"000010000",
  6342=>"000000111",
  6343=>"000001101",
  6344=>"001001001",
  6345=>"110000000",
  6346=>"000111111",
  6347=>"111111110",
  6348=>"110110110",
  6349=>"100100000",
  6350=>"111111100",
  6351=>"000000000",
  6352=>"010000000",
  6353=>"010110010",
  6354=>"000000000",
  6355=>"010110100",
  6356=>"111111000",
  6357=>"000000001",
  6358=>"010000000",
  6359=>"000001011",
  6360=>"111011000",
  6361=>"000000111",
  6362=>"111111111",
  6363=>"111000000",
  6364=>"011001111",
  6365=>"111111111",
  6366=>"010011001",
  6367=>"111000000",
  6368=>"111000000",
  6369=>"001000000",
  6370=>"101000100",
  6371=>"000110111",
  6372=>"000000000",
  6373=>"111110110",
  6374=>"111100001",
  6375=>"000000000",
  6376=>"111011000",
  6377=>"110110110",
  6378=>"111000000",
  6379=>"111000000",
  6380=>"011011001",
  6381=>"000110111",
  6382=>"110111111",
  6383=>"110111111",
  6384=>"001001111",
  6385=>"000111001",
  6386=>"111000000",
  6387=>"111001000",
  6388=>"111000000",
  6389=>"001011000",
  6390=>"000000110",
  6391=>"100111111",
  6392=>"000111111",
  6393=>"111100100",
  6394=>"110111111",
  6395=>"010000000",
  6396=>"011111111",
  6397=>"110111000",
  6398=>"000000110",
  6399=>"100111111",
  6400=>"000000100",
  6401=>"110110000",
  6402=>"000000000",
  6403=>"111110010",
  6404=>"000000111",
  6405=>"000000110",
  6406=>"000000111",
  6407=>"000011100",
  6408=>"000111111",
  6409=>"111111001",
  6410=>"111111100",
  6411=>"000001001",
  6412=>"000000111",
  6413=>"000110111",
  6414=>"100111111",
  6415=>"000000000",
  6416=>"000001000",
  6417=>"111111000",
  6418=>"111111111",
  6419=>"000000000",
  6420=>"001011000",
  6421=>"000001001",
  6422=>"111111101",
  6423=>"000000111",
  6424=>"010001001",
  6425=>"111110110",
  6426=>"100000110",
  6427=>"001001001",
  6428=>"111100111",
  6429=>"000100000",
  6430=>"000101000",
  6431=>"110000000",
  6432=>"111111001",
  6433=>"000000011",
  6434=>"001001000",
  6435=>"000000000",
  6436=>"000001011",
  6437=>"000000000",
  6438=>"111111011",
  6439=>"000111101",
  6440=>"111111000",
  6441=>"111111111",
  6442=>"110111001",
  6443=>"111111111",
  6444=>"111111011",
  6445=>"000001101",
  6446=>"000000000",
  6447=>"000000000",
  6448=>"110111111",
  6449=>"000000111",
  6450=>"011000001",
  6451=>"000000000",
  6452=>"111111111",
  6453=>"111000000",
  6454=>"000000111",
  6455=>"111101000",
  6456=>"111111000",
  6457=>"111100111",
  6458=>"000000111",
  6459=>"000000000",
  6460=>"000000000",
  6461=>"100100100",
  6462=>"000100110",
  6463=>"000000000",
  6464=>"000001000",
  6465=>"111111011",
  6466=>"000000000",
  6467=>"110100100",
  6468=>"111000111",
  6469=>"111111001",
  6470=>"000000000",
  6471=>"111111111",
  6472=>"111111111",
  6473=>"111111011",
  6474=>"000100001",
  6475=>"110100000",
  6476=>"000000000",
  6477=>"001000000",
  6478=>"110011111",
  6479=>"110110010",
  6480=>"110110111",
  6481=>"000101111",
  6482=>"001011001",
  6483=>"111111111",
  6484=>"000111110",
  6485=>"001100111",
  6486=>"000000000",
  6487=>"110111111",
  6488=>"111111111",
  6489=>"000000000",
  6490=>"011111111",
  6491=>"000000000",
  6492=>"000111111",
  6493=>"111111111",
  6494=>"000000000",
  6495=>"100000000",
  6496=>"111011000",
  6497=>"001101111",
  6498=>"000100001",
  6499=>"000001111",
  6500=>"010111111",
  6501=>"111000000",
  6502=>"101000000",
  6503=>"100101111",
  6504=>"001011111",
  6505=>"111000000",
  6506=>"000111111",
  6507=>"000000000",
  6508=>"000010111",
  6509=>"110110110",
  6510=>"000000000",
  6511=>"111011001",
  6512=>"000000000",
  6513=>"001101111",
  6514=>"010000000",
  6515=>"000000000",
  6516=>"111110111",
  6517=>"000111111",
  6518=>"000110111",
  6519=>"000000111",
  6520=>"111111111",
  6521=>"000000000",
  6522=>"111000000",
  6523=>"000000000",
  6524=>"100100000",
  6525=>"010100000",
  6526=>"111111000",
  6527=>"111000000",
  6528=>"000110110",
  6529=>"000000000",
  6530=>"110110110",
  6531=>"000100111",
  6532=>"111000000",
  6533=>"111111010",
  6534=>"001000000",
  6535=>"110000000",
  6536=>"001001011",
  6537=>"010000000",
  6538=>"100100110",
  6539=>"111111111",
  6540=>"111001111",
  6541=>"000000000",
  6542=>"000111111",
  6543=>"000000000",
  6544=>"000000001",
  6545=>"000000001",
  6546=>"101101100",
  6547=>"110111111",
  6548=>"111111111",
  6549=>"000000000",
  6550=>"000000000",
  6551=>"111111111",
  6552=>"111111111",
  6553=>"011001000",
  6554=>"111111111",
  6555=>"111000000",
  6556=>"000000000",
  6557=>"011010111",
  6558=>"111110110",
  6559=>"111111011",
  6560=>"001111111",
  6561=>"010110110",
  6562=>"011001011",
  6563=>"111111111",
  6564=>"001000000",
  6565=>"111111111",
  6566=>"000000000",
  6567=>"010111111",
  6568=>"010110010",
  6569=>"100100111",
  6570=>"000000001",
  6571=>"111000001",
  6572=>"000000000",
  6573=>"000111111",
  6574=>"100111111",
  6575=>"000001011",
  6576=>"111011111",
  6577=>"011011000",
  6578=>"010001000",
  6579=>"011111111",
  6580=>"110000111",
  6581=>"100100000",
  6582=>"000000001",
  6583=>"000000111",
  6584=>"111111111",
  6585=>"011111001",
  6586=>"000000000",
  6587=>"111000100",
  6588=>"000010000",
  6589=>"000110100",
  6590=>"111111000",
  6591=>"110101101",
  6592=>"001001111",
  6593=>"000000010",
  6594=>"010110111",
  6595=>"000000100",
  6596=>"000001100",
  6597=>"010111111",
  6598=>"001000111",
  6599=>"000000000",
  6600=>"100000011",
  6601=>"111111111",
  6602=>"101001100",
  6603=>"111111000",
  6604=>"111111010",
  6605=>"111010111",
  6606=>"000000000",
  6607=>"001001000",
  6608=>"000000000",
  6609=>"111010000",
  6610=>"000000001",
  6611=>"000000000",
  6612=>"000000100",
  6613=>"001101111",
  6614=>"010011111",
  6615=>"110111111",
  6616=>"100000110",
  6617=>"111111111",
  6618=>"110110000",
  6619=>"000000111",
  6620=>"000000000",
  6621=>"110111000",
  6622=>"001000000",
  6623=>"000100110",
  6624=>"000101000",
  6625=>"111101111",
  6626=>"010110000",
  6627=>"010000000",
  6628=>"111011111",
  6629=>"001000001",
  6630=>"111111000",
  6631=>"100110111",
  6632=>"111111000",
  6633=>"100110111",
  6634=>"110110111",
  6635=>"111111010",
  6636=>"110111110",
  6637=>"111111101",
  6638=>"000000000",
  6639=>"111111111",
  6640=>"111111111",
  6641=>"011011111",
  6642=>"000000000",
  6643=>"000001000",
  6644=>"111111000",
  6645=>"111001000",
  6646=>"000000000",
  6647=>"111110000",
  6648=>"000000000",
  6649=>"110111011",
  6650=>"000000001",
  6651=>"101100000",
  6652=>"010000010",
  6653=>"000000001",
  6654=>"111110111",
  6655=>"000000110",
  6656=>"000111101",
  6657=>"000000000",
  6658=>"111111111",
  6659=>"000000000",
  6660=>"111011111",
  6661=>"011111111",
  6662=>"000000000",
  6663=>"111111111",
  6664=>"111111111",
  6665=>"111111000",
  6666=>"000000000",
  6667=>"000000011",
  6668=>"000001011",
  6669=>"000000000",
  6670=>"111111111",
  6671=>"111111111",
  6672=>"110110110",
  6673=>"000000001",
  6674=>"000011111",
  6675=>"110000000",
  6676=>"111111100",
  6677=>"000000100",
  6678=>"010110000",
  6679=>"111111011",
  6680=>"000000000",
  6681=>"011000001",
  6682=>"111101111",
  6683=>"111111111",
  6684=>"111111111",
  6685=>"111110110",
  6686=>"000000000",
  6687=>"000001001",
  6688=>"000000000",
  6689=>"110111000",
  6690=>"000000111",
  6691=>"011011111",
  6692=>"111111111",
  6693=>"000000000",
  6694=>"000000000",
  6695=>"000000100",
  6696=>"000011000",
  6697=>"000110000",
  6698=>"111111111",
  6699=>"111000000",
  6700=>"000000000",
  6701=>"000000111",
  6702=>"111111011",
  6703=>"000000000",
  6704=>"000000011",
  6705=>"110000000",
  6706=>"011111101",
  6707=>"011111111",
  6708=>"000000010",
  6709=>"000010110",
  6710=>"000000000",
  6711=>"111011110",
  6712=>"000000100",
  6713=>"110100110",
  6714=>"100100110",
  6715=>"110100000",
  6716=>"000000101",
  6717=>"111111111",
  6718=>"010111110",
  6719=>"000000000",
  6720=>"110110110",
  6721=>"100000101",
  6722=>"110111111",
  6723=>"111110111",
  6724=>"010010111",
  6725=>"000000100",
  6726=>"000000000",
  6727=>"111111101",
  6728=>"111111010",
  6729=>"000000101",
  6730=>"111111111",
  6731=>"000000000",
  6732=>"111111000",
  6733=>"110100000",
  6734=>"000000001",
  6735=>"110000111",
  6736=>"000010110",
  6737=>"111001011",
  6738=>"000000001",
  6739=>"000000000",
  6740=>"000000000",
  6741=>"000000000",
  6742=>"001001111",
  6743=>"000000000",
  6744=>"000000000",
  6745=>"111111111",
  6746=>"111111111",
  6747=>"000100100",
  6748=>"001111111",
  6749=>"000000000",
  6750=>"101101110",
  6751=>"110000000",
  6752=>"000000000",
  6753=>"001001111",
  6754=>"111111111",
  6755=>"001000000",
  6756=>"000000110",
  6757=>"100100111",
  6758=>"111111111",
  6759=>"000000000",
  6760=>"011111111",
  6761=>"101101111",
  6762=>"111100100",
  6763=>"111110000",
  6764=>"001011011",
  6765=>"000000000",
  6766=>"010000010",
  6767=>"000000100",
  6768=>"001011101",
  6769=>"011000100",
  6770=>"000000000",
  6771=>"110111111",
  6772=>"111111111",
  6773=>"110100100",
  6774=>"000000000",
  6775=>"110101111",
  6776=>"011011111",
  6777=>"000010011",
  6778=>"000000110",
  6779=>"000100110",
  6780=>"111000100",
  6781=>"010011000",
  6782=>"001011111",
  6783=>"110111111",
  6784=>"000000010",
  6785=>"000000000",
  6786=>"000000000",
  6787=>"011001100",
  6788=>"111111111",
  6789=>"111110111",
  6790=>"010010110",
  6791=>"101101000",
  6792=>"111111111",
  6793=>"111011001",
  6794=>"111111011",
  6795=>"000000000",
  6796=>"111111100",
  6797=>"000011111",
  6798=>"111110000",
  6799=>"111111001",
  6800=>"010000000",
  6801=>"011001000",
  6802=>"000110110",
  6803=>"010011111",
  6804=>"000000000",
  6805=>"110110000",
  6806=>"100100110",
  6807=>"000000000",
  6808=>"000000000",
  6809=>"001011111",
  6810=>"111111001",
  6811=>"000000000",
  6812=>"110111110",
  6813=>"100000000",
  6814=>"001000000",
  6815=>"111111111",
  6816=>"111111111",
  6817=>"000000100",
  6818=>"001001011",
  6819=>"000001111",
  6820=>"000000000",
  6821=>"100000100",
  6822=>"111111111",
  6823=>"011111011",
  6824=>"000000000",
  6825=>"001001001",
  6826=>"100000000",
  6827=>"111100000",
  6828=>"000000100",
  6829=>"000011011",
  6830=>"011011001",
  6831=>"011001001",
  6832=>"111111011",
  6833=>"111111111",
  6834=>"111111111",
  6835=>"001000101",
  6836=>"000000000",
  6837=>"110011001",
  6838=>"011011011",
  6839=>"111110111",
  6840=>"011001001",
  6841=>"000000000",
  6842=>"000000000",
  6843=>"110110111",
  6844=>"111111111",
  6845=>"000100110",
  6846=>"000000000",
  6847=>"000101111",
  6848=>"011111111",
  6849=>"011111111",
  6850=>"000000100",
  6851=>"111011111",
  6852=>"000000000",
  6853=>"000000000",
  6854=>"000000000",
  6855=>"100000000",
  6856=>"010010000",
  6857=>"111001001",
  6858=>"110100101",
  6859=>"110110010",
  6860=>"001001111",
  6861=>"000000000",
  6862=>"111011011",
  6863=>"000000000",
  6864=>"000100000",
  6865=>"011011010",
  6866=>"111111000",
  6867=>"000000000",
  6868=>"000111001",
  6869=>"000000000",
  6870=>"000000000",
  6871=>"001000000",
  6872=>"100000000",
  6873=>"011011110",
  6874=>"111110111",
  6875=>"100111111",
  6876=>"001111111",
  6877=>"000000110",
  6878=>"111111001",
  6879=>"000000000",
  6880=>"111001001",
  6881=>"001000000",
  6882=>"000000000",
  6883=>"111111111",
  6884=>"000000000",
  6885=>"000000000",
  6886=>"000000000",
  6887=>"000000000",
  6888=>"111111000",
  6889=>"001000000",
  6890=>"000000101",
  6891=>"100111111",
  6892=>"101111001",
  6893=>"000100111",
  6894=>"011001000",
  6895=>"111001011",
  6896=>"111111111",
  6897=>"100111011",
  6898=>"111111111",
  6899=>"000000000",
  6900=>"100110110",
  6901=>"110000000",
  6902=>"111111111",
  6903=>"001001000",
  6904=>"000000100",
  6905=>"111101001",
  6906=>"100000111",
  6907=>"011111010",
  6908=>"000000000",
  6909=>"111001001",
  6910=>"110111000",
  6911=>"111111110",
  6912=>"111011001",
  6913=>"000001000",
  6914=>"000000100",
  6915=>"000001000",
  6916=>"000000000",
  6917=>"111111111",
  6918=>"000000000",
  6919=>"111100111",
  6920=>"011001100",
  6921=>"000000000",
  6922=>"111011001",
  6923=>"000000000",
  6924=>"101000000",
  6925=>"010010000",
  6926=>"011011111",
  6927=>"000000000",
  6928=>"111000000",
  6929=>"110000000",
  6930=>"110110110",
  6931=>"111111111",
  6932=>"101001000",
  6933=>"101000011",
  6934=>"001000000",
  6935=>"000000000",
  6936=>"111111100",
  6937=>"000000000",
  6938=>"110011000",
  6939=>"111110100",
  6940=>"000000000",
  6941=>"001000001",
  6942=>"000111111",
  6943=>"011101100",
  6944=>"100100111",
  6945=>"000000000",
  6946=>"000100000",
  6947=>"001011111",
  6948=>"000000000",
  6949=>"000000001",
  6950=>"000000000",
  6951=>"100100111",
  6952=>"000001000",
  6953=>"000000000",
  6954=>"010110111",
  6955=>"000100110",
  6956=>"000000000",
  6957=>"000100100",
  6958=>"110111001",
  6959=>"001001001",
  6960=>"111000011",
  6961=>"100000000",
  6962=>"000000000",
  6963=>"100000010",
  6964=>"000000111",
  6965=>"011001000",
  6966=>"110110110",
  6967=>"000000000",
  6968=>"000000100",
  6969=>"111100111",
  6970=>"110110111",
  6971=>"111111111",
  6972=>"010110110",
  6973=>"111111111",
  6974=>"101001001",
  6975=>"000100000",
  6976=>"111111111",
  6977=>"000011000",
  6978=>"111101111",
  6979=>"101001000",
  6980=>"000000100",
  6981=>"000111000",
  6982=>"111111000",
  6983=>"000000111",
  6984=>"110100001",
  6985=>"000001011",
  6986=>"000001111",
  6987=>"111111000",
  6988=>"000000100",
  6989=>"001110111",
  6990=>"100000000",
  6991=>"010000000",
  6992=>"100111011",
  6993=>"000000000",
  6994=>"110000000",
  6995=>"100111011",
  6996=>"000000000",
  6997=>"011011011",
  6998=>"000000000",
  6999=>"111111111",
  7000=>"111111111",
  7001=>"110111111",
  7002=>"000000000",
  7003=>"110100111",
  7004=>"111100100",
  7005=>"111111111",
  7006=>"000000000",
  7007=>"000000000",
  7008=>"001111100",
  7009=>"111111111",
  7010=>"111011001",
  7011=>"000000000",
  7012=>"000000000",
  7013=>"111111111",
  7014=>"000111111",
  7015=>"110010000",
  7016=>"001000001",
  7017=>"110010000",
  7018=>"111100000",
  7019=>"111111011",
  7020=>"000000000",
  7021=>"110110110",
  7022=>"100101100",
  7023=>"111001000",
  7024=>"100110110",
  7025=>"100100101",
  7026=>"111111101",
  7027=>"111000000",
  7028=>"111110111",
  7029=>"000000000",
  7030=>"111111111",
  7031=>"000000000",
  7032=>"110000111",
  7033=>"111101000",
  7034=>"110111010",
  7035=>"111111111",
  7036=>"000000000",
  7037=>"111111010",
  7038=>"110000010",
  7039=>"011111011",
  7040=>"011111111",
  7041=>"001001011",
  7042=>"000000001",
  7043=>"111111110",
  7044=>"110111111",
  7045=>"000111111",
  7046=>"100100100",
  7047=>"101111111",
  7048=>"000010111",
  7049=>"101001000",
  7050=>"001000000",
  7051=>"011000000",
  7052=>"001001111",
  7053=>"111111100",
  7054=>"011000111",
  7055=>"000000010",
  7056=>"000001001",
  7057=>"011111111",
  7058=>"000000110",
  7059=>"000000001",
  7060=>"111110000",
  7061=>"000000011",
  7062=>"111011011",
  7063=>"000000000",
  7064=>"000001000",
  7065=>"000100110",
  7066=>"000000001",
  7067=>"011111111",
  7068=>"000000000",
  7069=>"000000000",
  7070=>"000000000",
  7071=>"111111111",
  7072=>"111111111",
  7073=>"001011111",
  7074=>"010000100",
  7075=>"111111111",
  7076=>"111111111",
  7077=>"100101000",
  7078=>"000000001",
  7079=>"111111111",
  7080=>"001011111",
  7081=>"111111110",
  7082=>"111111111",
  7083=>"000000000",
  7084=>"000000000",
  7085=>"000000000",
  7086=>"000000000",
  7087=>"000111111",
  7088=>"000000000",
  7089=>"111111011",
  7090=>"111111111",
  7091=>"111000000",
  7092=>"111111111",
  7093=>"110111110",
  7094=>"111111011",
  7095=>"111101000",
  7096=>"110111111",
  7097=>"000000000",
  7098=>"111111100",
  7099=>"000000111",
  7100=>"111111111",
  7101=>"000000000",
  7102=>"000000100",
  7103=>"000000100",
  7104=>"000000111",
  7105=>"110000010",
  7106=>"101001101",
  7107=>"111111111",
  7108=>"001111111",
  7109=>"001110111",
  7110=>"000000000",
  7111=>"011001001",
  7112=>"000000000",
  7113=>"101011111",
  7114=>"011110110",
  7115=>"000000011",
  7116=>"100000000",
  7117=>"101000000",
  7118=>"000001000",
  7119=>"000000000",
  7120=>"001001011",
  7121=>"001000000",
  7122=>"111111111",
  7123=>"111111111",
  7124=>"011011000",
  7125=>"000111011",
  7126=>"111111110",
  7127=>"000000111",
  7128=>"001001000",
  7129=>"111111111",
  7130=>"110110111",
  7131=>"100110111",
  7132=>"111100010",
  7133=>"111111111",
  7134=>"111001001",
  7135=>"000001010",
  7136=>"111000001",
  7137=>"000000000",
  7138=>"000000000",
  7139=>"111100100",
  7140=>"001001010",
  7141=>"110110111",
  7142=>"000000000",
  7143=>"100110111",
  7144=>"001000001",
  7145=>"111001000",
  7146=>"000000000",
  7147=>"111000000",
  7148=>"111111111",
  7149=>"111011000",
  7150=>"011111110",
  7151=>"111111101",
  7152=>"000000000",
  7153=>"000000000",
  7154=>"111111111",
  7155=>"000000000",
  7156=>"000000000",
  7157=>"111111111",
  7158=>"000000000",
  7159=>"011001000",
  7160=>"000000000",
  7161=>"011011011",
  7162=>"000111011",
  7163=>"111101100",
  7164=>"101111111",
  7165=>"000000000",
  7166=>"111100111",
  7167=>"000000000",
  7168=>"000000000",
  7169=>"111111110",
  7170=>"011000000",
  7171=>"001001101",
  7172=>"010100100",
  7173=>"010010001",
  7174=>"100000000",
  7175=>"000000011",
  7176=>"001011011",
  7177=>"010011000",
  7178=>"111111110",
  7179=>"111111110",
  7180=>"100110110",
  7181=>"101111111",
  7182=>"000010101",
  7183=>"111111111",
  7184=>"000000000",
  7185=>"111111111",
  7186=>"000100110",
  7187=>"000000000",
  7188=>"001001000",
  7189=>"000000111",
  7190=>"111011001",
  7191=>"001000000",
  7192=>"110110110",
  7193=>"111100110",
  7194=>"111100111",
  7195=>"111111010",
  7196=>"111111011",
  7197=>"110100000",
  7198=>"000000001",
  7199=>"111000001",
  7200=>"100000010",
  7201=>"111111111",
  7202=>"001001001",
  7203=>"000001000",
  7204=>"000000000",
  7205=>"001010000",
  7206=>"000000111",
  7207=>"000000001",
  7208=>"110011000",
  7209=>"000001111",
  7210=>"000000000",
  7211=>"111111000",
  7212=>"000111111",
  7213=>"010000000",
  7214=>"001100100",
  7215=>"011110100",
  7216=>"000000000",
  7217=>"111111001",
  7218=>"001011011",
  7219=>"000001011",
  7220=>"000110110",
  7221=>"111001001",
  7222=>"100000000",
  7223=>"101101111",
  7224=>"011111111",
  7225=>"001111111",
  7226=>"000000000",
  7227=>"000000100",
  7228=>"000000000",
  7229=>"100000000",
  7230=>"110100000",
  7231=>"111100100",
  7232=>"001101001",
  7233=>"000000000",
  7234=>"001100101",
  7235=>"011001000",
  7236=>"111001000",
  7237=>"111011001",
  7238=>"111110000",
  7239=>"111111000",
  7240=>"000000001",
  7241=>"100000000",
  7242=>"010111111",
  7243=>"000000000",
  7244=>"101101000",
  7245=>"100000000",
  7246=>"000000100",
  7247=>"000000000",
  7248=>"000001000",
  7249=>"010111111",
  7250=>"111111110",
  7251=>"001001101",
  7252=>"101111111",
  7253=>"111001101",
  7254=>"111001111",
  7255=>"000000000",
  7256=>"010110110",
  7257=>"111111111",
  7258=>"111111111",
  7259=>"100000000",
  7260=>"111010000",
  7261=>"011000000",
  7262=>"000000000",
  7263=>"001111111",
  7264=>"111000110",
  7265=>"011011011",
  7266=>"011011000",
  7267=>"000000000",
  7268=>"111111111",
  7269=>"111111111",
  7270=>"011011111",
  7271=>"100100110",
  7272=>"000000000",
  7273=>"111111111",
  7274=>"111111111",
  7275=>"111001001",
  7276=>"010000000",
  7277=>"011001000",
  7278=>"110000000",
  7279=>"111000000",
  7280=>"111000000",
  7281=>"000010011",
  7282=>"001111011",
  7283=>"111101111",
  7284=>"111110100",
  7285=>"111111111",
  7286=>"011101111",
  7287=>"000111000",
  7288=>"000000001",
  7289=>"110110100",
  7290=>"000000101",
  7291=>"111111111",
  7292=>"011111111",
  7293=>"001101111",
  7294=>"100100110",
  7295=>"011011011",
  7296=>"011111111",
  7297=>"111111001",
  7298=>"000100111",
  7299=>"000000001",
  7300=>"111011111",
  7301=>"111011111",
  7302=>"000111111",
  7303=>"000100000",
  7304=>"000000000",
  7305=>"100110111",
  7306=>"000000000",
  7307=>"001001001",
  7308=>"111111111",
  7309=>"111111111",
  7310=>"111111111",
  7311=>"111010000",
  7312=>"001011001",
  7313=>"100110000",
  7314=>"111111111",
  7315=>"111001101",
  7316=>"010011010",
  7317=>"110110000",
  7318=>"011011111",
  7319=>"000000000",
  7320=>"010010010",
  7321=>"000000000",
  7322=>"111111100",
  7323=>"111000000",
  7324=>"111011011",
  7325=>"101100100",
  7326=>"111111111",
  7327=>"100001001",
  7328=>"000000000",
  7329=>"111011000",
  7330=>"111000110",
  7331=>"111111111",
  7332=>"101101001",
  7333=>"111111111",
  7334=>"010110111",
  7335=>"001001111",
  7336=>"111111100",
  7337=>"110111111",
  7338=>"111011011",
  7339=>"001001000",
  7340=>"111001011",
  7341=>"000000000",
  7342=>"111111111",
  7343=>"000110111",
  7344=>"000000000",
  7345=>"001001001",
  7346=>"100000000",
  7347=>"000000000",
  7348=>"100100111",
  7349=>"000000101",
  7350=>"000000000",
  7351=>"101001001",
  7352=>"000000000",
  7353=>"000000000",
  7354=>"100100000",
  7355=>"000000000",
  7356=>"111000000",
  7357=>"000001111",
  7358=>"111011110",
  7359=>"001001000",
  7360=>"110111000",
  7361=>"000000000",
  7362=>"000001001",
  7363=>"000000000",
  7364=>"000000000",
  7365=>"010000000",
  7366=>"000000000",
  7367=>"000000000",
  7368=>"110111010",
  7369=>"000000000",
  7370=>"011111011",
  7371=>"100111111",
  7372=>"000000100",
  7373=>"100111111",
  7374=>"000000000",
  7375=>"111001101",
  7376=>"011111111",
  7377=>"000000000",
  7378=>"111111000",
  7379=>"111111011",
  7380=>"111101001",
  7381=>"001001111",
  7382=>"111011000",
  7383=>"110111011",
  7384=>"001000000",
  7385=>"100100011",
  7386=>"000000000",
  7387=>"101100100",
  7388=>"000100000",
  7389=>"001000111",
  7390=>"000000000",
  7391=>"000000000",
  7392=>"000000000",
  7393=>"011011011",
  7394=>"111111111",
  7395=>"001110100",
  7396=>"111111111",
  7397=>"000000000",
  7398=>"111011001",
  7399=>"000000000",
  7400=>"111111111",
  7401=>"000000000",
  7402=>"111111111",
  7403=>"111011011",
  7404=>"111111111",
  7405=>"111111111",
  7406=>"001000111",
  7407=>"111011011",
  7408=>"111111110",
  7409=>"110011111",
  7410=>"111011001",
  7411=>"111111000",
  7412=>"000000000",
  7413=>"111111100",
  7414=>"000000000",
  7415=>"111111111",
  7416=>"111000010",
  7417=>"000000000",
  7418=>"111111111",
  7419=>"010000000",
  7420=>"000000011",
  7421=>"111111001",
  7422=>"101000000",
  7423=>"100111110",
  7424=>"001000000",
  7425=>"001001001",
  7426=>"111111111",
  7427=>"111101101",
  7428=>"011011000",
  7429=>"111111000",
  7430=>"000000000",
  7431=>"000001000",
  7432=>"000000000",
  7433=>"000000000",
  7434=>"000000000",
  7435=>"001010011",
  7436=>"110000000",
  7437=>"000000000",
  7438=>"111111000",
  7439=>"000011000",
  7440=>"111110111",
  7441=>"111111111",
  7442=>"000000111",
  7443=>"011011100",
  7444=>"000000000",
  7445=>"000000110",
  7446=>"111111111",
  7447=>"111110111",
  7448=>"000000001",
  7449=>"111100111",
  7450=>"000000101",
  7451=>"001011000",
  7452=>"011011001",
  7453=>"111111111",
  7454=>"000000000",
  7455=>"111001110",
  7456=>"101001000",
  7457=>"000000000",
  7458=>"011011001",
  7459=>"111111111",
  7460=>"101111111",
  7461=>"111111100",
  7462=>"100000000",
  7463=>"111111111",
  7464=>"100100100",
  7465=>"111111111",
  7466=>"101011001",
  7467=>"000010111",
  7468=>"111001001",
  7469=>"000000000",
  7470=>"000000000",
  7471=>"000100111",
  7472=>"100111111",
  7473=>"000000000",
  7474=>"111111111",
  7475=>"010000000",
  7476=>"011111000",
  7477=>"111111111",
  7478=>"001011000",
  7479=>"100000010",
  7480=>"000000000",
  7481=>"011011111",
  7482=>"111111111",
  7483=>"000110110",
  7484=>"001001001",
  7485=>"011000111",
  7486=>"111001111",
  7487=>"000000101",
  7488=>"111000001",
  7489=>"111111111",
  7490=>"000000000",
  7491=>"000000000",
  7492=>"000000001",
  7493=>"000001001",
  7494=>"100000000",
  7495=>"110110111",
  7496=>"000111111",
  7497=>"000000000",
  7498=>"000000000",
  7499=>"000110011",
  7500=>"001001000",
  7501=>"010010111",
  7502=>"000010111",
  7503=>"000000100",
  7504=>"010010101",
  7505=>"001000011",
  7506=>"111111111",
  7507=>"111111100",
  7508=>"000000000",
  7509=>"111101111",
  7510=>"010000000",
  7511=>"111111111",
  7512=>"000000001",
  7513=>"000000000",
  7514=>"001001000",
  7515=>"000000000",
  7516=>"111110000",
  7517=>"000000000",
  7518=>"001000111",
  7519=>"001000000",
  7520=>"100100110",
  7521=>"111111111",
  7522=>"000000011",
  7523=>"000000000",
  7524=>"110111011",
  7525=>"000111111",
  7526=>"000100000",
  7527=>"111011000",
  7528=>"000000000",
  7529=>"011111111",
  7530=>"000000000",
  7531=>"101101111",
  7532=>"000000000",
  7533=>"100000000",
  7534=>"111100111",
  7535=>"000001000",
  7536=>"110110000",
  7537=>"011011111",
  7538=>"000000000",
  7539=>"111101100",
  7540=>"111101101",
  7541=>"111100000",
  7542=>"111111111",
  7543=>"000110000",
  7544=>"000000000",
  7545=>"000000000",
  7546=>"001001001",
  7547=>"010110111",
  7548=>"111111011",
  7549=>"000000000",
  7550=>"111111001",
  7551=>"000001000",
  7552=>"000110111",
  7553=>"000110110",
  7554=>"111110110",
  7555=>"000000000",
  7556=>"111111000",
  7557=>"111111111",
  7558=>"111111111",
  7559=>"000000000",
  7560=>"000001000",
  7561=>"100110110",
  7562=>"011011011",
  7563=>"010110111",
  7564=>"000000000",
  7565=>"111111001",
  7566=>"111111111",
  7567=>"111111110",
  7568=>"000011000",
  7569=>"111111111",
  7570=>"111111111",
  7571=>"110110100",
  7572=>"000000000",
  7573=>"111111111",
  7574=>"110110000",
  7575=>"000000111",
  7576=>"111111111",
  7577=>"101101101",
  7578=>"000011011",
  7579=>"000000111",
  7580=>"101000101",
  7581=>"101111111",
  7582=>"101001011",
  7583=>"000000000",
  7584=>"101000001",
  7585=>"110111111",
  7586=>"000110110",
  7587=>"011001000",
  7588=>"010010000",
  7589=>"011111111",
  7590=>"000110000",
  7591=>"111111111",
  7592=>"111110000",
  7593=>"000000001",
  7594=>"111111111",
  7595=>"111111011",
  7596=>"000000000",
  7597=>"111111001",
  7598=>"101001001",
  7599=>"001000000",
  7600=>"111011000",
  7601=>"000000000",
  7602=>"000000000",
  7603=>"001011111",
  7604=>"111000000",
  7605=>"000000011",
  7606=>"000000000",
  7607=>"000011001",
  7608=>"111011000",
  7609=>"111111101",
  7610=>"110100001",
  7611=>"011001000",
  7612=>"000000000",
  7613=>"111000000",
  7614=>"011011000",
  7615=>"000001001",
  7616=>"101111110",
  7617=>"000000000",
  7618=>"011111011",
  7619=>"000000000",
  7620=>"000010110",
  7621=>"100001001",
  7622=>"000000000",
  7623=>"111111111",
  7624=>"111110100",
  7625=>"010000100",
  7626=>"000001111",
  7627=>"110111111",
  7628=>"110101111",
  7629=>"111111111",
  7630=>"000010000",
  7631=>"111111100",
  7632=>"011000000",
  7633=>"000000000",
  7634=>"000000001",
  7635=>"111000001",
  7636=>"110110100",
  7637=>"000010011",
  7638=>"011001001",
  7639=>"110001011",
  7640=>"001000000",
  7641=>"000000001",
  7642=>"100000100",
  7643=>"111111111",
  7644=>"111111111",
  7645=>"100000000",
  7646=>"000000000",
  7647=>"100111011",
  7648=>"000000000",
  7649=>"111111111",
  7650=>"000000100",
  7651=>"000010010",
  7652=>"000000000",
  7653=>"100111101",
  7654=>"000100000",
  7655=>"000000000",
  7656=>"011111111",
  7657=>"101001000",
  7658=>"110110100",
  7659=>"111111111",
  7660=>"000000000",
  7661=>"111000001",
  7662=>"000000000",
  7663=>"111110110",
  7664=>"111111111",
  7665=>"110110111",
  7666=>"001011011",
  7667=>"000000000",
  7668=>"111111111",
  7669=>"001001101",
  7670=>"110111111",
  7671=>"001101101",
  7672=>"111111011",
  7673=>"010110100",
  7674=>"100110000",
  7675=>"111010111",
  7676=>"101101100",
  7677=>"000000000",
  7678=>"111000000",
  7679=>"000000000",
  7680=>"111111110",
  7681=>"110111011",
  7682=>"101100000",
  7683=>"111111111",
  7684=>"111011110",
  7685=>"101101101",
  7686=>"100100011",
  7687=>"000000000",
  7688=>"000100000",
  7689=>"111110000",
  7690=>"111111111",
  7691=>"000000000",
  7692=>"000100100",
  7693=>"111111000",
  7694=>"111111111",
  7695=>"000001000",
  7696=>"000100111",
  7697=>"111110010",
  7698=>"000000000",
  7699=>"110110000",
  7700=>"111111111",
  7701=>"000000000",
  7702=>"100000000",
  7703=>"011000000",
  7704=>"000000111",
  7705=>"000100100",
  7706=>"000000000",
  7707=>"100000000",
  7708=>"100111011",
  7709=>"000000000",
  7710=>"011011010",
  7711=>"111111111",
  7712=>"111101000",
  7713=>"000000000",
  7714=>"100100000",
  7715=>"111111110",
  7716=>"111111111",
  7717=>"111011001",
  7718=>"000000000",
  7719=>"000001000",
  7720=>"111111111",
  7721=>"110010010",
  7722=>"000011011",
  7723=>"111001001",
  7724=>"001000000",
  7725=>"111110000",
  7726=>"000000000",
  7727=>"111111111",
  7728=>"000000000",
  7729=>"000000100",
  7730=>"000000000",
  7731=>"100000000",
  7732=>"011000000",
  7733=>"111011111",
  7734=>"001000110",
  7735=>"000111111",
  7736=>"111111111",
  7737=>"000000010",
  7738=>"000000111",
  7739=>"111110010",
  7740=>"000000000",
  7741=>"111111101",
  7742=>"100111111",
  7743=>"011001000",
  7744=>"001001111",
  7745=>"111001001",
  7746=>"000111111",
  7747=>"100100111",
  7748=>"100000000",
  7749=>"000000111",
  7750=>"000000000",
  7751=>"101100000",
  7752=>"001101110",
  7753=>"111000000",
  7754=>"100100111",
  7755=>"111111101",
  7756=>"111111111",
  7757=>"000000000",
  7758=>"000000000",
  7759=>"111110110",
  7760=>"000000000",
  7761=>"111111000",
  7762=>"001111111",
  7763=>"111110111",
  7764=>"000000000",
  7765=>"111010110",
  7766=>"111111111",
  7767=>"111111100",
  7768=>"001011011",
  7769=>"100000000",
  7770=>"101111111",
  7771=>"011001101",
  7772=>"111111111",
  7773=>"000011000",
  7774=>"000000000",
  7775=>"111111111",
  7776=>"111111111",
  7777=>"111111111",
  7778=>"001111111",
  7779=>"111100111",
  7780=>"011011111",
  7781=>"000000000",
  7782=>"111111111",
  7783=>"111111111",
  7784=>"000001001",
  7785=>"000000000",
  7786=>"111000110",
  7787=>"110111111",
  7788=>"111111111",
  7789=>"000001111",
  7790=>"000000000",
  7791=>"111111000",
  7792=>"000000000",
  7793=>"010010000",
  7794=>"111011111",
  7795=>"001001001",
  7796=>"001011111",
  7797=>"101111001",
  7798=>"000000000",
  7799=>"100111111",
  7800=>"000000000",
  7801=>"000000100",
  7802=>"110111000",
  7803=>"000000000",
  7804=>"001001000",
  7805=>"111111110",
  7806=>"100100100",
  7807=>"001000000",
  7808=>"110111111",
  7809=>"000101101",
  7810=>"111111000",
  7811=>"100000110",
  7812=>"101101001",
  7813=>"000000000",
  7814=>"001000000",
  7815=>"000010011",
  7816=>"111111100",
  7817=>"000001111",
  7818=>"000000000",
  7819=>"000000011",
  7820=>"100111000",
  7821=>"001000100",
  7822=>"100111111",
  7823=>"011011111",
  7824=>"111111000",
  7825=>"111111111",
  7826=>"001001001",
  7827=>"100111111",
  7828=>"000011000",
  7829=>"000001000",
  7830=>"011000000",
  7831=>"111111000",
  7832=>"111111111",
  7833=>"100111111",
  7834=>"111011000",
  7835=>"010011011",
  7836=>"000001001",
  7837=>"111000000",
  7838=>"111111000",
  7839=>"111001000",
  7840=>"101000000",
  7841=>"101001111",
  7842=>"000000000",
  7843=>"000000110",
  7844=>"111100110",
  7845=>"000010111",
  7846=>"111111111",
  7847=>"110110100",
  7848=>"000000001",
  7849=>"000000000",
  7850=>"111111000",
  7851=>"000000000",
  7852=>"111111111",
  7853=>"111111111",
  7854=>"111111111",
  7855=>"101000000",
  7856=>"000110111",
  7857=>"001101000",
  7858=>"010111111",
  7859=>"111100000",
  7860=>"111101111",
  7861=>"000000000",
  7862=>"111111111",
  7863=>"000100000",
  7864=>"101100000",
  7865=>"111111000",
  7866=>"000000000",
  7867=>"000000001",
  7868=>"111111100",
  7869=>"111111111",
  7870=>"000000000",
  7871=>"000001000",
  7872=>"110111111",
  7873=>"111111111",
  7874=>"111111000",
  7875=>"101100100",
  7876=>"000000000",
  7877=>"111111000",
  7878=>"100000011",
  7879=>"001101001",
  7880=>"001101000",
  7881=>"000100000",
  7882=>"000000100",
  7883=>"110110000",
  7884=>"000000010",
  7885=>"000110111",
  7886=>"110110100",
  7887=>"111111100",
  7888=>"111111101",
  7889=>"001000000",
  7890=>"000111111",
  7891=>"111111111",
  7892=>"000000000",
  7893=>"000000000",
  7894=>"111011111",
  7895=>"000000011",
  7896=>"000000000",
  7897=>"001111111",
  7898=>"000000000",
  7899=>"000000000",
  7900=>"001000111",
  7901=>"100000100",
  7902=>"100110111",
  7903=>"001101100",
  7904=>"011011011",
  7905=>"111000000",
  7906=>"000000000",
  7907=>"000000000",
  7908=>"100000100",
  7909=>"100110111",
  7910=>"111111100",
  7911=>"000111101",
  7912=>"100100111",
  7913=>"111111111",
  7914=>"001001010",
  7915=>"100000000",
  7916=>"011111111",
  7917=>"111111101",
  7918=>"111111000",
  7919=>"000000000",
  7920=>"000000110",
  7921=>"000000000",
  7922=>"000000000",
  7923=>"011011010",
  7924=>"000010111",
  7925=>"011111111",
  7926=>"011100001",
  7927=>"101101111",
  7928=>"000000000",
  7929=>"111111111",
  7930=>"000011110",
  7931=>"000000000",
  7932=>"110110110",
  7933=>"011011011",
  7934=>"000101100",
  7935=>"000100111",
  7936=>"000000000",
  7937=>"000000000",
  7938=>"000000000",
  7939=>"001000000",
  7940=>"000000000",
  7941=>"101111111",
  7942=>"111111111",
  7943=>"111111101",
  7944=>"110111110",
  7945=>"000000000",
  7946=>"000000000",
  7947=>"001111111",
  7948=>"111110111",
  7949=>"000000000",
  7950=>"000000000",
  7951=>"111111111",
  7952=>"110111111",
  7953=>"000000001",
  7954=>"001000000",
  7955=>"010000000",
  7956=>"111111101",
  7957=>"000000000",
  7958=>"111110000",
  7959=>"111110100",
  7960=>"111111111",
  7961=>"111111111",
  7962=>"111000000",
  7963=>"110111111",
  7964=>"110100000",
  7965=>"000000111",
  7966=>"001110110",
  7967=>"110000000",
  7968=>"111110111",
  7969=>"011010000",
  7970=>"000000100",
  7971=>"111100100",
  7972=>"000010011",
  7973=>"000000000",
  7974=>"111111111",
  7975=>"111111111",
  7976=>"000000000",
  7977=>"001000000",
  7978=>"000011011",
  7979=>"111001001",
  7980=>"000000100",
  7981=>"000000000",
  7982=>"000000000",
  7983=>"000111111",
  7984=>"111110111",
  7985=>"000000000",
  7986=>"111111110",
  7987=>"000000000",
  7988=>"000000000",
  7989=>"001000000",
  7990=>"000000000",
  7991=>"000000000",
  7992=>"111111000",
  7993=>"111111111",
  7994=>"111111101",
  7995=>"111111111",
  7996=>"000111100",
  7997=>"001001111",
  7998=>"000111111",
  7999=>"100111111",
  8000=>"000000000",
  8001=>"101101111",
  8002=>"011011111",
  8003=>"111111111",
  8004=>"011011000",
  8005=>"100111001",
  8006=>"111011011",
  8007=>"001000000",
  8008=>"000000000",
  8009=>"111111111",
  8010=>"111111011",
  8011=>"111100000",
  8012=>"100101111",
  8013=>"100000111",
  8014=>"000001111",
  8015=>"110000010",
  8016=>"110110000",
  8017=>"101001100",
  8018=>"111000000",
  8019=>"111000000",
  8020=>"111111111",
  8021=>"110000001",
  8022=>"000000000",
  8023=>"000000000",
  8024=>"000000000",
  8025=>"010000000",
  8026=>"111111011",
  8027=>"000001111",
  8028=>"000000000",
  8029=>"011111111",
  8030=>"000000000",
  8031=>"111100100",
  8032=>"000010000",
  8033=>"000000011",
  8034=>"111100000",
  8035=>"000000000",
  8036=>"111111111",
  8037=>"000000010",
  8038=>"111000101",
  8039=>"011001001",
  8040=>"000000000",
  8041=>"111111111",
  8042=>"110000000",
  8043=>"000110110",
  8044=>"011011111",
  8045=>"100110111",
  8046=>"111111100",
  8047=>"000100111",
  8048=>"101111011",
  8049=>"000000000",
  8050=>"111000000",
  8051=>"111110111",
  8052=>"111110110",
  8053=>"111011111",
  8054=>"000000000",
  8055=>"100101001",
  8056=>"110110110",
  8057=>"011111010",
  8058=>"100000000",
  8059=>"011111111",
  8060=>"101101001",
  8061=>"111000000",
  8062=>"000000001",
  8063=>"000000000",
  8064=>"001001001",
  8065=>"101011000",
  8066=>"000000101",
  8067=>"000000000",
  8068=>"000000111",
  8069=>"000000000",
  8070=>"000001001",
  8071=>"111111111",
  8072=>"111111011",
  8073=>"000111111",
  8074=>"101001000",
  8075=>"000011011",
  8076=>"111000000",
  8077=>"011111111",
  8078=>"010110110",
  8079=>"111100111",
  8080=>"000000000",
  8081=>"111111111",
  8082=>"111000000",
  8083=>"000101000",
  8084=>"000000000",
  8085=>"000001001",
  8086=>"111111100",
  8087=>"111111111",
  8088=>"111011111",
  8089=>"111111111",
  8090=>"111111010",
  8091=>"000000000",
  8092=>"100110111",
  8093=>"111111000",
  8094=>"000000111",
  8095=>"100101000",
  8096=>"000000000",
  8097=>"011011001",
  8098=>"011111111",
  8099=>"110110110",
  8100=>"000000000",
  8101=>"000000000",
  8102=>"000111000",
  8103=>"111110010",
  8104=>"010000000",
  8105=>"000000101",
  8106=>"111100000",
  8107=>"000000000",
  8108=>"000000000",
  8109=>"111111011",
  8110=>"000100101",
  8111=>"000111111",
  8112=>"110111111",
  8113=>"000000000",
  8114=>"111111111",
  8115=>"000000000",
  8116=>"000000000",
  8117=>"001000100",
  8118=>"111111111",
  8119=>"110000000",
  8120=>"000000100",
  8121=>"111111111",
  8122=>"001011011",
  8123=>"001011011",
  8124=>"111110000",
  8125=>"011011111",
  8126=>"011000000",
  8127=>"001001000",
  8128=>"011011111",
  8129=>"000000000",
  8130=>"111111111",
  8131=>"111111111",
  8132=>"111110000",
  8133=>"000000000",
  8134=>"111011000",
  8135=>"111111000",
  8136=>"000000000",
  8137=>"110000000",
  8138=>"000000000",
  8139=>"000111011",
  8140=>"111010111",
  8141=>"000000000",
  8142=>"111000000",
  8143=>"000000111",
  8144=>"000110110",
  8145=>"000000000",
  8146=>"000000000",
  8147=>"111001000",
  8148=>"011111111",
  8149=>"000100101",
  8150=>"001000011",
  8151=>"001001000",
  8152=>"000010110",
  8153=>"111111100",
  8154=>"111111111",
  8155=>"111111100",
  8156=>"011111011",
  8157=>"000111111",
  8158=>"000000000",
  8159=>"111110111",
  8160=>"111111111",
  8161=>"111111111",
  8162=>"011011000",
  8163=>"000010111",
  8164=>"111010000",
  8165=>"111111111",
  8166=>"000000111",
  8167=>"000000010",
  8168=>"000101111",
  8169=>"100110001",
  8170=>"010000000",
  8171=>"100100000",
  8172=>"100111111",
  8173=>"111111111",
  8174=>"111111111",
  8175=>"111111111",
  8176=>"100111111",
  8177=>"010111111",
  8178=>"000110100",
  8179=>"111111110",
  8180=>"000111111",
  8181=>"000000000",
  8182=>"000000111",
  8183=>"000000000",
  8184=>"000100110",
  8185=>"000000001",
  8186=>"111111111",
  8187=>"100000010",
  8188=>"100111011",
  8189=>"000000000",
  8190=>"011000001",
  8191=>"000001000",
  8192=>"100100110",
  8193=>"111110000",
  8194=>"000000111",
  8195=>"000111111",
  8196=>"000000001",
  8197=>"000000111",
  8198=>"000001001",
  8199=>"111111111",
  8200=>"001000000",
  8201=>"000000001",
  8202=>"000000011",
  8203=>"001111100",
  8204=>"111111111",
  8205=>"111111111",
  8206=>"000000100",
  8207=>"111111111",
  8208=>"111111000",
  8209=>"010010000",
  8210=>"001000111",
  8211=>"111111000",
  8212=>"000000111",
  8213=>"001000000",
  8214=>"111110000",
  8215=>"110101101",
  8216=>"000100100",
  8217=>"111011000",
  8218=>"111111111",
  8219=>"111101111",
  8220=>"000100111",
  8221=>"000000011",
  8222=>"111111111",
  8223=>"000000000",
  8224=>"010111111",
  8225=>"111000000",
  8226=>"000000111",
  8227=>"111111111",
  8228=>"000000111",
  8229=>"111101000",
  8230=>"111011011",
  8231=>"000001111",
  8232=>"111111111",
  8233=>"111001111",
  8234=>"000000111",
  8235=>"000101000",
  8236=>"111111000",
  8237=>"000101000",
  8238=>"000000010",
  8239=>"111000000",
  8240=>"000000010",
  8241=>"111111000",
  8242=>"000100110",
  8243=>"111111110",
  8244=>"000110100",
  8245=>"111111000",
  8246=>"100111111",
  8247=>"000111111",
  8248=>"000001111",
  8249=>"000000111",
  8250=>"000011010",
  8251=>"111111000",
  8252=>"000100111",
  8253=>"111000000",
  8254=>"110111111",
  8255=>"000111111",
  8256=>"011000000",
  8257=>"000100111",
  8258=>"001011010",
  8259=>"000011111",
  8260=>"000001111",
  8261=>"111001000",
  8262=>"111000000",
  8263=>"000110111",
  8264=>"000000011",
  8265=>"000000000",
  8266=>"000111000",
  8267=>"010110110",
  8268=>"110110000",
  8269=>"111001001",
  8270=>"111000000",
  8271=>"000000111",
  8272=>"000110011",
  8273=>"111111000",
  8274=>"111110000",
  8275=>"100100111",
  8276=>"000000000",
  8277=>"001000000",
  8278=>"111111111",
  8279=>"000010111",
  8280=>"001000100",
  8281=>"000000100",
  8282=>"000000011",
  8283=>"111110110",
  8284=>"010000000",
  8285=>"111111010",
  8286=>"000000000",
  8287=>"000000111",
  8288=>"110100110",
  8289=>"000000010",
  8290=>"000000000",
  8291=>"110100000",
  8292=>"010110000",
  8293=>"000000100",
  8294=>"000000111",
  8295=>"111011111",
  8296=>"111000000",
  8297=>"000000000",
  8298=>"011001000",
  8299=>"111111011",
  8300=>"010111110",
  8301=>"000000111",
  8302=>"110110111",
  8303=>"111000001",
  8304=>"111110010",
  8305=>"100111111",
  8306=>"001100110",
  8307=>"110001111",
  8308=>"111000000",
  8309=>"000101111",
  8310=>"111000111",
  8311=>"110111010",
  8312=>"000011111",
  8313=>"000000000",
  8314=>"000000000",
  8315=>"000000111",
  8316=>"000010111",
  8317=>"001111111",
  8318=>"001101000",
  8319=>"011001000",
  8320=>"000000000",
  8321=>"111111111",
  8322=>"111000000",
  8323=>"011000000",
  8324=>"000111111",
  8325=>"111000000",
  8326=>"000111100",
  8327=>"000000100",
  8328=>"111111000",
  8329=>"010000100",
  8330=>"000000000",
  8331=>"111111000",
  8332=>"000000111",
  8333=>"111001000",
  8334=>"111111000",
  8335=>"000111000",
  8336=>"000000000",
  8337=>"000000000",
  8338=>"000000111",
  8339=>"110111110",
  8340=>"000000000",
  8341=>"101000000",
  8342=>"111111001",
  8343=>"000000111",
  8344=>"000001001",
  8345=>"111000000",
  8346=>"111101110",
  8347=>"000100100",
  8348=>"000001101",
  8349=>"000000000",
  8350=>"111111101",
  8351=>"111111100",
  8352=>"111111111",
  8353=>"111111111",
  8354=>"111000000",
  8355=>"000111111",
  8356=>"000000000",
  8357=>"001000101",
  8358=>"111111111",
  8359=>"111000011",
  8360=>"000111111",
  8361=>"111111011",
  8362=>"001111001",
  8363=>"111100110",
  8364=>"111010000",
  8365=>"000000000",
  8366=>"101001001",
  8367=>"000010000",
  8368=>"000000100",
  8369=>"111010000",
  8370=>"111111110",
  8371=>"010000000",
  8372=>"110111010",
  8373=>"001111001",
  8374=>"000000000",
  8375=>"111111111",
  8376=>"000000000",
  8377=>"000000110",
  8378=>"000000000",
  8379=>"001000000",
  8380=>"000000111",
  8381=>"011011010",
  8382=>"100111000",
  8383=>"001101111",
  8384=>"000000000",
  8385=>"000000000",
  8386=>"000001011",
  8387=>"111101000",
  8388=>"111111111",
  8389=>"000000111",
  8390=>"000000010",
  8391=>"000111111",
  8392=>"110010000",
  8393=>"000101111",
  8394=>"000000000",
  8395=>"011001000",
  8396=>"000000111",
  8397=>"101111111",
  8398=>"010111111",
  8399=>"111111010",
  8400=>"111011110",
  8401=>"000000110",
  8402=>"000000000",
  8403=>"000000111",
  8404=>"000100010",
  8405=>"111111000",
  8406=>"000000110",
  8407=>"000111111",
  8408=>"000000100",
  8409=>"111111000",
  8410=>"000000101",
  8411=>"111110100",
  8412=>"111111001",
  8413=>"111111111",
  8414=>"111111110",
  8415=>"111111111",
  8416=>"000000100",
  8417=>"000111111",
  8418=>"011001111",
  8419=>"111111010",
  8420=>"101111000",
  8421=>"111111111",
  8422=>"111111000",
  8423=>"000111001",
  8424=>"111111000",
  8425=>"111100000",
  8426=>"101111111",
  8427=>"111111111",
  8428=>"111111111",
  8429=>"000000101",
  8430=>"111011000",
  8431=>"001000000",
  8432=>"100110100",
  8433=>"101100001",
  8434=>"001001101",
  8435=>"000000001",
  8436=>"011111000",
  8437=>"000000111",
  8438=>"110100000",
  8439=>"000000111",
  8440=>"111110100",
  8441=>"110110000",
  8442=>"001001000",
  8443=>"011010000",
  8444=>"111111001",
  8445=>"000000000",
  8446=>"011000000",
  8447=>"111001000",
  8448=>"000000111",
  8449=>"110111111",
  8450=>"000110111",
  8451=>"011111000",
  8452=>"111111100",
  8453=>"000000000",
  8454=>"000000111",
  8455=>"011111000",
  8456=>"000000001",
  8457=>"011000000",
  8458=>"000000001",
  8459=>"000000000",
  8460=>"110110000",
  8461=>"111111110",
  8462=>"010110000",
  8463=>"000110110",
  8464=>"101000000",
  8465=>"000000101",
  8466=>"000000000",
  8467=>"000000111",
  8468=>"110111111",
  8469=>"000100111",
  8470=>"000110111",
  8471=>"000000011",
  8472=>"110000000",
  8473=>"000000000",
  8474=>"111000000",
  8475=>"000000010",
  8476=>"000000100",
  8477=>"101111111",
  8478=>"000111111",
  8479=>"111000000",
  8480=>"000111111",
  8481=>"000000101",
  8482=>"000000111",
  8483=>"111111000",
  8484=>"000111111",
  8485=>"100000000",
  8486=>"111111111",
  8487=>"000011111",
  8488=>"000000000",
  8489=>"000111011",
  8490=>"000001111",
  8491=>"111000000",
  8492=>"000000001",
  8493=>"000111111",
  8494=>"101000000",
  8495=>"110000110",
  8496=>"011010011",
  8497=>"000000000",
  8498=>"111111111",
  8499=>"010000101",
  8500=>"111000000",
  8501=>"010111110",
  8502=>"111000000",
  8503=>"000011111",
  8504=>"000001000",
  8505=>"111110111",
  8506=>"100000111",
  8507=>"111111000",
  8508=>"000111111",
  8509=>"011111110",
  8510=>"111111000",
  8511=>"111000000",
  8512=>"000001111",
  8513=>"110010100",
  8514=>"001000111",
  8515=>"000100111",
  8516=>"001000000",
  8517=>"111111001",
  8518=>"000010111",
  8519=>"110110000",
  8520=>"110010111",
  8521=>"000000000",
  8522=>"111000000",
  8523=>"000000111",
  8524=>"110111111",
  8525=>"111111111",
  8526=>"001111111",
  8527=>"000000011",
  8528=>"001001110",
  8529=>"000000111",
  8530=>"000000111",
  8531=>"111101000",
  8532=>"111111000",
  8533=>"001111111",
  8534=>"011010000",
  8535=>"111000000",
  8536=>"111111111",
  8537=>"000000000",
  8538=>"111010010",
  8539=>"000100100",
  8540=>"001001111",
  8541=>"000000000",
  8542=>"111010000",
  8543=>"111111011",
  8544=>"000001001",
  8545=>"111010110",
  8546=>"100111110",
  8547=>"110111110",
  8548=>"111111110",
  8549=>"000111111",
  8550=>"000000000",
  8551=>"000000111",
  8552=>"100100110",
  8553=>"000000000",
  8554=>"000000000",
  8555=>"111111001",
  8556=>"101000001",
  8557=>"011111111",
  8558=>"110000000",
  8559=>"000000000",
  8560=>"111011110",
  8561=>"111010000",
  8562=>"000111111",
  8563=>"001000000",
  8564=>"000111000",
  8565=>"100100111",
  8566=>"000000100",
  8567=>"111111101",
  8568=>"100000001",
  8569=>"111111111",
  8570=>"000000000",
  8571=>"111101111",
  8572=>"000001000",
  8573=>"110000000",
  8574=>"111111000",
  8575=>"111111000",
  8576=>"110110000",
  8577=>"001000000",
  8578=>"111000000",
  8579=>"000111111",
  8580=>"011000110",
  8581=>"011011001",
  8582=>"000100010",
  8583=>"110110111",
  8584=>"000000000",
  8585=>"111111111",
  8586=>"000000000",
  8587=>"000000100",
  8588=>"110000111",
  8589=>"111111111",
  8590=>"000000000",
  8591=>"111000000",
  8592=>"000000110",
  8593=>"100111111",
  8594=>"000001111",
  8595=>"110111011",
  8596=>"000000000",
  8597=>"000000000",
  8598=>"100111011",
  8599=>"111111100",
  8600=>"011000000",
  8601=>"111111010",
  8602=>"111001000",
  8603=>"100000000",
  8604=>"000011011",
  8605=>"100000011",
  8606=>"000000000",
  8607=>"000000111",
  8608=>"111111000",
  8609=>"110100110",
  8610=>"111111101",
  8611=>"011111011",
  8612=>"100111100",
  8613=>"001110000",
  8614=>"000000000",
  8615=>"111010000",
  8616=>"000100110",
  8617=>"000000111",
  8618=>"100110111",
  8619=>"100110110",
  8620=>"000000101",
  8621=>"111111000",
  8622=>"111101000",
  8623=>"111000011",
  8624=>"000000111",
  8625=>"111111111",
  8626=>"001111111",
  8627=>"111111011",
  8628=>"000010110",
  8629=>"111100000",
  8630=>"111111111",
  8631=>"110100000",
  8632=>"111100000",
  8633=>"000000000",
  8634=>"111111000",
  8635=>"000111011",
  8636=>"111111111",
  8637=>"111111000",
  8638=>"111000000",
  8639=>"000000111",
  8640=>"000111000",
  8641=>"110000111",
  8642=>"011000010",
  8643=>"000000000",
  8644=>"011111111",
  8645=>"000010100",
  8646=>"111011111",
  8647=>"011011000",
  8648=>"001000100",
  8649=>"111000000",
  8650=>"000000111",
  8651=>"000000000",
  8652=>"000000000",
  8653=>"000000000",
  8654=>"000100100",
  8655=>"000101001",
  8656=>"110100000",
  8657=>"000100111",
  8658=>"111111001",
  8659=>"000000111",
  8660=>"101111111",
  8661=>"011111011",
  8662=>"000011111",
  8663=>"110000111",
  8664=>"000000100",
  8665=>"011000000",
  8666=>"000110111",
  8667=>"101000000",
  8668=>"111001000",
  8669=>"011111010",
  8670=>"000011000",
  8671=>"100000011",
  8672=>"000010111",
  8673=>"000000000",
  8674=>"111000000",
  8675=>"111111111",
  8676=>"000011111",
  8677=>"000101100",
  8678=>"000111000",
  8679=>"000000000",
  8680=>"000100111",
  8681=>"111111000",
  8682=>"100100000",
  8683=>"000000011",
  8684=>"111111111",
  8685=>"111000100",
  8686=>"001111000",
  8687=>"000000000",
  8688=>"000010000",
  8689=>"111001111",
  8690=>"101100111",
  8691=>"000000110",
  8692=>"100100000",
  8693=>"000100000",
  8694=>"110110110",
  8695=>"000111111",
  8696=>"000100111",
  8697=>"000000110",
  8698=>"111010110",
  8699=>"000000000",
  8700=>"000000111",
  8701=>"101101111",
  8702=>"111111000",
  8703=>"000000111",
  8704=>"111111110",
  8705=>"011011000",
  8706=>"111011001",
  8707=>"111110010",
  8708=>"110111110",
  8709=>"111000000",
  8710=>"111101101",
  8711=>"111111111",
  8712=>"111000001",
  8713=>"100101001",
  8714=>"000000000",
  8715=>"111101011",
  8716=>"110100000",
  8717=>"000111111",
  8718=>"000000000",
  8719=>"001000000",
  8720=>"000010000",
  8721=>"111100000",
  8722=>"111111001",
  8723=>"000000000",
  8724=>"000000000",
  8725=>"011011111",
  8726=>"111111111",
  8727=>"111011001",
  8728=>"110110110",
  8729=>"110100000",
  8730=>"101001000",
  8731=>"111100000",
  8732=>"111100100",
  8733=>"111111111",
  8734=>"100111001",
  8735=>"000000111",
  8736=>"111111111",
  8737=>"111000111",
  8738=>"001111100",
  8739=>"101111011",
  8740=>"111111110",
  8741=>"000010010",
  8742=>"111110111",
  8743=>"110100100",
  8744=>"111111000",
  8745=>"111111000",
  8746=>"111111111",
  8747=>"111111111",
  8748=>"101111110",
  8749=>"110000000",
  8750=>"001100000",
  8751=>"100000000",
  8752=>"000000000",
  8753=>"111111111",
  8754=>"001000000",
  8755=>"000000001",
  8756=>"000000000",
  8757=>"111111001",
  8758=>"111111111",
  8759=>"011111011",
  8760=>"011101100",
  8761=>"000000100",
  8762=>"000000000",
  8763=>"000111111",
  8764=>"111101111",
  8765=>"000000000",
  8766=>"001000111",
  8767=>"111111110",
  8768=>"000001001",
  8769=>"000000011",
  8770=>"000000100",
  8771=>"101100110",
  8772=>"000000111",
  8773=>"001000000",
  8774=>"111011010",
  8775=>"111111111",
  8776=>"001000001",
  8777=>"000000000",
  8778=>"000000110",
  8779=>"001000111",
  8780=>"000000000",
  8781=>"011111111",
  8782=>"111000011",
  8783=>"000000000",
  8784=>"110111110",
  8785=>"101101101",
  8786=>"000000000",
  8787=>"111111111",
  8788=>"000000000",
  8789=>"011100111",
  8790=>"001000100",
  8791=>"001001001",
  8792=>"001111111",
  8793=>"000000000",
  8794=>"000000111",
  8795=>"001011001",
  8796=>"111111111",
  8797=>"000000000",
  8798=>"111000000",
  8799=>"001010010",
  8800=>"110111111",
  8801=>"000000000",
  8802=>"111000000",
  8803=>"111111111",
  8804=>"100000000",
  8805=>"001111111",
  8806=>"010010000",
  8807=>"111111111",
  8808=>"000000000",
  8809=>"001000000",
  8810=>"111111010",
  8811=>"000000101",
  8812=>"000011001",
  8813=>"111111111",
  8814=>"000000000",
  8815=>"000001000",
  8816=>"101111111",
  8817=>"000000110",
  8818=>"000000000",
  8819=>"110100110",
  8820=>"000000110",
  8821=>"111111111",
  8822=>"111111111",
  8823=>"000000000",
  8824=>"000100100",
  8825=>"111100110",
  8826=>"111000001",
  8827=>"111111111",
  8828=>"110111000",
  8829=>"111111111",
  8830=>"111111001",
  8831=>"000000000",
  8832=>"001000000",
  8833=>"101111111",
  8834=>"011010000",
  8835=>"111111111",
  8836=>"101111111",
  8837=>"000000111",
  8838=>"010010000",
  8839=>"000000000",
  8840=>"110100101",
  8841=>"000111111",
  8842=>"101100100",
  8843=>"111110001",
  8844=>"001000100",
  8845=>"000000000",
  8846=>"111111000",
  8847=>"000000000",
  8848=>"111111111",
  8849=>"111010111",
  8850=>"011011000",
  8851=>"000000100",
  8852=>"111111010",
  8853=>"000000000",
  8854=>"000000000",
  8855=>"000000000",
  8856=>"000000000",
  8857=>"111111111",
  8858=>"000100000",
  8859=>"000000110",
  8860=>"111111111",
  8861=>"000000000",
  8862=>"111111111",
  8863=>"000000000",
  8864=>"000111111",
  8865=>"000000000",
  8866=>"111111111",
  8867=>"000000000",
  8868=>"111101001",
  8869=>"111010100",
  8870=>"111111111",
  8871=>"111111111",
  8872=>"000000000",
  8873=>"111111111",
  8874=>"111111111",
  8875=>"000000000",
  8876=>"000000000",
  8877=>"001001001",
  8878=>"000000000",
  8879=>"000000110",
  8880=>"000111101",
  8881=>"111001000",
  8882=>"101100100",
  8883=>"111111010",
  8884=>"000000000",
  8885=>"000111111",
  8886=>"000000000",
  8887=>"111110111",
  8888=>"000111111",
  8889=>"000000111",
  8890=>"001100100",
  8891=>"101001101",
  8892=>"000000000",
  8893=>"111100111",
  8894=>"111111111",
  8895=>"011011111",
  8896=>"111111110",
  8897=>"111111000",
  8898=>"110000000",
  8899=>"111111111",
  8900=>"000000000",
  8901=>"000000000",
  8902=>"111000000",
  8903=>"000000000",
  8904=>"111111011",
  8905=>"100000000",
  8906=>"011001111",
  8907=>"101111111",
  8908=>"000000000",
  8909=>"000111011",
  8910=>"000000000",
  8911=>"111000000",
  8912=>"111111110",
  8913=>"111011111",
  8914=>"111111111",
  8915=>"111010010",
  8916=>"111111100",
  8917=>"001001111",
  8918=>"000001000",
  8919=>"000010111",
  8920=>"101111000",
  8921=>"011111011",
  8922=>"000000000",
  8923=>"000000000",
  8924=>"111111111",
  8925=>"111111111",
  8926=>"110111110",
  8927=>"111111110",
  8928=>"000000000",
  8929=>"000000000",
  8930=>"000000100",
  8931=>"111111111",
  8932=>"011111111",
  8933=>"100010110",
  8934=>"000000000",
  8935=>"111111001",
  8936=>"000000000",
  8937=>"101100110",
  8938=>"111111111",
  8939=>"001001000",
  8940=>"110111111",
  8941=>"000110000",
  8942=>"110000001",
  8943=>"111001111",
  8944=>"000111000",
  8945=>"000000100",
  8946=>"111111101",
  8947=>"110000000",
  8948=>"011011100",
  8949=>"000000100",
  8950=>"110100100",
  8951=>"111111111",
  8952=>"111111111",
  8953=>"000000000",
  8954=>"111111111",
  8955=>"000000000",
  8956=>"110110110",
  8957=>"100100000",
  8958=>"111000000",
  8959=>"011011111",
  8960=>"111111000",
  8961=>"000100100",
  8962=>"111111111",
  8963=>"111111111",
  8964=>"111111100",
  8965=>"111001000",
  8966=>"000100111",
  8967=>"110110110",
  8968=>"111111111",
  8969=>"000000000",
  8970=>"001001010",
  8971=>"000011111",
  8972=>"000000000",
  8973=>"000000000",
  8974=>"111111111",
  8975=>"000000000",
  8976=>"000010000",
  8977=>"001111111",
  8978=>"000000000",
  8979=>"000111111",
  8980=>"000000001",
  8981=>"000000100",
  8982=>"011010110",
  8983=>"000000000",
  8984=>"000000000",
  8985=>"111111111",
  8986=>"111000000",
  8987=>"000110111",
  8988=>"110100000",
  8989=>"000010111",
  8990=>"111111111",
  8991=>"111111111",
  8992=>"011011111",
  8993=>"110111111",
  8994=>"111111111",
  8995=>"010111011",
  8996=>"011001000",
  8997=>"111111001",
  8998=>"011001001",
  8999=>"000000000",
  9000=>"101101000",
  9001=>"000000000",
  9002=>"111011000",
  9003=>"011000000",
  9004=>"101000000",
  9005=>"110110100",
  9006=>"111000111",
  9007=>"101000000",
  9008=>"110110111",
  9009=>"000000000",
  9010=>"001000000",
  9011=>"000000101",
  9012=>"000000101",
  9013=>"000000111",
  9014=>"001000000",
  9015=>"111111111",
  9016=>"000000000",
  9017=>"011011111",
  9018=>"001001000",
  9019=>"111111001",
  9020=>"000000100",
  9021=>"000000111",
  9022=>"000000000",
  9023=>"111111111",
  9024=>"111111111",
  9025=>"111110000",
  9026=>"000000000",
  9027=>"000000000",
  9028=>"000111100",
  9029=>"111111111",
  9030=>"111111111",
  9031=>"001111111",
  9032=>"000000000",
  9033=>"111111000",
  9034=>"110000110",
  9035=>"000000000",
  9036=>"011001101",
  9037=>"111111111",
  9038=>"000000001",
  9039=>"000000000",
  9040=>"111111111",
  9041=>"010000100",
  9042=>"111111110",
  9043=>"000101111",
  9044=>"000000111",
  9045=>"111111111",
  9046=>"111111000",
  9047=>"000111011",
  9048=>"111111111",
  9049=>"000011111",
  9050=>"110100111",
  9051=>"000000000",
  9052=>"000010010",
  9053=>"000000000",
  9054=>"010110110",
  9055=>"000000000",
  9056=>"000000000",
  9057=>"111111111",
  9058=>"111100110",
  9059=>"111111111",
  9060=>"111111001",
  9061=>"000000000",
  9062=>"111111000",
  9063=>"011011011",
  9064=>"000000000",
  9065=>"100101111",
  9066=>"110110100",
  9067=>"000001000",
  9068=>"011111100",
  9069=>"011111000",
  9070=>"110100110",
  9071=>"000000000",
  9072=>"000000000",
  9073=>"111111000",
  9074=>"010111111",
  9075=>"100100110",
  9076=>"111111001",
  9077=>"000000000",
  9078=>"101111111",
  9079=>"000000000",
  9080=>"111111000",
  9081=>"000001111",
  9082=>"100111111",
  9083=>"000000110",
  9084=>"110000100",
  9085=>"111111111",
  9086=>"001001111",
  9087=>"111101111",
  9088=>"011011011",
  9089=>"000000000",
  9090=>"110110110",
  9091=>"000000000",
  9092=>"111000011",
  9093=>"000000000",
  9094=>"000000000",
  9095=>"111111110",
  9096=>"000000000",
  9097=>"001000001",
  9098=>"111111111",
  9099=>"111111011",
  9100=>"111111111",
  9101=>"111111110",
  9102=>"111111110",
  9103=>"000000000",
  9104=>"111111100",
  9105=>"100000000",
  9106=>"111111111",
  9107=>"011011111",
  9108=>"111111111",
  9109=>"000000000",
  9110=>"111111111",
  9111=>"111000000",
  9112=>"100000111",
  9113=>"000001111",
  9114=>"111111111",
  9115=>"001101111",
  9116=>"111111111",
  9117=>"001000000",
  9118=>"000000000",
  9119=>"110000000",
  9120=>"011111011",
  9121=>"111111011",
  9122=>"010000000",
  9123=>"000000001",
  9124=>"111000000",
  9125=>"100111111",
  9126=>"111111111",
  9127=>"000000000",
  9128=>"000000000",
  9129=>"000000000",
  9130=>"111111111",
  9131=>"111011100",
  9132=>"111100000",
  9133=>"000000000",
  9134=>"100000000",
  9135=>"111111111",
  9136=>"111111000",
  9137=>"000000000",
  9138=>"000000000",
  9139=>"000000000",
  9140=>"111111100",
  9141=>"111111111",
  9142=>"111111111",
  9143=>"000100000",
  9144=>"011111111",
  9145=>"111111111",
  9146=>"111101001",
  9147=>"000000000",
  9148=>"000000000",
  9149=>"000000000",
  9150=>"000000000",
  9151=>"000000100",
  9152=>"101101000",
  9153=>"000000000",
  9154=>"111111111",
  9155=>"000000000",
  9156=>"100000000",
  9157=>"100100110",
  9158=>"111111111",
  9159=>"000111111",
  9160=>"100110001",
  9161=>"000000010",
  9162=>"001001111",
  9163=>"000000111",
  9164=>"100000101",
  9165=>"111111111",
  9166=>"000000001",
  9167=>"111111111",
  9168=>"000000000",
  9169=>"100100111",
  9170=>"111111111",
  9171=>"001001111",
  9172=>"000000100",
  9173=>"010000000",
  9174=>"000001000",
  9175=>"110101101",
  9176=>"000100000",
  9177=>"011000000",
  9178=>"000000100",
  9179=>"111111111",
  9180=>"111100100",
  9181=>"000110110",
  9182=>"001001111",
  9183=>"011111000",
  9184=>"000000000",
  9185=>"011011111",
  9186=>"111111111",
  9187=>"111011001",
  9188=>"000000000",
  9189=>"001111111",
  9190=>"000010001",
  9191=>"000000000",
  9192=>"111000000",
  9193=>"000111000",
  9194=>"000000000",
  9195=>"000000000",
  9196=>"000000000",
  9197=>"110000000",
  9198=>"111000001",
  9199=>"110100000",
  9200=>"000100111",
  9201=>"001000111",
  9202=>"111011011",
  9203=>"000010011",
  9204=>"011011011",
  9205=>"000111111",
  9206=>"000000000",
  9207=>"111111111",
  9208=>"111111101",
  9209=>"000000000",
  9210=>"111111111",
  9211=>"000000001",
  9212=>"000000000",
  9213=>"101011111",
  9214=>"000000011",
  9215=>"001000011",
  9216=>"000000000",
  9217=>"000110110",
  9218=>"011111111",
  9219=>"000000000",
  9220=>"000000000",
  9221=>"001000000",
  9222=>"000000001",
  9223=>"000111111",
  9224=>"000000000",
  9225=>"111001000",
  9226=>"000000000",
  9227=>"000000111",
  9228=>"000000000",
  9229=>"111111000",
  9230=>"101111000",
  9231=>"111111110",
  9232=>"101000000",
  9233=>"101111111",
  9234=>"001011011",
  9235=>"111111111",
  9236=>"111111111",
  9237=>"111001000",
  9238=>"111111101",
  9239=>"001000111",
  9240=>"100100000",
  9241=>"111111111",
  9242=>"011110111",
  9243=>"111111111",
  9244=>"000000000",
  9245=>"111011111",
  9246=>"000000100",
  9247=>"110110000",
  9248=>"111111110",
  9249=>"000101111",
  9250=>"010000000",
  9251=>"111111110",
  9252=>"000000000",
  9253=>"100111111",
  9254=>"011111000",
  9255=>"111000000",
  9256=>"111001111",
  9257=>"111110010",
  9258=>"110111011",
  9259=>"000000111",
  9260=>"111111111",
  9261=>"111111111",
  9262=>"000000000",
  9263=>"000000000",
  9264=>"111001010",
  9265=>"000000100",
  9266=>"000000000",
  9267=>"011001111",
  9268=>"000101111",
  9269=>"000000011",
  9270=>"111101111",
  9271=>"000000001",
  9272=>"101000000",
  9273=>"000000111",
  9274=>"000000000",
  9275=>"000110111",
  9276=>"101111111",
  9277=>"000000000",
  9278=>"000000000",
  9279=>"000000101",
  9280=>"111010110",
  9281=>"001000111",
  9282=>"000000100",
  9283=>"111111110",
  9284=>"000000000",
  9285=>"111111111",
  9286=>"111110100",
  9287=>"010010000",
  9288=>"111111111",
  9289=>"000000111",
  9290=>"111101000",
  9291=>"111001111",
  9292=>"001111111",
  9293=>"010111110",
  9294=>"111001000",
  9295=>"111111111",
  9296=>"000000111",
  9297=>"101000000",
  9298=>"110111111",
  9299=>"000011111",
  9300=>"000010111",
  9301=>"000100011",
  9302=>"001100101",
  9303=>"000000001",
  9304=>"000000000",
  9305=>"000000000",
  9306=>"000100111",
  9307=>"110111110",
  9308=>"101101111",
  9309=>"111111111",
  9310=>"011000000",
  9311=>"111111111",
  9312=>"001001111",
  9313=>"001000000",
  9314=>"001111111",
  9315=>"100100000",
  9316=>"000000111",
  9317=>"111111111",
  9318=>"100100110",
  9319=>"000000100",
  9320=>"000000000",
  9321=>"111101111",
  9322=>"000000000",
  9323=>"111111000",
  9324=>"000000000",
  9325=>"000000001",
  9326=>"000111111",
  9327=>"011011000",
  9328=>"000000000",
  9329=>"101111111",
  9330=>"000110111",
  9331=>"111111000",
  9332=>"000000000",
  9333=>"000000000",
  9334=>"000111111",
  9335=>"000000000",
  9336=>"111111111",
  9337=>"111100111",
  9338=>"000000000",
  9339=>"000000000",
  9340=>"100110100",
  9341=>"000000000",
  9342=>"000000000",
  9343=>"000000000",
  9344=>"001000000",
  9345=>"000000100",
  9346=>"111000000",
  9347=>"110111111",
  9348=>"000000010",
  9349=>"111101111",
  9350=>"111111111",
  9351=>"111011000",
  9352=>"111111111",
  9353=>"001000000",
  9354=>"000100110",
  9355=>"011111111",
  9356=>"000001101",
  9357=>"111111111",
  9358=>"111000000",
  9359=>"000000000",
  9360=>"111111111",
  9361=>"000001001",
  9362=>"000000100",
  9363=>"000110110",
  9364=>"010010000",
  9365=>"000000101",
  9366=>"111111111",
  9367=>"111000000",
  9368=>"000000000",
  9369=>"111111111",
  9370=>"000000000",
  9371=>"000110110",
  9372=>"000000110",
  9373=>"001001000",
  9374=>"000111111",
  9375=>"000000000",
  9376=>"011011001",
  9377=>"111111011",
  9378=>"000001001",
  9379=>"100110110",
  9380=>"000000000",
  9381=>"011111000",
  9382=>"111110111",
  9383=>"000110111",
  9384=>"000000000",
  9385=>"111101101",
  9386=>"000000000",
  9387=>"000000000",
  9388=>"111100000",
  9389=>"111011000",
  9390=>"000000000",
  9391=>"001000111",
  9392=>"111111111",
  9393=>"001110110",
  9394=>"111111111",
  9395=>"000000000",
  9396=>"111110110",
  9397=>"000000111",
  9398=>"000011001",
  9399=>"111111111",
  9400=>"111111001",
  9401=>"000000000",
  9402=>"000000000",
  9403=>"111100101",
  9404=>"111111111",
  9405=>"001001111",
  9406=>"011010000",
  9407=>"001101111",
  9408=>"000000000",
  9409=>"110111111",
  9410=>"000000011",
  9411=>"000001000",
  9412=>"001110111",
  9413=>"011111111",
  9414=>"000000000",
  9415=>"101111100",
  9416=>"111111111",
  9417=>"001000000",
  9418=>"010011000",
  9419=>"001000000",
  9420=>"101101101",
  9421=>"011111111",
  9422=>"000000000",
  9423=>"000000000",
  9424=>"000111110",
  9425=>"001001011",
  9426=>"001011000",
  9427=>"000111111",
  9428=>"111100000",
  9429=>"110110110",
  9430=>"111111010",
  9431=>"111111111",
  9432=>"011111110",
  9433=>"000000011",
  9434=>"011001000",
  9435=>"111111111",
  9436=>"000000100",
  9437=>"111111111",
  9438=>"001000000",
  9439=>"000000111",
  9440=>"111111111",
  9441=>"000011011",
  9442=>"111111111",
  9443=>"111111111",
  9444=>"000011111",
  9445=>"111111111",
  9446=>"111111111",
  9447=>"111011000",
  9448=>"001001000",
  9449=>"100000101",
  9450=>"111111110",
  9451=>"111111100",
  9452=>"000000100",
  9453=>"110111011",
  9454=>"011000000",
  9455=>"011111001",
  9456=>"011011011",
  9457=>"000000000",
  9458=>"000000001",
  9459=>"000000000",
  9460=>"011001000",
  9461=>"111111111",
  9462=>"111111111",
  9463=>"111011111",
  9464=>"000111111",
  9465=>"000000000",
  9466=>"111000000",
  9467=>"000000011",
  9468=>"011001001",
  9469=>"111100111",
  9470=>"111000110",
  9471=>"011000000",
  9472=>"111111111",
  9473=>"000000011",
  9474=>"100000000",
  9475=>"001111111",
  9476=>"111111001",
  9477=>"001001111",
  9478=>"000000000",
  9479=>"000000111",
  9480=>"111101111",
  9481=>"110110111",
  9482=>"011000000",
  9483=>"010000000",
  9484=>"111001001",
  9485=>"011101111",
  9486=>"001000101",
  9487=>"111111000",
  9488=>"111111111",
  9489=>"001000000",
  9490=>"111000000",
  9491=>"111111111",
  9492=>"000000000",
  9493=>"000010000",
  9494=>"111000000",
  9495=>"100000000",
  9496=>"111111111",
  9497=>"000000000",
  9498=>"111111111",
  9499=>"000000000",
  9500=>"001011111",
  9501=>"111111111",
  9502=>"111111111",
  9503=>"000000001",
  9504=>"100001000",
  9505=>"111111111",
  9506=>"111111111",
  9507=>"111111111",
  9508=>"000100100",
  9509=>"111111111",
  9510=>"000000000",
  9511=>"000000000",
  9512=>"010010111",
  9513=>"011011000",
  9514=>"001000000",
  9515=>"000000000",
  9516=>"000000000",
  9517=>"100000000",
  9518=>"000000000",
  9519=>"000000011",
  9520=>"111111111",
  9521=>"000000000",
  9522=>"000000000",
  9523=>"111111110",
  9524=>"000000000",
  9525=>"100000000",
  9526=>"010011111",
  9527=>"111111111",
  9528=>"111111000",
  9529=>"111111000",
  9530=>"000110111",
  9531=>"110110000",
  9532=>"110111111",
  9533=>"001001001",
  9534=>"000010000",
  9535=>"111111111",
  9536=>"111000000",
  9537=>"000000000",
  9538=>"000000111",
  9539=>"100111111",
  9540=>"111111111",
  9541=>"111111111",
  9542=>"000000101",
  9543=>"001000000",
  9544=>"111100111",
  9545=>"010000000",
  9546=>"101000001",
  9547=>"000101111",
  9548=>"000000000",
  9549=>"111111110",
  9550=>"000000000",
  9551=>"000111111",
  9552=>"000000000",
  9553=>"000100111",
  9554=>"001100111",
  9555=>"111000101",
  9556=>"111100100",
  9557=>"011011011",
  9558=>"000000001",
  9559=>"111111111",
  9560=>"000000000",
  9561=>"111111111",
  9562=>"111111111",
  9563=>"001000001",
  9564=>"111111110",
  9565=>"000000000",
  9566=>"101000001",
  9567=>"001001001",
  9568=>"101111111",
  9569=>"111111111",
  9570=>"100100110",
  9571=>"111110000",
  9572=>"000000000",
  9573=>"100000101",
  9574=>"110010111",
  9575=>"011011001",
  9576=>"110110111",
  9577=>"110110110",
  9578=>"000000000",
  9579=>"011001000",
  9580=>"011011111",
  9581=>"111111111",
  9582=>"000000000",
  9583=>"111111000",
  9584=>"010000000",
  9585=>"000000000",
  9586=>"101111111",
  9587=>"000110010",
  9588=>"010000000",
  9589=>"000111011",
  9590=>"111111111",
  9591=>"000000010",
  9592=>"111001111",
  9593=>"000000000",
  9594=>"111001000",
  9595=>"000000000",
  9596=>"100100000",
  9597=>"001000001",
  9598=>"011000101",
  9599=>"000000000",
  9600=>"111011001",
  9601=>"011111111",
  9602=>"111111001",
  9603=>"000000110",
  9604=>"010000000",
  9605=>"000000110",
  9606=>"111111001",
  9607=>"111111111",
  9608=>"111111111",
  9609=>"110100000",
  9610=>"111111000",
  9611=>"100100100",
  9612=>"000000001",
  9613=>"111111111",
  9614=>"000111111",
  9615=>"000000000",
  9616=>"111111010",
  9617=>"110111111",
  9618=>"101111011",
  9619=>"011111111",
  9620=>"111001000",
  9621=>"000000000",
  9622=>"011001000",
  9623=>"110110110",
  9624=>"111111000",
  9625=>"000100100",
  9626=>"000011000",
  9627=>"111111111",
  9628=>"000000000",
  9629=>"111111111",
  9630=>"000001001",
  9631=>"000000000",
  9632=>"000000000",
  9633=>"100110111",
  9634=>"001101011",
  9635=>"000000001",
  9636=>"100100001",
  9637=>"000110111",
  9638=>"000000000",
  9639=>"111111111",
  9640=>"001011111",
  9641=>"111111111",
  9642=>"001111111",
  9643=>"000000000",
  9644=>"000000000",
  9645=>"111111111",
  9646=>"111100000",
  9647=>"111000100",
  9648=>"111111111",
  9649=>"000000110",
  9650=>"111111001",
  9651=>"000000000",
  9652=>"111111111",
  9653=>"011111111",
  9654=>"111001000",
  9655=>"000000000",
  9656=>"100000000",
  9657=>"010000000",
  9658=>"111111111",
  9659=>"111111111",
  9660=>"011111011",
  9661=>"111111011",
  9662=>"101000000",
  9663=>"011001001",
  9664=>"000010011",
  9665=>"001011010",
  9666=>"111101111",
  9667=>"011011011",
  9668=>"001001000",
  9669=>"001001001",
  9670=>"000000000",
  9671=>"001011000",
  9672=>"010000000",
  9673=>"000000111",
  9674=>"100000111",
  9675=>"111111111",
  9676=>"111001000",
  9677=>"100000000",
  9678=>"001001011",
  9679=>"111010000",
  9680=>"100000000",
  9681=>"000000001",
  9682=>"111111111",
  9683=>"110010111",
  9684=>"001000111",
  9685=>"000000111",
  9686=>"001001111",
  9687=>"000000000",
  9688=>"111111111",
  9689=>"111000110",
  9690=>"000111111",
  9691=>"001001011",
  9692=>"000000111",
  9693=>"000000111",
  9694=>"000010011",
  9695=>"000000001",
  9696=>"000000000",
  9697=>"000001000",
  9698=>"000000000",
  9699=>"000000000",
  9700=>"111111111",
  9701=>"111111111",
  9702=>"111000000",
  9703=>"110111111",
  9704=>"001001000",
  9705=>"000000000",
  9706=>"010000000",
  9707=>"111111111",
  9708=>"111001000",
  9709=>"000100111",
  9710=>"111111000",
  9711=>"000000111",
  9712=>"000000000",
  9713=>"000000000",
  9714=>"000101100",
  9715=>"111111010",
  9716=>"000000000",
  9717=>"000000000",
  9718=>"111100000",
  9719=>"100001000",
  9720=>"000000111",
  9721=>"110101111",
  9722=>"000000000",
  9723=>"111111000",
  9724=>"000000000",
  9725=>"111101100",
  9726=>"111111111",
  9727=>"000000000",
  9728=>"100100100",
  9729=>"010010010",
  9730=>"000000000",
  9731=>"111111111",
  9732=>"111011011",
  9733=>"101100000",
  9734=>"000000000",
  9735=>"000000111",
  9736=>"111011001",
  9737=>"111000000",
  9738=>"000011111",
  9739=>"000000011",
  9740=>"000001101",
  9741=>"001011111",
  9742=>"101111111",
  9743=>"110111111",
  9744=>"111101111",
  9745=>"001111111",
  9746=>"000100100",
  9747=>"000000111",
  9748=>"000000000",
  9749=>"001100111",
  9750=>"000000000",
  9751=>"000000100",
  9752=>"000000101",
  9753=>"110000000",
  9754=>"111111111",
  9755=>"110111011",
  9756=>"000010010",
  9757=>"111111111",
  9758=>"111111111",
  9759=>"110011111",
  9760=>"000000000",
  9761=>"001001110",
  9762=>"111101001",
  9763=>"111111011",
  9764=>"111111111",
  9765=>"001000000",
  9766=>"000000000",
  9767=>"111111101",
  9768=>"111111100",
  9769=>"110111111",
  9770=>"011011011",
  9771=>"111100000",
  9772=>"111011011",
  9773=>"111111111",
  9774=>"000000000",
  9775=>"000000011",
  9776=>"111111111",
  9777=>"110010000",
  9778=>"011011011",
  9779=>"110000000",
  9780=>"001000000",
  9781=>"111111111",
  9782=>"000011011",
  9783=>"000000000",
  9784=>"000000000",
  9785=>"000000110",
  9786=>"111111000",
  9787=>"010000000",
  9788=>"000000111",
  9789=>"110111000",
  9790=>"011001110",
  9791=>"000000000",
  9792=>"110000010",
  9793=>"000000000",
  9794=>"111111111",
  9795=>"000000000",
  9796=>"001001001",
  9797=>"111010000",
  9798=>"000000000",
  9799=>"111111111",
  9800=>"110110110",
  9801=>"000000000",
  9802=>"000000011",
  9803=>"011111110",
  9804=>"000000001",
  9805=>"001001110",
  9806=>"100100000",
  9807=>"111111111",
  9808=>"000000000",
  9809=>"111111111",
  9810=>"000011010",
  9811=>"111111111",
  9812=>"101101111",
  9813=>"000000000",
  9814=>"111111000",
  9815=>"011011011",
  9816=>"000001000",
  9817=>"000000000",
  9818=>"111011011",
  9819=>"011001001",
  9820=>"011111111",
  9821=>"110000000",
  9822=>"000000000",
  9823=>"001000001",
  9824=>"000000000",
  9825=>"110110000",
  9826=>"000000010",
  9827=>"000000000",
  9828=>"111011110",
  9829=>"111000000",
  9830=>"111111011",
  9831=>"000000110",
  9832=>"000001001",
  9833=>"000000000",
  9834=>"000000000",
  9835=>"111011000",
  9836=>"000100001",
  9837=>"000000000",
  9838=>"111111111",
  9839=>"000100100",
  9840=>"111010000",
  9841=>"011000000",
  9842=>"111110100",
  9843=>"111111111",
  9844=>"110110110",
  9845=>"001000111",
  9846=>"111111001",
  9847=>"000000000",
  9848=>"111111111",
  9849=>"000001000",
  9850=>"000000001",
  9851=>"100000000",
  9852=>"111001011",
  9853=>"111111011",
  9854=>"000011011",
  9855=>"001000000",
  9856=>"000000000",
  9857=>"111111111",
  9858=>"100000000",
  9859=>"111111111",
  9860=>"111111111",
  9861=>"000000000",
  9862=>"001011011",
  9863=>"111111111",
  9864=>"111111111",
  9865=>"000000001",
  9866=>"000000000",
  9867=>"000000001",
  9868=>"111111111",
  9869=>"110100001",
  9870=>"000000000",
  9871=>"001101111",
  9872=>"000000000",
  9873=>"111111111",
  9874=>"110110000",
  9875=>"100110010",
  9876=>"010011111",
  9877=>"111111111",
  9878=>"011000000",
  9879=>"110111000",
  9880=>"011111000",
  9881=>"000000111",
  9882=>"000101000",
  9883=>"000000000",
  9884=>"100111110",
  9885=>"010111010",
  9886=>"100000011",
  9887=>"000110111",
  9888=>"000000000",
  9889=>"100000000",
  9890=>"011001011",
  9891=>"100100000",
  9892=>"001011001",
  9893=>"000010111",
  9894=>"001001111",
  9895=>"110110110",
  9896=>"010000000",
  9897=>"000000000",
  9898=>"111011001",
  9899=>"111001000",
  9900=>"100011111",
  9901=>"111111010",
  9902=>"010111000",
  9903=>"101101000",
  9904=>"000000000",
  9905=>"111011111",
  9906=>"111111111",
  9907=>"001101111",
  9908=>"001000000",
  9909=>"110110010",
  9910=>"000000000",
  9911=>"111111000",
  9912=>"000111111",
  9913=>"111011111",
  9914=>"000000000",
  9915=>"111111010",
  9916=>"000000000",
  9917=>"111011000",
  9918=>"111111000",
  9919=>"000000000",
  9920=>"000000000",
  9921=>"100110010",
  9922=>"011011011",
  9923=>"000001111",
  9924=>"111111100",
  9925=>"111111011",
  9926=>"000000100",
  9927=>"000000000",
  9928=>"110000100",
  9929=>"100100100",
  9930=>"111101001",
  9931=>"111110111",
  9932=>"000000100",
  9933=>"000100100",
  9934=>"000000000",
  9935=>"000111011",
  9936=>"000000000",
  9937=>"111111000",
  9938=>"011011000",
  9939=>"000000000",
  9940=>"111111111",
  9941=>"000000001",
  9942=>"000000000",
  9943=>"000111111",
  9944=>"111111111",
  9945=>"000110010",
  9946=>"111111000",
  9947=>"111111111",
  9948=>"000110111",
  9949=>"000000000",
  9950=>"100000000",
  9951=>"000000000",
  9952=>"100100100",
  9953=>"000000000",
  9954=>"111111100",
  9955=>"111011001",
  9956=>"000000000",
  9957=>"100110100",
  9958=>"000000111",
  9959=>"000000011",
  9960=>"000000011",
  9961=>"000000001",
  9962=>"110111001",
  9963=>"000111111",
  9964=>"011111111",
  9965=>"111110111",
  9966=>"000110110",
  9967=>"011111011",
  9968=>"111111111",
  9969=>"111000000",
  9970=>"111111111",
  9971=>"000000000",
  9972=>"011000000",
  9973=>"110000000",
  9974=>"000000100",
  9975=>"000000000",
  9976=>"011011001",
  9977=>"111001111",
  9978=>"000000000",
  9979=>"110000000",
  9980=>"001000110",
  9981=>"000001111",
  9982=>"111111111",
  9983=>"000110111",
  9984=>"000000000",
  9985=>"001000000",
  9986=>"111111111",
  9987=>"100000000",
  9988=>"000111111",
  9989=>"111011000",
  9990=>"000110000",
  9991=>"000000000",
  9992=>"100111010",
  9993=>"000000000",
  9994=>"111111011",
  9995=>"111110110",
  9996=>"000010110",
  9997=>"111111111",
  9998=>"111111011",
  9999=>"111111100",
  10000=>"011000110",
  10001=>"000110111",
  10002=>"111111111",
  10003=>"000000000",
  10004=>"111111000",
  10005=>"001111011",
  10006=>"001000000",
  10007=>"011111111",
  10008=>"111111111",
  10009=>"010000011",
  10010=>"110111111",
  10011=>"100101101",
  10012=>"110100000",
  10013=>"000000001",
  10014=>"000000001",
  10015=>"100111111",
  10016=>"000000111",
  10017=>"111111011",
  10018=>"000110100",
  10019=>"000000001",
  10020=>"001001001",
  10021=>"100110000",
  10022=>"110110111",
  10023=>"000000000",
  10024=>"111111111",
  10025=>"110000111",
  10026=>"111111110",
  10027=>"000000111",
  10028=>"011001111",
  10029=>"000001001",
  10030=>"000000000",
  10031=>"111111111",
  10032=>"001001011",
  10033=>"100000111",
  10034=>"000001011",
  10035=>"111001000",
  10036=>"100000000",
  10037=>"000000000",
  10038=>"000000111",
  10039=>"000001001",
  10040=>"000000000",
  10041=>"000000111",
  10042=>"111111111",
  10043=>"000000000",
  10044=>"001000000",
  10045=>"000000100",
  10046=>"111111011",
  10047=>"001111111",
  10048=>"010011111",
  10049=>"111111111",
  10050=>"110100000",
  10051=>"110100000",
  10052=>"111110000",
  10053=>"100110111",
  10054=>"001000000",
  10055=>"000110110",
  10056=>"111111110",
  10057=>"010000000",
  10058=>"111111110",
  10059=>"000000100",
  10060=>"000000011",
  10061=>"000000011",
  10062=>"011111011",
  10063=>"001011001",
  10064=>"000001011",
  10065=>"110010011",
  10066=>"000000000",
  10067=>"111111111",
  10068=>"000111011",
  10069=>"111111111",
  10070=>"000001111",
  10071=>"000001111",
  10072=>"000000000",
  10073=>"111111111",
  10074=>"111101000",
  10075=>"000000000",
  10076=>"000000000",
  10077=>"111111111",
  10078=>"000000000",
  10079=>"011000000",
  10080=>"000000011",
  10081=>"111111111",
  10082=>"011011101",
  10083=>"000000001",
  10084=>"111111010",
  10085=>"100000000",
  10086=>"111111110",
  10087=>"111110111",
  10088=>"000010000",
  10089=>"111001000",
  10090=>"111111111",
  10091=>"001000010",
  10092=>"110100110",
  10093=>"000000100",
  10094=>"000000111",
  10095=>"000000000",
  10096=>"000000000",
  10097=>"011011111",
  10098=>"111111111",
  10099=>"000000000",
  10100=>"101111111",
  10101=>"000010010",
  10102=>"010010010",
  10103=>"111000010",
  10104=>"000000001",
  10105=>"000000000",
  10106=>"111100001",
  10107=>"010110110",
  10108=>"000001111",
  10109=>"000000011",
  10110=>"111111100",
  10111=>"000000000",
  10112=>"000000000",
  10113=>"101110010",
  10114=>"111111111",
  10115=>"000000000",
  10116=>"000000000",
  10117=>"111111111",
  10118=>"110110110",
  10119=>"001001001",
  10120=>"111111111",
  10121=>"001011011",
  10122=>"100100100",
  10123=>"111001000",
  10124=>"111001000",
  10125=>"000000000",
  10126=>"011111000",
  10127=>"111111111",
  10128=>"000000111",
  10129=>"111111001",
  10130=>"111111111",
  10131=>"011011011",
  10132=>"001100100",
  10133=>"101000000",
  10134=>"001100000",
  10135=>"111111111",
  10136=>"111101111",
  10137=>"111111011",
  10138=>"000000000",
  10139=>"111111111",
  10140=>"011011001",
  10141=>"100111000",
  10142=>"000000011",
  10143=>"000000000",
  10144=>"000011011",
  10145=>"011111110",
  10146=>"111111110",
  10147=>"111111111",
  10148=>"111111111",
  10149=>"111101101",
  10150=>"111111111",
  10151=>"111111111",
  10152=>"000000000",
  10153=>"000000100",
  10154=>"100000000",
  10155=>"000000001",
  10156=>"011000011",
  10157=>"000000000",
  10158=>"111111111",
  10159=>"001111100",
  10160=>"111111111",
  10161=>"111101000",
  10162=>"000000000",
  10163=>"000000001",
  10164=>"000001001",
  10165=>"100110111",
  10166=>"100111000",
  10167=>"111110110",
  10168=>"000000000",
  10169=>"000000000",
  10170=>"000001001",
  10171=>"111111000",
  10172=>"100101111",
  10173=>"000000011",
  10174=>"000000000",
  10175=>"011011110",
  10176=>"111010000",
  10177=>"000000000",
  10178=>"111011010",
  10179=>"110000000",
  10180=>"000110110",
  10181=>"010011011",
  10182=>"000000100",
  10183=>"111000000",
  10184=>"000011000",
  10185=>"011111110",
  10186=>"100000000",
  10187=>"000100100",
  10188=>"111111111",
  10189=>"000110111",
  10190=>"010010000",
  10191=>"111111111",
  10192=>"000000000",
  10193=>"100111111",
  10194=>"001101111",
  10195=>"111111111",
  10196=>"001111100",
  10197=>"000111111",
  10198=>"100100100",
  10199=>"100100111",
  10200=>"111111111",
  10201=>"111100001",
  10202=>"111111110",
  10203=>"111111000",
  10204=>"111101101",
  10205=>"000111001",
  10206=>"000110100",
  10207=>"011111111",
  10208=>"100100110",
  10209=>"100110111",
  10210=>"000000000",
  10211=>"000000000",
  10212=>"000010010",
  10213=>"001011111",
  10214=>"110101111",
  10215=>"111000000",
  10216=>"111110110",
  10217=>"111001000",
  10218=>"110000000",
  10219=>"111111111",
  10220=>"110111011",
  10221=>"100000000",
  10222=>"000000000",
  10223=>"100000101",
  10224=>"011011011",
  10225=>"000001110",
  10226=>"110110010",
  10227=>"111010000",
  10228=>"001001001",
  10229=>"111111111",
  10230=>"110001001",
  10231=>"110000100",
  10232=>"000100111",
  10233=>"000010000",
  10234=>"000010110",
  10235=>"111111001",
  10236=>"000000111",
  10237=>"101111111",
  10238=>"001000000",
  10239=>"000000000",
  10240=>"001000000",
  10241=>"001000000",
  10242=>"111101111",
  10243=>"111111000",
  10244=>"000000100",
  10245=>"111111111",
  10246=>"000000000",
  10247=>"111011111",
  10248=>"111101111",
  10249=>"111001001",
  10250=>"000000111",
  10251=>"000000111",
  10252=>"100100000",
  10253=>"111110100",
  10254=>"111101000",
  10255=>"000001000",
  10256=>"111111111",
  10257=>"110110001",
  10258=>"000010111",
  10259=>"111111111",
  10260=>"111000000",
  10261=>"101111111",
  10262=>"110111111",
  10263=>"001011011",
  10264=>"111111111",
  10265=>"111111001",
  10266=>"001000001",
  10267=>"111010010",
  10268=>"000000110",
  10269=>"000100111",
  10270=>"011011111",
  10271=>"111111111",
  10272=>"000001111",
  10273=>"000001000",
  10274=>"000000000",
  10275=>"000000010",
  10276=>"000000000",
  10277=>"000000000",
  10278=>"111111100",
  10279=>"001000000",
  10280=>"111100111",
  10281=>"111111000",
  10282=>"000000100",
  10283=>"111110111",
  10284=>"111011000",
  10285=>"111111101",
  10286=>"111111111",
  10287=>"110110011",
  10288=>"101001000",
  10289=>"000000000",
  10290=>"001001000",
  10291=>"100100000",
  10292=>"000111111",
  10293=>"000001101",
  10294=>"111011100",
  10295=>"011000100",
  10296=>"111111111",
  10297=>"011011111",
  10298=>"000110000",
  10299=>"000001001",
  10300=>"000111111",
  10301=>"010000000",
  10302=>"001011100",
  10303=>"111100000",
  10304=>"000000111",
  10305=>"000110000",
  10306=>"011111010",
  10307=>"111010000",
  10308=>"110110000",
  10309=>"000000011",
  10310=>"111000000",
  10311=>"111111111",
  10312=>"011011000",
  10313=>"000000111",
  10314=>"000000111",
  10315=>"111000000",
  10316=>"000000100",
  10317=>"000000111",
  10318=>"011010000",
  10319=>"111110000",
  10320=>"000000110",
  10321=>"000111111",
  10322=>"010110000",
  10323=>"100100000",
  10324=>"000111100",
  10325=>"111111011",
  10326=>"001001001",
  10327=>"000000101",
  10328=>"111110010",
  10329=>"101000000",
  10330=>"111111000",
  10331=>"111001001",
  10332=>"111000000",
  10333=>"000101011",
  10334=>"111111000",
  10335=>"001000000",
  10336=>"000000000",
  10337=>"001000101",
  10338=>"000000110",
  10339=>"000000000",
  10340=>"000010000",
  10341=>"100000101",
  10342=>"111111111",
  10343=>"000000000",
  10344=>"000111111",
  10345=>"111000110",
  10346=>"100000111",
  10347=>"110111111",
  10348=>"111000000",
  10349=>"001001111",
  10350=>"000101111",
  10351=>"111111011",
  10352=>"011011000",
  10353=>"111110111",
  10354=>"000011001",
  10355=>"101001001",
  10356=>"101101111",
  10357=>"111111100",
  10358=>"000000111",
  10359=>"001011010",
  10360=>"000101111",
  10361=>"000111111",
  10362=>"111111000",
  10363=>"000000111",
  10364=>"011010010",
  10365=>"111111101",
  10366=>"111111000",
  10367=>"111001001",
  10368=>"000100111",
  10369=>"000001111",
  10370=>"000011111",
  10371=>"001011000",
  10372=>"111000000",
  10373=>"111111111",
  10374=>"000010110",
  10375=>"000011000",
  10376=>"001111111",
  10377=>"111111110",
  10378=>"000010000",
  10379=>"001000010",
  10380=>"001001111",
  10381=>"010010100",
  10382=>"000000111",
  10383=>"110111110",
  10384=>"001001000",
  10385=>"100101111",
  10386=>"110010000",
  10387=>"001011001",
  10388=>"111111010",
  10389=>"000101111",
  10390=>"000000000",
  10391=>"011111111",
  10392=>"100111111",
  10393=>"111111111",
  10394=>"000000010",
  10395=>"000111111",
  10396=>"001111000",
  10397=>"100111111",
  10398=>"000111111",
  10399=>"111111000",
  10400=>"000000000",
  10401=>"000000010",
  10402=>"001000110",
  10403=>"000000110",
  10404=>"101101000",
  10405=>"100001101",
  10406=>"001111000",
  10407=>"001011111",
  10408=>"000000000",
  10409=>"000000000",
  10410=>"100000000",
  10411=>"000000000",
  10412=>"111111111",
  10413=>"011000011",
  10414=>"000110111",
  10415=>"111000000",
  10416=>"111111111",
  10417=>"011111100",
  10418=>"001101000",
  10419=>"111111111",
  10420=>"000000000",
  10421=>"101000001",
  10422=>"001011000",
  10423=>"100110111",
  10424=>"111111111",
  10425=>"000111111",
  10426=>"100100000",
  10427=>"100000111",
  10428=>"111000001",
  10429=>"100000000",
  10430=>"110111111",
  10431=>"000000111",
  10432=>"100000000",
  10433=>"000000000",
  10434=>"111111000",
  10435=>"111111000",
  10436=>"000000000",
  10437=>"001001111",
  10438=>"011111111",
  10439=>"000101111",
  10440=>"100111111",
  10441=>"111001111",
  10442=>"000000000",
  10443=>"000111111",
  10444=>"000000000",
  10445=>"111111111",
  10446=>"111111110",
  10447=>"111111111",
  10448=>"000000000",
  10449=>"000010000",
  10450=>"111100100",
  10451=>"111011000",
  10452=>"000001111",
  10453=>"000100100",
  10454=>"111111011",
  10455=>"000000000",
  10456=>"101111000",
  10457=>"111110000",
  10458=>"011001001",
  10459=>"111111000",
  10460=>"111110111",
  10461=>"111111111",
  10462=>"000111111",
  10463=>"000000001",
  10464=>"000010111",
  10465=>"111000000",
  10466=>"111111111",
  10467=>"111111010",
  10468=>"100111111",
  10469=>"011001100",
  10470=>"111110000",
  10471=>"000000000",
  10472=>"000000110",
  10473=>"001111101",
  10474=>"111111011",
  10475=>"111000000",
  10476=>"000000000",
  10477=>"000000110",
  10478=>"111010000",
  10479=>"111111000",
  10480=>"111111000",
  10481=>"000000101",
  10482=>"000000001",
  10483=>"110010000",
  10484=>"111111000",
  10485=>"111100000",
  10486=>"100110111",
  10487=>"111101111",
  10488=>"110000000",
  10489=>"111000000",
  10490=>"110110111",
  10491=>"000001011",
  10492=>"111111111",
  10493=>"000000000",
  10494=>"111101111",
  10495=>"110110111",
  10496=>"111111000",
  10497=>"001011000",
  10498=>"000000000",
  10499=>"110000111",
  10500=>"111011000",
  10501=>"111110000",
  10502=>"000011111",
  10503=>"110000000",
  10504=>"111101000",
  10505=>"000110110",
  10506=>"110000000",
  10507=>"100000111",
  10508=>"000000000",
  10509=>"111111111",
  10510=>"101100000",
  10511=>"110110111",
  10512=>"100000111",
  10513=>"001000000",
  10514=>"111111111",
  10515=>"001000001",
  10516=>"110000000",
  10517=>"000011000",
  10518=>"010110000",
  10519=>"000011011",
  10520=>"111111111",
  10521=>"111011010",
  10522=>"111111000",
  10523=>"000000000",
  10524=>"011010010",
  10525=>"010000000",
  10526=>"111000000",
  10527=>"111011010",
  10528=>"001101111",
  10529=>"111000000",
  10530=>"111000111",
  10531=>"110110111",
  10532=>"111100111",
  10533=>"001011111",
  10534=>"001011001",
  10535=>"001000100",
  10536=>"000000000",
  10537=>"011010000",
  10538=>"111111000",
  10539=>"000000000",
  10540=>"111111111",
  10541=>"001111111",
  10542=>"111111000",
  10543=>"111110000",
  10544=>"001111111",
  10545=>"111100110",
  10546=>"011011111",
  10547=>"001111000",
  10548=>"000001000",
  10549=>"111101000",
  10550=>"111000000",
  10551=>"111111111",
  10552=>"000000101",
  10553=>"001000001",
  10554=>"111111111",
  10555=>"101001111",
  10556=>"001001000",
  10557=>"111111111",
  10558=>"000000000",
  10559=>"111111111",
  10560=>"000000111",
  10561=>"000101111",
  10562=>"000000000",
  10563=>"000000110",
  10564=>"111111111",
  10565=>"001101111",
  10566=>"000000100",
  10567=>"010000011",
  10568=>"111111110",
  10569=>"111000000",
  10570=>"000000000",
  10571=>"000000000",
  10572=>"101111111",
  10573=>"000111111",
  10574=>"111111000",
  10575=>"100111111",
  10576=>"011011111",
  10577=>"110000011",
  10578=>"100000111",
  10579=>"111001001",
  10580=>"000000000",
  10581=>"001000001",
  10582=>"000000111",
  10583=>"111000011",
  10584=>"111000000",
  10585=>"111111000",
  10586=>"000000001",
  10587=>"110010000",
  10588=>"110111000",
  10589=>"000000110",
  10590=>"000110100",
  10591=>"000001111",
  10592=>"000111101",
  10593=>"000000111",
  10594=>"100110111",
  10595=>"000000000",
  10596=>"000010000",
  10597=>"011000000",
  10598=>"011000000",
  10599=>"111111111",
  10600=>"010010011",
  10601=>"000011000",
  10602=>"000000000",
  10603=>"101111011",
  10604=>"111111110",
  10605=>"110111001",
  10606=>"000000000",
  10607=>"000000000",
  10608=>"000000000",
  10609=>"000000011",
  10610=>"001000000",
  10611=>"101011001",
  10612=>"100111111",
  10613=>"000111011",
  10614=>"000000011",
  10615=>"001100000",
  10616=>"000000000",
  10617=>"010010000",
  10618=>"011000000",
  10619=>"111000000",
  10620=>"111000100",
  10621=>"100000000",
  10622=>"000000000",
  10623=>"000000000",
  10624=>"111110110",
  10625=>"000101111",
  10626=>"100100110",
  10627=>"000000110",
  10628=>"111001111",
  10629=>"000000000",
  10630=>"000100000",
  10631=>"111110111",
  10632=>"001011000",
  10633=>"010000111",
  10634=>"000011111",
  10635=>"011000000",
  10636=>"000000001",
  10637=>"100110111",
  10638=>"000000000",
  10639=>"000100111",
  10640=>"111111000",
  10641=>"111110111",
  10642=>"001000110",
  10643=>"110100000",
  10644=>"001000111",
  10645=>"010110110",
  10646=>"000000000",
  10647=>"000010110",
  10648=>"000000111",
  10649=>"111001111",
  10650=>"111111111",
  10651=>"111111111",
  10652=>"101111111",
  10653=>"111111001",
  10654=>"000000111",
  10655=>"010011111",
  10656=>"110101111",
  10657=>"011111111",
  10658=>"100000001",
  10659=>"101101111",
  10660=>"100000000",
  10661=>"111111000",
  10662=>"001000000",
  10663=>"000000001",
  10664=>"000000000",
  10665=>"111000000",
  10666=>"111010000",
  10667=>"001111001",
  10668=>"111111000",
  10669=>"001000000",
  10670=>"111100111",
  10671=>"111111111",
  10672=>"000000000",
  10673=>"000000000",
  10674=>"100110000",
  10675=>"110000000",
  10676=>"110110000",
  10677=>"000000111",
  10678=>"011001011",
  10679=>"111110001",
  10680=>"111111000",
  10681=>"010000111",
  10682=>"111000000",
  10683=>"110110111",
  10684=>"111111111",
  10685=>"001000110",
  10686=>"000001100",
  10687=>"010010010",
  10688=>"000000000",
  10689=>"111111001",
  10690=>"000000000",
  10691=>"010000000",
  10692=>"000000100",
  10693=>"111001001",
  10694=>"011000101",
  10695=>"000111111",
  10696=>"110000001",
  10697=>"000011000",
  10698=>"001001111",
  10699=>"111111000",
  10700=>"010011000",
  10701=>"010001111",
  10702=>"011001111",
  10703=>"000001111",
  10704=>"000000100",
  10705=>"110111111",
  10706=>"111111000",
  10707=>"111111000",
  10708=>"101101111",
  10709=>"111111000",
  10710=>"000001001",
  10711=>"011001011",
  10712=>"000000000",
  10713=>"111011011",
  10714=>"111000000",
  10715=>"001011111",
  10716=>"100100111",
  10717=>"111000011",
  10718=>"111111001",
  10719=>"011001111",
  10720=>"011011011",
  10721=>"111000010",
  10722=>"000000000",
  10723=>"001011111",
  10724=>"000000101",
  10725=>"110101111",
  10726=>"111000100",
  10727=>"111100000",
  10728=>"101111111",
  10729=>"111111111",
  10730=>"111000000",
  10731=>"111010011",
  10732=>"000111000",
  10733=>"110010000",
  10734=>"000000110",
  10735=>"000000000",
  10736=>"000000000",
  10737=>"000000000",
  10738=>"111000111",
  10739=>"011000111",
  10740=>"111111000",
  10741=>"101100111",
  10742=>"000011001",
  10743=>"000011011",
  10744=>"001011001",
  10745=>"011011000",
  10746=>"010110110",
  10747=>"000000111",
  10748=>"100000000",
  10749=>"011000000",
  10750=>"111111000",
  10751=>"000001011",
  10752=>"111111111",
  10753=>"000100111",
  10754=>"000000000",
  10755=>"001011000",
  10756=>"001000000",
  10757=>"001000000",
  10758=>"000000000",
  10759=>"111000011",
  10760=>"000000111",
  10761=>"000001000",
  10762=>"000000000",
  10763=>"000101111",
  10764=>"000000000",
  10765=>"011000000",
  10766=>"110000100",
  10767=>"111001011",
  10768=>"000000000",
  10769=>"111011111",
  10770=>"001000101",
  10771=>"000000011",
  10772=>"000000000",
  10773=>"000000000",
  10774=>"111000000",
  10775=>"100101011",
  10776=>"001001001",
  10777=>"101100100",
  10778=>"000000000",
  10779=>"000000000",
  10780=>"110111111",
  10781=>"000000000",
  10782=>"011111111",
  10783=>"100100000",
  10784=>"000000000",
  10785=>"110110100",
  10786=>"111110000",
  10787=>"110000001",
  10788=>"000000011",
  10789=>"111001000",
  10790=>"001000101",
  10791=>"000111000",
  10792=>"111111111",
  10793=>"000000000",
  10794=>"101111011",
  10795=>"111000000",
  10796=>"111001001",
  10797=>"000000001",
  10798=>"000010000",
  10799=>"111111101",
  10800=>"000000100",
  10801=>"001000000",
  10802=>"111111111",
  10803=>"000000100",
  10804=>"111111111",
  10805=>"111000000",
  10806=>"111111111",
  10807=>"111111100",
  10808=>"111111111",
  10809=>"000000001",
  10810=>"000000000",
  10811=>"100100000",
  10812=>"000111111",
  10813=>"100000000",
  10814=>"011010010",
  10815=>"100100100",
  10816=>"111011011",
  10817=>"000000000",
  10818=>"000111111",
  10819=>"000000111",
  10820=>"001000000",
  10821=>"001001000",
  10822=>"001111111",
  10823=>"000000000",
  10824=>"111111001",
  10825=>"000000000",
  10826=>"111111001",
  10827=>"000000111",
  10828=>"111111000",
  10829=>"000000100",
  10830=>"011000001",
  10831=>"000000110",
  10832=>"100100100",
  10833=>"111111011",
  10834=>"111000000",
  10835=>"000001111",
  10836=>"000000110",
  10837=>"000000000",
  10838=>"101110110",
  10839=>"101111111",
  10840=>"000100000",
  10841=>"100100100",
  10842=>"000000101",
  10843=>"000010111",
  10844=>"110010110",
  10845=>"001001000",
  10846=>"000001001",
  10847=>"011000001",
  10848=>"000000111",
  10849=>"001000111",
  10850=>"111011101",
  10851=>"010011111",
  10852=>"000001000",
  10853=>"000000011",
  10854=>"101000000",
  10855=>"111001001",
  10856=>"000000000",
  10857=>"110111111",
  10858=>"000111101",
  10859=>"000000000",
  10860=>"100000000",
  10861=>"011000111",
  10862=>"001101111",
  10863=>"001001000",
  10864=>"111111111",
  10865=>"111111111",
  10866=>"111111000",
  10867=>"011001001",
  10868=>"000111111",
  10869=>"000000100",
  10870=>"000000110",
  10871=>"000010111",
  10872=>"000000001",
  10873=>"000000000",
  10874=>"000000000",
  10875=>"000000111",
  10876=>"110111111",
  10877=>"111000000",
  10878=>"000000000",
  10879=>"111111111",
  10880=>"110111111",
  10881=>"100111111",
  10882=>"000000111",
  10883=>"000000111",
  10884=>"111111111",
  10885=>"000000111",
  10886=>"111001000",
  10887=>"000011000",
  10888=>"000000000",
  10889=>"111000000",
  10890=>"000000000",
  10891=>"000000000",
  10892=>"010110101",
  10893=>"110111111",
  10894=>"111111111",
  10895=>"111110100",
  10896=>"111111111",
  10897=>"000000000",
  10898=>"111110000",
  10899=>"001011111",
  10900=>"111101000",
  10901=>"011011111",
  10902=>"111111111",
  10903=>"111111111",
  10904=>"000000111",
  10905=>"111111111",
  10906=>"000110011",
  10907=>"011000111",
  10908=>"111100000",
  10909=>"000111111",
  10910=>"101101101",
  10911=>"000100111",
  10912=>"111111110",
  10913=>"111111111",
  10914=>"000000111",
  10915=>"111111100",
  10916=>"000000000",
  10917=>"111000001",
  10918=>"000001000",
  10919=>"101111011",
  10920=>"000100111",
  10921=>"000101111",
  10922=>"000000000",
  10923=>"000000000",
  10924=>"001111111",
  10925=>"000101111",
  10926=>"101100000",
  10927=>"111111100",
  10928=>"000011111",
  10929=>"100000001",
  10930=>"111111010",
  10931=>"111111011",
  10932=>"101000000",
  10933=>"000000000",
  10934=>"011010000",
  10935=>"111111111",
  10936=>"111111111",
  10937=>"111110000",
  10938=>"010000100",
  10939=>"000100101",
  10940=>"111011000",
  10941=>"111111000",
  10942=>"111001011",
  10943=>"100111111",
  10944=>"111111000",
  10945=>"001111111",
  10946=>"111111001",
  10947=>"000110011",
  10948=>"000010011",
  10949=>"000000000",
  10950=>"111111000",
  10951=>"001111111",
  10952=>"111111111",
  10953=>"111111111",
  10954=>"111111111",
  10955=>"111111111",
  10956=>"000000111",
  10957=>"000111111",
  10958=>"000000000",
  10959=>"010010000",
  10960=>"000001111",
  10961=>"111111111",
  10962=>"001001111",
  10963=>"000000000",
  10964=>"111111000",
  10965=>"111000100",
  10966=>"001111101",
  10967=>"000000000",
  10968=>"110100000",
  10969=>"010111111",
  10970=>"000000000",
  10971=>"000000000",
  10972=>"001101001",
  10973=>"000100111",
  10974=>"111111100",
  10975=>"000000000",
  10976=>"000000000",
  10977=>"010011011",
  10978=>"111100000",
  10979=>"111111111",
  10980=>"001111111",
  10981=>"000000000",
  10982=>"001011011",
  10983=>"011111111",
  10984=>"000001000",
  10985=>"000000000",
  10986=>"000000001",
  10987=>"000000000",
  10988=>"000000000",
  10989=>"111110000",
  10990=>"110010111",
  10991=>"101111111",
  10992=>"000111111",
  10993=>"110110111",
  10994=>"111111111",
  10995=>"111111000",
  10996=>"000000000",
  10997=>"101111111",
  10998=>"100111111",
  10999=>"000000000",
  11000=>"000000000",
  11001=>"001000000",
  11002=>"100100111",
  11003=>"000000011",
  11004=>"111111111",
  11005=>"011111111",
  11006=>"000000110",
  11007=>"111111111",
  11008=>"101100110",
  11009=>"001111011",
  11010=>"111111111",
  11011=>"000000001",
  11012=>"111111101",
  11013=>"100001101",
  11014=>"111100110",
  11015=>"100100111",
  11016=>"000000111",
  11017=>"000010110",
  11018=>"111000000",
  11019=>"000000100",
  11020=>"000000111",
  11021=>"000000000",
  11022=>"001001101",
  11023=>"100100000",
  11024=>"111111111",
  11025=>"001000100",
  11026=>"000001011",
  11027=>"000000011",
  11028=>"000000111",
  11029=>"110111111",
  11030=>"111111101",
  11031=>"011111111",
  11032=>"000001111",
  11033=>"000100101",
  11034=>"001011000",
  11035=>"000011000",
  11036=>"111111111",
  11037=>"111111000",
  11038=>"111111111",
  11039=>"000000001",
  11040=>"111100000",
  11041=>"000100110",
  11042=>"000111111",
  11043=>"000000011",
  11044=>"111111111",
  11045=>"111011000",
  11046=>"000001001",
  11047=>"110000000",
  11048=>"111111111",
  11049=>"111111111",
  11050=>"000101101",
  11051=>"000111111",
  11052=>"111111001",
  11053=>"000101100",
  11054=>"101011111",
  11055=>"000000000",
  11056=>"001011111",
  11057=>"000000100",
  11058=>"000000000",
  11059=>"000000000",
  11060=>"000000000",
  11061=>"000010111",
  11062=>"111111111",
  11063=>"010000000",
  11064=>"010000000",
  11065=>"111000000",
  11066=>"111111111",
  11067=>"010010000",
  11068=>"001000101",
  11069=>"001000001",
  11070=>"111000000",
  11071=>"000000000",
  11072=>"111100000",
  11073=>"111100110",
  11074=>"100111111",
  11075=>"000111111",
  11076=>"000000111",
  11077=>"111111111",
  11078=>"010000111",
  11079=>"000000000",
  11080=>"011111111",
  11081=>"000000000",
  11082=>"000100111",
  11083=>"010010111",
  11084=>"010000000",
  11085=>"001111111",
  11086=>"000000111",
  11087=>"000001001",
  11088=>"001101000",
  11089=>"000100111",
  11090=>"111110111",
  11091=>"000100111",
  11092=>"000000001",
  11093=>"001001001",
  11094=>"000000000",
  11095=>"000000111",
  11096=>"000110110",
  11097=>"000000000",
  11098=>"111001000",
  11099=>"100001001",
  11100=>"000000101",
  11101=>"101101100",
  11102=>"000000000",
  11103=>"001000000",
  11104=>"000001111",
  11105=>"000000000",
  11106=>"111011011",
  11107=>"000000000",
  11108=>"110111100",
  11109=>"001111111",
  11110=>"000000000",
  11111=>"000011111",
  11112=>"110110101",
  11113=>"000010111",
  11114=>"000000000",
  11115=>"000111011",
  11116=>"000000001",
  11117=>"010000000",
  11118=>"000000000",
  11119=>"001000000",
  11120=>"000000000",
  11121=>"011110111",
  11122=>"111010000",
  11123=>"111000000",
  11124=>"111111110",
  11125=>"111000110",
  11126=>"111111111",
  11127=>"010111111",
  11128=>"111111111",
  11129=>"000000000",
  11130=>"000000000",
  11131=>"001001100",
  11132=>"111111111",
  11133=>"110000110",
  11134=>"000101001",
  11135=>"000000000",
  11136=>"111001111",
  11137=>"110110110",
  11138=>"000100000",
  11139=>"000000000",
  11140=>"000011111",
  11141=>"000000000",
  11142=>"000000011",
  11143=>"111111000",
  11144=>"000000001",
  11145=>"111011001",
  11146=>"111111111",
  11147=>"111111000",
  11148=>"100000000",
  11149=>"000000000",
  11150=>"000000111",
  11151=>"100000110",
  11152=>"001000000",
  11153=>"111110100",
  11154=>"011111111",
  11155=>"000000000",
  11156=>"110110111",
  11157=>"011011000",
  11158=>"000100001",
  11159=>"100100000",
  11160=>"110000100",
  11161=>"001000010",
  11162=>"111111111",
  11163=>"111101101",
  11164=>"111100111",
  11165=>"110110111",
  11166=>"000000000",
  11167=>"100100110",
  11168=>"000000000",
  11169=>"110111111",
  11170=>"101100000",
  11171=>"000000011",
  11172=>"111001011",
  11173=>"000000011",
  11174=>"000000000",
  11175=>"111011000",
  11176=>"001001000",
  11177=>"000000001",
  11178=>"111111111",
  11179=>"111000000",
  11180=>"111111110",
  11181=>"000001000",
  11182=>"000000111",
  11183=>"111111111",
  11184=>"111111110",
  11185=>"111111110",
  11186=>"010111111",
  11187=>"000101111",
  11188=>"110111101",
  11189=>"111111001",
  11190=>"111111001",
  11191=>"000000000",
  11192=>"000000000",
  11193=>"000000000",
  11194=>"111000000",
  11195=>"111111100",
  11196=>"111001011",
  11197=>"101001001",
  11198=>"110110111",
  11199=>"111110100",
  11200=>"000000000",
  11201=>"111111000",
  11202=>"000111111",
  11203=>"110111110",
  11204=>"110111111",
  11205=>"001000110",
  11206=>"111111110",
  11207=>"111111111",
  11208=>"000000000",
  11209=>"111011000",
  11210=>"000000001",
  11211=>"001000000",
  11212=>"111100000",
  11213=>"010110110",
  11214=>"111111001",
  11215=>"000010011",
  11216=>"000111111",
  11217=>"001000000",
  11218=>"011011111",
  11219=>"000111111",
  11220=>"111111100",
  11221=>"111111111",
  11222=>"001111111",
  11223=>"110000000",
  11224=>"111111111",
  11225=>"001111000",
  11226=>"000110111",
  11227=>"001011011",
  11228=>"000111111",
  11229=>"111001100",
  11230=>"000000000",
  11231=>"000100100",
  11232=>"011011111",
  11233=>"000100110",
  11234=>"111111000",
  11235=>"111011000",
  11236=>"101100000",
  11237=>"001111111",
  11238=>"000001001",
  11239=>"010110010",
  11240=>"010111111",
  11241=>"011110000",
  11242=>"000110111",
  11243=>"100000000",
  11244=>"000111111",
  11245=>"000000000",
  11246=>"111111111",
  11247=>"100000000",
  11248=>"111111000",
  11249=>"000111111",
  11250=>"100000011",
  11251=>"110000111",
  11252=>"110111111",
  11253=>"001001001",
  11254=>"111001000",
  11255=>"011011011",
  11256=>"111111111",
  11257=>"001101110",
  11258=>"001001101",
  11259=>"111111000",
  11260=>"001011001",
  11261=>"110000000",
  11262=>"001101111",
  11263=>"111110100",
  11264=>"100000000",
  11265=>"001000000",
  11266=>"111101101",
  11267=>"000000001",
  11268=>"001100100",
  11269=>"010000100",
  11270=>"111011000",
  11271=>"000000000",
  11272=>"111111000",
  11273=>"111111111",
  11274=>"000001111",
  11275=>"111111111",
  11276=>"110111111",
  11277=>"011110111",
  11278=>"100000000",
  11279=>"011011000",
  11280=>"000100001",
  11281=>"100111111",
  11282=>"010000001",
  11283=>"010000000",
  11284=>"110000000",
  11285=>"111000101",
  11286=>"110111000",
  11287=>"001001011",
  11288=>"110100100",
  11289=>"001001001",
  11290=>"000000000",
  11291=>"001000000",
  11292=>"111111111",
  11293=>"100111111",
  11294=>"010001001",
  11295=>"100100101",
  11296=>"000010011",
  11297=>"000000010",
  11298=>"100111110",
  11299=>"111111011",
  11300=>"111111110",
  11301=>"000000111",
  11302=>"000001111",
  11303=>"101101000",
  11304=>"000000000",
  11305=>"000111010",
  11306=>"000000100",
  11307=>"010111110",
  11308=>"000000000",
  11309=>"000111110",
  11310=>"000001111",
  11311=>"000000000",
  11312=>"100111101",
  11313=>"000011011",
  11314=>"011101101",
  11315=>"111101011",
  11316=>"000001000",
  11317=>"011000000",
  11318=>"111111110",
  11319=>"000000000",
  11320=>"111010011",
  11321=>"000000100",
  11322=>"011111111",
  11323=>"000111111",
  11324=>"111111000",
  11325=>"111001001",
  11326=>"110110000",
  11327=>"001000001",
  11328=>"000000000",
  11329=>"000110000",
  11330=>"111111111",
  11331=>"111010001",
  11332=>"110110110",
  11333=>"011111111",
  11334=>"111000000",
  11335=>"111111001",
  11336=>"011111001",
  11337=>"111000000",
  11338=>"000111010",
  11339=>"000000001",
  11340=>"111111110",
  11341=>"010010001",
  11342=>"001011111",
  11343=>"000000000",
  11344=>"000000110",
  11345=>"000100111",
  11346=>"111111111",
  11347=>"000100100",
  11348=>"001111101",
  11349=>"111111000",
  11350=>"111110000",
  11351=>"100110000",
  11352=>"101111111",
  11353=>"111101101",
  11354=>"010000000",
  11355=>"001000000",
  11356=>"111000000",
  11357=>"100100111",
  11358=>"111100000",
  11359=>"011011011",
  11360=>"100111111",
  11361=>"000000000",
  11362=>"010110111",
  11363=>"000000000",
  11364=>"111111000",
  11365=>"000000001",
  11366=>"111001100",
  11367=>"110100100",
  11368=>"000111111",
  11369=>"000000000",
  11370=>"111111010",
  11371=>"000000000",
  11372=>"011111111",
  11373=>"000110010",
  11374=>"100000101",
  11375=>"011111100",
  11376=>"111111011",
  11377=>"101100111",
  11378=>"101001000",
  11379=>"000000000",
  11380=>"001001000",
  11381=>"000000110",
  11382=>"000000111",
  11383=>"001001101",
  11384=>"100111111",
  11385=>"011111110",
  11386=>"110100100",
  11387=>"111000000",
  11388=>"111110100",
  11389=>"111111111",
  11390=>"100100000",
  11391=>"001001001",
  11392=>"011111111",
  11393=>"000000110",
  11394=>"110000000",
  11395=>"110111000",
  11396=>"001000011",
  11397=>"111100000",
  11398=>"110000011",
  11399=>"101100101",
  11400=>"000000000",
  11401=>"000001111",
  11402=>"111111111",
  11403=>"001001011",
  11404=>"000110100",
  11405=>"101000000",
  11406=>"000000000",
  11407=>"001000011",
  11408=>"000000100",
  11409=>"011111011",
  11410=>"000011111",
  11411=>"111111111",
  11412=>"001011110",
  11413=>"000000110",
  11414=>"010111111",
  11415=>"000000000",
  11416=>"001000000",
  11417=>"100000000",
  11418=>"111100000",
  11419=>"111111111",
  11420=>"110000000",
  11421=>"000000000",
  11422=>"111111111",
  11423=>"000111000",
  11424=>"000001001",
  11425=>"000001001",
  11426=>"000111111",
  11427=>"111000001",
  11428=>"001001001",
  11429=>"111111111",
  11430=>"000000000",
  11431=>"000101111",
  11432=>"000000000",
  11433=>"000000000",
  11434=>"000000000",
  11435=>"011111111",
  11436=>"111111111",
  11437=>"111110100",
  11438=>"111100000",
  11439=>"000000101",
  11440=>"000000111",
  11441=>"111001001",
  11442=>"000111111",
  11443=>"101111111",
  11444=>"100101111",
  11445=>"110111111",
  11446=>"010001100",
  11447=>"101000011",
  11448=>"001011101",
  11449=>"000000000",
  11450=>"110100000",
  11451=>"001001101",
  11452=>"111110100",
  11453=>"000000001",
  11454=>"111100010",
  11455=>"111101000",
  11456=>"100000000",
  11457=>"001000001",
  11458=>"001100101",
  11459=>"001100000",
  11460=>"001000111",
  11461=>"000000000",
  11462=>"000000000",
  11463=>"110100100",
  11464=>"000001011",
  11465=>"111111111",
  11466=>"000100100",
  11467=>"001000000",
  11468=>"110111100",
  11469=>"000001000",
  11470=>"111101111",
  11471=>"001000101",
  11472=>"011011111",
  11473=>"001000111",
  11474=>"000001011",
  11475=>"001011000",
  11476=>"000001001",
  11477=>"000000000",
  11478=>"000000000",
  11479=>"000000001",
  11480=>"011001111",
  11481=>"111111111",
  11482=>"000110110",
  11483=>"000000000",
  11484=>"001000111",
  11485=>"100111111",
  11486=>"000000000",
  11487=>"111010010",
  11488=>"000000011",
  11489=>"000000000",
  11490=>"000110110",
  11491=>"110100110",
  11492=>"100110111",
  11493=>"000000000",
  11494=>"110011000",
  11495=>"111000101",
  11496=>"111111000",
  11497=>"111111011",
  11498=>"001111000",
  11499=>"001000011",
  11500=>"001001111",
  11501=>"000000000",
  11502=>"111011111",
  11503=>"001000101",
  11504=>"000000000",
  11505=>"011000000",
  11506=>"011111111",
  11507=>"000001001",
  11508=>"111111111",
  11509=>"000100100",
  11510=>"001001011",
  11511=>"000100000",
  11512=>"000110010",
  11513=>"000000101",
  11514=>"111111111",
  11515=>"000010000",
  11516=>"000000000",
  11517=>"111000000",
  11518=>"000000100",
  11519=>"000111111",
  11520=>"100100111",
  11521=>"111100101",
  11522=>"111111111",
  11523=>"000000000",
  11524=>"010000000",
  11525=>"011000000",
  11526=>"111111000",
  11527=>"001000001",
  11528=>"001001000",
  11529=>"100100111",
  11530=>"000000001",
  11531=>"111111001",
  11532=>"100000000",
  11533=>"000000000",
  11534=>"000000000",
  11535=>"000000000",
  11536=>"011111110",
  11537=>"000000000",
  11538=>"000010111",
  11539=>"000010000",
  11540=>"000000010",
  11541=>"000100111",
  11542=>"000100100",
  11543=>"111111100",
  11544=>"000000001",
  11545=>"111111111",
  11546=>"011000100",
  11547=>"111000000",
  11548=>"110111101",
  11549=>"000000000",
  11550=>"000000000",
  11551=>"000000100",
  11552=>"001000000",
  11553=>"100000100",
  11554=>"110111111",
  11555=>"001001000",
  11556=>"010000000",
  11557=>"110111111",
  11558=>"000001111",
  11559=>"101000000",
  11560=>"000000100",
  11561=>"111111010",
  11562=>"000000111",
  11563=>"000010001",
  11564=>"001000000",
  11565=>"110000000",
  11566=>"111111111",
  11567=>"111110111",
  11568=>"111111111",
  11569=>"111100100",
  11570=>"111111110",
  11571=>"011011000",
  11572=>"111001000",
  11573=>"011001000",
  11574=>"000000000",
  11575=>"101000100",
  11576=>"010010000",
  11577=>"000000011",
  11578=>"000000101",
  11579=>"000000000",
  11580=>"110110111",
  11581=>"111111111",
  11582=>"100100101",
  11583=>"001011111",
  11584=>"100111111",
  11585=>"000000000",
  11586=>"001000110",
  11587=>"000001101",
  11588=>"000000000",
  11589=>"000000011",
  11590=>"110110010",
  11591=>"110111110",
  11592=>"111111100",
  11593=>"010011111",
  11594=>"010111111",
  11595=>"010100010",
  11596=>"000000111",
  11597=>"011001000",
  11598=>"100111111",
  11599=>"000000000",
  11600=>"011010111",
  11601=>"000000111",
  11602=>"011011011",
  11603=>"000000111",
  11604=>"100100100",
  11605=>"011011000",
  11606=>"000000000",
  11607=>"011001111",
  11608=>"000000000",
  11609=>"001001111",
  11610=>"111111111",
  11611=>"000000000",
  11612=>"000000000",
  11613=>"000000100",
  11614=>"011111111",
  11615=>"111011001",
  11616=>"111011000",
  11617=>"011000001",
  11618=>"000011011",
  11619=>"111101000",
  11620=>"000000000",
  11621=>"011000000",
  11622=>"000000000",
  11623=>"111111110",
  11624=>"001101101",
  11625=>"000011111",
  11626=>"000001111",
  11627=>"010011111",
  11628=>"001001000",
  11629=>"110111011",
  11630=>"010111111",
  11631=>"100111111",
  11632=>"000000100",
  11633=>"111000000",
  11634=>"000000111",
  11635=>"111101100",
  11636=>"010011011",
  11637=>"111111111",
  11638=>"111111100",
  11639=>"000000000",
  11640=>"111011000",
  11641=>"111101111",
  11642=>"001000000",
  11643=>"111010010",
  11644=>"010000011",
  11645=>"101000000",
  11646=>"011000000",
  11647=>"101000000",
  11648=>"110111110",
  11649=>"000000000",
  11650=>"111111011",
  11651=>"000000000",
  11652=>"111111111",
  11653=>"111111111",
  11654=>"011010000",
  11655=>"011011111",
  11656=>"110000000",
  11657=>"110000111",
  11658=>"000101111",
  11659=>"000111111",
  11660=>"011000001",
  11661=>"110100100",
  11662=>"101101110",
  11663=>"100000000",
  11664=>"000000000",
  11665=>"111111111",
  11666=>"000000100",
  11667=>"001001010",
  11668=>"111100111",
  11669=>"000011000",
  11670=>"111111011",
  11671=>"111001001",
  11672=>"000000101",
  11673=>"010111111",
  11674=>"111111001",
  11675=>"111111111",
  11676=>"111111111",
  11677=>"100100100",
  11678=>"100000000",
  11679=>"111111000",
  11680=>"000000000",
  11681=>"101000000",
  11682=>"100000000",
  11683=>"010111000",
  11684=>"100111010",
  11685=>"000100000",
  11686=>"101111111",
  11687=>"011111111",
  11688=>"111001101",
  11689=>"000110000",
  11690=>"111111111",
  11691=>"111111111",
  11692=>"000000000",
  11693=>"111111111",
  11694=>"000000001",
  11695=>"000011111",
  11696=>"001000111",
  11697=>"000000111",
  11698=>"011111110",
  11699=>"001101000",
  11700=>"111101111",
  11701=>"000000001",
  11702=>"011011111",
  11703=>"010010010",
  11704=>"000000000",
  11705=>"111111101",
  11706=>"111111111",
  11707=>"011111111",
  11708=>"000000110",
  11709=>"111011111",
  11710=>"000000000",
  11711=>"000100100",
  11712=>"111111111",
  11713=>"100101101",
  11714=>"111001111",
  11715=>"100101111",
  11716=>"111011001",
  11717=>"000000000",
  11718=>"000000000",
  11719=>"000000000",
  11720=>"110000000",
  11721=>"000000000",
  11722=>"001000000",
  11723=>"000111011",
  11724=>"100110000",
  11725=>"111111111",
  11726=>"001001111",
  11727=>"000000000",
  11728=>"011011000",
  11729=>"100001001",
  11730=>"000000000",
  11731=>"100100111",
  11732=>"110111100",
  11733=>"111111010",
  11734=>"000111111",
  11735=>"111111001",
  11736=>"101111101",
  11737=>"111111111",
  11738=>"111000001",
  11739=>"011010011",
  11740=>"011100111",
  11741=>"001000000",
  11742=>"111111000",
  11743=>"111111001",
  11744=>"000100100",
  11745=>"000000111",
  11746=>"000011111",
  11747=>"000000111",
  11748=>"000010111",
  11749=>"111001000",
  11750=>"011000000",
  11751=>"111110110",
  11752=>"110110111",
  11753=>"111111001",
  11754=>"110000000",
  11755=>"111101111",
  11756=>"001000101",
  11757=>"111011001",
  11758=>"100100101",
  11759=>"101001000",
  11760=>"110100001",
  11761=>"010110111",
  11762=>"001001111",
  11763=>"111000001",
  11764=>"111100110",
  11765=>"000000001",
  11766=>"111100000",
  11767=>"111111110",
  11768=>"001111011",
  11769=>"000001001",
  11770=>"111111111",
  11771=>"011000101",
  11772=>"111110000",
  11773=>"001000000",
  11774=>"100101101",
  11775=>"001000101",
  11776=>"010010010",
  11777=>"111111111",
  11778=>"000111111",
  11779=>"000000111",
  11780=>"000000110",
  11781=>"101111111",
  11782=>"000000000",
  11783=>"010000111",
  11784=>"111000000",
  11785=>"000000000",
  11786=>"000000000",
  11787=>"001000000",
  11788=>"111100000",
  11789=>"111110111",
  11790=>"001000000",
  11791=>"000000000",
  11792=>"111010000",
  11793=>"000000001",
  11794=>"111011000",
  11795=>"001000000",
  11796=>"000000001",
  11797=>"110111111",
  11798=>"000000000",
  11799=>"111111111",
  11800=>"100111111",
  11801=>"011000000",
  11802=>"100000000",
  11803=>"111111111",
  11804=>"111110000",
  11805=>"000111111",
  11806=>"111011011",
  11807=>"000000000",
  11808=>"111000000",
  11809=>"111110011",
  11810=>"111111000",
  11811=>"000000101",
  11812=>"111111000",
  11813=>"000000011",
  11814=>"111001000",
  11815=>"111111111",
  11816=>"011001001",
  11817=>"111001000",
  11818=>"000000000",
  11819=>"000111111",
  11820=>"111111000",
  11821=>"000101111",
  11822=>"111001000",
  11823=>"110110111",
  11824=>"111000111",
  11825=>"000000000",
  11826=>"011111111",
  11827=>"000000000",
  11828=>"100111000",
  11829=>"011011011",
  11830=>"000001011",
  11831=>"111000000",
  11832=>"111000000",
  11833=>"001101000",
  11834=>"111000000",
  11835=>"000000000",
  11836=>"100000000",
  11837=>"100111011",
  11838=>"000001111",
  11839=>"111000000",
  11840=>"011011000",
  11841=>"111111111",
  11842=>"000111111",
  11843=>"000000000",
  11844=>"000000000",
  11845=>"111110110",
  11846=>"000000001",
  11847=>"111111111",
  11848=>"011110000",
  11849=>"000000111",
  11850=>"000100100",
  11851=>"000000110",
  11852=>"100100111",
  11853=>"111110000",
  11854=>"000000000",
  11855=>"111111111",
  11856=>"111111111",
  11857=>"000011000",
  11858=>"111111111",
  11859=>"111111111",
  11860=>"000000000",
  11861=>"000000000",
  11862=>"100000011",
  11863=>"100100000",
  11864=>"111111111",
  11865=>"100100111",
  11866=>"000010110",
  11867=>"010000001",
  11868=>"000000111",
  11869=>"000000100",
  11870=>"110110111",
  11871=>"100111111",
  11872=>"100100001",
  11873=>"100000000",
  11874=>"111000000",
  11875=>"110001001",
  11876=>"000000000",
  11877=>"000000110",
  11878=>"110111111",
  11879=>"000101111",
  11880=>"000100100",
  11881=>"000100100",
  11882=>"111111010",
  11883=>"000010000",
  11884=>"000110111",
  11885=>"000000000",
  11886=>"111000000",
  11887=>"111111011",
  11888=>"111001000",
  11889=>"000000111",
  11890=>"100101001",
  11891=>"001011000",
  11892=>"110000000",
  11893=>"111111110",
  11894=>"000000001",
  11895=>"000000000",
  11896=>"000000000",
  11897=>"111111111",
  11898=>"000000000",
  11899=>"000000100",
  11900=>"111111110",
  11901=>"011111000",
  11902=>"011100000",
  11903=>"000000000",
  11904=>"000000000",
  11905=>"111111111",
  11906=>"111110000",
  11907=>"001111000",
  11908=>"111100000",
  11909=>"000000111",
  11910=>"110110110",
  11911=>"100000110",
  11912=>"110110100",
  11913=>"110110111",
  11914=>"111100101",
  11915=>"011111111",
  11916=>"111111011",
  11917=>"000000000",
  11918=>"110110000",
  11919=>"000000000",
  11920=>"000111111",
  11921=>"000000001",
  11922=>"110010000",
  11923=>"111000000",
  11924=>"000110110",
  11925=>"111111101",
  11926=>"110010010",
  11927=>"111111100",
  11928=>"001111111",
  11929=>"100111111",
  11930=>"000000000",
  11931=>"000000000",
  11932=>"111111000",
  11933=>"000110110",
  11934=>"000000110",
  11935=>"011111111",
  11936=>"000111001",
  11937=>"000000000",
  11938=>"000000111",
  11939=>"111111001",
  11940=>"000001011",
  11941=>"100000101",
  11942=>"111111111",
  11943=>"010111110",
  11944=>"111111110",
  11945=>"010110111",
  11946=>"001000000",
  11947=>"000000000",
  11948=>"010111110",
  11949=>"111111001",
  11950=>"111111000",
  11951=>"000000000",
  11952=>"000000000",
  11953=>"110110011",
  11954=>"111111011",
  11955=>"111000000",
  11956=>"111111111",
  11957=>"011011000",
  11958=>"111001000",
  11959=>"111111111",
  11960=>"000000001",
  11961=>"111111111",
  11962=>"000000000",
  11963=>"011010010",
  11964=>"000000000",
  11965=>"111111101",
  11966=>"000000000",
  11967=>"111010000",
  11968=>"000000000",
  11969=>"000000001",
  11970=>"000000000",
  11971=>"000001111",
  11972=>"000111111",
  11973=>"111101000",
  11974=>"000001001",
  11975=>"111101000",
  11976=>"011011110",
  11977=>"111111001",
  11978=>"101111001",
  11979=>"111111110",
  11980=>"111100000",
  11981=>"000100111",
  11982=>"111111111",
  11983=>"000000100",
  11984=>"111000000",
  11985=>"000001111",
  11986=>"111110111",
  11987=>"000000100",
  11988=>"000111111",
  11989=>"111111111",
  11990=>"000010111",
  11991=>"001000010",
  11992=>"101101111",
  11993=>"001101111",
  11994=>"111001111",
  11995=>"111111111",
  11996=>"100100111",
  11997=>"001000001",
  11998=>"000000011",
  11999=>"110111000",
  12000=>"111000000",
  12001=>"110000000",
  12002=>"010000000",
  12003=>"111111000",
  12004=>"011000000",
  12005=>"111111111",
  12006=>"000100110",
  12007=>"111101101",
  12008=>"000000000",
  12009=>"111110000",
  12010=>"111011001",
  12011=>"100000000",
  12012=>"111111111",
  12013=>"101100111",
  12014=>"111110010",
  12015=>"000000111",
  12016=>"110111111",
  12017=>"000000011",
  12018=>"000000000",
  12019=>"000001101",
  12020=>"110111111",
  12021=>"100111111",
  12022=>"100100100",
  12023=>"111111111",
  12024=>"000100111",
  12025=>"111111000",
  12026=>"000000000",
  12027=>"000011101",
  12028=>"111101101",
  12029=>"111011000",
  12030=>"001000000",
  12031=>"000000100",
  12032=>"000111000",
  12033=>"111101011",
  12034=>"000000001",
  12035=>"000000101",
  12036=>"111101101",
  12037=>"110111111",
  12038=>"000000000",
  12039=>"000000110",
  12040=>"101001001",
  12041=>"110000000",
  12042=>"101100000",
  12043=>"001001000",
  12044=>"111111000",
  12045=>"111000000",
  12046=>"000000111",
  12047=>"000000000",
  12048=>"101111111",
  12049=>"000000001",
  12050=>"111011000",
  12051=>"000000000",
  12052=>"000000000",
  12053=>"001000000",
  12054=>"111111101",
  12055=>"110111110",
  12056=>"000000000",
  12057=>"000000000",
  12058=>"000100111",
  12059=>"110111111",
  12060=>"100111111",
  12061=>"111111111",
  12062=>"001001011",
  12063=>"011001101",
  12064=>"000000000",
  12065=>"000000011",
  12066=>"000000111",
  12067=>"111111111",
  12068=>"111001000",
  12069=>"111111011",
  12070=>"011111111",
  12071=>"000000100",
  12072=>"110111111",
  12073=>"011011000",
  12074=>"111101000",
  12075=>"000000000",
  12076=>"001000000",
  12077=>"001001001",
  12078=>"101000011",
  12079=>"000000011",
  12080=>"111111111",
  12081=>"111111111",
  12082=>"000000000",
  12083=>"111000000",
  12084=>"000000111",
  12085=>"000000000",
  12086=>"101001101",
  12087=>"000000000",
  12088=>"111111100",
  12089=>"111110000",
  12090=>"000000000",
  12091=>"000000000",
  12092=>"000000000",
  12093=>"000100111",
  12094=>"000111111",
  12095=>"111111111",
  12096=>"000010011",
  12097=>"111111111",
  12098=>"001000000",
  12099=>"111111111",
  12100=>"000000000",
  12101=>"000000111",
  12102=>"000000111",
  12103=>"010011010",
  12104=>"000000000",
  12105=>"111011001",
  12106=>"111101101",
  12107=>"111011000",
  12108=>"000000000",
  12109=>"110011111",
  12110=>"111111111",
  12111=>"111111111",
  12112=>"110111010",
  12113=>"001000000",
  12114=>"000000000",
  12115=>"111111110",
  12116=>"100111111",
  12117=>"111011001",
  12118=>"111000000",
  12119=>"011011011",
  12120=>"111111111",
  12121=>"100000111",
  12122=>"100000000",
  12123=>"111111000",
  12124=>"000000111",
  12125=>"111111001",
  12126=>"100101101",
  12127=>"111111111",
  12128=>"001100111",
  12129=>"111111101",
  12130=>"110100100",
  12131=>"111111111",
  12132=>"100110110",
  12133=>"000000101",
  12134=>"000000001",
  12135=>"111111111",
  12136=>"110100111",
  12137=>"110000000",
  12138=>"111111111",
  12139=>"000011111",
  12140=>"011111111",
  12141=>"010111101",
  12142=>"100000000",
  12143=>"010000110",
  12144=>"010010111",
  12145=>"111111111",
  12146=>"111110000",
  12147=>"111110000",
  12148=>"000000001",
  12149=>"111111111",
  12150=>"011111011",
  12151=>"110100100",
  12152=>"000111111",
  12153=>"000011111",
  12154=>"100101101",
  12155=>"111111111",
  12156=>"111001111",
  12157=>"101111011",
  12158=>"001001001",
  12159=>"000110111",
  12160=>"011011111",
  12161=>"111111001",
  12162=>"011011011",
  12163=>"110000000",
  12164=>"111110000",
  12165=>"000110111",
  12166=>"011010000",
  12167=>"111100000",
  12168=>"111111111",
  12169=>"110000000",
  12170=>"111111111",
  12171=>"111000000",
  12172=>"111111111",
  12173=>"101100111",
  12174=>"111111111",
  12175=>"111111111",
  12176=>"000010011",
  12177=>"111111111",
  12178=>"111111100",
  12179=>"001000001",
  12180=>"111111000",
  12181=>"000000000",
  12182=>"001001011",
  12183=>"011001000",
  12184=>"000000001",
  12185=>"110010011",
  12186=>"000000000",
  12187=>"001000000",
  12188=>"001001000",
  12189=>"000000001",
  12190=>"110110110",
  12191=>"000000000",
  12192=>"001111000",
  12193=>"111100110",
  12194=>"101101111",
  12195=>"000010111",
  12196=>"111101000",
  12197=>"111111111",
  12198=>"111011111",
  12199=>"000111111",
  12200=>"111000000",
  12201=>"000000111",
  12202=>"000000110",
  12203=>"000100101",
  12204=>"111111001",
  12205=>"000000011",
  12206=>"000000000",
  12207=>"000000000",
  12208=>"000000000",
  12209=>"101100100",
  12210=>"000000111",
  12211=>"110110111",
  12212=>"000000000",
  12213=>"110010111",
  12214=>"111111111",
  12215=>"000000000",
  12216=>"111111000",
  12217=>"111011000",
  12218=>"000000111",
  12219=>"001000000",
  12220=>"010000000",
  12221=>"111111111",
  12222=>"101111101",
  12223=>"111001011",
  12224=>"000000000",
  12225=>"000001111",
  12226=>"011011111",
  12227=>"010110111",
  12228=>"100000000",
  12229=>"110110111",
  12230=>"001101111",
  12231=>"000001111",
  12232=>"001001111",
  12233=>"001101111",
  12234=>"101101111",
  12235=>"000000000",
  12236=>"000000000",
  12237=>"111101100",
  12238=>"111111111",
  12239=>"000011111",
  12240=>"000101111",
  12241=>"110111111",
  12242=>"001111111",
  12243=>"000000000",
  12244=>"111011000",
  12245=>"111011000",
  12246=>"000000011",
  12247=>"001101000",
  12248=>"111111111",
  12249=>"000000100",
  12250=>"000001001",
  12251=>"111001000",
  12252=>"111111011",
  12253=>"111111111",
  12254=>"011111111",
  12255=>"000001000",
  12256=>"110111111",
  12257=>"000001001",
  12258=>"100000000",
  12259=>"011000000",
  12260=>"111111110",
  12261=>"011111000",
  12262=>"000000000",
  12263=>"000001011",
  12264=>"101000000",
  12265=>"000000111",
  12266=>"111111101",
  12267=>"111111111",
  12268=>"000000111",
  12269=>"111110100",
  12270=>"111000000",
  12271=>"100111111",
  12272=>"000010011",
  12273=>"111111000",
  12274=>"001000000",
  12275=>"001101101",
  12276=>"111111000",
  12277=>"110000001",
  12278=>"111111001",
  12279=>"111111111",
  12280=>"001111011",
  12281=>"110000000",
  12282=>"110111101",
  12283=>"001001001",
  12284=>"111111000",
  12285=>"111001001",
  12286=>"001000000",
  12287=>"000100111",
  12288=>"111111111",
  12289=>"110000000",
  12290=>"111111010",
  12291=>"010110111",
  12292=>"111111110",
  12293=>"011000000",
  12294=>"011111000",
  12295=>"111001000",
  12296=>"011000000",
  12297=>"110111111",
  12298=>"001000000",
  12299=>"111000000",
  12300=>"111111111",
  12301=>"000000111",
  12302=>"100100111",
  12303=>"010111010",
  12304=>"000001100",
  12305=>"000010000",
  12306=>"000000000",
  12307=>"000000000",
  12308=>"000000111",
  12309=>"111111111",
  12310=>"000000101",
  12311=>"000100100",
  12312=>"111111111",
  12313=>"111011011",
  12314=>"000100111",
  12315=>"000001000",
  12316=>"101101111",
  12317=>"011111000",
  12318=>"000000000",
  12319=>"100111111",
  12320=>"111111111",
  12321=>"010111111",
  12322=>"111111110",
  12323=>"000000000",
  12324=>"111001000",
  12325=>"000000111",
  12326=>"001000000",
  12327=>"000000111",
  12328=>"111101111",
  12329=>"111111111",
  12330=>"111111000",
  12331=>"100100010",
  12332=>"000000000",
  12333=>"000000100",
  12334=>"001000100",
  12335=>"000011011",
  12336=>"111111110",
  12337=>"111001000",
  12338=>"101100100",
  12339=>"000000111",
  12340=>"000000000",
  12341=>"111111000",
  12342=>"111001000",
  12343=>"111111111",
  12344=>"100111100",
  12345=>"000000000",
  12346=>"111101111",
  12347=>"111101111",
  12348=>"101001000",
  12349=>"001000000",
  12350=>"111000000",
  12351=>"111001000",
  12352=>"000000000",
  12353=>"000100100",
  12354=>"000000000",
  12355=>"000000001",
  12356=>"110111111",
  12357=>"001001111",
  12358=>"100111111",
  12359=>"001000000",
  12360=>"011111111",
  12361=>"111101111",
  12362=>"010111111",
  12363=>"000000001",
  12364=>"011000000",
  12365=>"110111000",
  12366=>"001001000",
  12367=>"001001000",
  12368=>"000000000",
  12369=>"010010000",
  12370=>"111111110",
  12371=>"011011100",
  12372=>"111110000",
  12373=>"000000000",
  12374=>"111000100",
  12375=>"101111111",
  12376=>"011000111",
  12377=>"111000011",
  12378=>"110010000",
  12379=>"000110111",
  12380=>"101000111",
  12381=>"111000000",
  12382=>"110000101",
  12383=>"000010010",
  12384=>"111100111",
  12385=>"001001111",
  12386=>"000000000",
  12387=>"100101100",
  12388=>"111110000",
  12389=>"111111100",
  12390=>"000000100",
  12391=>"111000000",
  12392=>"111011111",
  12393=>"000000000",
  12394=>"111011000",
  12395=>"111000000",
  12396=>"000010111",
  12397=>"000000000",
  12398=>"000001111",
  12399=>"111110000",
  12400=>"111000000",
  12401=>"111111000",
  12402=>"000000000",
  12403=>"111011000",
  12404=>"000000000",
  12405=>"100110111",
  12406=>"100110111",
  12407=>"010010000",
  12408=>"000000000",
  12409=>"001000000",
  12410=>"000000000",
  12411=>"100100100",
  12412=>"000000000",
  12413=>"011111111",
  12414=>"000000000",
  12415=>"111111000",
  12416=>"000111111",
  12417=>"000000110",
  12418=>"001000000",
  12419=>"011001001",
  12420=>"000000101",
  12421=>"000000000",
  12422=>"000000101",
  12423=>"000000000",
  12424=>"000000000",
  12425=>"000000000",
  12426=>"001100101",
  12427=>"000000110",
  12428=>"000001111",
  12429=>"111111100",
  12430=>"000000000",
  12431=>"000000000",
  12432=>"000000000",
  12433=>"000000000",
  12434=>"011000000",
  12435=>"000000001",
  12436=>"010000000",
  12437=>"001001111",
  12438=>"000110111",
  12439=>"000000000",
  12440=>"111000000",
  12441=>"111111111",
  12442=>"100100101",
  12443=>"111111001",
  12444=>"111111111",
  12445=>"111001000",
  12446=>"001000000",
  12447=>"000000111",
  12448=>"110111000",
  12449=>"011001000",
  12450=>"111111100",
  12451=>"111111011",
  12452=>"000000000",
  12453=>"111111111",
  12454=>"111111100",
  12455=>"101000000",
  12456=>"010111111",
  12457=>"000111111",
  12458=>"111110100",
  12459=>"111101000",
  12460=>"000000000",
  12461=>"000000001",
  12462=>"001000101",
  12463=>"111101000",
  12464=>"010111001",
  12465=>"111111010",
  12466=>"111111011",
  12467=>"111111000",
  12468=>"111111111",
  12469=>"001001010",
  12470=>"000000100",
  12471=>"000000010",
  12472=>"000010111",
  12473=>"001000011",
  12474=>"000000000",
  12475=>"110110010",
  12476=>"100100111",
  12477=>"000000111",
  12478=>"111111111",
  12479=>"001111111",
  12480=>"111101111",
  12481=>"000000000",
  12482=>"000000000",
  12483=>"110110100",
  12484=>"111101111",
  12485=>"000000000",
  12486=>"000000000",
  12487=>"111111111",
  12488=>"000011011",
  12489=>"000001111",
  12490=>"000000100",
  12491=>"011011011",
  12492=>"111111111",
  12493=>"110000000",
  12494=>"111110110",
  12495=>"000000101",
  12496=>"000011111",
  12497=>"010000000",
  12498=>"111111111",
  12499=>"000000000",
  12500=>"101000000",
  12501=>"110111111",
  12502=>"000000000",
  12503=>"111111100",
  12504=>"001101110",
  12505=>"111111111",
  12506=>"101101101",
  12507=>"111111111",
  12508=>"000110111",
  12509=>"101101111",
  12510=>"100000000",
  12511=>"000000000",
  12512=>"111100111",
  12513=>"010010000",
  12514=>"000000100",
  12515=>"001000000",
  12516=>"000000000",
  12517=>"001111111",
  12518=>"000000111",
  12519=>"111111111",
  12520=>"111010010",
  12521=>"011111111",
  12522=>"111111100",
  12523=>"110000100",
  12524=>"000000110",
  12525=>"111000001",
  12526=>"000000011",
  12527=>"000000000",
  12528=>"110100000",
  12529=>"000000011",
  12530=>"000111111",
  12531=>"000000111",
  12532=>"111111000",
  12533=>"000000010",
  12534=>"111111001",
  12535=>"111111000",
  12536=>"000000000",
  12537=>"111111111",
  12538=>"000000000",
  12539=>"111000000",
  12540=>"011011011",
  12541=>"000000000",
  12542=>"111000001",
  12543=>"000000000",
  12544=>"000100100",
  12545=>"100000001",
  12546=>"000000001",
  12547=>"111111110",
  12548=>"000001111",
  12549=>"000000111",
  12550=>"111111111",
  12551=>"111111011",
  12552=>"000000000",
  12553=>"000000000",
  12554=>"111111111",
  12555=>"011000011",
  12556=>"000000000",
  12557=>"101001000",
  12558=>"000000000",
  12559=>"000000000",
  12560=>"110111100",
  12561=>"000000000",
  12562=>"000000111",
  12563=>"111111111",
  12564=>"111101111",
  12565=>"000001000",
  12566=>"000000100",
  12567=>"000001001",
  12568=>"001111000",
  12569=>"110010000",
  12570=>"111111100",
  12571=>"000000000",
  12572=>"111111001",
  12573=>"000000111",
  12574=>"000000000",
  12575=>"101101111",
  12576=>"000110001",
  12577=>"010001111",
  12578=>"111111000",
  12579=>"111111111",
  12580=>"110110000",
  12581=>"100111111",
  12582=>"001000001",
  12583=>"000111001",
  12584=>"101101111",
  12585=>"111111100",
  12586=>"111111111",
  12587=>"111100100",
  12588=>"000111111",
  12589=>"000000001",
  12590=>"111000111",
  12591=>"000000111",
  12592=>"111111100",
  12593=>"111111000",
  12594=>"111101011",
  12595=>"111010000",
  12596=>"000001000",
  12597=>"001001101",
  12598=>"000011011",
  12599=>"001011111",
  12600=>"000011111",
  12601=>"001001111",
  12602=>"000000000",
  12603=>"000000101",
  12604=>"000000001",
  12605=>"000111111",
  12606=>"000001000",
  12607=>"000000100",
  12608=>"011111111",
  12609=>"111111000",
  12610=>"111111111",
  12611=>"111101001",
  12612=>"101111110",
  12613=>"001000000",
  12614=>"101110110",
  12615=>"000000000",
  12616=>"000000000",
  12617=>"011010111",
  12618=>"011101111",
  12619=>"000000000",
  12620=>"111011011",
  12621=>"111100000",
  12622=>"101100110",
  12623=>"000110100",
  12624=>"011111001",
  12625=>"000000110",
  12626=>"001000000",
  12627=>"100000100",
  12628=>"111011000",
  12629=>"011011001",
  12630=>"000000111",
  12631=>"111000100",
  12632=>"000000001",
  12633=>"000000000",
  12634=>"000000100",
  12635=>"111011110",
  12636=>"011011000",
  12637=>"000000111",
  12638=>"111111110",
  12639=>"011111011",
  12640=>"000000000",
  12641=>"111111000",
  12642=>"001000010",
  12643=>"111111011",
  12644=>"101111111",
  12645=>"000000000",
  12646=>"000000000",
  12647=>"000110101",
  12648=>"000000110",
  12649=>"110111111",
  12650=>"000000100",
  12651=>"000010110",
  12652=>"110111110",
  12653=>"001000000",
  12654=>"000001001",
  12655=>"001011000",
  12656=>"000000001",
  12657=>"110011011",
  12658=>"111000000",
  12659=>"001001001",
  12660=>"111111000",
  12661=>"110110111",
  12662=>"111111111",
  12663=>"110100000",
  12664=>"000000000",
  12665=>"101000111",
  12666=>"000011111",
  12667=>"100010010",
  12668=>"110111000",
  12669=>"001000111",
  12670=>"110000000",
  12671=>"001001011",
  12672=>"111001111",
  12673=>"000000000",
  12674=>"100111111",
  12675=>"000001101",
  12676=>"001001011",
  12677=>"010111110",
  12678=>"000001000",
  12679=>"111111111",
  12680=>"001000111",
  12681=>"000000001",
  12682=>"000000000",
  12683=>"010111000",
  12684=>"000000100",
  12685=>"111111000",
  12686=>"000000000",
  12687=>"000000000",
  12688=>"000000000",
  12689=>"111111011",
  12690=>"001000110",
  12691=>"001000000",
  12692=>"011011111",
  12693=>"010010010",
  12694=>"111110100",
  12695=>"000000000",
  12696=>"000000000",
  12697=>"100000000",
  12698=>"111111111",
  12699=>"001001111",
  12700=>"001000111",
  12701=>"111101000",
  12702=>"000000000",
  12703=>"110110000",
  12704=>"000111111",
  12705=>"011001011",
  12706=>"111100000",
  12707=>"000111111",
  12708=>"111111000",
  12709=>"111110000",
  12710=>"111111111",
  12711=>"111111011",
  12712=>"111110100",
  12713=>"111111101",
  12714=>"111000100",
  12715=>"000000000",
  12716=>"100000111",
  12717=>"110010111",
  12718=>"010000000",
  12719=>"000000000",
  12720=>"111111101",
  12721=>"000000011",
  12722=>"000000000",
  12723=>"111111011",
  12724=>"001001011",
  12725=>"000000001",
  12726=>"000111111",
  12727=>"000000101",
  12728=>"000000000",
  12729=>"010000000",
  12730=>"001000011",
  12731=>"001001101",
  12732=>"000000111",
  12733=>"111001000",
  12734=>"001000000",
  12735=>"000000011",
  12736=>"111110000",
  12737=>"001001000",
  12738=>"010010111",
  12739=>"111000000",
  12740=>"111111111",
  12741=>"000000000",
  12742=>"000000001",
  12743=>"111111111",
  12744=>"000000100",
  12745=>"101000000",
  12746=>"000000100",
  12747=>"000001111",
  12748=>"000111111",
  12749=>"000000001",
  12750=>"000000101",
  12751=>"000000010",
  12752=>"000000000",
  12753=>"111001000",
  12754=>"000000000",
  12755=>"101000000",
  12756=>"001000101",
  12757=>"000010000",
  12758=>"100000110",
  12759=>"011111111",
  12760=>"000000000",
  12761=>"000000000",
  12762=>"111111100",
  12763=>"111111111",
  12764=>"000011111",
  12765=>"111000100",
  12766=>"111111000",
  12767=>"101111111",
  12768=>"100001000",
  12769=>"000000001",
  12770=>"110011111",
  12771=>"000000111",
  12772=>"011111111",
  12773=>"110111000",
  12774=>"000100111",
  12775=>"000000111",
  12776=>"000000101",
  12777=>"111111010",
  12778=>"110100000",
  12779=>"111111010",
  12780=>"111111011",
  12781=>"000000100",
  12782=>"000000000",
  12783=>"100111111",
  12784=>"000000000",
  12785=>"111111111",
  12786=>"111111111",
  12787=>"000000110",
  12788=>"001001111",
  12789=>"110110011",
  12790=>"000001000",
  12791=>"000000000",
  12792=>"011111000",
  12793=>"001001000",
  12794=>"000000000",
  12795=>"111001000",
  12796=>"111000000",
  12797=>"111111111",
  12798=>"110000000",
  12799=>"011011001",
  12800=>"100000111",
  12801=>"011110000",
  12802=>"111101111",
  12803=>"111110000",
  12804=>"001000001",
  12805=>"100101001",
  12806=>"101101111",
  12807=>"001000000",
  12808=>"000000000",
  12809=>"111001000",
  12810=>"000000000",
  12811=>"000000000",
  12812=>"001111111",
  12813=>"000000000",
  12814=>"111111111",
  12815=>"000110110",
  12816=>"000000000",
  12817=>"000111111",
  12818=>"100101111",
  12819=>"000000101",
  12820=>"100000001",
  12821=>"000000000",
  12822=>"001011000",
  12823=>"000000000",
  12824=>"110110110",
  12825=>"111111000",
  12826=>"111111110",
  12827=>"111111111",
  12828=>"000000000",
  12829=>"111111101",
  12830=>"011001000",
  12831=>"111011001",
  12832=>"111111110",
  12833=>"010010010",
  12834=>"001010011",
  12835=>"000010000",
  12836=>"110000000",
  12837=>"100101101",
  12838=>"111111111",
  12839=>"000000001",
  12840=>"111111111",
  12841=>"111111111",
  12842=>"010010000",
  12843=>"000000010",
  12844=>"001000111",
  12845=>"000000010",
  12846=>"111111100",
  12847=>"111111111",
  12848=>"110111110",
  12849=>"000110110",
  12850=>"000000000",
  12851=>"010111111",
  12852=>"111111101",
  12853=>"111111010",
  12854=>"000100110",
  12855=>"111111010",
  12856=>"000000001",
  12857=>"000000000",
  12858=>"000111011",
  12859=>"111111111",
  12860=>"111111101",
  12861=>"111111111",
  12862=>"111111111",
  12863=>"000000000",
  12864=>"000000001",
  12865=>"011111111",
  12866=>"000000000",
  12867=>"000111111",
  12868=>"100110110",
  12869=>"111111111",
  12870=>"000000011",
  12871=>"111110111",
  12872=>"100110111",
  12873=>"111111111",
  12874=>"111111111",
  12875=>"110111111",
  12876=>"110010110",
  12877=>"001011111",
  12878=>"000000000",
  12879=>"000000000",
  12880=>"011011011",
  12881=>"000000000",
  12882=>"111111111",
  12883=>"100110111",
  12884=>"101111111",
  12885=>"111000000",
  12886=>"000000000",
  12887=>"111111111",
  12888=>"101111111",
  12889=>"001000111",
  12890=>"000111111",
  12891=>"110110000",
  12892=>"101000000",
  12893=>"000000000",
  12894=>"111110010",
  12895=>"001011000",
  12896=>"111111111",
  12897=>"000000000",
  12898=>"111111111",
  12899=>"100111111",
  12900=>"000011111",
  12901=>"000000000",
  12902=>"111111000",
  12903=>"110000000",
  12904=>"001001111",
  12905=>"111111111",
  12906=>"000000000",
  12907=>"110111111",
  12908=>"101100100",
  12909=>"000101001",
  12910=>"000000100",
  12911=>"111111111",
  12912=>"010111111",
  12913=>"111111110",
  12914=>"000000000",
  12915=>"110111000",
  12916=>"111111111",
  12917=>"101000000",
  12918=>"011000100",
  12919=>"011111111",
  12920=>"000100101",
  12921=>"101000000",
  12922=>"110100100",
  12923=>"000010000",
  12924=>"110110110",
  12925=>"000000011",
  12926=>"101100000",
  12927=>"000000000",
  12928=>"000000000",
  12929=>"000000000",
  12930=>"000000000",
  12931=>"000000000",
  12932=>"000000000",
  12933=>"111001111",
  12934=>"111111110",
  12935=>"000000000",
  12936=>"000101111",
  12937=>"000000110",
  12938=>"000100111",
  12939=>"000101111",
  12940=>"000000000",
  12941=>"001001111",
  12942=>"011000000",
  12943=>"000000000",
  12944=>"100100100",
  12945=>"000000000",
  12946=>"000000001",
  12947=>"000000000",
  12948=>"101111111",
  12949=>"000000000",
  12950=>"000000000",
  12951=>"110000000",
  12952=>"000000100",
  12953=>"111111111",
  12954=>"111111111",
  12955=>"001000000",
  12956=>"000000000",
  12957=>"000011011",
  12958=>"100000100",
  12959=>"000000000",
  12960=>"000000100",
  12961=>"000000000",
  12962=>"110111111",
  12963=>"111111111",
  12964=>"011001001",
  12965=>"111111111",
  12966=>"101101111",
  12967=>"011011011",
  12968=>"111111111",
  12969=>"111000000",
  12970=>"111000000",
  12971=>"111111000",
  12972=>"000000000",
  12973=>"110110100",
  12974=>"001000101",
  12975=>"111111001",
  12976=>"111111110",
  12977=>"111111111",
  12978=>"111111111",
  12979=>"000000000",
  12980=>"111110110",
  12981=>"111111011",
  12982=>"100101001",
  12983=>"100000001",
  12984=>"111111111",
  12985=>"000000000",
  12986=>"000000000",
  12987=>"001011000",
  12988=>"111111111",
  12989=>"110011011",
  12990=>"000000000",
  12991=>"000000000",
  12992=>"010111010",
  12993=>"101001111",
  12994=>"000000000",
  12995=>"100000000",
  12996=>"111010011",
  12997=>"001000000",
  12998=>"111110100",
  12999=>"100000000",
  13000=>"000000000",
  13001=>"000000000",
  13002=>"100000001",
  13003=>"100000000",
  13004=>"000000000",
  13005=>"000000000",
  13006=>"011010000",
  13007=>"000000000",
  13008=>"001101111",
  13009=>"000110011",
  13010=>"000000000",
  13011=>"000001000",
  13012=>"001001011",
  13013=>"000000100",
  13014=>"000000000",
  13015=>"000000001",
  13016=>"111111111",
  13017=>"100111111",
  13018=>"000000000",
  13019=>"111111111",
  13020=>"000000000",
  13021=>"110011011",
  13022=>"110010011",
  13023=>"000000000",
  13024=>"111111111",
  13025=>"000000000",
  13026=>"111111111",
  13027=>"111111111",
  13028=>"111111010",
  13029=>"000011001",
  13030=>"011000000",
  13031=>"000000110",
  13032=>"111111000",
  13033=>"111111000",
  13034=>"101111111",
  13035=>"000000110",
  13036=>"000111111",
  13037=>"111111111",
  13038=>"111000110",
  13039=>"000100110",
  13040=>"011011010",
  13041=>"000000000",
  13042=>"111111111",
  13043=>"001001001",
  13044=>"010000000",
  13045=>"110110010",
  13046=>"011111011",
  13047=>"111111111",
  13048=>"000000000",
  13049=>"111101100",
  13050=>"000000000",
  13051=>"111111011",
  13052=>"111111000",
  13053=>"000000000",
  13054=>"100000000",
  13055=>"111111111",
  13056=>"110100001",
  13057=>"000000000",
  13058=>"011000000",
  13059=>"000000000",
  13060=>"111100101",
  13061=>"000000000",
  13062=>"111000101",
  13063=>"000000001",
  13064=>"100110111",
  13065=>"000000000",
  13066=>"111111111",
  13067=>"000000111",
  13068=>"111111011",
  13069=>"000000000",
  13070=>"000001000",
  13071=>"000000000",
  13072=>"001111111",
  13073=>"001001000",
  13074=>"000000000",
  13075=>"110111111",
  13076=>"000001111",
  13077=>"000000000",
  13078=>"110100010",
  13079=>"111001000",
  13080=>"100100100",
  13081=>"111111111",
  13082=>"111111111",
  13083=>"000000000",
  13084=>"110110100",
  13085=>"000000001",
  13086=>"000000000",
  13087=>"111111111",
  13088=>"010110100",
  13089=>"111000001",
  13090=>"100011000",
  13091=>"101100110",
  13092=>"011000000",
  13093=>"110111111",
  13094=>"011011011",
  13095=>"000000001",
  13096=>"111111010",
  13097=>"001000000",
  13098=>"101100110",
  13099=>"000000000",
  13100=>"111111011",
  13101=>"000000001",
  13102=>"111011011",
  13103=>"110000110",
  13104=>"111111110",
  13105=>"000000000",
  13106=>"111000001",
  13107=>"111111110",
  13108=>"000001000",
  13109=>"000100100",
  13110=>"000000111",
  13111=>"111111011",
  13112=>"000000000",
  13113=>"101111111",
  13114=>"000000000",
  13115=>"000111111",
  13116=>"000000111",
  13117=>"110011111",
  13118=>"011011011",
  13119=>"111011011",
  13120=>"110111111",
  13121=>"111111000",
  13122=>"000000011",
  13123=>"000000000",
  13124=>"000101001",
  13125=>"000100111",
  13126=>"111111110",
  13127=>"000000100",
  13128=>"111111111",
  13129=>"010000000",
  13130=>"000000000",
  13131=>"110111000",
  13132=>"000000000",
  13133=>"101110110",
  13134=>"000000101",
  13135=>"000000000",
  13136=>"100000010",
  13137=>"111101111",
  13138=>"000000111",
  13139=>"111111111",
  13140=>"101100000",
  13141=>"011011011",
  13142=>"001111111",
  13143=>"000000000",
  13144=>"101110111",
  13145=>"001110111",
  13146=>"111111111",
  13147=>"000000001",
  13148=>"000110011",
  13149=>"111111000",
  13150=>"111111111",
  13151=>"000000000",
  13152=>"100100100",
  13153=>"111111011",
  13154=>"001111000",
  13155=>"000101100",
  13156=>"000001011",
  13157=>"101001011",
  13158=>"000000000",
  13159=>"100000000",
  13160=>"111111001",
  13161=>"100100111",
  13162=>"000111000",
  13163=>"111001000",
  13164=>"110111111",
  13165=>"000000110",
  13166=>"000000111",
  13167=>"000010000",
  13168=>"000000000",
  13169=>"111111111",
  13170=>"000111111",
  13171=>"100000000",
  13172=>"110010000",
  13173=>"111100100",
  13174=>"000000000",
  13175=>"111110000",
  13176=>"110111111",
  13177=>"000000001",
  13178=>"000000111",
  13179=>"000000000",
  13180=>"111111111",
  13181=>"111111111",
  13182=>"100101111",
  13183=>"000000000",
  13184=>"101110111",
  13185=>"000000000",
  13186=>"111111110",
  13187=>"111111111",
  13188=>"000000000",
  13189=>"010100100",
  13190=>"000000000",
  13191=>"000000000",
  13192=>"000000000",
  13193=>"111111111",
  13194=>"011111111",
  13195=>"110011111",
  13196=>"111111111",
  13197=>"000111000",
  13198=>"010000000",
  13199=>"000010010",
  13200=>"011000000",
  13201=>"101111111",
  13202=>"000000000",
  13203=>"000000011",
  13204=>"100111111",
  13205=>"000000000",
  13206=>"000100111",
  13207=>"000001101",
  13208=>"111111000",
  13209=>"010111111",
  13210=>"011111111",
  13211=>"000000000",
  13212=>"111010000",
  13213=>"000000000",
  13214=>"011011011",
  13215=>"010111111",
  13216=>"000000000",
  13217=>"111111111",
  13218=>"111100100",
  13219=>"010111000",
  13220=>"111111111",
  13221=>"000000000",
  13222=>"111111111",
  13223=>"010111111",
  13224=>"000000100",
  13225=>"000000100",
  13226=>"111111111",
  13227=>"000000000",
  13228=>"000000000",
  13229=>"011010000",
  13230=>"010110000",
  13231=>"000011111",
  13232=>"010011000",
  13233=>"000000111",
  13234=>"001011111",
  13235=>"000000000",
  13236=>"001001000",
  13237=>"111001000",
  13238=>"111101000",
  13239=>"100100000",
  13240=>"011111111",
  13241=>"000000000",
  13242=>"111111111",
  13243=>"000000101",
  13244=>"001100100",
  13245=>"000000001",
  13246=>"100101111",
  13247=>"001111111",
  13248=>"111111011",
  13249=>"111111111",
  13250=>"000100111",
  13251=>"111101111",
  13252=>"100001111",
  13253=>"000101111",
  13254=>"100110000",
  13255=>"111111111",
  13256=>"001101111",
  13257=>"000000000",
  13258=>"111111111",
  13259=>"111111000",
  13260=>"111111011",
  13261=>"101111111",
  13262=>"100100001",
  13263=>"111111010",
  13264=>"111011000",
  13265=>"000000000",
  13266=>"110000000",
  13267=>"000000000",
  13268=>"011000000",
  13269=>"000110111",
  13270=>"000000000",
  13271=>"111111110",
  13272=>"111111010",
  13273=>"100100000",
  13274=>"001000000",
  13275=>"111000000",
  13276=>"000000000",
  13277=>"111101101",
  13278=>"111111100",
  13279=>"000011110",
  13280=>"111110110",
  13281=>"000101111",
  13282=>"000000000",
  13283=>"111111001",
  13284=>"000000000",
  13285=>"110110110",
  13286=>"000000001",
  13287=>"000001011",
  13288=>"111111111",
  13289=>"111111101",
  13290=>"111101001",
  13291=>"111111111",
  13292=>"111111000",
  13293=>"000000000",
  13294=>"001110111",
  13295=>"100000111",
  13296=>"000101111",
  13297=>"000110110",
  13298=>"000110110",
  13299=>"000100000",
  13300=>"101111111",
  13301=>"000000110",
  13302=>"010010010",
  13303=>"011011000",
  13304=>"000111111",
  13305=>"100000001",
  13306=>"110100100",
  13307=>"000000101",
  13308=>"000000000",
  13309=>"110111111",
  13310=>"000000000",
  13311=>"111111000",
  13312=>"000100111",
  13313=>"000000000",
  13314=>"111111110",
  13315=>"000001011",
  13316=>"011111111",
  13317=>"101111111",
  13318=>"000000001",
  13319=>"011111111",
  13320=>"100000000",
  13321=>"000001011",
  13322=>"001111111",
  13323=>"000111101",
  13324=>"000110000",
  13325=>"111000100",
  13326=>"000000000",
  13327=>"100000100",
  13328=>"111011000",
  13329=>"000011011",
  13330=>"000011000",
  13331=>"000000111",
  13332=>"111111111",
  13333=>"100000000",
  13334=>"100000000",
  13335=>"111000000",
  13336=>"100110110",
  13337=>"000110000",
  13338=>"110000001",
  13339=>"011101111",
  13340=>"111111100",
  13341=>"011111000",
  13342=>"001111111",
  13343=>"111111111",
  13344=>"000000000",
  13345=>"010111111",
  13346=>"111000000",
  13347=>"001000001",
  13348=>"010000111",
  13349=>"000000000",
  13350=>"000001111",
  13351=>"100000000",
  13352=>"000000111",
  13353=>"100000111",
  13354=>"000000100",
  13355=>"000000000",
  13356=>"111111000",
  13357=>"000000000",
  13358=>"111111111",
  13359=>"111111110",
  13360=>"001111111",
  13361=>"111111000",
  13362=>"000000111",
  13363=>"111011111",
  13364=>"110000000",
  13365=>"000111111",
  13366=>"111000000",
  13367=>"111001110",
  13368=>"000000000",
  13369=>"100000111",
  13370=>"000000000",
  13371=>"111000000",
  13372=>"111111111",
  13373=>"000000100",
  13374=>"000101111",
  13375=>"000101111",
  13376=>"000000100",
  13377=>"011011111",
  13378=>"111111111",
  13379=>"111111000",
  13380=>"000000110",
  13381=>"100100100",
  13382=>"111000000",
  13383=>"011111111",
  13384=>"001011011",
  13385=>"000111111",
  13386=>"000000110",
  13387=>"111101000",
  13388=>"001011111",
  13389=>"111111000",
  13390=>"000010110",
  13391=>"000000011",
  13392=>"000000001",
  13393=>"000000000",
  13394=>"000010111",
  13395=>"111100100",
  13396=>"111111000",
  13397=>"000000110",
  13398=>"000000111",
  13399=>"000000000",
  13400=>"111110111",
  13401=>"111000000",
  13402=>"000000000",
  13403=>"110010000",
  13404=>"100000000",
  13405=>"000100100",
  13406=>"111100111",
  13407=>"000110010",
  13408=>"111101111",
  13409=>"100000000",
  13410=>"111011111",
  13411=>"111111111",
  13412=>"001000000",
  13413=>"000001111",
  13414=>"111000111",
  13415=>"000000000",
  13416=>"010000101",
  13417=>"000111010",
  13418=>"111111111",
  13419=>"000000000",
  13420=>"111111111",
  13421=>"000000000",
  13422=>"111111001",
  13423=>"000000111",
  13424=>"000001111",
  13425=>"111101111",
  13426=>"001000001",
  13427=>"111101100",
  13428=>"000000000",
  13429=>"100110000",
  13430=>"000110110",
  13431=>"000001000",
  13432=>"000000000",
  13433=>"011001001",
  13434=>"011001000",
  13435=>"000000111",
  13436=>"111011000",
  13437=>"110011000",
  13438=>"001000000",
  13439=>"000000000",
  13440=>"111111111",
  13441=>"000000001",
  13442=>"111000000",
  13443=>"011111110",
  13444=>"001000001",
  13445=>"111000000",
  13446=>"100101111",
  13447=>"111110000",
  13448=>"111000000",
  13449=>"111000110",
  13450=>"001000000",
  13451=>"000111000",
  13452=>"001000111",
  13453=>"000000111",
  13454=>"111110111",
  13455=>"000000000",
  13456=>"011111111",
  13457=>"111111111",
  13458=>"000000001",
  13459=>"111100000",
  13460=>"001000000",
  13461=>"000000000",
  13462=>"110000000",
  13463=>"000000000",
  13464=>"100111111",
  13465=>"000001111",
  13466=>"001000000",
  13467=>"011011110",
  13468=>"111001001",
  13469=>"011011111",
  13470=>"111111111",
  13471=>"111111001",
  13472=>"111111100",
  13473=>"101111001",
  13474=>"000010110",
  13475=>"111111101",
  13476=>"000000000",
  13477=>"111111111",
  13478=>"111111100",
  13479=>"111111111",
  13480=>"000000100",
  13481=>"111111110",
  13482=>"000111111",
  13483=>"111111111",
  13484=>"110111111",
  13485=>"100100000",
  13486=>"000000001",
  13487=>"111111000",
  13488=>"000000000",
  13489=>"001111111",
  13490=>"000000110",
  13491=>"011000000",
  13492=>"000111111",
  13493=>"100000000",
  13494=>"000000111",
  13495=>"000000001",
  13496=>"011000110",
  13497=>"111111000",
  13498=>"000000100",
  13499=>"111111100",
  13500=>"000110000",
  13501=>"000000101",
  13502=>"000011000",
  13503=>"000011111",
  13504=>"111000000",
  13505=>"000000110",
  13506=>"111111111",
  13507=>"111111111",
  13508=>"000000000",
  13509=>"111111111",
  13510=>"111111111",
  13511=>"000000111",
  13512=>"000000000",
  13513=>"111111111",
  13514=>"000000000",
  13515=>"000000011",
  13516=>"000100101",
  13517=>"100100000",
  13518=>"111100000",
  13519=>"000000100",
  13520=>"000011000",
  13521=>"111011111",
  13522=>"000000110",
  13523=>"100000000",
  13524=>"111111111",
  13525=>"101111011",
  13526=>"000000011",
  13527=>"111110110",
  13528=>"011111111",
  13529=>"000000000",
  13530=>"000000010",
  13531=>"001111111",
  13532=>"111000000",
  13533=>"101101000",
  13534=>"000010001",
  13535=>"111110111",
  13536=>"000000111",
  13537=>"011001000",
  13538=>"000010000",
  13539=>"111111000",
  13540=>"000111111",
  13541=>"111111000",
  13542=>"000000111",
  13543=>"101001111",
  13544=>"000000000",
  13545=>"011111001",
  13546=>"000000111",
  13547=>"000000000",
  13548=>"111000000",
  13549=>"000000110",
  13550=>"111111111",
  13551=>"001001000",
  13552=>"111111000",
  13553=>"010110110",
  13554=>"011111111",
  13555=>"000000111",
  13556=>"111111000",
  13557=>"011011000",
  13558=>"001000100",
  13559=>"011111111",
  13560=>"011001000",
  13561=>"110000000",
  13562=>"000001000",
  13563=>"111111010",
  13564=>"000000000",
  13565=>"100000100",
  13566=>"100111111",
  13567=>"000000001",
  13568=>"110110000",
  13569=>"000000100",
  13570=>"111111000",
  13571=>"000000100",
  13572=>"000011011",
  13573=>"000000111",
  13574=>"001111000",
  13575=>"111110100",
  13576=>"111111111",
  13577=>"000000000",
  13578=>"111111110",
  13579=>"101000000",
  13580=>"111101000",
  13581=>"111001111",
  13582=>"000000000",
  13583=>"111010000",
  13584=>"111111000",
  13585=>"001000000",
  13586=>"100100110",
  13587=>"000010000",
  13588=>"000111111",
  13589=>"000001111",
  13590=>"011111110",
  13591=>"000000000",
  13592=>"111110000",
  13593=>"000111111",
  13594=>"111111111",
  13595=>"110000001",
  13596=>"000111100",
  13597=>"000000111",
  13598=>"111001111",
  13599=>"000000000",
  13600=>"001000000",
  13601=>"010011111",
  13602=>"000000111",
  13603=>"000000110",
  13604=>"111111111",
  13605=>"011111111",
  13606=>"111111111",
  13607=>"111000110",
  13608=>"111111111",
  13609=>"000000111",
  13610=>"111001000",
  13611=>"000000001",
  13612=>"000000000",
  13613=>"110100000",
  13614=>"000110111",
  13615=>"111000000",
  13616=>"110001111",
  13617=>"000111111",
  13618=>"111111110",
  13619=>"111111111",
  13620=>"010000111",
  13621=>"111000000",
  13622=>"000000000",
  13623=>"001100111",
  13624=>"101000000",
  13625=>"111000101",
  13626=>"111111000",
  13627=>"111110000",
  13628=>"101100100",
  13629=>"000000000",
  13630=>"100111111",
  13631=>"111111110",
  13632=>"011111111",
  13633=>"011111100",
  13634=>"100000111",
  13635=>"101000001",
  13636=>"000100111",
  13637=>"100000000",
  13638=>"000000000",
  13639=>"000000001",
  13640=>"110110100",
  13641=>"000000000",
  13642=>"011111111",
  13643=>"010010010",
  13644=>"010000000",
  13645=>"111000000",
  13646=>"000000001",
  13647=>"000000100",
  13648=>"111111000",
  13649=>"000000101",
  13650=>"111111111",
  13651=>"000000011",
  13652=>"000000001",
  13653=>"001000000",
  13654=>"111000000",
  13655=>"101000000",
  13656=>"111111111",
  13657=>"000000000",
  13658=>"101101001",
  13659=>"011111110",
  13660=>"100000111",
  13661=>"111111111",
  13662=>"111100110",
  13663=>"000111111",
  13664=>"000000000",
  13665=>"000000111",
  13666=>"011111111",
  13667=>"111111000",
  13668=>"000000111",
  13669=>"110000110",
  13670=>"000000111",
  13671=>"111000110",
  13672=>"101101101",
  13673=>"111010000",
  13674=>"100010111",
  13675=>"000011111",
  13676=>"000000000",
  13677=>"000001111",
  13678=>"000000011",
  13679=>"111111110",
  13680=>"111111110",
  13681=>"111111000",
  13682=>"111111000",
  13683=>"010100000",
  13684=>"111111000",
  13685=>"111111111",
  13686=>"001111011",
  13687=>"000111111",
  13688=>"111111000",
  13689=>"000000000",
  13690=>"111000000",
  13691=>"100000000",
  13692=>"111111111",
  13693=>"100000110",
  13694=>"100111001",
  13695=>"111001000",
  13696=>"001000001",
  13697=>"000100000",
  13698=>"000000001",
  13699=>"111100000",
  13700=>"111111000",
  13701=>"000111011",
  13702=>"110000000",
  13703=>"000000000",
  13704=>"100100110",
  13705=>"111001001",
  13706=>"111101111",
  13707=>"000100111",
  13708=>"011000000",
  13709=>"011111100",
  13710=>"111100111",
  13711=>"010111111",
  13712=>"000111111",
  13713=>"000100100",
  13714=>"111111000",
  13715=>"110011011",
  13716=>"111111111",
  13717=>"000011010",
  13718=>"011001100",
  13719=>"000100100",
  13720=>"011111100",
  13721=>"100011000",
  13722=>"000100101",
  13723=>"111000001",
  13724=>"000000000",
  13725=>"111110000",
  13726=>"000000111",
  13727=>"000100010",
  13728=>"000111111",
  13729=>"100101101",
  13730=>"001111101",
  13731=>"000000111",
  13732=>"111000100",
  13733=>"111111111",
  13734=>"100100111",
  13735=>"000010111",
  13736=>"111111000",
  13737=>"011010000",
  13738=>"001110110",
  13739=>"000000100",
  13740=>"000000000",
  13741=>"100000101",
  13742=>"000000101",
  13743=>"000000111",
  13744=>"000000000",
  13745=>"000000001",
  13746=>"000000000",
  13747=>"000011111",
  13748=>"000001111",
  13749=>"000000000",
  13750=>"001111111",
  13751=>"000111111",
  13752=>"110000110",
  13753=>"001011111",
  13754=>"000101111",
  13755=>"111110110",
  13756=>"001000001",
  13757=>"111111111",
  13758=>"111010000",
  13759=>"111111110",
  13760=>"111010010",
  13761=>"000000001",
  13762=>"111111111",
  13763=>"111111000",
  13764=>"111111110",
  13765=>"101000000",
  13766=>"011011101",
  13767=>"001100110",
  13768=>"000001001",
  13769=>"111111111",
  13770=>"000100100",
  13771=>"000011001",
  13772=>"000100111",
  13773=>"111101000",
  13774=>"111111110",
  13775=>"100111111",
  13776=>"111010111",
  13777=>"111111111",
  13778=>"011000111",
  13779=>"111111111",
  13780=>"001111111",
  13781=>"000000101",
  13782=>"000000111",
  13783=>"001001001",
  13784=>"000000111",
  13785=>"000111111",
  13786=>"010111111",
  13787=>"101001001",
  13788=>"000000101",
  13789=>"000000000",
  13790=>"000000111",
  13791=>"111111001",
  13792=>"001001111",
  13793=>"100001111",
  13794=>"000100000",
  13795=>"101000000",
  13796=>"111111111",
  13797=>"011001000",
  13798=>"111011111",
  13799=>"000000111",
  13800=>"000000000",
  13801=>"111111111",
  13802=>"110100111",
  13803=>"000000111",
  13804=>"000000001",
  13805=>"001001000",
  13806=>"001001001",
  13807=>"011111111",
  13808=>"000000000",
  13809=>"000111110",
  13810=>"001111111",
  13811=>"000000010",
  13812=>"001001011",
  13813=>"000101111",
  13814=>"111111111",
  13815=>"011111111",
  13816=>"000000001",
  13817=>"111111100",
  13818=>"000000111",
  13819=>"011111111",
  13820=>"011111111",
  13821=>"111111111",
  13822=>"000001111",
  13823=>"000000000",
  13824=>"011000000",
  13825=>"000000000",
  13826=>"101000111",
  13827=>"000000000",
  13828=>"000000110",
  13829=>"001000000",
  13830=>"000000000",
  13831=>"000111111",
  13832=>"111111111",
  13833=>"000000000",
  13834=>"001000001",
  13835=>"111111110",
  13836=>"100000000",
  13837=>"111111111",
  13838=>"011011001",
  13839=>"111101101",
  13840=>"111111111",
  13841=>"010111111",
  13842=>"000000011",
  13843=>"000000000",
  13844=>"000000000",
  13845=>"111010010",
  13846=>"111111011",
  13847=>"011111110",
  13848=>"101101000",
  13849=>"000000000",
  13850=>"101001111",
  13851=>"000000000",
  13852=>"101111111",
  13853=>"111111111",
  13854=>"000111001",
  13855=>"111111111",
  13856=>"111111111",
  13857=>"000000000",
  13858=>"101101111",
  13859=>"100000111",
  13860=>"111011111",
  13861=>"001011011",
  13862=>"000000000",
  13863=>"000000110",
  13864=>"111000000",
  13865=>"000000111",
  13866=>"000000111",
  13867=>"100011011",
  13868=>"100000111",
  13869=>"000000000",
  13870=>"000001111",
  13871=>"111000000",
  13872=>"001000000",
  13873=>"000000000",
  13874=>"111111100",
  13875=>"110000101",
  13876=>"111111111",
  13877=>"110100110",
  13878=>"111111111",
  13879=>"100110110",
  13880=>"000000000",
  13881=>"111111000",
  13882=>"000000001",
  13883=>"100111111",
  13884=>"111111110",
  13885=>"000111111",
  13886=>"111111001",
  13887=>"101101111",
  13888=>"111111000",
  13889=>"111111111",
  13890=>"000000000",
  13891=>"000000000",
  13892=>"110110111",
  13893=>"000000000",
  13894=>"001011000",
  13895=>"111111011",
  13896=>"011011111",
  13897=>"111111111",
  13898=>"001010111",
  13899=>"011010000",
  13900=>"000000110",
  13901=>"000000110",
  13902=>"110111100",
  13903=>"111111111",
  13904=>"011011101",
  13905=>"000111111",
  13906=>"001001010",
  13907=>"000000000",
  13908=>"111110000",
  13909=>"000100000",
  13910=>"111000000",
  13911=>"011111111",
  13912=>"100100000",
  13913=>"111101101",
  13914=>"000000001",
  13915=>"111100100",
  13916=>"000000000",
  13917=>"111111111",
  13918=>"111111111",
  13919=>"111111111",
  13920=>"000111111",
  13921=>"111110111",
  13922=>"011010011",
  13923=>"000000000",
  13924=>"000000101",
  13925=>"111111000",
  13926=>"100000000",
  13927=>"000000001",
  13928=>"000000000",
  13929=>"000111110",
  13930=>"111111111",
  13931=>"111101000",
  13932=>"000000000",
  13933=>"011001001",
  13934=>"111111111",
  13935=>"110111111",
  13936=>"111111111",
  13937=>"100100111",
  13938=>"110111111",
  13939=>"000000111",
  13940=>"111101101",
  13941=>"000000110",
  13942=>"001000000",
  13943=>"000000000",
  13944=>"000000000",
  13945=>"111111111",
  13946=>"000000000",
  13947=>"011011111",
  13948=>"110110000",
  13949=>"111110000",
  13950=>"000000000",
  13951=>"000011111",
  13952=>"100111111",
  13953=>"000110111",
  13954=>"111101111",
  13955=>"001000000",
  13956=>"101000000",
  13957=>"101001101",
  13958=>"100000100",
  13959=>"111111110",
  13960=>"101000000",
  13961=>"111000000",
  13962=>"000110000",
  13963=>"110111111",
  13964=>"000000000",
  13965=>"000000110",
  13966=>"000110110",
  13967=>"110110110",
  13968=>"000000000",
  13969=>"000000001",
  13970=>"000000000",
  13971=>"011111000",
  13972=>"101001111",
  13973=>"111110110",
  13974=>"111111111",
  13975=>"001000101",
  13976=>"011111111",
  13977=>"000000111",
  13978=>"111111111",
  13979=>"001000000",
  13980=>"111111111",
  13981=>"000000000",
  13982=>"111010011",
  13983=>"111110111",
  13984=>"111101001",
  13985=>"000000000",
  13986=>"000000000",
  13987=>"111011000",
  13988=>"100110110",
  13989=>"000000000",
  13990=>"110111111",
  13991=>"011000010",
  13992=>"110111111",
  13993=>"100000000",
  13994=>"000000000",
  13995=>"111001000",
  13996=>"000000001",
  13997=>"001011111",
  13998=>"010110111",
  13999=>"111000000",
  14000=>"000000100",
  14001=>"001010010",
  14002=>"110110111",
  14003=>"111111111",
  14004=>"111000000",
  14005=>"000100000",
  14006=>"000100111",
  14007=>"001011111",
  14008=>"000100111",
  14009=>"011011011",
  14010=>"000110000",
  14011=>"000110110",
  14012=>"111101111",
  14013=>"000111111",
  14014=>"000000000",
  14015=>"111110010",
  14016=>"110111111",
  14017=>"111111111",
  14018=>"000000000",
  14019=>"001101000",
  14020=>"110011111",
  14021=>"111111111",
  14022=>"111111111",
  14023=>"000000000",
  14024=>"000010010",
  14025=>"111111111",
  14026=>"111111100",
  14027=>"011111111",
  14028=>"111001100",
  14029=>"000000000",
  14030=>"000000000",
  14031=>"011011111",
  14032=>"111111110",
  14033=>"000111111",
  14034=>"000000010",
  14035=>"101000111",
  14036=>"000000000",
  14037=>"001000011",
  14038=>"111011001",
  14039=>"111001011",
  14040=>"100000100",
  14041=>"000000010",
  14042=>"111111111",
  14043=>"111111111",
  14044=>"111111110",
  14045=>"100111111",
  14046=>"100101111",
  14047=>"111111111",
  14048=>"000100110",
  14049=>"100000000",
  14050=>"011001001",
  14051=>"111000111",
  14052=>"111111111",
  14053=>"001000101",
  14054=>"000100110",
  14055=>"100110111",
  14056=>"000000111",
  14057=>"000111111",
  14058=>"100000111",
  14059=>"111101111",
  14060=>"001011010",
  14061=>"000000000",
  14062=>"111111101",
  14063=>"111000000",
  14064=>"000000011",
  14065=>"010111111",
  14066=>"111111111",
  14067=>"111101100",
  14068=>"111110010",
  14069=>"111111111",
  14070=>"000110110",
  14071=>"111111111",
  14072=>"000000001",
  14073=>"111000000",
  14074=>"100000100",
  14075=>"000110111",
  14076=>"100100111",
  14077=>"000000001",
  14078=>"000010011",
  14079=>"000110110",
  14080=>"110110111",
  14081=>"111100110",
  14082=>"111110000",
  14083=>"111101000",
  14084=>"111111111",
  14085=>"100100111",
  14086=>"011111111",
  14087=>"000000001",
  14088=>"101011111",
  14089=>"111001000",
  14090=>"100001111",
  14091=>"110001101",
  14092=>"001000000",
  14093=>"000000000",
  14094=>"100100000",
  14095=>"010111111",
  14096=>"111001000",
  14097=>"111111111",
  14098=>"000000111",
  14099=>"111011000",
  14100=>"111110000",
  14101=>"111111111",
  14102=>"001001001",
  14103=>"110111110",
  14104=>"100110000",
  14105=>"000000000",
  14106=>"001000001",
  14107=>"111111111",
  14108=>"111111111",
  14109=>"011011111",
  14110=>"000100100",
  14111=>"111111111",
  14112=>"000100110",
  14113=>"000000000",
  14114=>"011110110",
  14115=>"000000000",
  14116=>"000000111",
  14117=>"001000000",
  14118=>"011011001",
  14119=>"010011001",
  14120=>"111000110",
  14121=>"011001011",
  14122=>"100111111",
  14123=>"000000000",
  14124=>"000010111",
  14125=>"111000001",
  14126=>"000000000",
  14127=>"000000000",
  14128=>"100110111",
  14129=>"111111011",
  14130=>"111111000",
  14131=>"111111001",
  14132=>"010000000",
  14133=>"011111011",
  14134=>"011111100",
  14135=>"111111111",
  14136=>"111011000",
  14137=>"111010000",
  14138=>"000011000",
  14139=>"000000111",
  14140=>"111111000",
  14141=>"100100000",
  14142=>"111111111",
  14143=>"000000000",
  14144=>"100111000",
  14145=>"110111111",
  14146=>"100110111",
  14147=>"000000001",
  14148=>"111111111",
  14149=>"101001100",
  14150=>"111001001",
  14151=>"111000100",
  14152=>"111000000",
  14153=>"000000000",
  14154=>"101001000",
  14155=>"111111111",
  14156=>"000000000",
  14157=>"000000001",
  14158=>"000000011",
  14159=>"000001001",
  14160=>"111111111",
  14161=>"000000000",
  14162=>"101011011",
  14163=>"111111111",
  14164=>"100101111",
  14165=>"001011011",
  14166=>"000000101",
  14167=>"001101101",
  14168=>"111111111",
  14169=>"111111111",
  14170=>"000000000",
  14171=>"111110111",
  14172=>"011111111",
  14173=>"011010010",
  14174=>"100100100",
  14175=>"111110110",
  14176=>"000000000",
  14177=>"111010110",
  14178=>"100110100",
  14179=>"101101111",
  14180=>"111110110",
  14181=>"101000111",
  14182=>"000000001",
  14183=>"111110101",
  14184=>"110110111",
  14185=>"110100000",
  14186=>"000000000",
  14187=>"111001001",
  14188=>"100000000",
  14189=>"000111011",
  14190=>"000000000",
  14191=>"000110111",
  14192=>"000100111",
  14193=>"000000000",
  14194=>"111111111",
  14195=>"000001011",
  14196=>"010000000",
  14197=>"001000110",
  14198=>"111111111",
  14199=>"000100111",
  14200=>"000001001",
  14201=>"000000111",
  14202=>"111111111",
  14203=>"000000000",
  14204=>"101000000",
  14205=>"000000011",
  14206=>"000000001",
  14207=>"111111111",
  14208=>"111111111",
  14209=>"000000000",
  14210=>"000000000",
  14211=>"111101111",
  14212=>"111111111",
  14213=>"111111111",
  14214=>"000000000",
  14215=>"000000000",
  14216=>"001000001",
  14217=>"011111111",
  14218=>"110111111",
  14219=>"101101111",
  14220=>"101000000",
  14221=>"111001000",
  14222=>"000000011",
  14223=>"000000011",
  14224=>"000000000",
  14225=>"110100111",
  14226=>"000100100",
  14227=>"111111010",
  14228=>"000001000",
  14229=>"000000000",
  14230=>"000000000",
  14231=>"111011000",
  14232=>"111111111",
  14233=>"000001111",
  14234=>"000000011",
  14235=>"011111111",
  14236=>"000000011",
  14237=>"111110110",
  14238=>"000000000",
  14239=>"000011000",
  14240=>"000000111",
  14241=>"000000000",
  14242=>"011000001",
  14243=>"000000000",
  14244=>"011000000",
  14245=>"111111111",
  14246=>"111011111",
  14247=>"000000000",
  14248=>"111001000",
  14249=>"000000001",
  14250=>"000000111",
  14251=>"000100110",
  14252=>"001000000",
  14253=>"000001000",
  14254=>"111111111",
  14255=>"000000000",
  14256=>"111111111",
  14257=>"111111111",
  14258=>"000000000",
  14259=>"000000000",
  14260=>"000000011",
  14261=>"000000000",
  14262=>"000000111",
  14263=>"000011111",
  14264=>"100101000",
  14265=>"111111110",
  14266=>"000001111",
  14267=>"111111111",
  14268=>"000000110",
  14269=>"111110110",
  14270=>"111100100",
  14271=>"101111111",
  14272=>"100100111",
  14273=>"111111111",
  14274=>"111111111",
  14275=>"101101111",
  14276=>"110101101",
  14277=>"000001111",
  14278=>"010010000",
  14279=>"000001000",
  14280=>"000000000",
  14281=>"000111111",
  14282=>"111011001",
  14283=>"111111000",
  14284=>"100000000",
  14285=>"000000111",
  14286=>"100100110",
  14287=>"111111111",
  14288=>"110000000",
  14289=>"111111111",
  14290=>"011111111",
  14291=>"111011111",
  14292=>"001010011",
  14293=>"001111111",
  14294=>"000001111",
  14295=>"001111111",
  14296=>"001101111",
  14297=>"011000000",
  14298=>"010010000",
  14299=>"110100111",
  14300=>"010110000",
  14301=>"000100110",
  14302=>"111111111",
  14303=>"101000000",
  14304=>"001000000",
  14305=>"111111111",
  14306=>"100101111",
  14307=>"001000101",
  14308=>"100110000",
  14309=>"111000111",
  14310=>"000100111",
  14311=>"000000111",
  14312=>"101000000",
  14313=>"011111011",
  14314=>"111111111",
  14315=>"000000000",
  14316=>"001110111",
  14317=>"000100100",
  14318=>"000000000",
  14319=>"000000000",
  14320=>"010000000",
  14321=>"111111111",
  14322=>"111111101",
  14323=>"000110111",
  14324=>"111111111",
  14325=>"000000000",
  14326=>"111111111",
  14327=>"111111000",
  14328=>"111111111",
  14329=>"110100100",
  14330=>"111111111",
  14331=>"011000000",
  14332=>"000000111",
  14333=>"101101111",
  14334=>"000000000",
  14335=>"000100100",
  14336=>"000000000",
  14337=>"000000000",
  14338=>"111000000",
  14339=>"000000000",
  14340=>"001100110",
  14341=>"111000110",
  14342=>"100000001",
  14343=>"001001001",
  14344=>"000000000",
  14345=>"000000011",
  14346=>"000000000",
  14347=>"001000000",
  14348=>"110001001",
  14349=>"000000000",
  14350=>"011001001",
  14351=>"000000000",
  14352=>"000100100",
  14353=>"111111111",
  14354=>"100001101",
  14355=>"000000000",
  14356=>"000000001",
  14357=>"111111000",
  14358=>"110101001",
  14359=>"001001001",
  14360=>"001001101",
  14361=>"111111111",
  14362=>"000100000",
  14363=>"111111111",
  14364=>"010001011",
  14365=>"100000000",
  14366=>"011001110",
  14367=>"111110110",
  14368=>"010010000",
  14369=>"111111111",
  14370=>"001001001",
  14371=>"111101100",
  14372=>"111111111",
  14373=>"000000011",
  14374=>"101111111",
  14375=>"111111001",
  14376=>"001000111",
  14377=>"000000000",
  14378=>"000000000",
  14379=>"111111111",
  14380=>"000000000",
  14381=>"110110010",
  14382=>"111100100",
  14383=>"111101100",
  14384=>"001000000",
  14385=>"111111111",
  14386=>"100000001",
  14387=>"000010011",
  14388=>"110010000",
  14389=>"110111101",
  14390=>"111111111",
  14391=>"110111111",
  14392=>"000010111",
  14393=>"111001001",
  14394=>"000000001",
  14395=>"111110110",
  14396=>"000000000",
  14397=>"110111111",
  14398=>"111000000",
  14399=>"111011011",
  14400=>"101111101",
  14401=>"011111110",
  14402=>"011111111",
  14403=>"000000000",
  14404=>"101111111",
  14405=>"011101111",
  14406=>"110111111",
  14407=>"111111111",
  14408=>"111100100",
  14409=>"000000000",
  14410=>"111111111",
  14411=>"000001011",
  14412=>"110000000",
  14413=>"000000000",
  14414=>"111110111",
  14415=>"011111111",
  14416=>"111111111",
  14417=>"000100100",
  14418=>"110110110",
  14419=>"100101111",
  14420=>"000000000",
  14421=>"111001100",
  14422=>"000000110",
  14423=>"000100000",
  14424=>"001111011",
  14425=>"111111101",
  14426=>"000000111",
  14427=>"011111111",
  14428=>"110111111",
  14429=>"000000000",
  14430=>"011111000",
  14431=>"001001001",
  14432=>"111010000",
  14433=>"000000000",
  14434=>"000011111",
  14435=>"101111111",
  14436=>"001001001",
  14437=>"101111110",
  14438=>"111111111",
  14439=>"100100100",
  14440=>"110000000",
  14441=>"000100000",
  14442=>"110111011",
  14443=>"001000000",
  14444=>"100100000",
  14445=>"011011101",
  14446=>"100000100",
  14447=>"000000000",
  14448=>"110111111",
  14449=>"111111111",
  14450=>"011010010",
  14451=>"001111111",
  14452=>"000100111",
  14453=>"000000101",
  14454=>"011000011",
  14455=>"111011010",
  14456=>"001000000",
  14457=>"000000000",
  14458=>"110110110",
  14459=>"001000000",
  14460=>"100111101",
  14461=>"000000000",
  14462=>"111111111",
  14463=>"011000010",
  14464=>"000000000",
  14465=>"100000010",
  14466=>"111100000",
  14467=>"110110111",
  14468=>"000000111",
  14469=>"000000000",
  14470=>"000000011",
  14471=>"001110000",
  14472=>"000000000",
  14473=>"100101000",
  14474=>"110111111",
  14475=>"011011001",
  14476=>"111111011",
  14477=>"001001000",
  14478=>"001001111",
  14479=>"000000011",
  14480=>"000001011",
  14481=>"000000001",
  14482=>"000000000",
  14483=>"111111111",
  14484=>"001011111",
  14485=>"000100000",
  14486=>"000000000",
  14487=>"111111110",
  14488=>"000000000",
  14489=>"011111111",
  14490=>"111001011",
  14491=>"000011011",
  14492=>"111101100",
  14493=>"001000000",
  14494=>"111111010",
  14495=>"110000000",
  14496=>"000000000",
  14497=>"010000001",
  14498=>"111111101",
  14499=>"011000000",
  14500=>"000001111",
  14501=>"111111111",
  14502=>"000000000",
  14503=>"111111001",
  14504=>"000100000",
  14505=>"001001011",
  14506=>"000100100",
  14507=>"000000000",
  14508=>"000000001",
  14509=>"010110001",
  14510=>"101000011",
  14511=>"100111111",
  14512=>"000000001",
  14513=>"111111001",
  14514=>"101111111",
  14515=>"011111111",
  14516=>"111111111",
  14517=>"111100111",
  14518=>"000000000",
  14519=>"011011001",
  14520=>"000000000",
  14521=>"111011000",
  14522=>"000100101",
  14523=>"111101000",
  14524=>"111110100",
  14525=>"110111111",
  14526=>"111111111",
  14527=>"111111101",
  14528=>"100000000",
  14529=>"001000000",
  14530=>"111111110",
  14531=>"111101111",
  14532=>"111111111",
  14533=>"000000000",
  14534=>"101001000",
  14535=>"110111111",
  14536=>"000101111",
  14537=>"001101000",
  14538=>"000000100",
  14539=>"000000111",
  14540=>"000000000",
  14541=>"010111101",
  14542=>"111000001",
  14543=>"110000010",
  14544=>"111111111",
  14545=>"111111111",
  14546=>"000100110",
  14547=>"001000000",
  14548=>"011111111",
  14549=>"000000000",
  14550=>"000000010",
  14551=>"000000111",
  14552=>"000000000",
  14553=>"100100111",
  14554=>"110000000",
  14555=>"011011001",
  14556=>"001101111",
  14557=>"000000000",
  14558=>"111011000",
  14559=>"111110110",
  14560=>"000000000",
  14561=>"000000000",
  14562=>"011010000",
  14563=>"001001000",
  14564=>"100100010",
  14565=>"000100000",
  14566=>"111100111",
  14567=>"011111111",
  14568=>"111111111",
  14569=>"110110111",
  14570=>"000000011",
  14571=>"000010111",
  14572=>"100100111",
  14573=>"001001000",
  14574=>"111010001",
  14575=>"011111111",
  14576=>"011011011",
  14577=>"111011111",
  14578=>"000000000",
  14579=>"001011001",
  14580=>"011111011",
  14581=>"000100100",
  14582=>"010111111",
  14583=>"111110110",
  14584=>"110110110",
  14585=>"000000000",
  14586=>"100100110",
  14587=>"111111111",
  14588=>"110111110",
  14589=>"001110110",
  14590=>"111111111",
  14591=>"000000011",
  14592=>"101000000",
  14593=>"000000100",
  14594=>"000000000",
  14595=>"111111111",
  14596=>"000001111",
  14597=>"111011001",
  14598=>"000000000",
  14599=>"001001111",
  14600=>"100010110",
  14601=>"000000011",
  14602=>"001000000",
  14603=>"000000011",
  14604=>"000000000",
  14605=>"111101000",
  14606=>"000100000",
  14607=>"000000000",
  14608=>"001000110",
  14609=>"000000000",
  14610=>"000000000",
  14611=>"001000100",
  14612=>"000000000",
  14613=>"000000100",
  14614=>"111111110",
  14615=>"110000000",
  14616=>"001101111",
  14617=>"111111111",
  14618=>"111001001",
  14619=>"000001000",
  14620=>"000000000",
  14621=>"111111111",
  14622=>"000000000",
  14623=>"000010000",
  14624=>"000000000",
  14625=>"000000000",
  14626=>"000000110",
  14627=>"001111100",
  14628=>"001000111",
  14629=>"111110101",
  14630=>"111111111",
  14631=>"010010111",
  14632=>"000110110",
  14633=>"101000000",
  14634=>"000100001",
  14635=>"111111000",
  14636=>"111111011",
  14637=>"101101101",
  14638=>"111111111",
  14639=>"001001111",
  14640=>"111011000",
  14641=>"101100000",
  14642=>"110000000",
  14643=>"001000000",
  14644=>"000000000",
  14645=>"011110110",
  14646=>"100110110",
  14647=>"101000000",
  14648=>"111111100",
  14649=>"100100000",
  14650=>"101101001",
  14651=>"000000110",
  14652=>"000000100",
  14653=>"100100011",
  14654=>"000111110",
  14655=>"111111111",
  14656=>"001001001",
  14657=>"111111111",
  14658=>"001000011",
  14659=>"111110111",
  14660=>"001000000",
  14661=>"111111111",
  14662=>"000010110",
  14663=>"000000111",
  14664=>"111111111",
  14665=>"001100100",
  14666=>"011011111",
  14667=>"111101011",
  14668=>"000100100",
  14669=>"000100111",
  14670=>"011111011",
  14671=>"000000111",
  14672=>"000000001",
  14673=>"011110110",
  14674=>"000000111",
  14675=>"000100110",
  14676=>"000000100",
  14677=>"011111111",
  14678=>"001001000",
  14679=>"111111101",
  14680=>"111111111",
  14681=>"000000000",
  14682=>"111111111",
  14683=>"000000000",
  14684=>"100000000",
  14685=>"111101000",
  14686=>"000000001",
  14687=>"100111110",
  14688=>"000000011",
  14689=>"000000000",
  14690=>"000000001",
  14691=>"000111111",
  14692=>"000100100",
  14693=>"000110111",
  14694=>"000000000",
  14695=>"111111011",
  14696=>"001000000",
  14697=>"000000010",
  14698=>"000000000",
  14699=>"001001001",
  14700=>"000100100",
  14701=>"100111111",
  14702=>"011111111",
  14703=>"111111111",
  14704=>"000000000",
  14705=>"000000001",
  14706=>"101101110",
  14707=>"111111111",
  14708=>"111111111",
  14709=>"111011111",
  14710=>"001000000",
  14711=>"011100110",
  14712=>"111111111",
  14713=>"111111001",
  14714=>"011111111",
  14715=>"000000000",
  14716=>"000000111",
  14717=>"000111000",
  14718=>"001000010",
  14719=>"111111110",
  14720=>"101101111",
  14721=>"000000000",
  14722=>"100110110",
  14723=>"000000111",
  14724=>"111111000",
  14725=>"110110000",
  14726=>"000000001",
  14727=>"111000010",
  14728=>"100111111",
  14729=>"111000001",
  14730=>"000000110",
  14731=>"000000110",
  14732=>"111111111",
  14733=>"111111101",
  14734=>"111111111",
  14735=>"001000000",
  14736=>"000000000",
  14737=>"111110000",
  14738=>"000000000",
  14739=>"001000000",
  14740=>"111111101",
  14741=>"011111100",
  14742=>"000000100",
  14743=>"110110111",
  14744=>"110110001",
  14745=>"001000100",
  14746=>"000000001",
  14747=>"000000000",
  14748=>"000000000",
  14749=>"111111111",
  14750=>"000000001",
  14751=>"111111010",
  14752=>"000000000",
  14753=>"001000001",
  14754=>"101000111",
  14755=>"011000000",
  14756=>"000000011",
  14757=>"111111111",
  14758=>"111111111",
  14759=>"001101111",
  14760=>"000000100",
  14761=>"001001000",
  14762=>"011001000",
  14763=>"000000000",
  14764=>"000000000",
  14765=>"000000000",
  14766=>"001000101",
  14767=>"111101001",
  14768=>"111111111",
  14769=>"111101110",
  14770=>"000000000",
  14771=>"111111111",
  14772=>"110111111",
  14773=>"111000001",
  14774=>"001111111",
  14775=>"111111111",
  14776=>"101110111",
  14777=>"101101111",
  14778=>"111111111",
  14779=>"011110100",
  14780=>"110000100",
  14781=>"111111111",
  14782=>"111111111",
  14783=>"110110100",
  14784=>"011001101",
  14785=>"111111111",
  14786=>"000000000",
  14787=>"001111111",
  14788=>"011011001",
  14789=>"001001111",
  14790=>"010110110",
  14791=>"111110110",
  14792=>"101101111",
  14793=>"011011111",
  14794=>"111111011",
  14795=>"000011111",
  14796=>"111111111",
  14797=>"000000001",
  14798=>"111110000",
  14799=>"001001000",
  14800=>"111111111",
  14801=>"001111101",
  14802=>"100100100",
  14803=>"000000000",
  14804=>"100000001",
  14805=>"000000001",
  14806=>"000000000",
  14807=>"110100000",
  14808=>"011111111",
  14809=>"000000000",
  14810=>"000000111",
  14811=>"111111111",
  14812=>"111111100",
  14813=>"100111111",
  14814=>"000000000",
  14815=>"000000100",
  14816=>"001001001",
  14817=>"100000110",
  14818=>"011010110",
  14819=>"111101101",
  14820=>"001011111",
  14821=>"101110111",
  14822=>"010011011",
  14823=>"111111111",
  14824=>"001111111",
  14825=>"000100000",
  14826=>"001000000",
  14827=>"111101111",
  14828=>"001000000",
  14829=>"111111111",
  14830=>"010011001",
  14831=>"100100000",
  14832=>"100100101",
  14833=>"001001000",
  14834=>"000000110",
  14835=>"010000000",
  14836=>"111001001",
  14837=>"000000111",
  14838=>"111111000",
  14839=>"111111111",
  14840=>"000000000",
  14841=>"111111111",
  14842=>"001111111",
  14843=>"000000000",
  14844=>"011000000",
  14845=>"111011011",
  14846=>"001001111",
  14847=>"111011011",
  14848=>"001111101",
  14849=>"111110010",
  14850=>"101000011",
  14851=>"000000111",
  14852=>"000100100",
  14853=>"010010010",
  14854=>"000110100",
  14855=>"111111111",
  14856=>"000000110",
  14857=>"111000000",
  14858=>"000000000",
  14859=>"111011111",
  14860=>"100000000",
  14861=>"110110100",
  14862=>"000000001",
  14863=>"110110000",
  14864=>"101100111",
  14865=>"000000111",
  14866=>"111111111",
  14867=>"111001000",
  14868=>"110000000",
  14869=>"000000111",
  14870=>"111011011",
  14871=>"001101100",
  14872=>"111001111",
  14873=>"000001110",
  14874=>"000001001",
  14875=>"011011101",
  14876=>"100100100",
  14877=>"011111111",
  14878=>"011001111",
  14879=>"110111111",
  14880=>"111000001",
  14881=>"101000101",
  14882=>"000110111",
  14883=>"000001111",
  14884=>"111111000",
  14885=>"001000000",
  14886=>"000111000",
  14887=>"110000000",
  14888=>"111111110",
  14889=>"111011000",
  14890=>"001101111",
  14891=>"000110010",
  14892=>"000111111",
  14893=>"011111111",
  14894=>"000000000",
  14895=>"111111111",
  14896=>"111111000",
  14897=>"100101101",
  14898=>"100100101",
  14899=>"000101101",
  14900=>"111111000",
  14901=>"110001000",
  14902=>"111000000",
  14903=>"001110111",
  14904=>"001010110",
  14905=>"111000001",
  14906=>"011000000",
  14907=>"000000011",
  14908=>"111111111",
  14909=>"111111101",
  14910=>"110000111",
  14911=>"001000111",
  14912=>"001000011",
  14913=>"001000100",
  14914=>"101111111",
  14915=>"100000110",
  14916=>"000000001",
  14917=>"000000000",
  14918=>"000111111",
  14919=>"111111111",
  14920=>"100000000",
  14921=>"111000001",
  14922=>"111110111",
  14923=>"000011111",
  14924=>"111111111",
  14925=>"000110000",
  14926=>"000000000",
  14927=>"111111100",
  14928=>"001001000",
  14929=>"000000001",
  14930=>"101001111",
  14931=>"001001001",
  14932=>"000100000",
  14933=>"001000100",
  14934=>"110100100",
  14935=>"111111000",
  14936=>"000100100",
  14937=>"001000000",
  14938=>"000011000",
  14939=>"100001011",
  14940=>"000100111",
  14941=>"111101000",
  14942=>"000000000",
  14943=>"000000111",
  14944=>"111001111",
  14945=>"000001001",
  14946=>"001000000",
  14947=>"000000111",
  14948=>"000010111",
  14949=>"100000111",
  14950=>"110100111",
  14951=>"111000000",
  14952=>"111111001",
  14953=>"111111111",
  14954=>"000000000",
  14955=>"011000000",
  14956=>"010101000",
  14957=>"000111000",
  14958=>"110110110",
  14959=>"111110000",
  14960=>"111011000",
  14961=>"011101110",
  14962=>"101001001",
  14963=>"101101100",
  14964=>"111000000",
  14965=>"111111000",
  14966=>"000000111",
  14967=>"111111100",
  14968=>"001000000",
  14969=>"000000000",
  14970=>"100000001",
  14971=>"000000011",
  14972=>"111111000",
  14973=>"001001000",
  14974=>"111111111",
  14975=>"111111100",
  14976=>"011000000",
  14977=>"111000101",
  14978=>"000111000",
  14979=>"000100100",
  14980=>"001011110",
  14981=>"111110000",
  14982=>"111111111",
  14983=>"011111111",
  14984=>"100000000",
  14985=>"001000010",
  14986=>"000100000",
  14987=>"001100000",
  14988=>"000000001",
  14989=>"000100000",
  14990=>"111001001",
  14991=>"111111111",
  14992=>"100000110",
  14993=>"111111001",
  14994=>"000000111",
  14995=>"111101000",
  14996=>"011000000",
  14997=>"111000100",
  14998=>"111100000",
  14999=>"011011000",
  15000=>"111111000",
  15001=>"111000000",
  15002=>"110000000",
  15003=>"000110111",
  15004=>"000000000",
  15005=>"101000101",
  15006=>"111111001",
  15007=>"110100100",
  15008=>"000000011",
  15009=>"111111011",
  15010=>"000111111",
  15011=>"111111111",
  15012=>"111100111",
  15013=>"000000000",
  15014=>"000111010",
  15015=>"101101001",
  15016=>"000000000",
  15017=>"001001111",
  15018=>"001011000",
  15019=>"000111111",
  15020=>"111111000",
  15021=>"101100100",
  15022=>"110111111",
  15023=>"111111111",
  15024=>"000000000",
  15025=>"000000100",
  15026=>"111111111",
  15027=>"111000001",
  15028=>"111110110",
  15029=>"010011111",
  15030=>"000000000",
  15031=>"111111111",
  15032=>"000000000",
  15033=>"000000000",
  15034=>"110110000",
  15035=>"110000000",
  15036=>"110110000",
  15037=>"111111111",
  15038=>"011011011",
  15039=>"110111111",
  15040=>"000110111",
  15041=>"111110111",
  15042=>"001000111",
  15043=>"000001111",
  15044=>"111110011",
  15045=>"111011000",
  15046=>"101011000",
  15047=>"111111110",
  15048=>"000000000",
  15049=>"111010110",
  15050=>"110111011",
  15051=>"111111010",
  15052=>"000010110",
  15053=>"000000010",
  15054=>"000111111",
  15055=>"100110100",
  15056=>"111010000",
  15057=>"111000001",
  15058=>"100000110",
  15059=>"111111000",
  15060=>"110110100",
  15061=>"110111110",
  15062=>"110000000",
  15063=>"000000000",
  15064=>"000000111",
  15065=>"000101111",
  15066=>"000000001",
  15067=>"110000110",
  15068=>"111001000",
  15069=>"000000100",
  15070=>"010111111",
  15071=>"111100010",
  15072=>"000000000",
  15073=>"111001000",
  15074=>"111111001",
  15075=>"110000000",
  15076=>"111111111",
  15077=>"010010110",
  15078=>"110111011",
  15079=>"111000111",
  15080=>"000100111",
  15081=>"001001001",
  15082=>"011000110",
  15083=>"111111111",
  15084=>"100000000",
  15085=>"111010000",
  15086=>"110100100",
  15087=>"111101111",
  15088=>"111111000",
  15089=>"000000111",
  15090=>"111011000",
  15091=>"010111011",
  15092=>"000000000",
  15093=>"001001001",
  15094=>"101111011",
  15095=>"000000000",
  15096=>"111111111",
  15097=>"111000000",
  15098=>"000000110",
  15099=>"111111000",
  15100=>"100111110",
  15101=>"111010110",
  15102=>"110000000",
  15103=>"000010111",
  15104=>"000000000",
  15105=>"111001001",
  15106=>"111101100",
  15107=>"100100000",
  15108=>"000001110",
  15109=>"000000000",
  15110=>"101111111",
  15111=>"110000111",
  15112=>"000000001",
  15113=>"000000000",
  15114=>"111110111",
  15115=>"111000000",
  15116=>"000000001",
  15117=>"001001000",
  15118=>"100100110",
  15119=>"000001111",
  15120=>"001000100",
  15121=>"111111111",
  15122=>"000000000",
  15123=>"111000000",
  15124=>"011011000",
  15125=>"101001000",
  15126=>"111100000",
  15127=>"000110111",
  15128=>"000000000",
  15129=>"100000000",
  15130=>"001100000",
  15131=>"000010011",
  15132=>"000000000",
  15133=>"000000000",
  15134=>"000000000",
  15135=>"110111111",
  15136=>"111101111",
  15137=>"001111111",
  15138=>"000111111",
  15139=>"111111100",
  15140=>"011000000",
  15141=>"001101011",
  15142=>"111111110",
  15143=>"000000111",
  15144=>"000000000",
  15145=>"111000100",
  15146=>"000000000",
  15147=>"001111111",
  15148=>"110111011",
  15149=>"000010011",
  15150=>"000000111",
  15151=>"000000100",
  15152=>"000000000",
  15153=>"000000000",
  15154=>"000000111",
  15155=>"111110010",
  15156=>"111111111",
  15157=>"101111111",
  15158=>"000000011",
  15159=>"101000000",
  15160=>"001001001",
  15161=>"000000000",
  15162=>"111010000",
  15163=>"000001001",
  15164=>"100100000",
  15165=>"111110000",
  15166=>"110110110",
  15167=>"111111111",
  15168=>"101000001",
  15169=>"001111111",
  15170=>"000000100",
  15171=>"111110000",
  15172=>"000000000",
  15173=>"000000000",
  15174=>"000000000",
  15175=>"111111111",
  15176=>"001000000",
  15177=>"000000101",
  15178=>"100000100",
  15179=>"111011011",
  15180=>"010000010",
  15181=>"111110111",
  15182=>"010001000",
  15183=>"011111111",
  15184=>"000000000",
  15185=>"111110100",
  15186=>"001101000",
  15187=>"110110110",
  15188=>"001111111",
  15189=>"111111011",
  15190=>"010001001",
  15191=>"101111100",
  15192=>"110111111",
  15193=>"000001111",
  15194=>"111111111",
  15195=>"011000110",
  15196=>"000000111",
  15197=>"111111001",
  15198=>"001011111",
  15199=>"111100100",
  15200=>"100111110",
  15201=>"000100110",
  15202=>"100101011",
  15203=>"111111111",
  15204=>"110101100",
  15205=>"110000000",
  15206=>"000000000",
  15207=>"111111111",
  15208=>"111100000",
  15209=>"000111111",
  15210=>"110101001",
  15211=>"101001001",
  15212=>"000001000",
  15213=>"110111000",
  15214=>"000000000",
  15215=>"000000111",
  15216=>"010000000",
  15217=>"111111111",
  15218=>"001011111",
  15219=>"101111111",
  15220=>"000000110",
  15221=>"000111111",
  15222=>"000111111",
  15223=>"000111111",
  15224=>"011111011",
  15225=>"101111100",
  15226=>"111010000",
  15227=>"110110000",
  15228=>"001000100",
  15229=>"011111111",
  15230=>"111110110",
  15231=>"000000001",
  15232=>"000100100",
  15233=>"111111110",
  15234=>"111111110",
  15235=>"111010000",
  15236=>"000000000",
  15237=>"001001000",
  15238=>"000000111",
  15239=>"110110000",
  15240=>"000000111",
  15241=>"111000111",
  15242=>"111111111",
  15243=>"001001111",
  15244=>"001000011",
  15245=>"110111111",
  15246=>"000100000",
  15247=>"011111111",
  15248=>"000000000",
  15249=>"000111111",
  15250=>"001110000",
  15251=>"111111111",
  15252=>"111001101",
  15253=>"010010000",
  15254=>"000000111",
  15255=>"101100000",
  15256=>"110110111",
  15257=>"000110110",
  15258=>"000000000",
  15259=>"000000000",
  15260=>"000010111",
  15261=>"000000001",
  15262=>"000010000",
  15263=>"111000000",
  15264=>"000010110",
  15265=>"111101000",
  15266=>"000000000",
  15267=>"000000000",
  15268=>"010111101",
  15269=>"111111001",
  15270=>"100100001",
  15271=>"000000000",
  15272=>"111101001",
  15273=>"011010000",
  15274=>"000000000",
  15275=>"101000000",
  15276=>"000100111",
  15277=>"110111001",
  15278=>"000001011",
  15279=>"110100100",
  15280=>"000111111",
  15281=>"110100100",
  15282=>"000100111",
  15283=>"110111111",
  15284=>"111111111",
  15285=>"000000000",
  15286=>"101101111",
  15287=>"000000000",
  15288=>"110110110",
  15289=>"000000111",
  15290=>"011111110",
  15291=>"100100111",
  15292=>"000001111",
  15293=>"001010000",
  15294=>"111101000",
  15295=>"101100000",
  15296=>"111101100",
  15297=>"000000000",
  15298=>"000010111",
  15299=>"111111111",
  15300=>"110111111",
  15301=>"111111001",
  15302=>"111111001",
  15303=>"011001000",
  15304=>"010000100",
  15305=>"010000010",
  15306=>"110000000",
  15307=>"001011000",
  15308=>"100100111",
  15309=>"111010000",
  15310=>"000000111",
  15311=>"010111111",
  15312=>"110000000",
  15313=>"000000010",
  15314=>"000000000",
  15315=>"000001001",
  15316=>"111111001",
  15317=>"001001000",
  15318=>"000000111",
  15319=>"010000001",
  15320=>"100110100",
  15321=>"000000111",
  15322=>"011110111",
  15323=>"100100000",
  15324=>"110111111",
  15325=>"111001111",
  15326=>"111100111",
  15327=>"110000000",
  15328=>"001001000",
  15329=>"011001011",
  15330=>"100001100",
  15331=>"000000000",
  15332=>"110100110",
  15333=>"000100110",
  15334=>"001000000",
  15335=>"000000110",
  15336=>"000100110",
  15337=>"000111111",
  15338=>"111111111",
  15339=>"111110110",
  15340=>"000000111",
  15341=>"000000110",
  15342=>"011011000",
  15343=>"001000010",
  15344=>"111111110",
  15345=>"000111011",
  15346=>"011000000",
  15347=>"111001001",
  15348=>"111111110",
  15349=>"011001000",
  15350=>"110110110",
  15351=>"111000100",
  15352=>"011111011",
  15353=>"000000010",
  15354=>"110111111",
  15355=>"001011111",
  15356=>"001001100",
  15357=>"111101001",
  15358=>"000110111",
  15359=>"001011011",
  15360=>"101000111",
  15361=>"111111000",
  15362=>"101101111",
  15363=>"111110011",
  15364=>"001001001",
  15365=>"001000000",
  15366=>"010111111",
  15367=>"111111101",
  15368=>"001000001",
  15369=>"111011011",
  15370=>"101001101",
  15371=>"111111000",
  15372=>"110110010",
  15373=>"000000000",
  15374=>"110110010",
  15375=>"000010000",
  15376=>"000000000",
  15377=>"111111110",
  15378=>"000000000",
  15379=>"000000000",
  15380=>"000000001",
  15381=>"000001111",
  15382=>"000000000",
  15383=>"101100100",
  15384=>"000000001",
  15385=>"000000000",
  15386=>"111111111",
  15387=>"000000100",
  15388=>"111111111",
  15389=>"001111111",
  15390=>"110111111",
  15391=>"001101000",
  15392=>"010011111",
  15393=>"000000000",
  15394=>"000000111",
  15395=>"111000000",
  15396=>"111111111",
  15397=>"001000000",
  15398=>"000000000",
  15399=>"000000000",
  15400=>"001111111",
  15401=>"111000000",
  15402=>"000000011",
  15403=>"111111010",
  15404=>"111001000",
  15405=>"000000000",
  15406=>"000000111",
  15407=>"111110100",
  15408=>"111111111",
  15409=>"011010010",
  15410=>"111001001",
  15411=>"000000000",
  15412=>"000100011",
  15413=>"000000100",
  15414=>"000000000",
  15415=>"010110111",
  15416=>"000011110",
  15417=>"001111011",
  15418=>"000111111",
  15419=>"001001111",
  15420=>"001001000",
  15421=>"111111010",
  15422=>"111111111",
  15423=>"011011011",
  15424=>"111101111",
  15425=>"111111111",
  15426=>"000000001",
  15427=>"111101111",
  15428=>"001001111",
  15429=>"110011000",
  15430=>"000000100",
  15431=>"000000000",
  15432=>"011011001",
  15433=>"111101111",
  15434=>"111111101",
  15435=>"000000000",
  15436=>"111111111",
  15437=>"000000000",
  15438=>"001001111",
  15439=>"111000000",
  15440=>"000010011",
  15441=>"111101000",
  15442=>"001000101",
  15443=>"001001000",
  15444=>"111111111",
  15445=>"110100000",
  15446=>"000000001",
  15447=>"100000000",
  15448=>"110010010",
  15449=>"101000100",
  15450=>"000000000",
  15451=>"010110110",
  15452=>"000110110",
  15453=>"000000001",
  15454=>"000001001",
  15455=>"000001001",
  15456=>"001000000",
  15457=>"000011111",
  15458=>"111111011",
  15459=>"101101111",
  15460=>"111111000",
  15461=>"111111101",
  15462=>"000011111",
  15463=>"000000000",
  15464=>"111111111",
  15465=>"001001111",
  15466=>"111010000",
  15467=>"111000000",
  15468=>"111111101",
  15469=>"111111110",
  15470=>"000000001",
  15471=>"000110111",
  15472=>"111111111",
  15473=>"000100111",
  15474=>"010000000",
  15475=>"000000000",
  15476=>"000000100",
  15477=>"010111111",
  15478=>"111011101",
  15479=>"100111111",
  15480=>"000000111",
  15481=>"111000000",
  15482=>"000000000",
  15483=>"000111111",
  15484=>"111111000",
  15485=>"001001001",
  15486=>"000000000",
  15487=>"001111011",
  15488=>"000000001",
  15489=>"000000011",
  15490=>"111000000",
  15491=>"000111111",
  15492=>"000000000",
  15493=>"111100000",
  15494=>"111111111",
  15495=>"000000000",
  15496=>"000000011",
  15497=>"111111111",
  15498=>"111111111",
  15499=>"001001111",
  15500=>"111111111",
  15501=>"111111110",
  15502=>"111111111",
  15503=>"000000000",
  15504=>"000000101",
  15505=>"000000000",
  15506=>"000000000",
  15507=>"001001001",
  15508=>"000111011",
  15509=>"010000000",
  15510=>"000010011",
  15511=>"000000000",
  15512=>"000000000",
  15513=>"111111010",
  15514=>"000111111",
  15515=>"111011111",
  15516=>"111111111",
  15517=>"111111111",
  15518=>"111111101",
  15519=>"000100100",
  15520=>"111110110",
  15521=>"111111111",
  15522=>"000000000",
  15523=>"111111111",
  15524=>"111100000",
  15525=>"001000100",
  15526=>"000000111",
  15527=>"000011001",
  15528=>"101000100",
  15529=>"001100000",
  15530=>"111111010",
  15531=>"011011011",
  15532=>"000000100",
  15533=>"111011111",
  15534=>"111111111",
  15535=>"111101000",
  15536=>"111011010",
  15537=>"000001000",
  15538=>"111111111",
  15539=>"000000000",
  15540=>"000000001",
  15541=>"001111111",
  15542=>"001000000",
  15543=>"111111111",
  15544=>"000000100",
  15545=>"111111111",
  15546=>"100000000",
  15547=>"110000101",
  15548=>"000000111",
  15549=>"100100111",
  15550=>"000000000",
  15551=>"000111111",
  15552=>"100000100",
  15553=>"101101111",
  15554=>"000000000",
  15555=>"000000000",
  15556=>"111111011",
  15557=>"000000001",
  15558=>"010000110",
  15559=>"110001001",
  15560=>"110010000",
  15561=>"111111111",
  15562=>"001000001",
  15563=>"000011011",
  15564=>"111101101",
  15565=>"000001011",
  15566=>"111000000",
  15567=>"000000011",
  15568=>"000110111",
  15569=>"111110111",
  15570=>"111111110",
  15571=>"100111000",
  15572=>"111101111",
  15573=>"000111011",
  15574=>"000000000",
  15575=>"111111111",
  15576=>"000000000",
  15577=>"000001001",
  15578=>"111111111",
  15579=>"011001000",
  15580=>"111111111",
  15581=>"001001101",
  15582=>"000000000",
  15583=>"000000000",
  15584=>"111100111",
  15585=>"110110110",
  15586=>"110110111",
  15587=>"000000000",
  15588=>"000011100",
  15589=>"111111001",
  15590=>"000000111",
  15591=>"000000000",
  15592=>"111111010",
  15593=>"111111111",
  15594=>"000000001",
  15595=>"001001000",
  15596=>"111001001",
  15597=>"001000000",
  15598=>"000000111",
  15599=>"001000000",
  15600=>"100111111",
  15601=>"000000000",
  15602=>"111111111",
  15603=>"000000000",
  15604=>"000000001",
  15605=>"000000000",
  15606=>"000000011",
  15607=>"111111111",
  15608=>"111111101",
  15609=>"010111110",
  15610=>"000000000",
  15611=>"101000000",
  15612=>"011001001",
  15613=>"011011111",
  15614=>"111111111",
  15615=>"010111010",
  15616=>"000000000",
  15617=>"011011001",
  15618=>"000000000",
  15619=>"001011000",
  15620=>"000000000",
  15621=>"000110110",
  15622=>"111111000",
  15623=>"110010000",
  15624=>"000011000",
  15625=>"000000000",
  15626=>"100000100",
  15627=>"000111011",
  15628=>"111000111",
  15629=>"111111101",
  15630=>"000001000",
  15631=>"111111111",
  15632=>"000111111",
  15633=>"110111111",
  15634=>"111111111",
  15635=>"000110111",
  15636=>"111111111",
  15637=>"000001001",
  15638=>"000000001",
  15639=>"100100000",
  15640=>"111111110",
  15641=>"111111011",
  15642=>"111111010",
  15643=>"000000000",
  15644=>"001000000",
  15645=>"000000001",
  15646=>"000000000",
  15647=>"000000011",
  15648=>"000000000",
  15649=>"111101111",
  15650=>"100100101",
  15651=>"111111111",
  15652=>"111100000",
  15653=>"111101111",
  15654=>"000000000",
  15655=>"000001011",
  15656=>"111110110",
  15657=>"000000000",
  15658=>"100110010",
  15659=>"111101001",
  15660=>"000000000",
  15661=>"000100010",
  15662=>"111111000",
  15663=>"000000000",
  15664=>"010010000",
  15665=>"110000000",
  15666=>"001000111",
  15667=>"110110000",
  15668=>"000000000",
  15669=>"110110010",
  15670=>"111011001",
  15671=>"100110111",
  15672=>"111110000",
  15673=>"101101111",
  15674=>"010010000",
  15675=>"000100111",
  15676=>"000011011",
  15677=>"000000000",
  15678=>"110000000",
  15679=>"000000000",
  15680=>"110100111",
  15681=>"000000000",
  15682=>"111111110",
  15683=>"010111010",
  15684=>"000101111",
  15685=>"001111111",
  15686=>"010111111",
  15687=>"000001011",
  15688=>"000000000",
  15689=>"000000000",
  15690=>"000000001",
  15691=>"100000100",
  15692=>"111111110",
  15693=>"100000000",
  15694=>"111101100",
  15695=>"001000000",
  15696=>"111111000",
  15697=>"000000011",
  15698=>"000000001",
  15699=>"000000110",
  15700=>"000000000",
  15701=>"011001001",
  15702=>"000000001",
  15703=>"000000000",
  15704=>"000000001",
  15705=>"000000000",
  15706=>"001011011",
  15707=>"111000010",
  15708=>"111000000",
  15709=>"111000100",
  15710=>"001000000",
  15711=>"111111100",
  15712=>"110011000",
  15713=>"011011001",
  15714=>"011111100",
  15715=>"111111000",
  15716=>"110111111",
  15717=>"000000000",
  15718=>"000000000",
  15719=>"111111010",
  15720=>"011001111",
  15721=>"000000111",
  15722=>"111111111",
  15723=>"111111111",
  15724=>"110110110",
  15725=>"001111111",
  15726=>"111001001",
  15727=>"000000011",
  15728=>"000000000",
  15729=>"111111111",
  15730=>"111111110",
  15731=>"111111111",
  15732=>"111111111",
  15733=>"000000000",
  15734=>"001001001",
  15735=>"001000000",
  15736=>"111111000",
  15737=>"000000000",
  15738=>"000000000",
  15739=>"000111111",
  15740=>"001000000",
  15741=>"111111110",
  15742=>"000000000",
  15743=>"101111111",
  15744=>"111001000",
  15745=>"000000111",
  15746=>"111111111",
  15747=>"100001000",
  15748=>"000000000",
  15749=>"000010111",
  15750=>"011110010",
  15751=>"001111111",
  15752=>"111011001",
  15753=>"000000110",
  15754=>"111001001",
  15755=>"010010000",
  15756=>"111111111",
  15757=>"111011011",
  15758=>"000110010",
  15759=>"000000000",
  15760=>"001000000",
  15761=>"001011011",
  15762=>"000010011",
  15763=>"010110111",
  15764=>"011000000",
  15765=>"000000000",
  15766=>"111000000",
  15767=>"100010001",
  15768=>"000000000",
  15769=>"111111011",
  15770=>"000000010",
  15771=>"000111111",
  15772=>"000000001",
  15773=>"111001010",
  15774=>"000000000",
  15775=>"000110110",
  15776=>"110110111",
  15777=>"000001001",
  15778=>"001000001",
  15779=>"111100100",
  15780=>"111111111",
  15781=>"111111111",
  15782=>"001000001",
  15783=>"000000000",
  15784=>"111001101",
  15785=>"111111100",
  15786=>"111000111",
  15787=>"111110000",
  15788=>"101000000",
  15789=>"111110101",
  15790=>"000000001",
  15791=>"000100100",
  15792=>"001000101",
  15793=>"000000000",
  15794=>"000000000",
  15795=>"001001000",
  15796=>"000000100",
  15797=>"001001000",
  15798=>"000000000",
  15799=>"000001111",
  15800=>"011000000",
  15801=>"111001111",
  15802=>"000000011",
  15803=>"011011000",
  15804=>"000000000",
  15805=>"000000000",
  15806=>"000100000",
  15807=>"010111000",
  15808=>"001000001",
  15809=>"000000000",
  15810=>"111111011",
  15811=>"111111111",
  15812=>"111111111",
  15813=>"011111111",
  15814=>"110000000",
  15815=>"000000001",
  15816=>"000000000",
  15817=>"101000010",
  15818=>"101100111",
  15819=>"111011000",
  15820=>"000000000",
  15821=>"000000000",
  15822=>"100000000",
  15823=>"000111111",
  15824=>"111111000",
  15825=>"111111000",
  15826=>"001111111",
  15827=>"000000000",
  15828=>"001111111",
  15829=>"111111111",
  15830=>"111101100",
  15831=>"111110001",
  15832=>"001111111",
  15833=>"110110010",
  15834=>"000001001",
  15835=>"001001001",
  15836=>"111111111",
  15837=>"000000000",
  15838=>"101000011",
  15839=>"000111100",
  15840=>"010110111",
  15841=>"000111001",
  15842=>"111111111",
  15843=>"110110111",
  15844=>"110110111",
  15845=>"111000101",
  15846=>"001001011",
  15847=>"000000000",
  15848=>"000000000",
  15849=>"111000000",
  15850=>"100111000",
  15851=>"100000000",
  15852=>"101000000",
  15853=>"110111111",
  15854=>"111111111",
  15855=>"000000111",
  15856=>"000000011",
  15857=>"011001000",
  15858=>"111111111",
  15859=>"000000100",
  15860=>"111111111",
  15861=>"000110100",
  15862=>"111111000",
  15863=>"011010000",
  15864=>"111111111",
  15865=>"001001001",
  15866=>"110010000",
  15867=>"011001111",
  15868=>"000000000",
  15869=>"111111111",
  15870=>"111111111",
  15871=>"000000111",
  15872=>"000001001",
  15873=>"111000000",
  15874=>"111000001",
  15875=>"010010111",
  15876=>"001001011",
  15877=>"000000000",
  15878=>"000000001",
  15879=>"111001111",
  15880=>"110111000",
  15881=>"110111111",
  15882=>"000000011",
  15883=>"111111010",
  15884=>"110100100",
  15885=>"111000000",
  15886=>"111000100",
  15887=>"000111110",
  15888=>"000000001",
  15889=>"000000111",
  15890=>"000000000",
  15891=>"111001000",
  15892=>"000000000",
  15893=>"111000000",
  15894=>"111100100",
  15895=>"000000011",
  15896=>"000001100",
  15897=>"000000001",
  15898=>"000000111",
  15899=>"111111000",
  15900=>"110111111",
  15901=>"000000000",
  15902=>"101101000",
  15903=>"000111111",
  15904=>"000111111",
  15905=>"111100000",
  15906=>"000001111",
  15907=>"111111000",
  15908=>"111000000",
  15909=>"111111111",
  15910=>"111000000",
  15911=>"111111000",
  15912=>"111111111",
  15913=>"001111111",
  15914=>"111110000",
  15915=>"110111010",
  15916=>"111011011",
  15917=>"000000000",
  15918=>"111111111",
  15919=>"000000100",
  15920=>"111111000",
  15921=>"000000111",
  15922=>"111110011",
  15923=>"000001111",
  15924=>"111111001",
  15925=>"001011111",
  15926=>"011111011",
  15927=>"001000000",
  15928=>"000000000",
  15929=>"111000000",
  15930=>"111111011",
  15931=>"010101000",
  15932=>"000000000",
  15933=>"011000000",
  15934=>"111111110",
  15935=>"000000000",
  15936=>"011111111",
  15937=>"111001000",
  15938=>"110111011",
  15939=>"000000000",
  15940=>"111001000",
  15941=>"001111111",
  15942=>"111000000",
  15943=>"001000001",
  15944=>"111111011",
  15945=>"111110101",
  15946=>"000000000",
  15947=>"111111111",
  15948=>"111111000",
  15949=>"000000011",
  15950=>"111011000",
  15951=>"110110000",
  15952=>"000000001",
  15953=>"111000000",
  15954=>"111111000",
  15955=>"101001111",
  15956=>"000000000",
  15957=>"000000000",
  15958=>"111111000",
  15959=>"100110100",
  15960=>"111111000",
  15961=>"100111100",
  15962=>"010111110",
  15963=>"111000000",
  15964=>"000111111",
  15965=>"110111011",
  15966=>"111000000",
  15967=>"101111111",
  15968=>"010000111",
  15969=>"111011000",
  15970=>"110110000",
  15971=>"001001000",
  15972=>"111111111",
  15973=>"111111001",
  15974=>"011000110",
  15975=>"100101111",
  15976=>"110111111",
  15977=>"111000110",
  15978=>"111000000",
  15979=>"111110000",
  15980=>"011010000",
  15981=>"111000011",
  15982=>"110000000",
  15983=>"100110111",
  15984=>"001111111",
  15985=>"000000111",
  15986=>"011000111",
  15987=>"000000100",
  15988=>"110000000",
  15989=>"001000000",
  15990=>"000000000",
  15991=>"000000111",
  15992=>"000111111",
  15993=>"000000111",
  15994=>"111111111",
  15995=>"000000000",
  15996=>"010000100",
  15997=>"010011111",
  15998=>"000000011",
  15999=>"100111110",
  16000=>"000000000",
  16001=>"111111000",
  16002=>"111000100",
  16003=>"000111111",
  16004=>"000000000",
  16005=>"000100000",
  16006=>"000110111",
  16007=>"000000000",
  16008=>"110000000",
  16009=>"000000100",
  16010=>"111000111",
  16011=>"111111111",
  16012=>"100111110",
  16013=>"111111111",
  16014=>"111000000",
  16015=>"001001000",
  16016=>"000111111",
  16017=>"000000001",
  16018=>"111111111",
  16019=>"100000010",
  16020=>"111001000",
  16021=>"000000101",
  16022=>"000111000",
  16023=>"000000010",
  16024=>"001000001",
  16025=>"111111111",
  16026=>"011000000",
  16027=>"111001000",
  16028=>"011000000",
  16029=>"000101111",
  16030=>"111111010",
  16031=>"001000000",
  16032=>"101111111",
  16033=>"000010111",
  16034=>"000000111",
  16035=>"000111111",
  16036=>"011011010",
  16037=>"000000111",
  16038=>"100000111",
  16039=>"000000001",
  16040=>"111000000",
  16041=>"111111111",
  16042=>"001001111",
  16043=>"000000100",
  16044=>"111101101",
  16045=>"000000000",
  16046=>"000000000",
  16047=>"001000111",
  16048=>"000110000",
  16049=>"000111110",
  16050=>"111111010",
  16051=>"111000000",
  16052=>"000000011",
  16053=>"010111111",
  16054=>"000000000",
  16055=>"100000000",
  16056=>"101000000",
  16057=>"000100111",
  16058=>"111011111",
  16059=>"001000000",
  16060=>"100000001",
  16061=>"110000111",
  16062=>"111000100",
  16063=>"000000000",
  16064=>"111110000",
  16065=>"000000111",
  16066=>"110110111",
  16067=>"111111001",
  16068=>"000111111",
  16069=>"101000000",
  16070=>"011011000",
  16071=>"101100000",
  16072=>"000110111",
  16073=>"000001000",
  16074=>"111111000",
  16075=>"111111111",
  16076=>"000000111",
  16077=>"000111001",
  16078=>"111101111",
  16079=>"111111000",
  16080=>"111111000",
  16081=>"111111111",
  16082=>"001111111",
  16083=>"111111000",
  16084=>"000001111",
  16085=>"011111111",
  16086=>"000000000",
  16087=>"001000000",
  16088=>"000000000",
  16089=>"000111111",
  16090=>"111111111",
  16091=>"000000000",
  16092=>"111111000",
  16093=>"111111001",
  16094=>"000000111",
  16095=>"000000000",
  16096=>"000000000",
  16097=>"110000000",
  16098=>"010111100",
  16099=>"111111111",
  16100=>"000001001",
  16101=>"111000000",
  16102=>"110111111",
  16103=>"111111000",
  16104=>"111111000",
  16105=>"000000001",
  16106=>"000000001",
  16107=>"101111000",
  16108=>"111111100",
  16109=>"000000000",
  16110=>"000001000",
  16111=>"000001000",
  16112=>"001000000",
  16113=>"000111111",
  16114=>"011011011",
  16115=>"000000000",
  16116=>"000011111",
  16117=>"111111111",
  16118=>"000111111",
  16119=>"111111011",
  16120=>"100000000",
  16121=>"000000111",
  16122=>"011111111",
  16123=>"000111000",
  16124=>"011111000",
  16125=>"011000000",
  16126=>"000000000",
  16127=>"000000001",
  16128=>"011000000",
  16129=>"011011001",
  16130=>"111111111",
  16131=>"111000000",
  16132=>"110111011",
  16133=>"111000110",
  16134=>"111111111",
  16135=>"000000000",
  16136=>"011011000",
  16137=>"000000111",
  16138=>"000000111",
  16139=>"011000101",
  16140=>"110100000",
  16141=>"100111111",
  16142=>"100110111",
  16143=>"001000110",
  16144=>"000000000",
  16145=>"001001111",
  16146=>"000000000",
  16147=>"000000011",
  16148=>"111111111",
  16149=>"100101000",
  16150=>"001000000",
  16151=>"000101111",
  16152=>"000111111",
  16153=>"000111111",
  16154=>"000000000",
  16155=>"111111111",
  16156=>"111111100",
  16157=>"111000100",
  16158=>"011000000",
  16159=>"111111000",
  16160=>"000000001",
  16161=>"000000011",
  16162=>"111111111",
  16163=>"101000000",
  16164=>"111111000",
  16165=>"001011111",
  16166=>"111111111",
  16167=>"000000000",
  16168=>"100000000",
  16169=>"000011010",
  16170=>"000000111",
  16171=>"111111111",
  16172=>"000100110",
  16173=>"000001110",
  16174=>"001001100",
  16175=>"111111011",
  16176=>"000011010",
  16177=>"001000000",
  16178=>"111111000",
  16179=>"000000111",
  16180=>"111100000",
  16181=>"100001111",
  16182=>"111111010",
  16183=>"011010000",
  16184=>"100101000",
  16185=>"000000000",
  16186=>"000100100",
  16187=>"000001111",
  16188=>"100111111",
  16189=>"001000000",
  16190=>"111101000",
  16191=>"000000000",
  16192=>"111101100",
  16193=>"000111111",
  16194=>"111111111",
  16195=>"110000000",
  16196=>"000000001",
  16197=>"000110000",
  16198=>"000000000",
  16199=>"010011000",
  16200=>"000000000",
  16201=>"011000000",
  16202=>"000111111",
  16203=>"110111001",
  16204=>"000000101",
  16205=>"110111111",
  16206=>"111000001",
  16207=>"000000110",
  16208=>"100000001",
  16209=>"000000000",
  16210=>"001110000",
  16211=>"000001111",
  16212=>"000000011",
  16213=>"000001001",
  16214=>"000000000",
  16215=>"000111111",
  16216=>"000000000",
  16217=>"011011000",
  16218=>"001000000",
  16219=>"000000000",
  16220=>"111001000",
  16221=>"001111111",
  16222=>"001000100",
  16223=>"010000000",
  16224=>"000000111",
  16225=>"111111111",
  16226=>"000011010",
  16227=>"011000011",
  16228=>"110110100",
  16229=>"000000001",
  16230=>"000000000",
  16231=>"111110111",
  16232=>"111111100",
  16233=>"000000000",
  16234=>"101101111",
  16235=>"111000000",
  16236=>"001001000",
  16237=>"000010000",
  16238=>"010000110",
  16239=>"111000111",
  16240=>"010110111",
  16241=>"010000111",
  16242=>"000000000",
  16243=>"000100111",
  16244=>"000010011",
  16245=>"000000111",
  16246=>"111111000",
  16247=>"000000000",
  16248=>"000111110",
  16249=>"110111111",
  16250=>"100000110",
  16251=>"000111111",
  16252=>"100100111",
  16253=>"111001111",
  16254=>"001000000",
  16255=>"001000000",
  16256=>"000110110",
  16257=>"111001000",
  16258=>"011111111",
  16259=>"000001000",
  16260=>"000000000",
  16261=>"111111111",
  16262=>"011000000",
  16263=>"111000000",
  16264=>"111000000",
  16265=>"111000110",
  16266=>"000000011",
  16267=>"111110010",
  16268=>"111111000",
  16269=>"000100110",
  16270=>"111111000",
  16271=>"000000111",
  16272=>"000000000",
  16273=>"111000000",
  16274=>"000000111",
  16275=>"011001111",
  16276=>"000001000",
  16277=>"000000000",
  16278=>"101111111",
  16279=>"011111111",
  16280=>"000000001",
  16281=>"111011111",
  16282=>"101000001",
  16283=>"111101100",
  16284=>"000000000",
  16285=>"010010110",
  16286=>"000000000",
  16287=>"110000000",
  16288=>"000000000",
  16289=>"010010011",
  16290=>"001111100",
  16291=>"000000000",
  16292=>"000111110",
  16293=>"111000111",
  16294=>"111111110",
  16295=>"000011110",
  16296=>"111100000",
  16297=>"111111111",
  16298=>"000000111",
  16299=>"000000000",
  16300=>"111111001",
  16301=>"011010000",
  16302=>"000100100",
  16303=>"000000000",
  16304=>"000000000",
  16305=>"000001001",
  16306=>"111000000",
  16307=>"000000000",
  16308=>"000000111",
  16309=>"111111000",
  16310=>"001100111",
  16311=>"111101000",
  16312=>"000000000",
  16313=>"111111100",
  16314=>"000101111",
  16315=>"001000000",
  16316=>"000000000",
  16317=>"111111000",
  16318=>"000000000",
  16319=>"111000000",
  16320=>"111011011",
  16321=>"100111111",
  16322=>"011011111",
  16323=>"111001000",
  16324=>"001011001",
  16325=>"000000111",
  16326=>"111111100",
  16327=>"101101000",
  16328=>"011000000",
  16329=>"011000000",
  16330=>"111111110",
  16331=>"001111111",
  16332=>"100000011",
  16333=>"000000111",
  16334=>"110000000",
  16335=>"000000111",
  16336=>"010000010",
  16337=>"000000001",
  16338=>"111011001",
  16339=>"111111111",
  16340=>"110111111",
  16341=>"000111111",
  16342=>"000111000",
  16343=>"011011011",
  16344=>"000000001",
  16345=>"000000000",
  16346=>"110111111",
  16347=>"011110000",
  16348=>"111111001",
  16349=>"000000000",
  16350=>"011000000",
  16351=>"001011011",
  16352=>"111111101",
  16353=>"100000000",
  16354=>"000000000",
  16355=>"000000111",
  16356=>"111111111",
  16357=>"011011111",
  16358=>"111000000",
  16359=>"000000111",
  16360=>"111000001",
  16361=>"000000000",
  16362=>"000000011",
  16363=>"000111111",
  16364=>"111000000",
  16365=>"101000000",
  16366=>"010111000",
  16367=>"000000100",
  16368=>"111111111",
  16369=>"000000011",
  16370=>"001000000",
  16371=>"011011000",
  16372=>"011000000",
  16373=>"111111111",
  16374=>"111111111",
  16375=>"001001001",
  16376=>"111111011",
  16377=>"111011000",
  16378=>"000000001",
  16379=>"101000001",
  16380=>"111111000",
  16381=>"000000100",
  16382=>"000001111",
  16383=>"001000111",
  16384=>"000100000",
  16385=>"111111000",
  16386=>"111000000",
  16387=>"001111000",
  16388=>"000110110",
  16389=>"111111111",
  16390=>"000000000",
  16391=>"111111000",
  16392=>"100101101",
  16393=>"010111010",
  16394=>"000000000",
  16395=>"100000000",
  16396=>"000000100",
  16397=>"111111111",
  16398=>"000110110",
  16399=>"000000010",
  16400=>"000000111",
  16401=>"000000111",
  16402=>"000000000",
  16403=>"111111111",
  16404=>"001000000",
  16405=>"000010011",
  16406=>"111000000",
  16407=>"000001001",
  16408=>"111111111",
  16409=>"000000111",
  16410=>"111111111",
  16411=>"111111001",
  16412=>"000100110",
  16413=>"111111111",
  16414=>"000000111",
  16415=>"110111111",
  16416=>"000000000",
  16417=>"111111111",
  16418=>"000000011",
  16419=>"100000000",
  16420=>"000111111",
  16421=>"111111001",
  16422=>"111111100",
  16423=>"111101000",
  16424=>"000000000",
  16425=>"000000000",
  16426=>"011001000",
  16427=>"111000111",
  16428=>"000100111",
  16429=>"111111000",
  16430=>"100100000",
  16431=>"111000000",
  16432=>"111101000",
  16433=>"000000000",
  16434=>"000000000",
  16435=>"100000000",
  16436=>"000100000",
  16437=>"111111000",
  16438=>"000000011",
  16439=>"110011111",
  16440=>"000111111",
  16441=>"111110100",
  16442=>"000000000",
  16443=>"111001000",
  16444=>"111111000",
  16445=>"111000000",
  16446=>"000010011",
  16447=>"111010111",
  16448=>"000000000",
  16449=>"000000000",
  16450=>"111111000",
  16451=>"000000000",
  16452=>"110000000",
  16453=>"111001000",
  16454=>"111111000",
  16455=>"001011000",
  16456=>"000111111",
  16457=>"000000000",
  16458=>"001001001",
  16459=>"000000111",
  16460=>"111111111",
  16461=>"000000111",
  16462=>"100000000",
  16463=>"000010000",
  16464=>"111011000",
  16465=>"000010100",
  16466=>"100100111",
  16467=>"000000000",
  16468=>"000000000",
  16469=>"000000011",
  16470=>"111100100",
  16471=>"000000111",
  16472=>"111111000",
  16473=>"000000000",
  16474=>"110100100",
  16475=>"100100000",
  16476=>"000001011",
  16477=>"011011001",
  16478=>"110010000",
  16479=>"101011000",
  16480=>"111000000",
  16481=>"000111111",
  16482=>"111011011",
  16483=>"111000111",
  16484=>"111111011",
  16485=>"000001000",
  16486=>"000000000",
  16487=>"000000000",
  16488=>"000111111",
  16489=>"110100111",
  16490=>"111111011",
  16491=>"111110000",
  16492=>"000000000",
  16493=>"000111111",
  16494=>"001000011",
  16495=>"111011011",
  16496=>"111111000",
  16497=>"100000100",
  16498=>"011111111",
  16499=>"111001000",
  16500=>"000000111",
  16501=>"000000001",
  16502=>"000000000",
  16503=>"110000000",
  16504=>"000000000",
  16505=>"101011000",
  16506=>"000000000",
  16507=>"000010010",
  16508=>"111101101",
  16509=>"011111011",
  16510=>"010000011",
  16511=>"000000111",
  16512=>"000011010",
  16513=>"011001000",
  16514=>"100000000",
  16515=>"001001000",
  16516=>"111011000",
  16517=>"111110010",
  16518=>"000110111",
  16519=>"000100111",
  16520=>"111111000",
  16521=>"111000000",
  16522=>"100100100",
  16523=>"000000000",
  16524=>"011100001",
  16525=>"111111111",
  16526=>"000000111",
  16527=>"000000000",
  16528=>"000000111",
  16529=>"110111110",
  16530=>"000010111",
  16531=>"100111111",
  16532=>"000000000",
  16533=>"111000000",
  16534=>"000000111",
  16535=>"100100100",
  16536=>"000111001",
  16537=>"101100111",
  16538=>"110111100",
  16539=>"000010111",
  16540=>"011000000",
  16541=>"000010010",
  16542=>"000000000",
  16543=>"101111111",
  16544=>"111101010",
  16545=>"110000000",
  16546=>"100110111",
  16547=>"100111000",
  16548=>"110000000",
  16549=>"100111111",
  16550=>"111111011",
  16551=>"111111101",
  16552=>"111000000",
  16553=>"111100000",
  16554=>"000111000",
  16555=>"000001111",
  16556=>"111110110",
  16557=>"100001111",
  16558=>"100000000",
  16559=>"000100111",
  16560=>"101111000",
  16561=>"000011111",
  16562=>"011011111",
  16563=>"000100101",
  16564=>"111111000",
  16565=>"111001111",
  16566=>"000110110",
  16567=>"000000001",
  16568=>"111111111",
  16569=>"111111111",
  16570=>"110000000",
  16571=>"000001011",
  16572=>"111001001",
  16573=>"000000111",
  16574=>"111111111",
  16575=>"011000000",
  16576=>"000000000",
  16577=>"111000000",
  16578=>"000110111",
  16579=>"111111010",
  16580=>"000111111",
  16581=>"010111000",
  16582=>"000001011",
  16583=>"111111111",
  16584=>"010111110",
  16585=>"000000000",
  16586=>"110100000",
  16587=>"111111000",
  16588=>"111000000",
  16589=>"111111111",
  16590=>"111011000",
  16591=>"001000000",
  16592=>"101000000",
  16593=>"111001001",
  16594=>"000000000",
  16595=>"000000001",
  16596=>"000100000",
  16597=>"001000100",
  16598=>"011111000",
  16599=>"111111111",
  16600=>"000000111",
  16601=>"111111111",
  16602=>"000100111",
  16603=>"000000000",
  16604=>"111111110",
  16605=>"000000000",
  16606=>"000111111",
  16607=>"001111000",
  16608=>"010000000",
  16609=>"110111111",
  16610=>"000110111",
  16611=>"111111000",
  16612=>"000111011",
  16613=>"000000000",
  16614=>"000000000",
  16615=>"111111111",
  16616=>"100000000",
  16617=>"011001111",
  16618=>"001000000",
  16619=>"110111111",
  16620=>"000000011",
  16621=>"111010000",
  16622=>"000100110",
  16623=>"111111111",
  16624=>"111011000",
  16625=>"000000111",
  16626=>"000000111",
  16627=>"110111000",
  16628=>"111111111",
  16629=>"111000000",
  16630=>"001110111",
  16631=>"100000000",
  16632=>"110000000",
  16633=>"000000000",
  16634=>"111101111",
  16635=>"111111000",
  16636=>"001011111",
  16637=>"000000001",
  16638=>"000000001",
  16639=>"111001000",
  16640=>"000000000",
  16641=>"100110111",
  16642=>"011001001",
  16643=>"000100111",
  16644=>"001000000",
  16645=>"100011010",
  16646=>"111011011",
  16647=>"001100111",
  16648=>"111101100",
  16649=>"000000111",
  16650=>"111000000",
  16651=>"000111111",
  16652=>"111000000",
  16653=>"000000000",
  16654=>"000000000",
  16655=>"000000000",
  16656=>"111011011",
  16657=>"111110111",
  16658=>"111001000",
  16659=>"000000000",
  16660=>"111111110",
  16661=>"000110111",
  16662=>"011111011",
  16663=>"110011111",
  16664=>"111111111",
  16665=>"000111111",
  16666=>"111111111",
  16667=>"100110111",
  16668=>"011111001",
  16669=>"000000111",
  16670=>"101100111",
  16671=>"011010100",
  16672=>"110110111",
  16673=>"000000111",
  16674=>"000000000",
  16675=>"111111111",
  16676=>"111000000",
  16677=>"011000001",
  16678=>"000000000",
  16679=>"111111110",
  16680=>"100111110",
  16681=>"000000000",
  16682=>"100110111",
  16683=>"011010000",
  16684=>"111100000",
  16685=>"000111111",
  16686=>"111110111",
  16687=>"000010000",
  16688=>"111100100",
  16689=>"011111111",
  16690=>"111111111",
  16691=>"111000001",
  16692=>"000000000",
  16693=>"000001111",
  16694=>"111000111",
  16695=>"000111000",
  16696=>"000000100",
  16697=>"101111111",
  16698=>"000000001",
  16699=>"100111101",
  16700=>"001000000",
  16701=>"111111111",
  16702=>"000000111",
  16703=>"000000001",
  16704=>"000110111",
  16705=>"000100111",
  16706=>"111111000",
  16707=>"000000000",
  16708=>"111110111",
  16709=>"111111111",
  16710=>"000111110",
  16711=>"011010000",
  16712=>"000000111",
  16713=>"000000000",
  16714=>"110000001",
  16715=>"000000101",
  16716=>"000010011",
  16717=>"000001111",
  16718=>"111111111",
  16719=>"110111111",
  16720=>"101101111",
  16721=>"110111001",
  16722=>"000000111",
  16723=>"000000011",
  16724=>"000011111",
  16725=>"111011111",
  16726=>"000101100",
  16727=>"111000000",
  16728=>"000010111",
  16729=>"000000001",
  16730=>"000111111",
  16731=>"111111111",
  16732=>"100100110",
  16733=>"111111111",
  16734=>"111111000",
  16735=>"001011111",
  16736=>"000100100",
  16737=>"100000011",
  16738=>"000111111",
  16739=>"011111000",
  16740=>"001001000",
  16741=>"000000000",
  16742=>"000000111",
  16743=>"000000111",
  16744=>"000000000",
  16745=>"111000001",
  16746=>"011000010",
  16747=>"000000111",
  16748=>"110111001",
  16749=>"000000000",
  16750=>"000000111",
  16751=>"000000111",
  16752=>"011001000",
  16753=>"111111111",
  16754=>"011111000",
  16755=>"000000100",
  16756=>"000000000",
  16757=>"100111001",
  16758=>"010000101",
  16759=>"100000111",
  16760=>"111000000",
  16761=>"011000111",
  16762=>"111000001",
  16763=>"000111111",
  16764=>"000000001",
  16765=>"111111111",
  16766=>"011111001",
  16767=>"000000111",
  16768=>"110111011",
  16769=>"111111111",
  16770=>"111110001",
  16771=>"111000000",
  16772=>"111111111",
  16773=>"110110100",
  16774=>"100011111",
  16775=>"111111111",
  16776=>"111000111",
  16777=>"111111111",
  16778=>"111111000",
  16779=>"111100111",
  16780=>"111011111",
  16781=>"000000000",
  16782=>"000000011",
  16783=>"111000000",
  16784=>"111111110",
  16785=>"000111100",
  16786=>"100110000",
  16787=>"110000001",
  16788=>"111111111",
  16789=>"001011001",
  16790=>"101000001",
  16791=>"000001001",
  16792=>"000000011",
  16793=>"000110110",
  16794=>"000000100",
  16795=>"000001000",
  16796=>"101100000",
  16797=>"111100110",
  16798=>"011001000",
  16799=>"001000000",
  16800=>"111111000",
  16801=>"001110111",
  16802=>"000000000",
  16803=>"111000100",
  16804=>"101000101",
  16805=>"111111000",
  16806=>"100000001",
  16807=>"100000111",
  16808=>"111011001",
  16809=>"011011111",
  16810=>"111111111",
  16811=>"110110111",
  16812=>"111011010",
  16813=>"111111111",
  16814=>"111101110",
  16815=>"111111111",
  16816=>"111111000",
  16817=>"111111111",
  16818=>"001101000",
  16819=>"111110101",
  16820=>"000000000",
  16821=>"000000010",
  16822=>"000110111",
  16823=>"111011011",
  16824=>"000101111",
  16825=>"111011111",
  16826=>"100001101",
  16827=>"110111111",
  16828=>"000001000",
  16829=>"100111101",
  16830=>"000111111",
  16831=>"000000000",
  16832=>"000111011",
  16833=>"110010010",
  16834=>"000111111",
  16835=>"111111111",
  16836=>"010100101",
  16837=>"111000000",
  16838=>"000000000",
  16839=>"111100000",
  16840=>"000000011",
  16841=>"100000000",
  16842=>"100000000",
  16843=>"111000111",
  16844=>"000000111",
  16845=>"111111111",
  16846=>"110100111",
  16847=>"111100111",
  16848=>"000000111",
  16849=>"000000010",
  16850=>"000010000",
  16851=>"111111011",
  16852=>"010100100",
  16853=>"111010000",
  16854=>"000000000",
  16855=>"000000011",
  16856=>"111000000",
  16857=>"000000110",
  16858=>"010000000",
  16859=>"000000000",
  16860=>"000000111",
  16861=>"111001111",
  16862=>"001000000",
  16863=>"111111000",
  16864=>"110000000",
  16865=>"111111111",
  16866=>"000000000",
  16867=>"111111011",
  16868=>"011111111",
  16869=>"000000000",
  16870=>"111111110",
  16871=>"000000111",
  16872=>"000100110",
  16873=>"000000000",
  16874=>"011000111",
  16875=>"100111111",
  16876=>"000000111",
  16877=>"001101111",
  16878=>"000111000",
  16879=>"011011111",
  16880=>"110111111",
  16881=>"011111111",
  16882=>"110000000",
  16883=>"100101000",
  16884=>"100110010",
  16885=>"111111001",
  16886=>"111111101",
  16887=>"000000011",
  16888=>"010010000",
  16889=>"000001101",
  16890=>"111111000",
  16891=>"000000111",
  16892=>"111011111",
  16893=>"011111110",
  16894=>"001000000",
  16895=>"000000000",
  16896=>"000000001",
  16897=>"111111111",
  16898=>"001100000",
  16899=>"111111111",
  16900=>"100100100",
  16901=>"111111100",
  16902=>"111100111",
  16903=>"111111111",
  16904=>"111111111",
  16905=>"000000000",
  16906=>"010000000",
  16907=>"010000101",
  16908=>"001011111",
  16909=>"000000000",
  16910=>"100000000",
  16911=>"000000010",
  16912=>"000000001",
  16913=>"000000000",
  16914=>"110110000",
  16915=>"001111111",
  16916=>"000000000",
  16917=>"001001001",
  16918=>"111111111",
  16919=>"000000000",
  16920=>"000000000",
  16921=>"001111111",
  16922=>"000000000",
  16923=>"011111111",
  16924=>"111111111",
  16925=>"000000000",
  16926=>"110000000",
  16927=>"111111101",
  16928=>"001110111",
  16929=>"111111110",
  16930=>"000000110",
  16931=>"000000001",
  16932=>"000100111",
  16933=>"111111111",
  16934=>"110000100",
  16935=>"011000000",
  16936=>"111111111",
  16937=>"001000000",
  16938=>"011011111",
  16939=>"100111111",
  16940=>"000000111",
  16941=>"000000100",
  16942=>"111111111",
  16943=>"111111110",
  16944=>"000100100",
  16945=>"001011011",
  16946=>"001111111",
  16947=>"000000100",
  16948=>"000100100",
  16949=>"100100100",
  16950=>"111110111",
  16951=>"111111101",
  16952=>"111011111",
  16953=>"001010111",
  16954=>"111011011",
  16955=>"000100000",
  16956=>"001001111",
  16957=>"000000000",
  16958=>"000110101",
  16959=>"010110111",
  16960=>"000000000",
  16961=>"110110110",
  16962=>"010111111",
  16963=>"111111111",
  16964=>"001001001",
  16965=>"111111100",
  16966=>"111110111",
  16967=>"001000000",
  16968=>"111111111",
  16969=>"001001000",
  16970=>"101000000",
  16971=>"111000000",
  16972=>"111111111",
  16973=>"000000101",
  16974=>"001011000",
  16975=>"000000000",
  16976=>"000000000",
  16977=>"111111111",
  16978=>"000000000",
  16979=>"000000000",
  16980=>"000000000",
  16981=>"000011110",
  16982=>"101110111",
  16983=>"010110010",
  16984=>"111100000",
  16985=>"000000000",
  16986=>"111111111",
  16987=>"110110000",
  16988=>"111111111",
  16989=>"011111011",
  16990=>"111111111",
  16991=>"111111111",
  16992=>"000101001",
  16993=>"001110100",
  16994=>"111111111",
  16995=>"111111111",
  16996=>"000000100",
  16997=>"000011111",
  16998=>"111100000",
  16999=>"001110110",
  17000=>"111111111",
  17001=>"111111111",
  17002=>"111010111",
  17003=>"000000000",
  17004=>"100000001",
  17005=>"111111111",
  17006=>"111111111",
  17007=>"001110000",
  17008=>"111110110",
  17009=>"110000111",
  17010=>"001011011",
  17011=>"000000000",
  17012=>"001000000",
  17013=>"000000000",
  17014=>"000000000",
  17015=>"111000000",
  17016=>"000000000",
  17017=>"000000000",
  17018=>"011111101",
  17019=>"111111111",
  17020=>"000000000",
  17021=>"000000000",
  17022=>"111111111",
  17023=>"000000000",
  17024=>"111111111",
  17025=>"111000000",
  17026=>"000000000",
  17027=>"011011001",
  17028=>"000000000",
  17029=>"100000101",
  17030=>"111111111",
  17031=>"111111111",
  17032=>"000000000",
  17033=>"111110110",
  17034=>"111111111",
  17035=>"000000000",
  17036=>"111101100",
  17037=>"111111111",
  17038=>"101001000",
  17039=>"000000111",
  17040=>"001001011",
  17041=>"000110110",
  17042=>"000000000",
  17043=>"010111111",
  17044=>"000000000",
  17045=>"111111111",
  17046=>"000000000",
  17047=>"000000000",
  17048=>"111001111",
  17049=>"111111111",
  17050=>"110111110",
  17051=>"000000000",
  17052=>"111111110",
  17053=>"001000000",
  17054=>"000000000",
  17055=>"000000000",
  17056=>"101000000",
  17057=>"101110111",
  17058=>"111111111",
  17059=>"001000000",
  17060=>"000110111",
  17061=>"111011101",
  17062=>"000000111",
  17063=>"000011011",
  17064=>"000000101",
  17065=>"000000000",
  17066=>"110111111",
  17067=>"000000000",
  17068=>"000000000",
  17069=>"110100000",
  17070=>"000001101",
  17071=>"111111110",
  17072=>"000000000",
  17073=>"111111111",
  17074=>"111111111",
  17075=>"010101111",
  17076=>"110111111",
  17077=>"111000000",
  17078=>"000000010",
  17079=>"111111111",
  17080=>"011001111",
  17081=>"000000000",
  17082=>"000000000",
  17083=>"000000000",
  17084=>"111111111",
  17085=>"111111000",
  17086=>"111111111",
  17087=>"011011111",
  17088=>"000000000",
  17089=>"100000000",
  17090=>"111110000",
  17091=>"111111111",
  17092=>"000000000",
  17093=>"000100110",
  17094=>"000000000",
  17095=>"101000001",
  17096=>"011111010",
  17097=>"111111111",
  17098=>"000000000",
  17099=>"111111111",
  17100=>"110110111",
  17101=>"000001000",
  17102=>"100000000",
  17103=>"000000000",
  17104=>"111110000",
  17105=>"111111111",
  17106=>"010000111",
  17107=>"000000000",
  17108=>"000000000",
  17109=>"000000000",
  17110=>"000110110",
  17111=>"101111111",
  17112=>"111100110",
  17113=>"100000101",
  17114=>"111011011",
  17115=>"000000000",
  17116=>"111111111",
  17117=>"111110111",
  17118=>"000000000",
  17119=>"000010000",
  17120=>"000000000",
  17121=>"111111111",
  17122=>"010000000",
  17123=>"000000101",
  17124=>"111111111",
  17125=>"111000111",
  17126=>"111111000",
  17127=>"111111111",
  17128=>"111111111",
  17129=>"000000000",
  17130=>"111111111",
  17131=>"111111111",
  17132=>"000000010",
  17133=>"000000000",
  17134=>"000000000",
  17135=>"111111001",
  17136=>"100000000",
  17137=>"000000000",
  17138=>"000100001",
  17139=>"000000000",
  17140=>"111110111",
  17141=>"111111111",
  17142=>"111111001",
  17143=>"101000001",
  17144=>"000001101",
  17145=>"100000000",
  17146=>"111011111",
  17147=>"000000000",
  17148=>"111111111",
  17149=>"111111011",
  17150=>"000010011",
  17151=>"000000000",
  17152=>"000110111",
  17153=>"001011011",
  17154=>"001101000",
  17155=>"111111111",
  17156=>"000000000",
  17157=>"110110111",
  17158=>"111111111",
  17159=>"110100110",
  17160=>"111111111",
  17161=>"010000000",
  17162=>"100000000",
  17163=>"000000001",
  17164=>"111000000",
  17165=>"000000000",
  17166=>"000000000",
  17167=>"111101000",
  17168=>"110111111",
  17169=>"111111111",
  17170=>"000000000",
  17171=>"000000000",
  17172=>"000000000",
  17173=>"111101111",
  17174=>"000000000",
  17175=>"001011000",
  17176=>"111110111",
  17177=>"111111000",
  17178=>"000000000",
  17179=>"111001000",
  17180=>"111111111",
  17181=>"000111111",
  17182=>"010111111",
  17183=>"111111110",
  17184=>"000000000",
  17185=>"010111001",
  17186=>"110000000",
  17187=>"000000000",
  17188=>"110000000",
  17189=>"111000000",
  17190=>"111111111",
  17191=>"011000001",
  17192=>"010010000",
  17193=>"000000000",
  17194=>"111111110",
  17195=>"011010011",
  17196=>"111111111",
  17197=>"110100110",
  17198=>"111111111",
  17199=>"111001000",
  17200=>"000000000",
  17201=>"111111111",
  17202=>"010000110",
  17203=>"010000000",
  17204=>"100101111",
  17205=>"111111111",
  17206=>"110110000",
  17207=>"000000000",
  17208=>"001000000",
  17209=>"000000000",
  17210=>"110111111",
  17211=>"000000000",
  17212=>"101000101",
  17213=>"111111001",
  17214=>"000000000",
  17215=>"000000000",
  17216=>"111111000",
  17217=>"110111111",
  17218=>"000000000",
  17219=>"111100000",
  17220=>"000000110",
  17221=>"000000110",
  17222=>"000000000",
  17223=>"000000000",
  17224=>"000000001",
  17225=>"111100100",
  17226=>"011000000",
  17227=>"000000000",
  17228=>"000000000",
  17229=>"001000000",
  17230=>"111111111",
  17231=>"100000010",
  17232=>"000000001",
  17233=>"111111111",
  17234=>"000000000",
  17235=>"111111101",
  17236=>"111111111",
  17237=>"001000000",
  17238=>"000100111",
  17239=>"111111111",
  17240=>"111010000",
  17241=>"010011111",
  17242=>"000110111",
  17243=>"000001111",
  17244=>"000000000",
  17245=>"000000000",
  17246=>"000000000",
  17247=>"111111110",
  17248=>"000000000",
  17249=>"111111100",
  17250=>"001000000",
  17251=>"000000000",
  17252=>"000110000",
  17253=>"111001000",
  17254=>"000000000",
  17255=>"111001101",
  17256=>"000001000",
  17257=>"101111111",
  17258=>"000000111",
  17259=>"110110111",
  17260=>"000001000",
  17261=>"000000000",
  17262=>"000000000",
  17263=>"000001011",
  17264=>"101000100",
  17265=>"000000000",
  17266=>"111111000",
  17267=>"111111111",
  17268=>"000000000",
  17269=>"000000100",
  17270=>"000000000",
  17271=>"000000000",
  17272=>"111111111",
  17273=>"000000000",
  17274=>"000000110",
  17275=>"111001000",
  17276=>"000000000",
  17277=>"000000000",
  17278=>"111111111",
  17279=>"111111111",
  17280=>"000000010",
  17281=>"111111110",
  17282=>"110111111",
  17283=>"000000000",
  17284=>"000000011",
  17285=>"000000000",
  17286=>"111111111",
  17287=>"000100111",
  17288=>"000000000",
  17289=>"111111111",
  17290=>"111000111",
  17291=>"111111111",
  17292=>"000011000",
  17293=>"000000110",
  17294=>"010010000",
  17295=>"000100111",
  17296=>"000000001",
  17297=>"111000000",
  17298=>"000000000",
  17299=>"010111011",
  17300=>"000000001",
  17301=>"000000000",
  17302=>"000100101",
  17303=>"001000000",
  17304=>"011011111",
  17305=>"110111111",
  17306=>"111000000",
  17307=>"111110111",
  17308=>"000000001",
  17309=>"111010111",
  17310=>"111011011",
  17311=>"100100110",
  17312=>"000000000",
  17313=>"000000000",
  17314=>"100101001",
  17315=>"111111111",
  17316=>"000000111",
  17317=>"110100000",
  17318=>"011011111",
  17319=>"011111111",
  17320=>"000000001",
  17321=>"111000000",
  17322=>"101000000",
  17323=>"000000000",
  17324=>"101101101",
  17325=>"110000000",
  17326=>"000000011",
  17327=>"111111111",
  17328=>"111000010",
  17329=>"000000000",
  17330=>"000000111",
  17331=>"111001000",
  17332=>"000000000",
  17333=>"000000000",
  17334=>"000110000",
  17335=>"111110000",
  17336=>"010000000",
  17337=>"000010111",
  17338=>"000100000",
  17339=>"111111111",
  17340=>"111111111",
  17341=>"111111111",
  17342=>"100000000",
  17343=>"011011000",
  17344=>"000000111",
  17345=>"000000000",
  17346=>"111111111",
  17347=>"000111000",
  17348=>"111111001",
  17349=>"001000111",
  17350=>"111110011",
  17351=>"111001000",
  17352=>"111000101",
  17353=>"111111111",
  17354=>"111001000",
  17355=>"111100000",
  17356=>"000000000",
  17357=>"111110000",
  17358=>"111111110",
  17359=>"111011111",
  17360=>"000000010",
  17361=>"111111111",
  17362=>"111111111",
  17363=>"110111111",
  17364=>"111110110",
  17365=>"000000000",
  17366=>"001000110",
  17367=>"111111111",
  17368=>"000000000",
  17369=>"000110111",
  17370=>"000000000",
  17371=>"000001111",
  17372=>"000001111",
  17373=>"110000000",
  17374=>"000000001",
  17375=>"111110001",
  17376=>"110110000",
  17377=>"111000000",
  17378=>"000000000",
  17379=>"000000000",
  17380=>"000110110",
  17381=>"110100000",
  17382=>"111111100",
  17383=>"101111111",
  17384=>"111111111",
  17385=>"000000001",
  17386=>"000000000",
  17387=>"000000000",
  17388=>"101111111",
  17389=>"001000000",
  17390=>"000000110",
  17391=>"111111111",
  17392=>"011111000",
  17393=>"000000000",
  17394=>"101001000",
  17395=>"000000000",
  17396=>"111111111",
  17397=>"100111110",
  17398=>"000000000",
  17399=>"111110110",
  17400=>"111111111",
  17401=>"100110000",
  17402=>"000000000",
  17403=>"111110110",
  17404=>"111111111",
  17405=>"111111111",
  17406=>"110100111",
  17407=>"001000000",
  17408=>"100001011",
  17409=>"111111000",
  17410=>"101000111",
  17411=>"000011011",
  17412=>"000001001",
  17413=>"000110010",
  17414=>"110110110",
  17415=>"111111111",
  17416=>"000001011",
  17417=>"000010000",
  17418=>"111111001",
  17419=>"000110111",
  17420=>"111111110",
  17421=>"001000000",
  17422=>"101100000",
  17423=>"111111110",
  17424=>"101000100",
  17425=>"000111111",
  17426=>"010111111",
  17427=>"000000001",
  17428=>"000000011",
  17429=>"000000111",
  17430=>"111011010",
  17431=>"000000000",
  17432=>"110110111",
  17433=>"110001000",
  17434=>"000000000",
  17435=>"110110111",
  17436=>"000000000",
  17437=>"001111111",
  17438=>"001001001",
  17439=>"000001111",
  17440=>"001111100",
  17441=>"000111001",
  17442=>"111110000",
  17443=>"111110000",
  17444=>"110011010",
  17445=>"100000101",
  17446=>"010000000",
  17447=>"010111011",
  17448=>"001000111",
  17449=>"101000000",
  17450=>"111101111",
  17451=>"111000001",
  17452=>"000100111",
  17453=>"011011000",
  17454=>"000000000",
  17455=>"111111111",
  17456=>"110111111",
  17457=>"000011111",
  17458=>"100111111",
  17459=>"000000000",
  17460=>"010000000",
  17461=>"111111111",
  17462=>"111000000",
  17463=>"011000000",
  17464=>"111100000",
  17465=>"011101110",
  17466=>"100100000",
  17467=>"111111111",
  17468=>"000000000",
  17469=>"111111111",
  17470=>"111111111",
  17471=>"110000000",
  17472=>"000100100",
  17473=>"100000100",
  17474=>"000000001",
  17475=>"000000100",
  17476=>"101101000",
  17477=>"000010110",
  17478=>"000000100",
  17479=>"000000000",
  17480=>"100100000",
  17481=>"000000111",
  17482=>"000000000",
  17483=>"000000000",
  17484=>"111111100",
  17485=>"111111111",
  17486=>"111111111",
  17487=>"111111111",
  17488=>"111111111",
  17489=>"111111011",
  17490=>"111111111",
  17491=>"001001001",
  17492=>"000000000",
  17493=>"000100100",
  17494=>"110000001",
  17495=>"000000000",
  17496=>"000000101",
  17497=>"101100100",
  17498=>"000010111",
  17499=>"110010000",
  17500=>"111111111",
  17501=>"111111100",
  17502=>"000000000",
  17503=>"111000000",
  17504=>"000000000",
  17505=>"110110010",
  17506=>"000000000",
  17507=>"011001001",
  17508=>"001111000",
  17509=>"101001111",
  17510=>"110111111",
  17511=>"000000000",
  17512=>"000111111",
  17513=>"001001011",
  17514=>"011101111",
  17515=>"000100111",
  17516=>"111000011",
  17517=>"111111010",
  17518=>"000001111",
  17519=>"000000111",
  17520=>"100100000",
  17521=>"000000000",
  17522=>"001001001",
  17523=>"111111111",
  17524=>"000000000",
  17525=>"111111111",
  17526=>"001001000",
  17527=>"000110111",
  17528=>"000000101",
  17529=>"110111111",
  17530=>"000000000",
  17531=>"100000000",
  17532=>"100100000",
  17533=>"110110010",
  17534=>"000000000",
  17535=>"111111011",
  17536=>"000000000",
  17537=>"110111010",
  17538=>"111111111",
  17539=>"000100001",
  17540=>"110100100",
  17541=>"001000000",
  17542=>"110111000",
  17543=>"111011011",
  17544=>"000011111",
  17545=>"000000100",
  17546=>"100000000",
  17547=>"000000111",
  17548=>"000000100",
  17549=>"100000000",
  17550=>"001101001",
  17551=>"110111110",
  17552=>"000100111",
  17553=>"000000001",
  17554=>"100110100",
  17555=>"110111111",
  17556=>"000000000",
  17557=>"000100100",
  17558=>"001000000",
  17559=>"111111000",
  17560=>"000000000",
  17561=>"111111000",
  17562=>"010001000",
  17563=>"000000100",
  17564=>"001101111",
  17565=>"111100000",
  17566=>"111111111",
  17567=>"000000100",
  17568=>"000101101",
  17569=>"101000000",
  17570=>"111100100",
  17571=>"111000100",
  17572=>"111111111",
  17573=>"111111111",
  17574=>"000000101",
  17575=>"000011001",
  17576=>"000000000",
  17577=>"000100110",
  17578=>"000000000",
  17579=>"000001000",
  17580=>"111001101",
  17581=>"100001000",
  17582=>"111111010",
  17583=>"000000000",
  17584=>"000000111",
  17585=>"101110110",
  17586=>"010111111",
  17587=>"000111111",
  17588=>"111001000",
  17589=>"111111010",
  17590=>"110111111",
  17591=>"000000101",
  17592=>"111011001",
  17593=>"001011011",
  17594=>"001000111",
  17595=>"111111111",
  17596=>"000000000",
  17597=>"000000000",
  17598=>"000111101",
  17599=>"101001000",
  17600=>"000000001",
  17601=>"111000000",
  17602=>"111111001",
  17603=>"001001000",
  17604=>"110111111",
  17605=>"111001001",
  17606=>"000100001",
  17607=>"000000000",
  17608=>"000111111",
  17609=>"110000000",
  17610=>"000000000",
  17611=>"111111111",
  17612=>"100100000",
  17613=>"000000000",
  17614=>"111111111",
  17615=>"110111111",
  17616=>"111101101",
  17617=>"000110000",
  17618=>"100000000",
  17619=>"001000000",
  17620=>"111100111",
  17621=>"100000000",
  17622=>"000000000",
  17623=>"111111001",
  17624=>"111111010",
  17625=>"111111011",
  17626=>"111111011",
  17627=>"001000000",
  17628=>"110000000",
  17629=>"000000000",
  17630=>"000000000",
  17631=>"111001111",
  17632=>"111111111",
  17633=>"000000000",
  17634=>"000000000",
  17635=>"111111110",
  17636=>"000000000",
  17637=>"011110011",
  17638=>"000010010",
  17639=>"001000000",
  17640=>"000000000",
  17641=>"001000000",
  17642=>"000000000",
  17643=>"011001111",
  17644=>"111111111",
  17645=>"000000000",
  17646=>"001000100",
  17647=>"000000100",
  17648=>"000000000",
  17649=>"011010111",
  17650=>"111111010",
  17651=>"111001001",
  17652=>"000000101",
  17653=>"110110000",
  17654=>"000100100",
  17655=>"000000000",
  17656=>"001111111",
  17657=>"000000000",
  17658=>"111111000",
  17659=>"001101100",
  17660=>"000100111",
  17661=>"000100000",
  17662=>"111010111",
  17663=>"111111111",
  17664=>"111000000",
  17665=>"001001111",
  17666=>"000000000",
  17667=>"001000111",
  17668=>"001000000",
  17669=>"101101100",
  17670=>"100000000",
  17671=>"000000101",
  17672=>"101000000",
  17673=>"111111000",
  17674=>"000000000",
  17675=>"100000000",
  17676=>"101101111",
  17677=>"100100111",
  17678=>"000101111",
  17679=>"010000000",
  17680=>"000000000",
  17681=>"110111110",
  17682=>"110111111",
  17683=>"000110110",
  17684=>"000000000",
  17685=>"111111111",
  17686=>"110110010",
  17687=>"111111100",
  17688=>"111111111",
  17689=>"111111000",
  17690=>"000000000",
  17691=>"010010010",
  17692=>"000001110",
  17693=>"000000000",
  17694=>"000000000",
  17695=>"110100111",
  17696=>"111111110",
  17697=>"111111000",
  17698=>"111111101",
  17699=>"111111110",
  17700=>"100110110",
  17701=>"010011111",
  17702=>"111010000",
  17703=>"000100111",
  17704=>"111111111",
  17705=>"000111111",
  17706=>"111111000",
  17707=>"000000000",
  17708=>"000000100",
  17709=>"111111000",
  17710=>"111111111",
  17711=>"000000000",
  17712=>"101111110",
  17713=>"100000000",
  17714=>"111111111",
  17715=>"000000000",
  17716=>"111000001",
  17717=>"110111000",
  17718=>"001001000",
  17719=>"000000000",
  17720=>"111111111",
  17721=>"000000110",
  17722=>"011000000",
  17723=>"111111011",
  17724=>"000000000",
  17725=>"100100010",
  17726=>"001001001",
  17727=>"111111111",
  17728=>"111000100",
  17729=>"111111111",
  17730=>"111111110",
  17731=>"001001001",
  17732=>"000000000",
  17733=>"000000000",
  17734=>"000100100",
  17735=>"000000000",
  17736=>"000000001",
  17737=>"010111111",
  17738=>"111111000",
  17739=>"000010000",
  17740=>"000000000",
  17741=>"000010010",
  17742=>"000000100",
  17743=>"110110010",
  17744=>"100110110",
  17745=>"000100100",
  17746=>"000000000",
  17747=>"000000000",
  17748=>"000000011",
  17749=>"011011001",
  17750=>"111111110",
  17751=>"100100100",
  17752=>"000001000",
  17753=>"011011111",
  17754=>"111001000",
  17755=>"111011000",
  17756=>"000000001",
  17757=>"000010010",
  17758=>"111110000",
  17759=>"000110000",
  17760=>"111001000",
  17761=>"000000001",
  17762=>"100110110",
  17763=>"000000101",
  17764=>"111111000",
  17765=>"000000000",
  17766=>"111111111",
  17767=>"111111111",
  17768=>"000000001",
  17769=>"111111000",
  17770=>"001011111",
  17771=>"111110000",
  17772=>"111111000",
  17773=>"000000100",
  17774=>"000110000",
  17775=>"111100100",
  17776=>"110000111",
  17777=>"110111110",
  17778=>"011111111",
  17779=>"111111000",
  17780=>"110000000",
  17781=>"100000000",
  17782=>"110100101",
  17783=>"111111111",
  17784=>"101000101",
  17785=>"000000111",
  17786=>"000000111",
  17787=>"111000000",
  17788=>"001111111",
  17789=>"111111111",
  17790=>"000000000",
  17791=>"000000000",
  17792=>"000000100",
  17793=>"000100000",
  17794=>"000111111",
  17795=>"000000000",
  17796=>"000011111",
  17797=>"001001000",
  17798=>"000000111",
  17799=>"110110100",
  17800=>"111111111",
  17801=>"000000000",
  17802=>"001000000",
  17803=>"111111111",
  17804=>"111111111",
  17805=>"111110001",
  17806=>"111111111",
  17807=>"111011011",
  17808=>"000000000",
  17809=>"111111011",
  17810=>"000100101",
  17811=>"011000101",
  17812=>"111111111",
  17813=>"000000000",
  17814=>"110110110",
  17815=>"111111010",
  17816=>"001011001",
  17817=>"110110110",
  17818=>"000000000",
  17819=>"000000101",
  17820=>"000000001",
  17821=>"011001111",
  17822=>"001001101",
  17823=>"000110011",
  17824=>"111111010",
  17825=>"011111000",
  17826=>"011001000",
  17827=>"111111011",
  17828=>"011001111",
  17829=>"011001011",
  17830=>"100100111",
  17831=>"001000000",
  17832=>"000000000",
  17833=>"001000000",
  17834=>"111111111",
  17835=>"011011000",
  17836=>"000000000",
  17837=>"000000000",
  17838=>"111001111",
  17839=>"000000100",
  17840=>"000001111",
  17841=>"011111000",
  17842=>"111001000",
  17843=>"000000000",
  17844=>"001111001",
  17845=>"000000000",
  17846=>"110111111",
  17847=>"101111000",
  17848=>"111111111",
  17849=>"011010000",
  17850=>"000000000",
  17851=>"000100100",
  17852=>"000000000",
  17853=>"100110111",
  17854=>"011011000",
  17855=>"000001000",
  17856=>"001001000",
  17857=>"001101110",
  17858=>"101001111",
  17859=>"000010000",
  17860=>"001001000",
  17861=>"001001001",
  17862=>"001000101",
  17863=>"001001001",
  17864=>"111000000",
  17865=>"100100111",
  17866=>"111110100",
  17867=>"000000000",
  17868=>"000011000",
  17869=>"111111111",
  17870=>"000000000",
  17871=>"000000000",
  17872=>"001001011",
  17873=>"010111111",
  17874=>"011111001",
  17875=>"000000000",
  17876=>"001001001",
  17877=>"100111111",
  17878=>"000000111",
  17879=>"011011001",
  17880=>"000000111",
  17881=>"000000111",
  17882=>"000011011",
  17883=>"011000000",
  17884=>"000000000",
  17885=>"001011111",
  17886=>"111111011",
  17887=>"000100100",
  17888=>"001001001",
  17889=>"111000000",
  17890=>"000000111",
  17891=>"000000000",
  17892=>"111111110",
  17893=>"011111111",
  17894=>"011011000",
  17895=>"111000000",
  17896=>"110110100",
  17897=>"000000000",
  17898=>"100000000",
  17899=>"000000000",
  17900=>"000000101",
  17901=>"110110010",
  17902=>"001001001",
  17903=>"110100000",
  17904=>"101101100",
  17905=>"010111111",
  17906=>"111111111",
  17907=>"001000000",
  17908=>"111111000",
  17909=>"000000000",
  17910=>"000000000",
  17911=>"110110000",
  17912=>"000100111",
  17913=>"011011000",
  17914=>"000000000",
  17915=>"111101101",
  17916=>"001000001",
  17917=>"110100110",
  17918=>"000000100",
  17919=>"000000001",
  17920=>"110110010",
  17921=>"111111001",
  17922=>"000000101",
  17923=>"000000111",
  17924=>"111111011",
  17925=>"000001001",
  17926=>"110110111",
  17927=>"001111110",
  17928=>"111001111",
  17929=>"000000000",
  17930=>"111111111",
  17931=>"111110110",
  17932=>"100110111",
  17933=>"001001101",
  17934=>"000100000",
  17935=>"000000010",
  17936=>"001001111",
  17937=>"011111111",
  17938=>"111001001",
  17939=>"001000000",
  17940=>"001000001",
  17941=>"000000000",
  17942=>"000000101",
  17943=>"001100100",
  17944=>"000000100",
  17945=>"000100001",
  17946=>"000000000",
  17947=>"111111111",
  17948=>"000000000",
  17949=>"000000110",
  17950=>"111101000",
  17951=>"000000110",
  17952=>"101001000",
  17953=>"000000000",
  17954=>"110110010",
  17955=>"111111010",
  17956=>"111010000",
  17957=>"000000101",
  17958=>"111110110",
  17959=>"000010011",
  17960=>"111101000",
  17961=>"000000101",
  17962=>"100100000",
  17963=>"000000111",
  17964=>"001000000",
  17965=>"111011000",
  17966=>"001001011",
  17967=>"111110111",
  17968=>"110000111",
  17969=>"111011000",
  17970=>"000000000",
  17971=>"111111000",
  17972=>"000000000",
  17973=>"000100000",
  17974=>"111101100",
  17975=>"000000100",
  17976=>"010111010",
  17977=>"000111111",
  17978=>"001111111",
  17979=>"111110110",
  17980=>"000000000",
  17981=>"001000000",
  17982=>"001100000",
  17983=>"000101111",
  17984=>"000000000",
  17985=>"000010010",
  17986=>"000000111",
  17987=>"000000100",
  17988=>"000000010",
  17989=>"000000000",
  17990=>"111110110",
  17991=>"111001000",
  17992=>"000100111",
  17993=>"111111111",
  17994=>"101100111",
  17995=>"110111111",
  17996=>"110110000",
  17997=>"111111000",
  17998=>"000000000",
  17999=>"001001001",
  18000=>"111111011",
  18001=>"111001100",
  18002=>"110111000",
  18003=>"100100000",
  18004=>"110000000",
  18005=>"001000010",
  18006=>"000000010",
  18007=>"000001111",
  18008=>"110110000",
  18009=>"111111111",
  18010=>"000000000",
  18011=>"010010010",
  18012=>"100000000",
  18013=>"000000100",
  18014=>"010010000",
  18015=>"110110111",
  18016=>"111111110",
  18017=>"000000000",
  18018=>"110110000",
  18019=>"111100100",
  18020=>"000000000",
  18021=>"000000000",
  18022=>"000000000",
  18023=>"000101111",
  18024=>"111111001",
  18025=>"000000111",
  18026=>"111001011",
  18027=>"111100110",
  18028=>"000110110",
  18029=>"000000000",
  18030=>"110110000",
  18031=>"111001101",
  18032=>"111100111",
  18033=>"000000000",
  18034=>"000000011",
  18035=>"101111010",
  18036=>"011001001",
  18037=>"111110111",
  18038=>"000000000",
  18039=>"111011000",
  18040=>"000000110",
  18041=>"111111111",
  18042=>"001000001",
  18043=>"010010000",
  18044=>"110110100",
  18045=>"001010000",
  18046=>"001000100",
  18047=>"000000000",
  18048=>"000000000",
  18049=>"000111110",
  18050=>"111000100",
  18051=>"001010010",
  18052=>"000100111",
  18053=>"000000011",
  18054=>"000100100",
  18055=>"110111111",
  18056=>"011001100",
  18057=>"111111111",
  18058=>"111111000",
  18059=>"001000110",
  18060=>"111111110",
  18061=>"000000010",
  18062=>"101000101",
  18063=>"000000000",
  18064=>"001000101",
  18065=>"000000000",
  18066=>"000001011",
  18067=>"110111100",
  18068=>"001001101",
  18069=>"110000000",
  18070=>"101111111",
  18071=>"001001111",
  18072=>"001001111",
  18073=>"100000111",
  18074=>"000000111",
  18075=>"110110000",
  18076=>"001000000",
  18077=>"000000000",
  18078=>"001111100",
  18079=>"111111111",
  18080=>"111111111",
  18081=>"000111011",
  18082=>"110100101",
  18083=>"000000000",
  18084=>"110111110",
  18085=>"000110110",
  18086=>"011001001",
  18087=>"000011001",
  18088=>"000100011",
  18089=>"101001001",
  18090=>"111010011",
  18091=>"000100111",
  18092=>"000000000",
  18093=>"110110100",
  18094=>"000000000",
  18095=>"111100111",
  18096=>"110111000",
  18097=>"000001010",
  18098=>"111111010",
  18099=>"111111111",
  18100=>"000000000",
  18101=>"000001111",
  18102=>"001001011",
  18103=>"111111111",
  18104=>"111001001",
  18105=>"111111111",
  18106=>"111001001",
  18107=>"000000000",
  18108=>"010000000",
  18109=>"111000001",
  18110=>"101101111",
  18111=>"111110110",
  18112=>"111111011",
  18113=>"111111011",
  18114=>"111101000",
  18115=>"000100101",
  18116=>"001101111",
  18117=>"101111111",
  18118=>"000000000",
  18119=>"111111000",
  18120=>"000100000",
  18121=>"110111001",
  18122=>"111111010",
  18123=>"000000000",
  18124=>"111111111",
  18125=>"000111001",
  18126=>"001000000",
  18127=>"000000000",
  18128=>"000000011",
  18129=>"001001111",
  18130=>"000000000",
  18131=>"000000000",
  18132=>"000000000",
  18133=>"111111000",
  18134=>"111100000",
  18135=>"011110000",
  18136=>"111111111",
  18137=>"000001001",
  18138=>"000000000",
  18139=>"110000000",
  18140=>"111111111",
  18141=>"011111111",
  18142=>"111101000",
  18143=>"010110010",
  18144=>"010110000",
  18145=>"000010000",
  18146=>"000110111",
  18147=>"000000000",
  18148=>"110100000",
  18149=>"010110110",
  18150=>"010010010",
  18151=>"100110000",
  18152=>"111110111",
  18153=>"100000000",
  18154=>"000000000",
  18155=>"111011111",
  18156=>"101110111",
  18157=>"111111111",
  18158=>"111111111",
  18159=>"000111100",
  18160=>"110111111",
  18161=>"000000010",
  18162=>"111001000",
  18163=>"000000111",
  18164=>"000000000",
  18165=>"110100101",
  18166=>"000001001",
  18167=>"111111011",
  18168=>"111101000",
  18169=>"110111111",
  18170=>"000000000",
  18171=>"000000100",
  18172=>"000111100",
  18173=>"110110000",
  18174=>"111000111",
  18175=>"111111000",
  18176=>"000000111",
  18177=>"111001011",
  18178=>"000000100",
  18179=>"000000111",
  18180=>"111111000",
  18181=>"000000001",
  18182=>"001111111",
  18183=>"000000010",
  18184=>"110111111",
  18185=>"111001100",
  18186=>"110110010",
  18187=>"010000111",
  18188=>"000000000",
  18189=>"011000010",
  18190=>"000110000",
  18191=>"011011111",
  18192=>"100101111",
  18193=>"000000000",
  18194=>"000000000",
  18195=>"110000000",
  18196=>"111111111",
  18197=>"101000111",
  18198=>"111110110",
  18199=>"110000101",
  18200=>"110100000",
  18201=>"000000000",
  18202=>"000000000",
  18203=>"001000000",
  18204=>"110111110",
  18205=>"000000000",
  18206=>"101111111",
  18207=>"000000000",
  18208=>"111111000",
  18209=>"000000000",
  18210=>"000111000",
  18211=>"001001101",
  18212=>"111111100",
  18213=>"111111111",
  18214=>"010010010",
  18215=>"111000000",
  18216=>"001001111",
  18217=>"000000001",
  18218=>"111110111",
  18219=>"001000111",
  18220=>"000000000",
  18221=>"000000000",
  18222=>"111110111",
  18223=>"111111110",
  18224=>"000000101",
  18225=>"000111110",
  18226=>"001000110",
  18227=>"000000000",
  18228=>"000010010",
  18229=>"111000000",
  18230=>"000000111",
  18231=>"001000000",
  18232=>"111101111",
  18233=>"101101111",
  18234=>"111111111",
  18235=>"000001001",
  18236=>"000000111",
  18237=>"000000100",
  18238=>"110000111",
  18239=>"111111111",
  18240=>"111111111",
  18241=>"000001110",
  18242=>"110110001",
  18243=>"000000111",
  18244=>"111111111",
  18245=>"111101000",
  18246=>"001111101",
  18247=>"010100110",
  18248=>"111000111",
  18249=>"010011111",
  18250=>"111110100",
  18251=>"000110100",
  18252=>"000000101",
  18253=>"111111111",
  18254=>"000000000",
  18255=>"001011111",
  18256=>"000010110",
  18257=>"001101111",
  18258=>"111111111",
  18259=>"001001111",
  18260=>"101000101",
  18261=>"011011000",
  18262=>"000000000",
  18263=>"000000111",
  18264=>"000000000",
  18265=>"000000000",
  18266=>"111100000",
  18267=>"101000100",
  18268=>"110110110",
  18269=>"100001000",
  18270=>"111111110",
  18271=>"011010110",
  18272=>"101001101",
  18273=>"000000000",
  18274=>"000110011",
  18275=>"000111111",
  18276=>"111001000",
  18277=>"101001000",
  18278=>"000100111",
  18279=>"000100110",
  18280=>"001001111",
  18281=>"000111111",
  18282=>"000000010",
  18283=>"010110111",
  18284=>"110110110",
  18285=>"000001101",
  18286=>"001111111",
  18287=>"000000000",
  18288=>"000000110",
  18289=>"111111001",
  18290=>"100111110",
  18291=>"110110000",
  18292=>"010010010",
  18293=>"000000000",
  18294=>"011000000",
  18295=>"000000000",
  18296=>"001001111",
  18297=>"111110100",
  18298=>"001111111",
  18299=>"110111111",
  18300=>"000000000",
  18301=>"001000001",
  18302=>"100000000",
  18303=>"000110111",
  18304=>"110110100",
  18305=>"001000111",
  18306=>"001000000",
  18307=>"101000000",
  18308=>"000000110",
  18309=>"010000011",
  18310=>"111111111",
  18311=>"111111111",
  18312=>"111110000",
  18313=>"000000000",
  18314=>"010000000",
  18315=>"111000000",
  18316=>"111111111",
  18317=>"111111011",
  18318=>"111111111",
  18319=>"111110100",
  18320=>"111111111",
  18321=>"000100110",
  18322=>"000000000",
  18323=>"000000111",
  18324=>"110010010",
  18325=>"000001010",
  18326=>"100000101",
  18327=>"100000000",
  18328=>"110010111",
  18329=>"111110000",
  18330=>"000000001",
  18331=>"110110011",
  18332=>"000010110",
  18333=>"000000000",
  18334=>"111001001",
  18335=>"000001111",
  18336=>"000000000",
  18337=>"000110110",
  18338=>"000000000",
  18339=>"111111111",
  18340=>"000001111",
  18341=>"111111111",
  18342=>"111000000",
  18343=>"000001001",
  18344=>"101111110",
  18345=>"000000001",
  18346=>"111111001",
  18347=>"000000000",
  18348=>"111001000",
  18349=>"001100111",
  18350=>"101111111",
  18351=>"001011000",
  18352=>"111111100",
  18353=>"001001011",
  18354=>"110110000",
  18355=>"111101111",
  18356=>"000001000",
  18357=>"000000000",
  18358=>"001000111",
  18359=>"000000111",
  18360=>"010010111",
  18361=>"010001011",
  18362=>"001101000",
  18363=>"001000000",
  18364=>"000111011",
  18365=>"000000000",
  18366=>"111011000",
  18367=>"110111111",
  18368=>"111111000",
  18369=>"100111111",
  18370=>"111111111",
  18371=>"101101111",
  18372=>"000000010",
  18373=>"100100110",
  18374=>"000000001",
  18375=>"110000000",
  18376=>"111000000",
  18377=>"000000001",
  18378=>"000000010",
  18379=>"000000111",
  18380=>"110010010",
  18381=>"001111111",
  18382=>"111110111",
  18383=>"001111111",
  18384=>"010111111",
  18385=>"001001111",
  18386=>"000000000",
  18387=>"111001111",
  18388=>"011001001",
  18389=>"111000100",
  18390=>"000000000",
  18391=>"111111111",
  18392=>"110110000",
  18393=>"111011000",
  18394=>"000000000",
  18395=>"000000000",
  18396=>"111001101",
  18397=>"101000111",
  18398=>"111110010",
  18399=>"100000000",
  18400=>"111110110",
  18401=>"001011000",
  18402=>"111111111",
  18403=>"000000011",
  18404=>"111111111",
  18405=>"111111111",
  18406=>"000000000",
  18407=>"001001101",
  18408=>"111101111",
  18409=>"000000000",
  18410=>"011111111",
  18411=>"010110000",
  18412=>"001011000",
  18413=>"011111111",
  18414=>"100110000",
  18415=>"011011111",
  18416=>"000001111",
  18417=>"111110110",
  18418=>"001011111",
  18419=>"000000000",
  18420=>"001000000",
  18421=>"000000110",
  18422=>"111111111",
  18423=>"000010010",
  18424=>"111111111",
  18425=>"011111111",
  18426=>"111111111",
  18427=>"000000001",
  18428=>"111110001",
  18429=>"110110110",
  18430=>"111110110",
  18431=>"011001111",
  18432=>"011010110",
  18433=>"000000000",
  18434=>"101001000",
  18435=>"110100111",
  18436=>"001111111",
  18437=>"111011011",
  18438=>"111101111",
  18439=>"001011111",
  18440=>"001111111",
  18441=>"111111000",
  18442=>"111111101",
  18443=>"000000000",
  18444=>"000001000",
  18445=>"000010010",
  18446=>"111111111",
  18447=>"111111111",
  18448=>"111111111",
  18449=>"111111011",
  18450=>"000000000",
  18451=>"000110110",
  18452=>"111111111",
  18453=>"111111111",
  18454=>"000000000",
  18455=>"011111111",
  18456=>"000000110",
  18457=>"011111111",
  18458=>"111001111",
  18459=>"111001001",
  18460=>"000000000",
  18461=>"000000000",
  18462=>"000000010",
  18463=>"000000000",
  18464=>"010010111",
  18465=>"000000000",
  18466=>"100101001",
  18467=>"001001101",
  18468=>"111111111",
  18469=>"000100111",
  18470=>"000000000",
  18471=>"110100001",
  18472=>"111111111",
  18473=>"111111111",
  18474=>"001000000",
  18475=>"111111111",
  18476=>"000000001",
  18477=>"111111111",
  18478=>"000001100",
  18479=>"111111110",
  18480=>"000000000",
  18481=>"001000000",
  18482=>"110010010",
  18483=>"110000000",
  18484=>"111111111",
  18485=>"000011011",
  18486=>"010001000",
  18487=>"111111111",
  18488=>"000100000",
  18489=>"000010000",
  18490=>"100000000",
  18491=>"111111111",
  18492=>"001000000",
  18493=>"100000111",
  18494=>"111111011",
  18495=>"111101001",
  18496=>"000000000",
  18497=>"011000100",
  18498=>"101001001",
  18499=>"111111101",
  18500=>"011111111",
  18501=>"000000110",
  18502=>"111111110",
  18503=>"111111111",
  18504=>"000000000",
  18505=>"000000001",
  18506=>"100000100",
  18507=>"011000111",
  18508=>"000100111",
  18509=>"000000000",
  18510=>"111111111",
  18511=>"111101001",
  18512=>"100100111",
  18513=>"000000000",
  18514=>"001001000",
  18515=>"111001001",
  18516=>"000000000",
  18517=>"111111110",
  18518=>"000001110",
  18519=>"111111111",
  18520=>"000000100",
  18521=>"000000000",
  18522=>"010111111",
  18523=>"001001001",
  18524=>"000000000",
  18525=>"000000000",
  18526=>"100100000",
  18527=>"000000000",
  18528=>"000000000",
  18529=>"111111111",
  18530=>"100110110",
  18531=>"111000000",
  18532=>"000000010",
  18533=>"000000000",
  18534=>"110111111",
  18535=>"000110000",
  18536=>"000000111",
  18537=>"001000000",
  18538=>"111111111",
  18539=>"110010000",
  18540=>"101111111",
  18541=>"000000000",
  18542=>"000000000",
  18543=>"000000000",
  18544=>"000000000",
  18545=>"000000001",
  18546=>"011001001",
  18547=>"000000000",
  18548=>"111111100",
  18549=>"001001111",
  18550=>"111111010",
  18551=>"100101001",
  18552=>"001001001",
  18553=>"000000000",
  18554=>"001001011",
  18555=>"000000000",
  18556=>"000111111",
  18557=>"000000001",
  18558=>"000000000",
  18559=>"111000000",
  18560=>"111001000",
  18561=>"010110111",
  18562=>"000000000",
  18563=>"000000000",
  18564=>"110100000",
  18565=>"000000000",
  18566=>"000000000",
  18567=>"110000011",
  18568=>"110110100",
  18569=>"000000000",
  18570=>"111101111",
  18571=>"111000000",
  18572=>"110000000",
  18573=>"000000000",
  18574=>"111000011",
  18575=>"000000110",
  18576=>"000000111",
  18577=>"000001011",
  18578=>"110111110",
  18579=>"111111111",
  18580=>"010111000",
  18581=>"000110000",
  18582=>"000000000",
  18583=>"000000100",
  18584=>"111111111",
  18585=>"111111001",
  18586=>"111010000",
  18587=>"111111111",
  18588=>"111111111",
  18589=>"001101110",
  18590=>"000011011",
  18591=>"000000000",
  18592=>"011000000",
  18593=>"100110111",
  18594=>"000001000",
  18595=>"001111010",
  18596=>"111111111",
  18597=>"111111111",
  18598=>"111111111",
  18599=>"001001011",
  18600=>"000000000",
  18601=>"001001001",
  18602=>"000000000",
  18603=>"111111111",
  18604=>"000001100",
  18605=>"000000001",
  18606=>"000000000",
  18607=>"000000100",
  18608=>"000111111",
  18609=>"000000000",
  18610=>"100110110",
  18611=>"000101010",
  18612=>"111101000",
  18613=>"000000000",
  18614=>"000000000",
  18615=>"100100000",
  18616=>"100101111",
  18617=>"000000111",
  18618=>"100101101",
  18619=>"111111111",
  18620=>"111000000",
  18621=>"000111111",
  18622=>"111111000",
  18623=>"010000010",
  18624=>"111111111",
  18625=>"111111111",
  18626=>"000011111",
  18627=>"001001111",
  18628=>"111111111",
  18629=>"000000111",
  18630=>"000000101",
  18631=>"100101101",
  18632=>"000000000",
  18633=>"111111101",
  18634=>"110111101",
  18635=>"100000000",
  18636=>"101101001",
  18637=>"111111111",
  18638=>"111101000",
  18639=>"000111111",
  18640=>"111010001",
  18641=>"000000000",
  18642=>"000000000",
  18643=>"000000000",
  18644=>"100000000",
  18645=>"111111111",
  18646=>"011111111",
  18647=>"000000000",
  18648=>"111111000",
  18649=>"000000000",
  18650=>"110000000",
  18651=>"000000000",
  18652=>"010001111",
  18653=>"000111110",
  18654=>"111111000",
  18655=>"000000001",
  18656=>"000000000",
  18657=>"111111111",
  18658=>"000000000",
  18659=>"000000000",
  18660=>"111111011",
  18661=>"100110111",
  18662=>"111111111",
  18663=>"011111111",
  18664=>"111111111",
  18665=>"000000000",
  18666=>"101101111",
  18667=>"111111111",
  18668=>"000000000",
  18669=>"111111111",
  18670=>"111111000",
  18671=>"000000011",
  18672=>"111111000",
  18673=>"111111011",
  18674=>"111111111",
  18675=>"001001111",
  18676=>"100000000",
  18677=>"000000000",
  18678=>"101001000",
  18679=>"000000000",
  18680=>"111111110",
  18681=>"000001001",
  18682=>"011001111",
  18683=>"001001000",
  18684=>"000000000",
  18685=>"001001000",
  18686=>"000001111",
  18687=>"000110010",
  18688=>"111111111",
  18689=>"000010110",
  18690=>"000000000",
  18691=>"111110000",
  18692=>"110100000",
  18693=>"110100111",
  18694=>"111101101",
  18695=>"010100000",
  18696=>"111100110",
  18697=>"000000011",
  18698=>"111111111",
  18699=>"110101000",
  18700=>"000000000",
  18701=>"000100111",
  18702=>"111111110",
  18703=>"000000010",
  18704=>"000000000",
  18705=>"000000000",
  18706=>"111000000",
  18707=>"000000001",
  18708=>"000000000",
  18709=>"111100000",
  18710=>"011001001",
  18711=>"001001101",
  18712=>"001000110",
  18713=>"110111111",
  18714=>"110110110",
  18715=>"111111111",
  18716=>"001001011",
  18717=>"001001111",
  18718=>"110110100",
  18719=>"111111111",
  18720=>"000000011",
  18721=>"010111000",
  18722=>"011111111",
  18723=>"111111111",
  18724=>"000000000",
  18725=>"000000010",
  18726=>"111111111",
  18727=>"111101100",
  18728=>"000100110",
  18729=>"000000000",
  18730=>"110000000",
  18731=>"000000000",
  18732=>"000000000",
  18733=>"110000000",
  18734=>"000000000",
  18735=>"000000000",
  18736=>"000100011",
  18737=>"000100110",
  18738=>"011011011",
  18739=>"111111111",
  18740=>"000110000",
  18741=>"000000000",
  18742=>"010001111",
  18743=>"001001101",
  18744=>"010000000",
  18745=>"000000111",
  18746=>"000000110",
  18747=>"000000000",
  18748=>"111111110",
  18749=>"111101000",
  18750=>"000100111",
  18751=>"111011001",
  18752=>"001000000",
  18753=>"000000111",
  18754=>"111111111",
  18755=>"000000000",
  18756=>"000000000",
  18757=>"000000000",
  18758=>"111111001",
  18759=>"111111000",
  18760=>"000000000",
  18761=>"111111100",
  18762=>"110110110",
  18763=>"010011001",
  18764=>"110000000",
  18765=>"011001000",
  18766=>"111111111",
  18767=>"111111111",
  18768=>"000000000",
  18769=>"000000000",
  18770=>"111000000",
  18771=>"111111000",
  18772=>"000000000",
  18773=>"111111011",
  18774=>"001001000",
  18775=>"000000000",
  18776=>"111111111",
  18777=>"000001000",
  18778=>"111111111",
  18779=>"001000000",
  18780=>"111001000",
  18781=>"110000000",
  18782=>"000000000",
  18783=>"000000001",
  18784=>"010111111",
  18785=>"000011011",
  18786=>"000000000",
  18787=>"000000000",
  18788=>"000000000",
  18789=>"000000000",
  18790=>"111111111",
  18791=>"111011010",
  18792=>"000000000",
  18793=>"111011111",
  18794=>"011000000",
  18795=>"110111101",
  18796=>"000000000",
  18797=>"000100001",
  18798=>"010000000",
  18799=>"000100111",
  18800=>"011011010",
  18801=>"000000000",
  18802=>"110111111",
  18803=>"110111111",
  18804=>"100000010",
  18805=>"000001101",
  18806=>"000000001",
  18807=>"011000011",
  18808=>"000000000",
  18809=>"000011011",
  18810=>"111111111",
  18811=>"001000100",
  18812=>"000000100",
  18813=>"011001000",
  18814=>"000011010",
  18815=>"000000000",
  18816=>"000000000",
  18817=>"111001101",
  18818=>"011111001",
  18819=>"000000000",
  18820=>"001101100",
  18821=>"001000000",
  18822=>"111111111",
  18823=>"010000000",
  18824=>"010011111",
  18825=>"100100000",
  18826=>"111011111",
  18827=>"100101100",
  18828=>"111111111",
  18829=>"010010010",
  18830=>"000000000",
  18831=>"000000000",
  18832=>"000000010",
  18833=>"000000000",
  18834=>"011111111",
  18835=>"111111111",
  18836=>"000000000",
  18837=>"000010011",
  18838=>"100000000",
  18839=>"000000000",
  18840=>"001000000",
  18841=>"111111111",
  18842=>"111001100",
  18843=>"101111111",
  18844=>"001011011",
  18845=>"011111011",
  18846=>"101101111",
  18847=>"000000000",
  18848=>"000000000",
  18849=>"011111010",
  18850=>"001001111",
  18851=>"111111111",
  18852=>"110111000",
  18853=>"101001000",
  18854=>"101101111",
  18855=>"011011000",
  18856=>"000000000",
  18857=>"000000111",
  18858=>"111111111",
  18859=>"000100101",
  18860=>"111111111",
  18861=>"000000000",
  18862=>"000111000",
  18863=>"101111111",
  18864=>"100000000",
  18865=>"000000000",
  18866=>"011110110",
  18867=>"000000000",
  18868=>"110101111",
  18869=>"011001000",
  18870=>"111111011",
  18871=>"000000000",
  18872=>"000000000",
  18873=>"111111011",
  18874=>"000000110",
  18875=>"000000111",
  18876=>"000000000",
  18877=>"111111110",
  18878=>"101101101",
  18879=>"001011000",
  18880=>"100111111",
  18881=>"001000000",
  18882=>"100001001",
  18883=>"000000000",
  18884=>"000000000",
  18885=>"111111001",
  18886=>"000001100",
  18887=>"111011001",
  18888=>"000000000",
  18889=>"101000000",
  18890=>"000010111",
  18891=>"100100100",
  18892=>"101000101",
  18893=>"000000000",
  18894=>"110110000",
  18895=>"111111111",
  18896=>"000000000",
  18897=>"100100000",
  18898=>"111111010",
  18899=>"111001000",
  18900=>"011011000",
  18901=>"000000000",
  18902=>"000001111",
  18903=>"000000100",
  18904=>"000110111",
  18905=>"000010011",
  18906=>"101001001",
  18907=>"000001000",
  18908=>"100100011",
  18909=>"011100111",
  18910=>"111111111",
  18911=>"001001000",
  18912=>"010111101",
  18913=>"111110100",
  18914=>"111111111",
  18915=>"111111111",
  18916=>"111111000",
  18917=>"111111111",
  18918=>"111110000",
  18919=>"110110100",
  18920=>"111111111",
  18921=>"100100111",
  18922=>"000000111",
  18923=>"011001011",
  18924=>"111111111",
  18925=>"100100000",
  18926=>"000000000",
  18927=>"000100101",
  18928=>"101101101",
  18929=>"100100000",
  18930=>"101111111",
  18931=>"000011010",
  18932=>"000000000",
  18933=>"110110110",
  18934=>"000000000",
  18935=>"000110100",
  18936=>"101000000",
  18937=>"110110010",
  18938=>"000001000",
  18939=>"111111000",
  18940=>"000000110",
  18941=>"000000000",
  18942=>"000000000",
  18943=>"111001001",
  18944=>"000000100",
  18945=>"111001000",
  18946=>"111000111",
  18947=>"001000000",
  18948=>"110111111",
  18949=>"000000100",
  18950=>"010111010",
  18951=>"111111111",
  18952=>"111111111",
  18953=>"000000111",
  18954=>"000111111",
  18955=>"000000000",
  18956=>"000110110",
  18957=>"000000100",
  18958=>"000000000",
  18959=>"000000000",
  18960=>"111001011",
  18961=>"011010000",
  18962=>"000000000",
  18963=>"000000000",
  18964=>"111100000",
  18965=>"000111111",
  18966=>"111001000",
  18967=>"000001001",
  18968=>"000000000",
  18969=>"001001110",
  18970=>"000010111",
  18971=>"100010011",
  18972=>"000000101",
  18973=>"000000110",
  18974=>"111111111",
  18975=>"010110111",
  18976=>"111111110",
  18977=>"001011001",
  18978=>"110111111",
  18979=>"000000000",
  18980=>"111111111",
  18981=>"101000000",
  18982=>"111111111",
  18983=>"000111111",
  18984=>"110111110",
  18985=>"000100100",
  18986=>"111100100",
  18987=>"111000000",
  18988=>"000000000",
  18989=>"110100100",
  18990=>"101000000",
  18991=>"101000000",
  18992=>"100001001",
  18993=>"010111010",
  18994=>"000011011",
  18995=>"111101000",
  18996=>"101101111",
  18997=>"110010000",
  18998=>"000000000",
  18999=>"100000001",
  19000=>"111111111",
  19001=>"101111110",
  19002=>"111111111",
  19003=>"000000111",
  19004=>"101000101",
  19005=>"000110111",
  19006=>"001111010",
  19007=>"101111101",
  19008=>"001001011",
  19009=>"000100000",
  19010=>"111100001",
  19011=>"111110111",
  19012=>"000110111",
  19013=>"000001000",
  19014=>"111000000",
  19015=>"111001001",
  19016=>"000101001",
  19017=>"011001001",
  19018=>"110111111",
  19019=>"111111111",
  19020=>"000000000",
  19021=>"111101001",
  19022=>"011111111",
  19023=>"111100000",
  19024=>"000011000",
  19025=>"111111111",
  19026=>"110100100",
  19027=>"001000000",
  19028=>"000000001",
  19029=>"111111110",
  19030=>"000000011",
  19031=>"101111010",
  19032=>"001000111",
  19033=>"111111101",
  19034=>"111010000",
  19035=>"100100010",
  19036=>"000010000",
  19037=>"111001101",
  19038=>"000111111",
  19039=>"000000000",
  19040=>"011010000",
  19041=>"111111111",
  19042=>"001000000",
  19043=>"111000001",
  19044=>"111111110",
  19045=>"111000000",
  19046=>"001011000",
  19047=>"001000101",
  19048=>"111111111",
  19049=>"011011000",
  19050=>"111110111",
  19051=>"110111111",
  19052=>"000111011",
  19053=>"111100000",
  19054=>"111000001",
  19055=>"110111111",
  19056=>"000000000",
  19057=>"100101111",
  19058=>"001000000",
  19059=>"100010111",
  19060=>"111001000",
  19061=>"100100100",
  19062=>"000000000",
  19063=>"000000000",
  19064=>"101101111",
  19065=>"101101111",
  19066=>"000001001",
  19067=>"000001111",
  19068=>"100000111",
  19069=>"000000000",
  19070=>"000000000",
  19071=>"000111111",
  19072=>"000000000",
  19073=>"110110000",
  19074=>"111000100",
  19075=>"111111000",
  19076=>"111111111",
  19077=>"010010000",
  19078=>"111101000",
  19079=>"111001000",
  19080=>"001000000",
  19081=>"001000000",
  19082=>"001111111",
  19083=>"000000000",
  19084=>"111111111",
  19085=>"111101001",
  19086=>"000000100",
  19087=>"000000000",
  19088=>"101000000",
  19089=>"000000000",
  19090=>"000011000",
  19091=>"111110110",
  19092=>"111111111",
  19093=>"001111000",
  19094=>"111111111",
  19095=>"111000101",
  19096=>"000000000",
  19097=>"000001001",
  19098=>"111110010",
  19099=>"000000000",
  19100=>"110111111",
  19101=>"001000101",
  19102=>"111111100",
  19103=>"111111111",
  19104=>"111111110",
  19105=>"001111101",
  19106=>"111111111",
  19107=>"111001000",
  19108=>"000011011",
  19109=>"000000000",
  19110=>"111000100",
  19111=>"011111110",
  19112=>"111111111",
  19113=>"000000100",
  19114=>"000000000",
  19115=>"111111101",
  19116=>"111011111",
  19117=>"100000100",
  19118=>"111111110",
  19119=>"010111111",
  19120=>"000000000",
  19121=>"101100100",
  19122=>"010111011",
  19123=>"000101111",
  19124=>"111011000",
  19125=>"001000000",
  19126=>"000000000",
  19127=>"111100000",
  19128=>"000000100",
  19129=>"111111111",
  19130=>"101000000",
  19131=>"100000110",
  19132=>"101000000",
  19133=>"011011010",
  19134=>"101000000",
  19135=>"001111111",
  19136=>"001000000",
  19137=>"111011010",
  19138=>"000000111",
  19139=>"000000001",
  19140=>"111111111",
  19141=>"001000000",
  19142=>"111110111",
  19143=>"000000011",
  19144=>"100000001",
  19145=>"111101000",
  19146=>"001111011",
  19147=>"111111100",
  19148=>"000111111",
  19149=>"000100100",
  19150=>"110110111",
  19151=>"000011111",
  19152=>"010000110",
  19153=>"111001000",
  19154=>"111111001",
  19155=>"000000110",
  19156=>"101011000",
  19157=>"111000000",
  19158=>"001000000",
  19159=>"000000000",
  19160=>"111000000",
  19161=>"000000100",
  19162=>"011010000",
  19163=>"110111111",
  19164=>"111100100",
  19165=>"111011000",
  19166=>"110111111",
  19167=>"111011110",
  19168=>"000000111",
  19169=>"000000111",
  19170=>"111111100",
  19171=>"010000010",
  19172=>"001101000",
  19173=>"000111110",
  19174=>"101101111",
  19175=>"000000100",
  19176=>"111111011",
  19177=>"000000000",
  19178=>"000001110",
  19179=>"001111110",
  19180=>"111101101",
  19181=>"111111000",
  19182=>"111111111",
  19183=>"101000000",
  19184=>"101000000",
  19185=>"111110011",
  19186=>"011111011",
  19187=>"101000000",
  19188=>"110111111",
  19189=>"110000000",
  19190=>"000111111",
  19191=>"111111111",
  19192=>"111010000",
  19193=>"000000000",
  19194=>"111111111",
  19195=>"111111111",
  19196=>"001000111",
  19197=>"011011001",
  19198=>"000100000",
  19199=>"000000000",
  19200=>"101000000",
  19201=>"001011011",
  19202=>"010000000",
  19203=>"100000010",
  19204=>"000000000",
  19205=>"110110000",
  19206=>"111111111",
  19207=>"011001111",
  19208=>"100000000",
  19209=>"000000000",
  19210=>"000000000",
  19211=>"110111110",
  19212=>"001001001",
  19213=>"101001011",
  19214=>"111111111",
  19215=>"111111000",
  19216=>"000101110",
  19217=>"010111111",
  19218=>"001001001",
  19219=>"000000100",
  19220=>"111000000",
  19221=>"111111111",
  19222=>"001000000",
  19223=>"100101101",
  19224=>"001001001",
  19225=>"011011000",
  19226=>"000101101",
  19227=>"100000000",
  19228=>"000100101",
  19229=>"000111111",
  19230=>"000000000",
  19231=>"011111111",
  19232=>"100110000",
  19233=>"000000000",
  19234=>"000000000",
  19235=>"111110000",
  19236=>"000000000",
  19237=>"101000000",
  19238=>"000000000",
  19239=>"111111111",
  19240=>"111000000",
  19241=>"000111111",
  19242=>"000111111",
  19243=>"111111000",
  19244=>"000011111",
  19245=>"011001000",
  19246=>"000110111",
  19247=>"000010111",
  19248=>"000000000",
  19249=>"000000000",
  19250=>"011111101",
  19251=>"000000000",
  19252=>"000011111",
  19253=>"011011001",
  19254=>"111111101",
  19255=>"111111111",
  19256=>"110010000",
  19257=>"111100111",
  19258=>"000000001",
  19259=>"111000000",
  19260=>"000000100",
  19261=>"011001000",
  19262=>"000111111",
  19263=>"111111100",
  19264=>"001000000",
  19265=>"000000000",
  19266=>"000001001",
  19267=>"111000000",
  19268=>"000000000",
  19269=>"111100000",
  19270=>"000000111",
  19271=>"000000010",
  19272=>"111111111",
  19273=>"000001111",
  19274=>"000000000",
  19275=>"100011110",
  19276=>"110001000",
  19277=>"111111111",
  19278=>"100000000",
  19279=>"111010010",
  19280=>"011000000",
  19281=>"101000001",
  19282=>"000000000",
  19283=>"000000100",
  19284=>"000000000",
  19285=>"011011011",
  19286=>"101111111",
  19287=>"111111111",
  19288=>"111111011",
  19289=>"000000001",
  19290=>"111111111",
  19291=>"111011011",
  19292=>"000000000",
  19293=>"101101001",
  19294=>"101100100",
  19295=>"001000000",
  19296=>"000000000",
  19297=>"111100000",
  19298=>"111100111",
  19299=>"111001001",
  19300=>"110111110",
  19301=>"000000000",
  19302=>"111110111",
  19303=>"111001001",
  19304=>"111111111",
  19305=>"000000000",
  19306=>"000000000",
  19307=>"111001100",
  19308=>"000110111",
  19309=>"001000000",
  19310=>"010111111",
  19311=>"010000000",
  19312=>"000000000",
  19313=>"010010000",
  19314=>"001000000",
  19315=>"000111111",
  19316=>"110110110",
  19317=>"000000101",
  19318=>"111011111",
  19319=>"010010000",
  19320=>"111101101",
  19321=>"000000100",
  19322=>"000000000",
  19323=>"000000000",
  19324=>"000000101",
  19325=>"111100000",
  19326=>"000001000",
  19327=>"000111111",
  19328=>"010111111",
  19329=>"100111111",
  19330=>"100101001",
  19331=>"111111111",
  19332=>"010000011",
  19333=>"111101001",
  19334=>"101111111",
  19335=>"111111000",
  19336=>"000000000",
  19337=>"000000010",
  19338=>"001000001",
  19339=>"111111110",
  19340=>"111011111",
  19341=>"000110111",
  19342=>"010111111",
  19343=>"011000010",
  19344=>"000000111",
  19345=>"000000000",
  19346=>"111111111",
  19347=>"100000000",
  19348=>"111010011",
  19349=>"000000010",
  19350=>"000000000",
  19351=>"000000000",
  19352=>"100000000",
  19353=>"000000000",
  19354=>"110111111",
  19355=>"111110000",
  19356=>"000100000",
  19357=>"001000000",
  19358=>"101100000",
  19359=>"110111111",
  19360=>"000000000",
  19361=>"010111111",
  19362=>"000000010",
  19363=>"111000000",
  19364=>"111111110",
  19365=>"110111111",
  19366=>"001001001",
  19367=>"111111111",
  19368=>"000000000",
  19369=>"001000000",
  19370=>"010111010",
  19371=>"111001000",
  19372=>"000011111",
  19373=>"111101111",
  19374=>"111100000",
  19375=>"111111001",
  19376=>"111000111",
  19377=>"000011111",
  19378=>"000000000",
  19379=>"000000000",
  19380=>"001000000",
  19381=>"000000000",
  19382=>"000000110",
  19383=>"000111000",
  19384=>"111101001",
  19385=>"000011011",
  19386=>"111010110",
  19387=>"010111111",
  19388=>"000010000",
  19389=>"001000000",
  19390=>"111111100",
  19391=>"100110100",
  19392=>"000000000",
  19393=>"000000000",
  19394=>"001000000",
  19395=>"000000001",
  19396=>"001001110",
  19397=>"010011111",
  19398=>"000000000",
  19399=>"000000000",
  19400=>"000001000",
  19401=>"100000111",
  19402=>"001111111",
  19403=>"000000000",
  19404=>"000000000",
  19405=>"110111111",
  19406=>"000000000",
  19407=>"111101001",
  19408=>"111100000",
  19409=>"111111011",
  19410=>"100100000",
  19411=>"000000000",
  19412=>"011111111",
  19413=>"111101000",
  19414=>"111111001",
  19415=>"010111111",
  19416=>"101000000",
  19417=>"111101100",
  19418=>"111111000",
  19419=>"000000000",
  19420=>"011101100",
  19421=>"111111101",
  19422=>"000111111",
  19423=>"000100000",
  19424=>"101001000",
  19425=>"000100111",
  19426=>"000000000",
  19427=>"011000000",
  19428=>"111111111",
  19429=>"111100000",
  19430=>"000000110",
  19431=>"111011000",
  19432=>"111000000",
  19433=>"111000000",
  19434=>"110111110",
  19435=>"101001000",
  19436=>"111111010",
  19437=>"001000100",
  19438=>"101101101",
  19439=>"001001011",
  19440=>"000000000",
  19441=>"000111111",
  19442=>"000000000",
  19443=>"111111111",
  19444=>"111111111",
  19445=>"000000000",
  19446=>"111111111",
  19447=>"011000000",
  19448=>"110111011",
  19449=>"000001001",
  19450=>"111011000",
  19451=>"001000000",
  19452=>"000000000",
  19453=>"111111111",
  19454=>"111111000",
  19455=>"000000000",
  19456=>"110000100",
  19457=>"111000000",
  19458=>"000000000",
  19459=>"000110110",
  19460=>"111111111",
  19461=>"001001001",
  19462=>"111101101",
  19463=>"111001111",
  19464=>"000000000",
  19465=>"001111110",
  19466=>"010000000",
  19467=>"000000100",
  19468=>"001011011",
  19469=>"111000000",
  19470=>"001000000",
  19471=>"000110000",
  19472=>"000110110",
  19473=>"111111111",
  19474=>"111111110",
  19475=>"000000000",
  19476=>"111000000",
  19477=>"111111111",
  19478=>"000000100",
  19479=>"110110100",
  19480=>"000000000",
  19481=>"000000111",
  19482=>"110111111",
  19483=>"111111111",
  19484=>"100100111",
  19485=>"000011000",
  19486=>"000000000",
  19487=>"000000111",
  19488=>"111111111",
  19489=>"000000000",
  19490=>"110111111",
  19491=>"111111000",
  19492=>"111111110",
  19493=>"000000000",
  19494=>"111001000",
  19495=>"110100000",
  19496=>"111011110",
  19497=>"111111111",
  19498=>"000000000",
  19499=>"000000111",
  19500=>"000000000",
  19501=>"000000000",
  19502=>"011011011",
  19503=>"110010011",
  19504=>"000000110",
  19505=>"100000100",
  19506=>"000000000",
  19507=>"000111111",
  19508=>"111101000",
  19509=>"110110010",
  19510=>"000000100",
  19511=>"101100000",
  19512=>"000110111",
  19513=>"111111101",
  19514=>"111111111",
  19515=>"111111010",
  19516=>"000000100",
  19517=>"000111111",
  19518=>"000000000",
  19519=>"111011111",
  19520=>"111111111",
  19521=>"111111011",
  19522=>"011111000",
  19523=>"111111111",
  19524=>"111011011",
  19525=>"000000111",
  19526=>"111111010",
  19527=>"111000000",
  19528=>"100110111",
  19529=>"111111111",
  19530=>"111111111",
  19531=>"111111000",
  19532=>"000000011",
  19533=>"000000100",
  19534=>"000000000",
  19535=>"000000111",
  19536=>"111111000",
  19537=>"000001000",
  19538=>"110000000",
  19539=>"111010000",
  19540=>"000000000",
  19541=>"000000100",
  19542=>"110010000",
  19543=>"111111111",
  19544=>"001111110",
  19545=>"111000000",
  19546=>"001001111",
  19547=>"001000000",
  19548=>"111111111",
  19549=>"000000111",
  19550=>"000000110",
  19551=>"000000000",
  19552=>"111001000",
  19553=>"000110000",
  19554=>"111111000",
  19555=>"000000111",
  19556=>"110111010",
  19557=>"111111000",
  19558=>"101110111",
  19559=>"111100101",
  19560=>"001100000",
  19561=>"000000000",
  19562=>"111111111",
  19563=>"111111001",
  19564=>"000000000",
  19565=>"111111000",
  19566=>"000000100",
  19567=>"000000101",
  19568=>"100000000",
  19569=>"011000000",
  19570=>"001110000",
  19571=>"000000110",
  19572=>"111000000",
  19573=>"110111000",
  19574=>"111111111",
  19575=>"000000000",
  19576=>"000000000",
  19577=>"111111111",
  19578=>"111011011",
  19579=>"111111000",
  19580=>"100000000",
  19581=>"000000000",
  19582=>"111111011",
  19583=>"000000000",
  19584=>"110100111",
  19585=>"111111111",
  19586=>"000000000",
  19587=>"111111000",
  19588=>"111111111",
  19589=>"000000100",
  19590=>"000001001",
  19591=>"111110010",
  19592=>"011000111",
  19593=>"000010111",
  19594=>"111011001",
  19595=>"001000110",
  19596=>"101111111",
  19597=>"000100111",
  19598=>"111111000",
  19599=>"001101001",
  19600=>"111111111",
  19601=>"000000000",
  19602=>"000011111",
  19603=>"111111111",
  19604=>"001000001",
  19605=>"000000000",
  19606=>"111111111",
  19607=>"000000000",
  19608=>"111001110",
  19609=>"000000001",
  19610=>"000010110",
  19611=>"000000000",
  19612=>"000000000",
  19613=>"011011111",
  19614=>"111101000",
  19615=>"111111000",
  19616=>"111111101",
  19617=>"011111111",
  19618=>"000011110",
  19619=>"010000000",
  19620=>"111111111",
  19621=>"000000111",
  19622=>"000000000",
  19623=>"000000000",
  19624=>"111111111",
  19625=>"100000000",
  19626=>"100100111",
  19627=>"111010110",
  19628=>"000111111",
  19629=>"111111111",
  19630=>"111111000",
  19631=>"111001001",
  19632=>"111111100",
  19633=>"011010000",
  19634=>"111111111",
  19635=>"100000100",
  19636=>"000000000",
  19637=>"110111000",
  19638=>"000000000",
  19639=>"011111000",
  19640=>"000000000",
  19641=>"111000001",
  19642=>"111111111",
  19643=>"110111100",
  19644=>"000000000",
  19645=>"100000101",
  19646=>"100111000",
  19647=>"000000000",
  19648=>"111001011",
  19649=>"111111110",
  19650=>"111111111",
  19651=>"111111111",
  19652=>"001011111",
  19653=>"000000000",
  19654=>"110010001",
  19655=>"001001000",
  19656=>"000111111",
  19657=>"011111111",
  19658=>"000000111",
  19659=>"101101111",
  19660=>"000010000",
  19661=>"111111000",
  19662=>"000000000",
  19663=>"000011011",
  19664=>"111111111",
  19665=>"111111111",
  19666=>"111110000",
  19667=>"001111000",
  19668=>"100110110",
  19669=>"111111000",
  19670=>"000001001",
  19671=>"001000000",
  19672=>"111000000",
  19673=>"000000000",
  19674=>"111111111",
  19675=>"000000111",
  19676=>"111110000",
  19677=>"000110110",
  19678=>"001000000",
  19679=>"111111111",
  19680=>"111101100",
  19681=>"000000111",
  19682=>"000100111",
  19683=>"110111111",
  19684=>"000111111",
  19685=>"000000000",
  19686=>"011001000",
  19687=>"011111000",
  19688=>"010111110",
  19689=>"110111010",
  19690=>"111111110",
  19691=>"111111111",
  19692=>"000000001",
  19693=>"000000000",
  19694=>"000000101",
  19695=>"000000000",
  19696=>"101111110",
  19697=>"000111110",
  19698=>"111111111",
  19699=>"111111111",
  19700=>"000010110",
  19701=>"110011000",
  19702=>"011011001",
  19703=>"000110000",
  19704=>"111111111",
  19705=>"001111111",
  19706=>"000000000",
  19707=>"111111111",
  19708=>"111111111",
  19709=>"001001111",
  19710=>"111111111",
  19711=>"111000000",
  19712=>"000000101",
  19713=>"000010000",
  19714=>"111111011",
  19715=>"000000000",
  19716=>"111111000",
  19717=>"010000000",
  19718=>"111111000",
  19719=>"000011001",
  19720=>"000000000",
  19721=>"000000000",
  19722=>"000000000",
  19723=>"111111000",
  19724=>"111110110",
  19725=>"110111111",
  19726=>"000111000",
  19727=>"001101111",
  19728=>"000000000",
  19729=>"110111111",
  19730=>"100000000",
  19731=>"000000111",
  19732=>"111101111",
  19733=>"000000000",
  19734=>"000111001",
  19735=>"000000111",
  19736=>"000000000",
  19737=>"110110000",
  19738=>"000011011",
  19739=>"101111111",
  19740=>"000000000",
  19741=>"000000000",
  19742=>"111101111",
  19743=>"111001000",
  19744=>"000000000",
  19745=>"000000101",
  19746=>"111111011",
  19747=>"111011001",
  19748=>"000000000",
  19749=>"110111111",
  19750=>"000110111",
  19751=>"000000000",
  19752=>"111011000",
  19753=>"110111111",
  19754=>"111111011",
  19755=>"111111001",
  19756=>"000000000",
  19757=>"000100100",
  19758=>"000000000",
  19759=>"100000000",
  19760=>"111111000",
  19761=>"000011000",
  19762=>"111111111",
  19763=>"100101111",
  19764=>"000000000",
  19765=>"000000000",
  19766=>"000100000",
  19767=>"000000000",
  19768=>"000000001",
  19769=>"100000001",
  19770=>"000000000",
  19771=>"011111111",
  19772=>"000000000",
  19773=>"000010110",
  19774=>"100100111",
  19775=>"000000000",
  19776=>"011100101",
  19777=>"111111000",
  19778=>"000000111",
  19779=>"111111111",
  19780=>"000101000",
  19781=>"000000000",
  19782=>"111111111",
  19783=>"111111111",
  19784=>"000000000",
  19785=>"101000000",
  19786=>"000111111",
  19787=>"010111001",
  19788=>"110000000",
  19789=>"111111000",
  19790=>"111111101",
  19791=>"000111111",
  19792=>"000000100",
  19793=>"111111111",
  19794=>"110111110",
  19795=>"111110111",
  19796=>"111111111",
  19797=>"001011001",
  19798=>"111111000",
  19799=>"111110000",
  19800=>"011011111",
  19801=>"000000000",
  19802=>"000111110",
  19803=>"111111011",
  19804=>"000000000",
  19805=>"001111111",
  19806=>"011011111",
  19807=>"000000000",
  19808=>"000100100",
  19809=>"111000000",
  19810=>"011011111",
  19811=>"100000000",
  19812=>"111111111",
  19813=>"000000000",
  19814=>"100000100",
  19815=>"000000100",
  19816=>"011011000",
  19817=>"000111011",
  19818=>"000100111",
  19819=>"111111000",
  19820=>"111110110",
  19821=>"000010010",
  19822=>"111111000",
  19823=>"000000000",
  19824=>"000000000",
  19825=>"000000000",
  19826=>"101000000",
  19827=>"000000100",
  19828=>"111111111",
  19829=>"000000000",
  19830=>"000001000",
  19831=>"111110000",
  19832=>"000100100",
  19833=>"100110111",
  19834=>"001000000",
  19835=>"000010100",
  19836=>"100000000",
  19837=>"000000101",
  19838=>"000110000",
  19839=>"111111011",
  19840=>"001000000",
  19841=>"001000111",
  19842=>"000111111",
  19843=>"000000000",
  19844=>"100110110",
  19845=>"111111110",
  19846=>"100110111",
  19847=>"010010000",
  19848=>"000000000",
  19849=>"110111000",
  19850=>"011001010",
  19851=>"011101111",
  19852=>"111111111",
  19853=>"011011001",
  19854=>"010111111",
  19855=>"000111111",
  19856=>"111111001",
  19857=>"111111000",
  19858=>"111110001",
  19859=>"000000000",
  19860=>"000000111",
  19861=>"000100000",
  19862=>"000000000",
  19863=>"000000010",
  19864=>"111111111",
  19865=>"100110010",
  19866=>"001000000",
  19867=>"111111110",
  19868=>"000100100",
  19869=>"011111100",
  19870=>"000000000",
  19871=>"000111111",
  19872=>"000001011",
  19873=>"000000111",
  19874=>"111111111",
  19875=>"000000110",
  19876=>"011111100",
  19877=>"111011111",
  19878=>"001000000",
  19879=>"110111111",
  19880=>"110111111",
  19881=>"001000000",
  19882=>"110111111",
  19883=>"000000000",
  19884=>"000000100",
  19885=>"100111101",
  19886=>"000000010",
  19887=>"110111110",
  19888=>"111000011",
  19889=>"111111000",
  19890=>"000000001",
  19891=>"100001000",
  19892=>"000011110",
  19893=>"110111111",
  19894=>"111111111",
  19895=>"000000000",
  19896=>"000000010",
  19897=>"000001000",
  19898=>"010100110",
  19899=>"000000000",
  19900=>"011000000",
  19901=>"111111000",
  19902=>"111000000",
  19903=>"011000000",
  19904=>"000000111",
  19905=>"000000000",
  19906=>"000000001",
  19907=>"000000111",
  19908=>"000011111",
  19909=>"000110111",
  19910=>"011101100",
  19911=>"000001001",
  19912=>"000001101",
  19913=>"101000000",
  19914=>"111011011",
  19915=>"000100111",
  19916=>"111111000",
  19917=>"000000000",
  19918=>"110111101",
  19919=>"011111111",
  19920=>"110011000",
  19921=>"000010000",
  19922=>"101111111",
  19923=>"101000000",
  19924=>"101111111",
  19925=>"000000000",
  19926=>"111111110",
  19927=>"110110111",
  19928=>"000011111",
  19929=>"000000000",
  19930=>"000000000",
  19931=>"000000000",
  19932=>"101111111",
  19933=>"111111111",
  19934=>"000000000",
  19935=>"000110111",
  19936=>"100100111",
  19937=>"111000000",
  19938=>"111111111",
  19939=>"101001000",
  19940=>"000000000",
  19941=>"011000000",
  19942=>"100101100",
  19943=>"010010000",
  19944=>"010100111",
  19945=>"000010011",
  19946=>"111111100",
  19947=>"000011111",
  19948=>"000000000",
  19949=>"001111000",
  19950=>"000000111",
  19951=>"000000000",
  19952=>"000000100",
  19953=>"000000000",
  19954=>"011111111",
  19955=>"000111111",
  19956=>"111110111",
  19957=>"000000000",
  19958=>"000011111",
  19959=>"000100110",
  19960=>"110110110",
  19961=>"100110000",
  19962=>"001001001",
  19963=>"000100111",
  19964=>"001010111",
  19965=>"001000000",
  19966=>"111001001",
  19967=>"100110111",
  19968=>"111111111",
  19969=>"011000111",
  19970=>"111101111",
  19971=>"111111111",
  19972=>"001101111",
  19973=>"001000000",
  19974=>"111111111",
  19975=>"111111111",
  19976=>"111010100",
  19977=>"111100101",
  19978=>"101000100",
  19979=>"000000000",
  19980=>"110011001",
  19981=>"000000011",
  19982=>"111111111",
  19983=>"001111111",
  19984=>"000000000",
  19985=>"011000000",
  19986=>"001111111",
  19987=>"100000111",
  19988=>"000000000",
  19989=>"000000001",
  19990=>"111011111",
  19991=>"111101001",
  19992=>"000000000",
  19993=>"000000000",
  19994=>"110000010",
  19995=>"010000000",
  19996=>"110000000",
  19997=>"000011111",
  19998=>"110110110",
  19999=>"111111000",
  20000=>"111111000",
  20001=>"000000111",
  20002=>"111111111",
  20003=>"111110000",
  20004=>"000000111",
  20005=>"111110111",
  20006=>"111110111",
  20007=>"000000100",
  20008=>"111000000",
  20009=>"000010111",
  20010=>"000000000",
  20011=>"100111111",
  20012=>"110111111",
  20013=>"111111111",
  20014=>"100000101",
  20015=>"000000000",
  20016=>"000000000",
  20017=>"111111111",
  20018=>"000111000",
  20019=>"111100000",
  20020=>"001000000",
  20021=>"000000000",
  20022=>"000111111",
  20023=>"000000001",
  20024=>"110111111",
  20025=>"000000000",
  20026=>"111001000",
  20027=>"110110000",
  20028=>"111000000",
  20029=>"000111111",
  20030=>"111110010",
  20031=>"000000000",
  20032=>"000001000",
  20033=>"001001100",
  20034=>"000111111",
  20035=>"011111111",
  20036=>"111111111",
  20037=>"000000000",
  20038=>"000000111",
  20039=>"000000000",
  20040=>"111011000",
  20041=>"000000000",
  20042=>"111111111",
  20043=>"000000111",
  20044=>"100100000",
  20045=>"111010000",
  20046=>"110110111",
  20047=>"000111111",
  20048=>"000000000",
  20049=>"100111111",
  20050=>"000001111",
  20051=>"001001000",
  20052=>"000000000",
  20053=>"111011111",
  20054=>"000000000",
  20055=>"111001000",
  20056=>"111101001",
  20057=>"101000000",
  20058=>"000000110",
  20059=>"000000001",
  20060=>"000000111",
  20061=>"000010000",
  20062=>"111111111",
  20063=>"010110110",
  20064=>"111111111",
  20065=>"000000000",
  20066=>"111111011",
  20067=>"111111111",
  20068=>"001001111",
  20069=>"111100100",
  20070=>"111111111",
  20071=>"000000000",
  20072=>"000000000",
  20073=>"111001011",
  20074=>"001111111",
  20075=>"010010010",
  20076=>"111111011",
  20077=>"111111111",
  20078=>"001111111",
  20079=>"111111011",
  20080=>"000000000",
  20081=>"000100111",
  20082=>"000110110",
  20083=>"111110000",
  20084=>"000000000",
  20085=>"000111111",
  20086=>"000000000",
  20087=>"111111111",
  20088=>"100000000",
  20089=>"011001000",
  20090=>"000000010",
  20091=>"000111111",
  20092=>"001000000",
  20093=>"111111111",
  20094=>"110110111",
  20095=>"111111111",
  20096=>"000000111",
  20097=>"000000000",
  20098=>"000000000",
  20099=>"110110000",
  20100=>"111000000",
  20101=>"111110111",
  20102=>"000000001",
  20103=>"011000000",
  20104=>"110110000",
  20105=>"000011011",
  20106=>"111111111",
  20107=>"100100000",
  20108=>"111111111",
  20109=>"111000000",
  20110=>"100000000",
  20111=>"111111111",
  20112=>"111100101",
  20113=>"111111111",
  20114=>"110110111",
  20115=>"100000000",
  20116=>"000011111",
  20117=>"111011011",
  20118=>"000000000",
  20119=>"000000000",
  20120=>"111100000",
  20121=>"100101011",
  20122=>"000000000",
  20123=>"000000000",
  20124=>"111111111",
  20125=>"000000000",
  20126=>"110111011",
  20127=>"000000000",
  20128=>"111111111",
  20129=>"110010010",
  20130=>"111111111",
  20131=>"000000000",
  20132=>"111110100",
  20133=>"111111111",
  20134=>"111000000",
  20135=>"110100100",
  20136=>"000010011",
  20137=>"111110110",
  20138=>"101001101",
  20139=>"001000001",
  20140=>"111111111",
  20141=>"000110111",
  20142=>"000000000",
  20143=>"000110111",
  20144=>"111111111",
  20145=>"000000110",
  20146=>"111111111",
  20147=>"111000000",
  20148=>"111011100",
  20149=>"101000000",
  20150=>"011010111",
  20151=>"101111111",
  20152=>"111000111",
  20153=>"111111111",
  20154=>"110000000",
  20155=>"111000010",
  20156=>"111111000",
  20157=>"001000011",
  20158=>"111111011",
  20159=>"110000000",
  20160=>"111011001",
  20161=>"111111111",
  20162=>"001000000",
  20163=>"000000000",
  20164=>"100000000",
  20165=>"000000000",
  20166=>"000010000",
  20167=>"000011101",
  20168=>"000000010",
  20169=>"100000000",
  20170=>"000000000",
  20171=>"000000000",
  20172=>"100100110",
  20173=>"000100000",
  20174=>"011111111",
  20175=>"000000000",
  20176=>"111000111",
  20177=>"111000111",
  20178=>"111111111",
  20179=>"000011000",
  20180=>"111111111",
  20181=>"000000000",
  20182=>"110000000",
  20183=>"100001001",
  20184=>"101011111",
  20185=>"111111111",
  20186=>"000001101",
  20187=>"000010111",
  20188=>"000000000",
  20189=>"111111111",
  20190=>"111100100",
  20191=>"111111111",
  20192=>"001101000",
  20193=>"000000000",
  20194=>"111111110",
  20195=>"101100001",
  20196=>"000000011",
  20197=>"000000000",
  20198=>"001001000",
  20199=>"001000111",
  20200=>"001000000",
  20201=>"110000000",
  20202=>"111111111",
  20203=>"111011010",
  20204=>"100100111",
  20205=>"000000011",
  20206=>"111111011",
  20207=>"101000110",
  20208=>"100000000",
  20209=>"100100101",
  20210=>"111111111",
  20211=>"111110100",
  20212=>"111001111",
  20213=>"111111111",
  20214=>"110000101",
  20215=>"111111110",
  20216=>"000000000",
  20217=>"010000000",
  20218=>"111111000",
  20219=>"000100100",
  20220=>"000000000",
  20221=>"000000010",
  20222=>"110111111",
  20223=>"110111110",
  20224=>"100000000",
  20225=>"011111011",
  20226=>"111111111",
  20227=>"111000000",
  20228=>"101000000",
  20229=>"000111111",
  20230=>"111000000",
  20231=>"000000001",
  20232=>"110111110",
  20233=>"000000000",
  20234=>"001011001",
  20235=>"111111011",
  20236=>"110100000",
  20237=>"100101011",
  20238=>"110010101",
  20239=>"000000000",
  20240=>"000110111",
  20241=>"111001001",
  20242=>"000010111",
  20243=>"111100100",
  20244=>"111111111",
  20245=>"000000000",
  20246=>"001011111",
  20247=>"011111101",
  20248=>"000000000",
  20249=>"111111111",
  20250=>"111111111",
  20251=>"000001101",
  20252=>"000000100",
  20253=>"011010111",
  20254=>"000000000",
  20255=>"111000101",
  20256=>"000000000",
  20257=>"000000000",
  20258=>"110111111",
  20259=>"000000010",
  20260=>"111111111",
  20261=>"000111111",
  20262=>"101100101",
  20263=>"000000000",
  20264=>"000000011",
  20265=>"011110010",
  20266=>"000000000",
  20267=>"000000000",
  20268=>"000001000",
  20269=>"010110100",
  20270=>"000000111",
  20271=>"000000000",
  20272=>"000000000",
  20273=>"011111111",
  20274=>"001001011",
  20275=>"111111010",
  20276=>"110110111",
  20277=>"111111001",
  20278=>"000000000",
  20279=>"011110110",
  20280=>"110100000",
  20281=>"111110110",
  20282=>"100111011",
  20283=>"111111111",
  20284=>"111000100",
  20285=>"110111000",
  20286=>"001000000",
  20287=>"000000010",
  20288=>"111111100",
  20289=>"111111111",
  20290=>"111101111",
  20291=>"111111101",
  20292=>"000000001",
  20293=>"000000000",
  20294=>"100000000",
  20295=>"000111000",
  20296=>"000111111",
  20297=>"001000111",
  20298=>"110110111",
  20299=>"000001000",
  20300=>"000000111",
  20301=>"000000111",
  20302=>"000010111",
  20303=>"000111111",
  20304=>"010011000",
  20305=>"111111111",
  20306=>"000000000",
  20307=>"010011100",
  20308=>"011011000",
  20309=>"011011011",
  20310=>"011011010",
  20311=>"000000100",
  20312=>"111010000",
  20313=>"000000001",
  20314=>"000111111",
  20315=>"000000000",
  20316=>"000000100",
  20317=>"101111111",
  20318=>"000000000",
  20319=>"111111000",
  20320=>"111000111",
  20321=>"111111000",
  20322=>"011001100",
  20323=>"111111111",
  20324=>"011111111",
  20325=>"111111001",
  20326=>"111001001",
  20327=>"000000000",
  20328=>"000000000",
  20329=>"111111100",
  20330=>"000000111",
  20331=>"000000000",
  20332=>"110000000",
  20333=>"111110111",
  20334=>"000000001",
  20335=>"101100111",
  20336=>"111111111",
  20337=>"111111111",
  20338=>"011111111",
  20339=>"101100100",
  20340=>"110110010",
  20341=>"111111111",
  20342=>"100110000",
  20343=>"000001011",
  20344=>"111111111",
  20345=>"000000111",
  20346=>"000011111",
  20347=>"000000011",
  20348=>"111111011",
  20349=>"111111111",
  20350=>"000010111",
  20351=>"000000000",
  20352=>"001111111",
  20353=>"111111000",
  20354=>"000000110",
  20355=>"100000000",
  20356=>"000000001",
  20357=>"111110000",
  20358=>"111111111",
  20359=>"010011000",
  20360=>"011111111",
  20361=>"011111111",
  20362=>"000000000",
  20363=>"000000010",
  20364=>"000000001",
  20365=>"000000000",
  20366=>"111111010",
  20367=>"000000000",
  20368=>"000000000",
  20369=>"011011001",
  20370=>"000001101",
  20371=>"101001111",
  20372=>"110000111",
  20373=>"111110010",
  20374=>"000000000",
  20375=>"111011001",
  20376=>"100101101",
  20377=>"111111011",
  20378=>"010010010",
  20379=>"111000000",
  20380=>"010011011",
  20381=>"000000000",
  20382=>"111110000",
  20383=>"000000000",
  20384=>"100100000",
  20385=>"110110111",
  20386=>"111111111",
  20387=>"000001111",
  20388=>"111111000",
  20389=>"111111111",
  20390=>"000000111",
  20391=>"000000000",
  20392=>"111111110",
  20393=>"000000000",
  20394=>"111111111",
  20395=>"111001111",
  20396=>"010010000",
  20397=>"100000011",
  20398=>"000110011",
  20399=>"000011111",
  20400=>"010011111",
  20401=>"110100000",
  20402=>"111111111",
  20403=>"111111111",
  20404=>"110000110",
  20405=>"000000000",
  20406=>"101111111",
  20407=>"100101001",
  20408=>"111111111",
  20409=>"000010011",
  20410=>"111011111",
  20411=>"110000000",
  20412=>"001011000",
  20413=>"000011111",
  20414=>"110111111",
  20415=>"000000100",
  20416=>"110000000",
  20417=>"000000111",
  20418=>"111111111",
  20419=>"100100110",
  20420=>"000000000",
  20421=>"000100110",
  20422=>"000000000",
  20423=>"111111111",
  20424=>"000100000",
  20425=>"000111111",
  20426=>"000100110",
  20427=>"110111110",
  20428=>"101000000",
  20429=>"111111111",
  20430=>"000000111",
  20431=>"111111111",
  20432=>"111111111",
  20433=>"111111110",
  20434=>"000000011",
  20435=>"000000000",
  20436=>"111011001",
  20437=>"001001000",
  20438=>"111011000",
  20439=>"111111110",
  20440=>"000000000",
  20441=>"000000000",
  20442=>"000000111",
  20443=>"111100111",
  20444=>"000000111",
  20445=>"111111111",
  20446=>"001000000",
  20447=>"100110111",
  20448=>"101111111",
  20449=>"111111111",
  20450=>"111011111",
  20451=>"010100101",
  20452=>"101000000",
  20453=>"111111111",
  20454=>"000000000",
  20455=>"000001111",
  20456=>"111100000",
  20457=>"111000000",
  20458=>"001000000",
  20459=>"111000001",
  20460=>"000000111",
  20461=>"111100100",
  20462=>"000001011",
  20463=>"101100000",
  20464=>"111110110",
  20465=>"111111111",
  20466=>"000111111",
  20467=>"000000000",
  20468=>"111111000",
  20469=>"000000011",
  20470=>"001001000",
  20471=>"111011010",
  20472=>"111100000",
  20473=>"011001101",
  20474=>"001011011",
  20475=>"000111111",
  20476=>"000000111",
  20477=>"000000000",
  20478=>"000000000",
  20479=>"110111111",
  20480=>"101000000",
  20481=>"111000000",
  20482=>"110000100",
  20483=>"110111111",
  20484=>"000000111",
  20485=>"111100111",
  20486=>"000000000",
  20487=>"000000000",
  20488=>"011000001",
  20489=>"000111110",
  20490=>"001000001",
  20491=>"000001000",
  20492=>"000000001",
  20493=>"000000000",
  20494=>"000110111",
  20495=>"111111000",
  20496=>"000000001",
  20497=>"000000000",
  20498=>"001111001",
  20499=>"010110111",
  20500=>"000000100",
  20501=>"111111110",
  20502=>"110010110",
  20503=>"111100111",
  20504=>"111110000",
  20505=>"000001111",
  20506=>"111111111",
  20507=>"000000110",
  20508=>"111111111",
  20509=>"111110010",
  20510=>"000000110",
  20511=>"110111111",
  20512=>"000000011",
  20513=>"111111100",
  20514=>"000000000",
  20515=>"000000000",
  20516=>"111111111",
  20517=>"000000100",
  20518=>"110111111",
  20519=>"100100111",
  20520=>"000000000",
  20521=>"000000100",
  20522=>"101000001",
  20523=>"000000000",
  20524=>"000000000",
  20525=>"000101111",
  20526=>"001000001",
  20527=>"000000000",
  20528=>"000000000",
  20529=>"111111111",
  20530=>"001001001",
  20531=>"100000010",
  20532=>"000000001",
  20533=>"110011011",
  20534=>"000000011",
  20535=>"000010111",
  20536=>"111111111",
  20537=>"000000010",
  20538=>"000000000",
  20539=>"011011111",
  20540=>"111111111",
  20541=>"111111111",
  20542=>"011111111",
  20543=>"101000000",
  20544=>"011000000",
  20545=>"110010111",
  20546=>"001011011",
  20547=>"110100011",
  20548=>"011000000",
  20549=>"001001001",
  20550=>"000000000",
  20551=>"111111101",
  20552=>"001001001",
  20553=>"000000000",
  20554=>"111111001",
  20555=>"010010110",
  20556=>"000000111",
  20557=>"010010011",
  20558=>"111111000",
  20559=>"111111111",
  20560=>"001000000",
  20561=>"000011001",
  20562=>"000000000",
  20563=>"111111011",
  20564=>"000110111",
  20565=>"000000100",
  20566=>"011011011",
  20567=>"000000000",
  20568=>"111111011",
  20569=>"000000000",
  20570=>"111111000",
  20571=>"001001000",
  20572=>"111111111",
  20573=>"110000011",
  20574=>"000000000",
  20575=>"111111101",
  20576=>"111111101",
  20577=>"111111111",
  20578=>"111111011",
  20579=>"111111111",
  20580=>"100100000",
  20581=>"000001011",
  20582=>"000000000",
  20583=>"000000001",
  20584=>"000010010",
  20585=>"111111110",
  20586=>"011011000",
  20587=>"111111010",
  20588=>"111001001",
  20589=>"111111110",
  20590=>"111111111",
  20591=>"000010000",
  20592=>"110110010",
  20593=>"011011111",
  20594=>"111111110",
  20595=>"110100110",
  20596=>"000000111",
  20597=>"000001001",
  20598=>"111111111",
  20599=>"111000111",
  20600=>"000001001",
  20601=>"111111100",
  20602=>"001111111",
  20603=>"000011011",
  20604=>"111111110",
  20605=>"001001001",
  20606=>"011011000",
  20607=>"111101111",
  20608=>"000000000",
  20609=>"111111111",
  20610=>"001111111",
  20611=>"011111111",
  20612=>"111111111",
  20613=>"000000111",
  20614=>"110110110",
  20615=>"100000000",
  20616=>"001000010",
  20617=>"001001001",
  20618=>"111111111",
  20619=>"000000001",
  20620=>"111111111",
  20621=>"111010000",
  20622=>"000000000",
  20623=>"000000001",
  20624=>"111011011",
  20625=>"000100111",
  20626=>"000000011",
  20627=>"111101111",
  20628=>"000000000",
  20629=>"011011011",
  20630=>"111111111",
  20631=>"000000000",
  20632=>"111111110",
  20633=>"000100000",
  20634=>"000000010",
  20635=>"011111011",
  20636=>"011111110",
  20637=>"000000111",
  20638=>"000001111",
  20639=>"010000000",
  20640=>"110111111",
  20641=>"110110010",
  20642=>"000000000",
  20643=>"111111111",
  20644=>"001101000",
  20645=>"111111111",
  20646=>"111111111",
  20647=>"011111010",
  20648=>"000000000",
  20649=>"000000000",
  20650=>"000000100",
  20651=>"000000000",
  20652=>"000001101",
  20653=>"110111110",
  20654=>"000010010",
  20655=>"011011001",
  20656=>"111000000",
  20657=>"011111001",
  20658=>"111111111",
  20659=>"000000000",
  20660=>"111100000",
  20661=>"000001001",
  20662=>"000000000",
  20663=>"100000000",
  20664=>"000000000",
  20665=>"111111000",
  20666=>"001011011",
  20667=>"000000001",
  20668=>"111111111",
  20669=>"000000000",
  20670=>"110000010",
  20671=>"111111111",
  20672=>"111111111",
  20673=>"000000110",
  20674=>"001000000",
  20675=>"000000011",
  20676=>"000000000",
  20677=>"000000110",
  20678=>"000000000",
  20679=>"000000000",
  20680=>"000100000",
  20681=>"111100100",
  20682=>"111111111",
  20683=>"001001001",
  20684=>"111111000",
  20685=>"110100000",
  20686=>"011001101",
  20687=>"000000111",
  20688=>"000000000",
  20689=>"111111111",
  20690=>"001000000",
  20691=>"000000000",
  20692=>"111111011",
  20693=>"111111111",
  20694=>"101101101",
  20695=>"110000111",
  20696=>"100100111",
  20697=>"000000000",
  20698=>"000000000",
  20699=>"011100111",
  20700=>"111111111",
  20701=>"100000111",
  20702=>"111001111",
  20703=>"000000111",
  20704=>"101100000",
  20705=>"111110110",
  20706=>"000000000",
  20707=>"001000000",
  20708=>"111111111",
  20709=>"100000000",
  20710=>"001001000",
  20711=>"011001001",
  20712=>"000000000",
  20713=>"100101111",
  20714=>"111000000",
  20715=>"000001111",
  20716=>"111111111",
  20717=>"000000000",
  20718=>"001111101",
  20719=>"010000011",
  20720=>"000000000",
  20721=>"001000000",
  20722=>"111111111",
  20723=>"011010000",
  20724=>"011000001",
  20725=>"110110110",
  20726=>"111111111",
  20727=>"111000000",
  20728=>"000000000",
  20729=>"000000000",
  20730=>"110000000",
  20731=>"000000000",
  20732=>"111100000",
  20733=>"110000100",
  20734=>"001101111",
  20735=>"000111111",
  20736=>"111111100",
  20737=>"111100100",
  20738=>"111111100",
  20739=>"000010001",
  20740=>"111111111",
  20741=>"100000000",
  20742=>"111111111",
  20743=>"000010110",
  20744=>"001001111",
  20745=>"100100110",
  20746=>"111111111",
  20747=>"111111111",
  20748=>"111101001",
  20749=>"111111111",
  20750=>"111111010",
  20751=>"000011111",
  20752=>"000000000",
  20753=>"000000001",
  20754=>"000000111",
  20755=>"100100100",
  20756=>"000000101",
  20757=>"000000000",
  20758=>"010011011",
  20759=>"011001011",
  20760=>"100100110",
  20761=>"011111011",
  20762=>"000000001",
  20763=>"001111111",
  20764=>"100010000",
  20765=>"111111111",
  20766=>"000001111",
  20767=>"000000000",
  20768=>"000000010",
  20769=>"000000000",
  20770=>"100000000",
  20771=>"000000111",
  20772=>"000000100",
  20773=>"111111111",
  20774=>"011011011",
  20775=>"101111111",
  20776=>"111111101",
  20777=>"011000000",
  20778=>"000000000",
  20779=>"100100111",
  20780=>"000100000",
  20781=>"110100100",
  20782=>"010000111",
  20783=>"000000001",
  20784=>"010110110",
  20785=>"000111111",
  20786=>"100000000",
  20787=>"000000001",
  20788=>"111111110",
  20789=>"100100010",
  20790=>"000001011",
  20791=>"000001001",
  20792=>"100000000",
  20793=>"000000000",
  20794=>"000000000",
  20795=>"111111000",
  20796=>"111111111",
  20797=>"100000000",
  20798=>"111111111",
  20799=>"000010011",
  20800=>"000000000",
  20801=>"100001000",
  20802=>"111111111",
  20803=>"111111111",
  20804=>"111111111",
  20805=>"011001000",
  20806=>"100100100",
  20807=>"000011111",
  20808=>"000000000",
  20809=>"000100110",
  20810=>"111111111",
  20811=>"111111111",
  20812=>"001001000",
  20813=>"110000000",
  20814=>"000000000",
  20815=>"101111011",
  20816=>"001001001",
  20817=>"110110011",
  20818=>"111111111",
  20819=>"101101111",
  20820=>"101000000",
  20821=>"011011011",
  20822=>"000000000",
  20823=>"111011111",
  20824=>"000000000",
  20825=>"111111111",
  20826=>"111111111",
  20827=>"110100100",
  20828=>"111111111",
  20829=>"000000000",
  20830=>"000000000",
  20831=>"111111100",
  20832=>"100000000",
  20833=>"001001011",
  20834=>"110111111",
  20835=>"111110000",
  20836=>"000001111",
  20837=>"000000111",
  20838=>"000000111",
  20839=>"100100110",
  20840=>"111111111",
  20841=>"111000000",
  20842=>"101000000",
  20843=>"100000000",
  20844=>"011000000",
  20845=>"000010111",
  20846=>"000000000",
  20847=>"000000000",
  20848=>"011011111",
  20849=>"000000111",
  20850=>"111011001",
  20851=>"111001000",
  20852=>"010011001",
  20853=>"000000111",
  20854=>"000000001",
  20855=>"110100100",
  20856=>"111111111",
  20857=>"000000000",
  20858=>"111111111",
  20859=>"111110111",
  20860=>"000000111",
  20861=>"111111111",
  20862=>"010010111",
  20863=>"111111111",
  20864=>"111111000",
  20865=>"000000011",
  20866=>"000000000",
  20867=>"110000100",
  20868=>"000100110",
  20869=>"000100110",
  20870=>"001000000",
  20871=>"110110000",
  20872=>"100110000",
  20873=>"110111111",
  20874=>"111111110",
  20875=>"000000000",
  20876=>"101101111",
  20877=>"001110110",
  20878=>"011111010",
  20879=>"111111111",
  20880=>"001100000",
  20881=>"111000000",
  20882=>"000000000",
  20883=>"110110111",
  20884=>"000000000",
  20885=>"000010000",
  20886=>"111111111",
  20887=>"000000111",
  20888=>"111111111",
  20889=>"111111111",
  20890=>"000000000",
  20891=>"000111111",
  20892=>"111111111",
  20893=>"000000000",
  20894=>"001000000",
  20895=>"000000000",
  20896=>"011011000",
  20897=>"111111111",
  20898=>"110110110",
  20899=>"111101111",
  20900=>"110111111",
  20901=>"000111111",
  20902=>"000000000",
  20903=>"110000100",
  20904=>"000000000",
  20905=>"111100100",
  20906=>"001001111",
  20907=>"111111111",
  20908=>"000000000",
  20909=>"111111000",
  20910=>"111111000",
  20911=>"111111111",
  20912=>"000000000",
  20913=>"111111111",
  20914=>"000011000",
  20915=>"000001111",
  20916=>"101100000",
  20917=>"111111000",
  20918=>"110110110",
  20919=>"000000111",
  20920=>"100000000",
  20921=>"001000000",
  20922=>"011111111",
  20923=>"111111010",
  20924=>"100000000",
  20925=>"111111111",
  20926=>"000100000",
  20927=>"100110110",
  20928=>"000000000",
  20929=>"111100000",
  20930=>"000000000",
  20931=>"111100111",
  20932=>"111010111",
  20933=>"001011000",
  20934=>"000100111",
  20935=>"111111100",
  20936=>"011010000",
  20937=>"000000000",
  20938=>"010000000",
  20939=>"111100100",
  20940=>"000000011",
  20941=>"111111111",
  20942=>"000000000",
  20943=>"000000000",
  20944=>"000000000",
  20945=>"011111111",
  20946=>"111111011",
  20947=>"111111111",
  20948=>"001011111",
  20949=>"011110100",
  20950=>"000111111",
  20951=>"000000000",
  20952=>"111100101",
  20953=>"011111111",
  20954=>"001000011",
  20955=>"000000001",
  20956=>"000110111",
  20957=>"000000000",
  20958=>"111111111",
  20959=>"001000110",
  20960=>"000001000",
  20961=>"011000000",
  20962=>"000000111",
  20963=>"111111010",
  20964=>"000000000",
  20965=>"111111111",
  20966=>"000000001",
  20967=>"100100111",
  20968=>"000000000",
  20969=>"111001000",
  20970=>"010000001",
  20971=>"011000000",
  20972=>"011010000",
  20973=>"000001011",
  20974=>"000000000",
  20975=>"110000000",
  20976=>"000000101",
  20977=>"000000000",
  20978=>"111111111",
  20979=>"110010010",
  20980=>"111111111",
  20981=>"111111111",
  20982=>"000000000",
  20983=>"000000000",
  20984=>"000000000",
  20985=>"000100011",
  20986=>"001000100",
  20987=>"000000000",
  20988=>"000000000",
  20989=>"111111111",
  20990=>"001000000",
  20991=>"101111101",
  20992=>"100110110",
  20993=>"110000000",
  20994=>"000000100",
  20995=>"011111000",
  20996=>"000000000",
  20997=>"011111110",
  20998=>"001000000",
  20999=>"111111111",
  21000=>"111111000",
  21001=>"011000000",
  21002=>"100001001",
  21003=>"100000000",
  21004=>"001001001",
  21005=>"001010000",
  21006=>"000000110",
  21007=>"001111111",
  21008=>"110000111",
  21009=>"000010100",
  21010=>"111111111",
  21011=>"100100000",
  21012=>"000000000",
  21013=>"101000001",
  21014=>"011011111",
  21015=>"101100100",
  21016=>"101011000",
  21017=>"111111011",
  21018=>"000000000",
  21019=>"001011000",
  21020=>"111111011",
  21021=>"111111111",
  21022=>"111110110",
  21023=>"000000000",
  21024=>"000000111",
  21025=>"000110000",
  21026=>"111011001",
  21027=>"000110100",
  21028=>"000000000",
  21029=>"000000110",
  21030=>"010111111",
  21031=>"000111111",
  21032=>"001110000",
  21033=>"100000001",
  21034=>"000000100",
  21035=>"000010011",
  21036=>"001001101",
  21037=>"111101111",
  21038=>"011111111",
  21039=>"111110100",
  21040=>"001000000",
  21041=>"011010000",
  21042=>"101001101",
  21043=>"011001000",
  21044=>"111111111",
  21045=>"110100010",
  21046=>"001111010",
  21047=>"010010110",
  21048=>"111100000",
  21049=>"001001000",
  21050=>"001001011",
  21051=>"000000111",
  21052=>"111001001",
  21053=>"000000000",
  21054=>"001001011",
  21055=>"110111111",
  21056=>"111111111",
  21057=>"001011000",
  21058=>"111001001",
  21059=>"000000101",
  21060=>"110111011",
  21061=>"111111111",
  21062=>"000000111",
  21063=>"111111111",
  21064=>"101100100",
  21065=>"101001000",
  21066=>"101101111",
  21067=>"001000011",
  21068=>"000000000",
  21069=>"010010000",
  21070=>"001011011",
  21071=>"101001000",
  21072=>"000000000",
  21073=>"101111101",
  21074=>"111111111",
  21075=>"001101101",
  21076=>"011011010",
  21077=>"000000011",
  21078=>"010010000",
  21079=>"011001001",
  21080=>"000100110",
  21081=>"100100100",
  21082=>"111111111",
  21083=>"110110100",
  21084=>"111111111",
  21085=>"000000101",
  21086=>"010000101",
  21087=>"110110110",
  21088=>"001001000",
  21089=>"001011101",
  21090=>"000000000",
  21091=>"111100100",
  21092=>"100100000",
  21093=>"110111100",
  21094=>"011011000",
  21095=>"010011011",
  21096=>"000000000",
  21097=>"000001000",
  21098=>"000000000",
  21099=>"000000010",
  21100=>"111111111",
  21101=>"111111111",
  21102=>"111010010",
  21103=>"111111111",
  21104=>"011011010",
  21105=>"110110111",
  21106=>"110010100",
  21107=>"111000111",
  21108=>"011000000",
  21109=>"010010111",
  21110=>"000000000",
  21111=>"011011111",
  21112=>"001000001",
  21113=>"111011000",
  21114=>"010110000",
  21115=>"000000000",
  21116=>"110110110",
  21117=>"010111010",
  21118=>"110110011",
  21119=>"000000000",
  21120=>"000100100",
  21121=>"110010110",
  21122=>"000001001",
  21123=>"000010000",
  21124=>"111111000",
  21125=>"101101111",
  21126=>"110111111",
  21127=>"011111111",
  21128=>"000000101",
  21129=>"000100111",
  21130=>"000000000",
  21131=>"110000000",
  21132=>"000000000",
  21133=>"111011011",
  21134=>"001001000",
  21135=>"011000001",
  21136=>"000000000",
  21137=>"011000100",
  21138=>"110000011",
  21139=>"000000011",
  21140=>"011011011",
  21141=>"011010010",
  21142=>"100101111",
  21143=>"100100101",
  21144=>"001101101",
  21145=>"001101101",
  21146=>"111101011",
  21147=>"000000000",
  21148=>"001001111",
  21149=>"011000000",
  21150=>"011011011",
  21151=>"111101001",
  21152=>"000001101",
  21153=>"011111111",
  21154=>"011010000",
  21155=>"000011010",
  21156=>"010010110",
  21157=>"001011000",
  21158=>"000010000",
  21159=>"011011011",
  21160=>"000000000",
  21161=>"011011111",
  21162=>"100110110",
  21163=>"111000000",
  21164=>"100111111",
  21165=>"000110110",
  21166=>"100100111",
  21167=>"111111111",
  21168=>"000010000",
  21169=>"111111011",
  21170=>"010111011",
  21171=>"010001000",
  21172=>"011011001",
  21173=>"011011011",
  21174=>"010111111",
  21175=>"111111111",
  21176=>"001001111",
  21177=>"100111111",
  21178=>"011011011",
  21179=>"000010000",
  21180=>"000011111",
  21181=>"011000000",
  21182=>"111111101",
  21183=>"110111111",
  21184=>"000001101",
  21185=>"000010000",
  21186=>"000000111",
  21187=>"110111111",
  21188=>"111111111",
  21189=>"000001101",
  21190=>"110100010",
  21191=>"000000000",
  21192=>"111011011",
  21193=>"000010011",
  21194=>"000000000",
  21195=>"111110111",
  21196=>"001001001",
  21197=>"011001000",
  21198=>"000000000",
  21199=>"000000000",
  21200=>"001001000",
  21201=>"110010000",
  21202=>"000000011",
  21203=>"001100000",
  21204=>"111011011",
  21205=>"110111011",
  21206=>"000001101",
  21207=>"111111100",
  21208=>"111111111",
  21209=>"001101110",
  21210=>"100101101",
  21211=>"010011011",
  21212=>"111110010",
  21213=>"000100010",
  21214=>"000000000",
  21215=>"010011000",
  21216=>"000111110",
  21217=>"101000000",
  21218=>"100001011",
  21219=>"010111111",
  21220=>"011010010",
  21221=>"001011011",
  21222=>"111111111",
  21223=>"111111111",
  21224=>"000000000",
  21225=>"111111111",
  21226=>"011111111",
  21227=>"101101111",
  21228=>"011011111",
  21229=>"100100100",
  21230=>"111111110",
  21231=>"111100111",
  21232=>"111110010",
  21233=>"010000000",
  21234=>"000010011",
  21235=>"000100111",
  21236=>"110111111",
  21237=>"100000000",
  21238=>"001011001",
  21239=>"000000001",
  21240=>"111111101",
  21241=>"001000001",
  21242=>"000001011",
  21243=>"001001000",
  21244=>"011001001",
  21245=>"111101100",
  21246=>"010010000",
  21247=>"011111111",
  21248=>"011011001",
  21249=>"011001001",
  21250=>"000010010",
  21251=>"010000000",
  21252=>"010100100",
  21253=>"000000010",
  21254=>"101001101",
  21255=>"001011101",
  21256=>"010111111",
  21257=>"111111111",
  21258=>"000000101",
  21259=>"000110110",
  21260=>"101101101",
  21261=>"001001111",
  21262=>"000000110",
  21263=>"001001111",
  21264=>"011011000",
  21265=>"001111111",
  21266=>"011001001",
  21267=>"000000011",
  21268=>"011011011",
  21269=>"001000111",
  21270=>"111001001",
  21271=>"011110111",
  21272=>"110110110",
  21273=>"010010100",
  21274=>"110011011",
  21275=>"001000111",
  21276=>"110110100",
  21277=>"000011111",
  21278=>"000111011",
  21279=>"001010110",
  21280=>"111111111",
  21281=>"100100110",
  21282=>"100110111",
  21283=>"110100100",
  21284=>"000000000",
  21285=>"000011011",
  21286=>"111111111",
  21287=>"000111111",
  21288=>"000010010",
  21289=>"111011001",
  21290=>"001111010",
  21291=>"100100100",
  21292=>"011011011",
  21293=>"000111000",
  21294=>"000000010",
  21295=>"011011001",
  21296=>"000110111",
  21297=>"000000010",
  21298=>"000000000",
  21299=>"111100000",
  21300=>"000010111",
  21301=>"101011111",
  21302=>"011011101",
  21303=>"010110111",
  21304=>"111111110",
  21305=>"100000100",
  21306=>"011011011",
  21307=>"000000000",
  21308=>"010110111",
  21309=>"000010000",
  21310=>"010011000",
  21311=>"011000011",
  21312=>"000000000",
  21313=>"100110111",
  21314=>"000011010",
  21315=>"000000000",
  21316=>"111111111",
  21317=>"000110000",
  21318=>"110111011",
  21319=>"111000000",
  21320=>"001001101",
  21321=>"000000111",
  21322=>"011100110",
  21323=>"011011001",
  21324=>"000000011",
  21325=>"110010011",
  21326=>"000000001",
  21327=>"001001000",
  21328=>"011111011",
  21329=>"000000000",
  21330=>"000000101",
  21331=>"111001001",
  21332=>"110111111",
  21333=>"011011011",
  21334=>"011011000",
  21335=>"001000000",
  21336=>"111111110",
  21337=>"111111111",
  21338=>"011011011",
  21339=>"000100100",
  21340=>"000000100",
  21341=>"011001001",
  21342=>"111111111",
  21343=>"110110000",
  21344=>"111111111",
  21345=>"011011000",
  21346=>"011011111",
  21347=>"111100000",
  21348=>"110110110",
  21349=>"001001011",
  21350=>"111000000",
  21351=>"100000000",
  21352=>"000000110",
  21353=>"100000000",
  21354=>"001000001",
  21355=>"001011111",
  21356=>"111111111",
  21357=>"010111010",
  21358=>"111111111",
  21359=>"011111111",
  21360=>"011111111",
  21361=>"000111111",
  21362=>"110000111",
  21363=>"011001001",
  21364=>"011011000",
  21365=>"111110111",
  21366=>"011111010",
  21367=>"111111111",
  21368=>"111101101",
  21369=>"000010111",
  21370=>"100000000",
  21371=>"000001011",
  21372=>"000000000",
  21373=>"000000010",
  21374=>"011001000",
  21375=>"000000000",
  21376=>"110010010",
  21377=>"011111111",
  21378=>"011011001",
  21379=>"000000000",
  21380=>"001001001",
  21381=>"000000000",
  21382=>"110111011",
  21383=>"001100000",
  21384=>"001000000",
  21385=>"000100000",
  21386=>"010111111",
  21387=>"100100100",
  21388=>"000000000",
  21389=>"010000000",
  21390=>"011001000",
  21391=>"000000000",
  21392=>"000010010",
  21393=>"000000000",
  21394=>"111011001",
  21395=>"011001001",
  21396=>"000011111",
  21397=>"000011000",
  21398=>"000000000",
  21399=>"100110100",
  21400=>"000100110",
  21401=>"010011011",
  21402=>"000000001",
  21403=>"000101111",
  21404=>"100100100",
  21405=>"000100001",
  21406=>"110010011",
  21407=>"000101001",
  21408=>"010010010",
  21409=>"000000010",
  21410=>"000010000",
  21411=>"000000000",
  21412=>"111111000",
  21413=>"111111111",
  21414=>"111111111",
  21415=>"010010111",
  21416=>"000000000",
  21417=>"100100000",
  21418=>"000000000",
  21419=>"111000111",
  21420=>"000000000",
  21421=>"000000011",
  21422=>"000111010",
  21423=>"111111011",
  21424=>"111110110",
  21425=>"000001011",
  21426=>"111111111",
  21427=>"000000000",
  21428=>"110110111",
  21429=>"111110100",
  21430=>"110110100",
  21431=>"111110000",
  21432=>"001001000",
  21433=>"000110111",
  21434=>"000001001",
  21435=>"001011111",
  21436=>"111111111",
  21437=>"000000000",
  21438=>"111111111",
  21439=>"000010111",
  21440=>"111111111",
  21441=>"111111111",
  21442=>"111111111",
  21443=>"000000001",
  21444=>"110100000",
  21445=>"101101001",
  21446=>"000000000",
  21447=>"001001111",
  21448=>"000001101",
  21449=>"000011011",
  21450=>"011011001",
  21451=>"001101101",
  21452=>"111111000",
  21453=>"110110110",
  21454=>"010000001",
  21455=>"110011000",
  21456=>"110000000",
  21457=>"000001001",
  21458=>"110110010",
  21459=>"001111111",
  21460=>"011011001",
  21461=>"100110110",
  21462=>"001001000",
  21463=>"001001001",
  21464=>"010111111",
  21465=>"000011100",
  21466=>"001000010",
  21467=>"011010000",
  21468=>"000110110",
  21469=>"000100101",
  21470=>"111011111",
  21471=>"010000000",
  21472=>"101001100",
  21473=>"111111111",
  21474=>"000000000",
  21475=>"000111111",
  21476=>"010110000",
  21477=>"000000000",
  21478=>"001100100",
  21479=>"110111110",
  21480=>"011111011",
  21481=>"011011111",
  21482=>"100000110",
  21483=>"000000001",
  21484=>"000111111",
  21485=>"001001101",
  21486=>"100100110",
  21487=>"000011111",
  21488=>"011010000",
  21489=>"111111111",
  21490=>"000010100",
  21491=>"000000111",
  21492=>"100110110",
  21493=>"111010010",
  21494=>"000000111",
  21495=>"000000001",
  21496=>"111111110",
  21497=>"001101001",
  21498=>"011011111",
  21499=>"000000000",
  21500=>"000010001",
  21501=>"110111111",
  21502=>"110110110",
  21503=>"110110110",
  21504=>"111111111",
  21505=>"110110000",
  21506=>"000000111",
  21507=>"111111111",
  21508=>"111111111",
  21509=>"000000010",
  21510=>"111100100",
  21511=>"000000000",
  21512=>"011111111",
  21513=>"000000011",
  21514=>"000000000",
  21515=>"111100100",
  21516=>"110110110",
  21517=>"000000000",
  21518=>"000000000",
  21519=>"000000101",
  21520=>"000101001",
  21521=>"111111111",
  21522=>"111101101",
  21523=>"111101001",
  21524=>"001001001",
  21525=>"000011111",
  21526=>"000100111",
  21527=>"001000000",
  21528=>"111110010",
  21529=>"111111000",
  21530=>"001011001",
  21531=>"000100101",
  21532=>"111111111",
  21533=>"111101111",
  21534=>"111001011",
  21535=>"000111000",
  21536=>"111101101",
  21537=>"110110100",
  21538=>"111111111",
  21539=>"110111111",
  21540=>"111111000",
  21541=>"110011001",
  21542=>"000001000",
  21543=>"100111111",
  21544=>"000000000",
  21545=>"000000000",
  21546=>"111111111",
  21547=>"000000000",
  21548=>"000001001",
  21549=>"000001111",
  21550=>"000000000",
  21551=>"011000000",
  21552=>"010000000",
  21553=>"111111110",
  21554=>"001000100",
  21555=>"011111000",
  21556=>"110111111",
  21557=>"001010010",
  21558=>"100001001",
  21559=>"000111011",
  21560=>"111111111",
  21561=>"000000000",
  21562=>"000011111",
  21563=>"111001111",
  21564=>"111011000",
  21565=>"000100000",
  21566=>"110100000",
  21567=>"011011000",
  21568=>"011111111",
  21569=>"000000000",
  21570=>"011001000",
  21571=>"111111111",
  21572=>"011011011",
  21573=>"110100000",
  21574=>"000001101",
  21575=>"111111001",
  21576=>"001000011",
  21577=>"000000111",
  21578=>"000000000",
  21579=>"101111101",
  21580=>"001001000",
  21581=>"110000000",
  21582=>"111011111",
  21583=>"111111111",
  21584=>"000111011",
  21585=>"111111111",
  21586=>"111010110",
  21587=>"000010110",
  21588=>"000100111",
  21589=>"100110110",
  21590=>"000000001",
  21591=>"100100110",
  21592=>"000000000",
  21593=>"001000101",
  21594=>"011110110",
  21595=>"100000000",
  21596=>"000000000",
  21597=>"000000111",
  21598=>"111111111",
  21599=>"001000000",
  21600=>"110100000",
  21601=>"111111111",
  21602=>"100100111",
  21603=>"110100000",
  21604=>"101000000",
  21605=>"000000000",
  21606=>"000000111",
  21607=>"000000000",
  21608=>"000010111",
  21609=>"111111111",
  21610=>"001001111",
  21611=>"111111111",
  21612=>"010000000",
  21613=>"110110110",
  21614=>"000000000",
  21615=>"000000000",
  21616=>"111111111",
  21617=>"000000000",
  21618=>"011001000",
  21619=>"101111111",
  21620=>"111100101",
  21621=>"100101111",
  21622=>"111111110",
  21623=>"111000101",
  21624=>"000000100",
  21625=>"100111111",
  21626=>"000000000",
  21627=>"001000000",
  21628=>"001011011",
  21629=>"010111111",
  21630=>"000000000",
  21631=>"111111111",
  21632=>"000010000",
  21633=>"001001001",
  21634=>"011000000",
  21635=>"111111011",
  21636=>"110110111",
  21637=>"000000000",
  21638=>"000000000",
  21639=>"110000000",
  21640=>"011010011",
  21641=>"000000111",
  21642=>"010010000",
  21643=>"000000001",
  21644=>"111111111",
  21645=>"000000000",
  21646=>"111111110",
  21647=>"111111111",
  21648=>"000000000",
  21649=>"111111111",
  21650=>"000000000",
  21651=>"101111111",
  21652=>"000000000",
  21653=>"000000000",
  21654=>"100011011",
  21655=>"000000011",
  21656=>"100000101",
  21657=>"111111111",
  21658=>"000000000",
  21659=>"001001001",
  21660=>"011111111",
  21661=>"100101111",
  21662=>"111111111",
  21663=>"000000000",
  21664=>"111111011",
  21665=>"000001000",
  21666=>"000100000",
  21667=>"111111101",
  21668=>"100000000",
  21669=>"111111111",
  21670=>"101100000",
  21671=>"100100110",
  21672=>"000100000",
  21673=>"111111111",
  21674=>"000000000",
  21675=>"000000000",
  21676=>"011111111",
  21677=>"011111011",
  21678=>"111111110",
  21679=>"000000000",
  21680=>"110110111",
  21681=>"011101111",
  21682=>"111001000",
  21683=>"111111111",
  21684=>"100100100",
  21685=>"000000000",
  21686=>"111101000",
  21687=>"000000000",
  21688=>"000111111",
  21689=>"111111111",
  21690=>"111001100",
  21691=>"011111100",
  21692=>"000000000",
  21693=>"000000111",
  21694=>"000111111",
  21695=>"000000000",
  21696=>"000000000",
  21697=>"111111000",
  21698=>"111101111",
  21699=>"000000000",
  21700=>"001001111",
  21701=>"000000110",
  21702=>"000000111",
  21703=>"100001001",
  21704=>"110111111",
  21705=>"111000000",
  21706=>"001001001",
  21707=>"001011011",
  21708=>"001000000",
  21709=>"111111111",
  21710=>"111111001",
  21711=>"000000000",
  21712=>"110000011",
  21713=>"000000011",
  21714=>"001000100",
  21715=>"000000000",
  21716=>"111000000",
  21717=>"111111000",
  21718=>"000000000",
  21719=>"000001000",
  21720=>"011011011",
  21721=>"111110110",
  21722=>"111111111",
  21723=>"000111111",
  21724=>"000000000",
  21725=>"000000000",
  21726=>"000000000",
  21727=>"111111101",
  21728=>"000000000",
  21729=>"000000000",
  21730=>"000000000",
  21731=>"111111111",
  21732=>"001011111",
  21733=>"011011111",
  21734=>"010010011",
  21735=>"101001000",
  21736=>"000101111",
  21737=>"101001111",
  21738=>"111111111",
  21739=>"000000111",
  21740=>"111111111",
  21741=>"001001011",
  21742=>"111111111",
  21743=>"001011111",
  21744=>"110000000",
  21745=>"011011011",
  21746=>"100100011",
  21747=>"000000111",
  21748=>"110110110",
  21749=>"111000000",
  21750=>"000000000",
  21751=>"000100111",
  21752=>"000000000",
  21753=>"100000000",
  21754=>"000111000",
  21755=>"101000001",
  21756=>"111011001",
  21757=>"001011000",
  21758=>"011110110",
  21759=>"101101000",
  21760=>"000110011",
  21761=>"001000000",
  21762=>"111111111",
  21763=>"000000000",
  21764=>"000000000",
  21765=>"000000000",
  21766=>"111111111",
  21767=>"000000000",
  21768=>"110111001",
  21769=>"100100000",
  21770=>"000000001",
  21771=>"111111000",
  21772=>"000000000",
  21773=>"100011001",
  21774=>"000000100",
  21775=>"000000110",
  21776=>"001001101",
  21777=>"000100110",
  21778=>"000000000",
  21779=>"000000101",
  21780=>"101101111",
  21781=>"111100100",
  21782=>"110111111",
  21783=>"000000000",
  21784=>"000111111",
  21785=>"111111000",
  21786=>"000100101",
  21787=>"011001111",
  21788=>"000110000",
  21789=>"000000000",
  21790=>"000000000",
  21791=>"000000010",
  21792=>"111110110",
  21793=>"111111011",
  21794=>"011011000",
  21795=>"000000111",
  21796=>"001001111",
  21797=>"000100111",
  21798=>"111110110",
  21799=>"000000110",
  21800=>"111100101",
  21801=>"111111111",
  21802=>"000000000",
  21803=>"000000000",
  21804=>"000000000",
  21805=>"011011111",
  21806=>"101111111",
  21807=>"010010010",
  21808=>"111111111",
  21809=>"000001000",
  21810=>"001111111",
  21811=>"010010000",
  21812=>"111110000",
  21813=>"100110111",
  21814=>"110110100",
  21815=>"000100101",
  21816=>"111000000",
  21817=>"000000000",
  21818=>"001000100",
  21819=>"001001000",
  21820=>"000110110",
  21821=>"111111111",
  21822=>"110100000",
  21823=>"000000110",
  21824=>"000000000",
  21825=>"000101001",
  21826=>"111111111",
  21827=>"000000000",
  21828=>"001011000",
  21829=>"000000000",
  21830=>"111100000",
  21831=>"111111111",
  21832=>"000000000",
  21833=>"000000000",
  21834=>"000010111",
  21835=>"110110110",
  21836=>"000100110",
  21837=>"000000001",
  21838=>"000000000",
  21839=>"010110110",
  21840=>"001000110",
  21841=>"111111111",
  21842=>"111111111",
  21843=>"111000000",
  21844=>"000010000",
  21845=>"111110000",
  21846=>"111111111",
  21847=>"000000000",
  21848=>"000000000",
  21849=>"000000000",
  21850=>"111011110",
  21851=>"011111111",
  21852=>"000011001",
  21853=>"100000101",
  21854=>"010110111",
  21855=>"011011011",
  21856=>"000000000",
  21857=>"111100000",
  21858=>"110010011",
  21859=>"111111011",
  21860=>"000000001",
  21861=>"000111001",
  21862=>"000000000",
  21863=>"000000000",
  21864=>"111000000",
  21865=>"000110000",
  21866=>"101111111",
  21867=>"000000001",
  21868=>"000011001",
  21869=>"000111111",
  21870=>"011010000",
  21871=>"100100000",
  21872=>"111111111",
  21873=>"101000101",
  21874=>"000110111",
  21875=>"000011001",
  21876=>"100000000",
  21877=>"110100000",
  21878=>"011111001",
  21879=>"011010100",
  21880=>"111111111",
  21881=>"001001000",
  21882=>"111111001",
  21883=>"110110000",
  21884=>"111100100",
  21885=>"011111011",
  21886=>"101000000",
  21887=>"000010000",
  21888=>"000000000",
  21889=>"000111000",
  21890=>"111100001",
  21891=>"110100000",
  21892=>"011000110",
  21893=>"000010111",
  21894=>"111111111",
  21895=>"111110000",
  21896=>"101001101",
  21897=>"111111111",
  21898=>"001000000",
  21899=>"000000110",
  21900=>"000000000",
  21901=>"001000000",
  21902=>"000000011",
  21903=>"000011010",
  21904=>"001001000",
  21905=>"000001011",
  21906=>"000000100",
  21907=>"000000010",
  21908=>"111111111",
  21909=>"000000110",
  21910=>"000000000",
  21911=>"000110111",
  21912=>"110110110",
  21913=>"000000100",
  21914=>"111111111",
  21915=>"000101111",
  21916=>"010110100",
  21917=>"001001000",
  21918=>"011011001",
  21919=>"111111111",
  21920=>"111111111",
  21921=>"000000000",
  21922=>"000110111",
  21923=>"111111001",
  21924=>"000110111",
  21925=>"111011111",
  21926=>"100111111",
  21927=>"111111111",
  21928=>"000011011",
  21929=>"000110000",
  21930=>"111111111",
  21931=>"110111011",
  21932=>"001001001",
  21933=>"111000000",
  21934=>"001001100",
  21935=>"000000000",
  21936=>"001000000",
  21937=>"000000000",
  21938=>"111111111",
  21939=>"000000000",
  21940=>"001111111",
  21941=>"101101001",
  21942=>"110100100",
  21943=>"000010000",
  21944=>"000000001",
  21945=>"111011000",
  21946=>"111000000",
  21947=>"101101101",
  21948=>"011000000",
  21949=>"000000110",
  21950=>"000000000",
  21951=>"001011011",
  21952=>"001001011",
  21953=>"010111111",
  21954=>"010110110",
  21955=>"111111011",
  21956=>"011011001",
  21957=>"011001000",
  21958=>"000100111",
  21959=>"001111111",
  21960=>"111101000",
  21961=>"111111011",
  21962=>"001011011",
  21963=>"000100111",
  21964=>"000000000",
  21965=>"111001000",
  21966=>"000000000",
  21967=>"111111111",
  21968=>"111011011",
  21969=>"101111111",
  21970=>"000100100",
  21971=>"111111111",
  21972=>"000100001",
  21973=>"111111111",
  21974=>"011011011",
  21975=>"110111011",
  21976=>"000000000",
  21977=>"100101111",
  21978=>"111111111",
  21979=>"111111111",
  21980=>"011011011",
  21981=>"111111111",
  21982=>"110000001",
  21983=>"101101101",
  21984=>"111111111",
  21985=>"100111111",
  21986=>"111111011",
  21987=>"000000001",
  21988=>"000000000",
  21989=>"000111000",
  21990=>"000000111",
  21991=>"011000000",
  21992=>"111111111",
  21993=>"000010000",
  21994=>"000000001",
  21995=>"111100101",
  21996=>"000000000",
  21997=>"110110110",
  21998=>"011111011",
  21999=>"000000000",
  22000=>"111111110",
  22001=>"000000001",
  22002=>"111110100",
  22003=>"000000011",
  22004=>"000000000",
  22005=>"010111111",
  22006=>"100100000",
  22007=>"111111011",
  22008=>"010010011",
  22009=>"000110110",
  22010=>"111100000",
  22011=>"001001001",
  22012=>"111111111",
  22013=>"001001101",
  22014=>"000001000",
  22015=>"000010000",
  22016=>"011011011",
  22017=>"000000000",
  22018=>"000000111",
  22019=>"000111111",
  22020=>"000111111",
  22021=>"111111100",
  22022=>"111111111",
  22023=>"111111111",
  22024=>"000000000",
  22025=>"011011000",
  22026=>"111110000",
  22027=>"101101111",
  22028=>"001110110",
  22029=>"001001111",
  22030=>"011111111",
  22031=>"000001001",
  22032=>"111000000",
  22033=>"000100111",
  22034=>"111100100",
  22035=>"000100111",
  22036=>"000001101",
  22037=>"001000000",
  22038=>"000000000",
  22039=>"110100100",
  22040=>"000001111",
  22041=>"100110111",
  22042=>"101001011",
  22043=>"000000000",
  22044=>"000110111",
  22045=>"011111000",
  22046=>"000000000",
  22047=>"101000000",
  22048=>"001001000",
  22049=>"100110110",
  22050=>"111110000",
  22051=>"000000001",
  22052=>"000000000",
  22053=>"111011111",
  22054=>"111111111",
  22055=>"111111111",
  22056=>"111111111",
  22057=>"110000111",
  22058=>"111111111",
  22059=>"100000000",
  22060=>"110000000",
  22061=>"101111111",
  22062=>"000011011",
  22063=>"111110100",
  22064=>"111111111",
  22065=>"111111111",
  22066=>"000000001",
  22067=>"110111111",
  22068=>"000000000",
  22069=>"000110111",
  22070=>"111000000",
  22071=>"111111111",
  22072=>"011111110",
  22073=>"111110111",
  22074=>"111111111",
  22075=>"000000000",
  22076=>"001000111",
  22077=>"010011100",
  22078=>"111111111",
  22079=>"000000000",
  22080=>"111110111",
  22081=>"110000000",
  22082=>"111111101",
  22083=>"110100101",
  22084=>"011000010",
  22085=>"001001001",
  22086=>"111010000",
  22087=>"110111111",
  22088=>"111011011",
  22089=>"111101000",
  22090=>"000000011",
  22091=>"000000000",
  22092=>"111111111",
  22093=>"001000011",
  22094=>"111000000",
  22095=>"111000000",
  22096=>"011111111",
  22097=>"111000000",
  22098=>"001111000",
  22099=>"000000000",
  22100=>"111111011",
  22101=>"000000001",
  22102=>"000110111",
  22103=>"000000000",
  22104=>"011111111",
  22105=>"111000000",
  22106=>"000000000",
  22107=>"110010010",
  22108=>"000000000",
  22109=>"110000110",
  22110=>"000000001",
  22111=>"111011111",
  22112=>"000001000",
  22113=>"111101111",
  22114=>"001000000",
  22115=>"000000000",
  22116=>"010111110",
  22117=>"000001001",
  22118=>"111111111",
  22119=>"000000000",
  22120=>"111111100",
  22121=>"000000000",
  22122=>"100100000",
  22123=>"101000111",
  22124=>"000000000",
  22125=>"111100110",
  22126=>"111111011",
  22127=>"000000000",
  22128=>"101101111",
  22129=>"000000000",
  22130=>"010000000",
  22131=>"011001111",
  22132=>"011000000",
  22133=>"010001000",
  22134=>"111111100",
  22135=>"110000000",
  22136=>"111001101",
  22137=>"111111111",
  22138=>"000000000",
  22139=>"000000001",
  22140=>"110110110",
  22141=>"001101111",
  22142=>"000000000",
  22143=>"111001000",
  22144=>"111111111",
  22145=>"111111111",
  22146=>"000000000",
  22147=>"000110101",
  22148=>"000010111",
  22149=>"000100101",
  22150=>"111111111",
  22151=>"000000000",
  22152=>"101101001",
  22153=>"000000010",
  22154=>"000000000",
  22155=>"000000110",
  22156=>"011000000",
  22157=>"111010110",
  22158=>"110010111",
  22159=>"000000100",
  22160=>"111001000",
  22161=>"000000000",
  22162=>"011111111",
  22163=>"001001001",
  22164=>"000000001",
  22165=>"111111111",
  22166=>"100111111",
  22167=>"000000000",
  22168=>"000000000",
  22169=>"101111111",
  22170=>"000000110",
  22171=>"001001001",
  22172=>"000100110",
  22173=>"000001000",
  22174=>"000000001",
  22175=>"011111001",
  22176=>"101111111",
  22177=>"111111111",
  22178=>"111111110",
  22179=>"000000000",
  22180=>"000100110",
  22181=>"100111111",
  22182=>"111111111",
  22183=>"010111111",
  22184=>"011000110",
  22185=>"111111111",
  22186=>"111111111",
  22187=>"000000111",
  22188=>"111111111",
  22189=>"000110110",
  22190=>"000110110",
  22191=>"000000000",
  22192=>"011111000",
  22193=>"011010011",
  22194=>"111101000",
  22195=>"000000000",
  22196=>"100100111",
  22197=>"011000000",
  22198=>"111111111",
  22199=>"000111111",
  22200=>"100111111",
  22201=>"111111111",
  22202=>"000000000",
  22203=>"000110010",
  22204=>"000010111",
  22205=>"111110001",
  22206=>"011011011",
  22207=>"111111110",
  22208=>"000000000",
  22209=>"100110110",
  22210=>"001101101",
  22211=>"000000000",
  22212=>"000001000",
  22213=>"000000000",
  22214=>"000000110",
  22215=>"000110000",
  22216=>"101000000",
  22217=>"000000000",
  22218=>"001001111",
  22219=>"000010111",
  22220=>"000001111",
  22221=>"001000010",
  22222=>"100000001",
  22223=>"000000000",
  22224=>"011000000",
  22225=>"100100100",
  22226=>"000111100",
  22227=>"000000001",
  22228=>"001000000",
  22229=>"110111111",
  22230=>"000000000",
  22231=>"011000001",
  22232=>"010011000",
  22233=>"110110010",
  22234=>"000000000",
  22235=>"000000000",
  22236=>"000000001",
  22237=>"000000000",
  22238=>"111111111",
  22239=>"000110111",
  22240=>"000000000",
  22241=>"000110111",
  22242=>"000000100",
  22243=>"010100000",
  22244=>"111101101",
  22245=>"110110100",
  22246=>"111111000",
  22247=>"000000000",
  22248=>"000111000",
  22249=>"000000001",
  22250=>"000000000",
  22251=>"000000000",
  22252=>"011111111",
  22253=>"000000000",
  22254=>"000000111",
  22255=>"111110010",
  22256=>"110111111",
  22257=>"111111110",
  22258=>"110010000",
  22259=>"000000110",
  22260=>"000110000",
  22261=>"000000000",
  22262=>"011000001",
  22263=>"111111111",
  22264=>"110110111",
  22265=>"110111111",
  22266=>"000000000",
  22267=>"110110110",
  22268=>"001000000",
  22269=>"010111001",
  22270=>"000000101",
  22271=>"111000000",
  22272=>"000000000",
  22273=>"000000000",
  22274=>"000000001",
  22275=>"000000000",
  22276=>"000000000",
  22277=>"000000100",
  22278=>"000011111",
  22279=>"100101000",
  22280=>"001010000",
  22281=>"000000000",
  22282=>"001001101",
  22283=>"000000001",
  22284=>"000000000",
  22285=>"000000000",
  22286=>"001000000",
  22287=>"111000000",
  22288=>"000100111",
  22289=>"111111111",
  22290=>"111101101",
  22291=>"111111111",
  22292=>"111111111",
  22293=>"000000000",
  22294=>"110110000",
  22295=>"111011000",
  22296=>"000000101",
  22297=>"000000111",
  22298=>"111100101",
  22299=>"000001000",
  22300=>"111111110",
  22301=>"000011001",
  22302=>"100000000",
  22303=>"011001101",
  22304=>"010110000",
  22305=>"111111111",
  22306=>"000010011",
  22307=>"001001001",
  22308=>"000000000",
  22309=>"100000110",
  22310=>"110000000",
  22311=>"000111000",
  22312=>"000000000",
  22313=>"111111110",
  22314=>"000000000",
  22315=>"111011000",
  22316=>"111000000",
  22317=>"000111111",
  22318=>"000000000",
  22319=>"001000000",
  22320=>"110110111",
  22321=>"000000000",
  22322=>"000000000",
  22323=>"111000000",
  22324=>"111100100",
  22325=>"001011000",
  22326=>"100011111",
  22327=>"000000000",
  22328=>"100000000",
  22329=>"100100111",
  22330=>"000111111",
  22331=>"111110111",
  22332=>"000000001",
  22333=>"000110100",
  22334=>"000100110",
  22335=>"111111000",
  22336=>"111111111",
  22337=>"000000000",
  22338=>"111111110",
  22339=>"111111111",
  22340=>"111111010",
  22341=>"000111111",
  22342=>"111000000",
  22343=>"000000000",
  22344=>"000000000",
  22345=>"100000000",
  22346=>"001111111",
  22347=>"111011011",
  22348=>"101100010",
  22349=>"100000000",
  22350=>"001110000",
  22351=>"010000100",
  22352=>"001001111",
  22353=>"000000111",
  22354=>"000000000",
  22355=>"000000000",
  22356=>"000000000",
  22357=>"001011011",
  22358=>"000000100",
  22359=>"100111111",
  22360=>"111111111",
  22361=>"000000000",
  22362=>"000110000",
  22363=>"000000000",
  22364=>"000000001",
  22365=>"111001111",
  22366=>"111000000",
  22367=>"000000000",
  22368=>"111111111",
  22369=>"111111111",
  22370=>"011011011",
  22371=>"000000000",
  22372=>"001001001",
  22373=>"010111111",
  22374=>"000000111",
  22375=>"011110111",
  22376=>"110110111",
  22377=>"100000000",
  22378=>"011111011",
  22379=>"111111111",
  22380=>"110110110",
  22381=>"111110110",
  22382=>"111111111",
  22383=>"000111011",
  22384=>"000000000",
  22385=>"000100100",
  22386=>"011011001",
  22387=>"000010000",
  22388=>"000011001",
  22389=>"110010000",
  22390=>"010111110",
  22391=>"000000000",
  22392=>"000000111",
  22393=>"100000101",
  22394=>"110110111",
  22395=>"011010000",
  22396=>"111100000",
  22397=>"000000000",
  22398=>"111101101",
  22399=>"000000000",
  22400=>"000000110",
  22401=>"111110111",
  22402=>"000100101",
  22403=>"111111111",
  22404=>"111111111",
  22405=>"111111011",
  22406=>"111111111",
  22407=>"111111111",
  22408=>"111111111",
  22409=>"111111111",
  22410=>"011110110",
  22411=>"111110000",
  22412=>"100000001",
  22413=>"001011011",
  22414=>"111111011",
  22415=>"111111111",
  22416=>"000000000",
  22417=>"111111111",
  22418=>"101000001",
  22419=>"000000100",
  22420=>"000000000",
  22421=>"000001000",
  22422=>"000001000",
  22423=>"110100000",
  22424=>"111111111",
  22425=>"111000010",
  22426=>"001000000",
  22427=>"011111000",
  22428=>"011111111",
  22429=>"000000000",
  22430=>"000000000",
  22431=>"100000000",
  22432=>"000100100",
  22433=>"001000000",
  22434=>"000000001",
  22435=>"111111111",
  22436=>"111111111",
  22437=>"000000000",
  22438=>"110000000",
  22439=>"000100000",
  22440=>"000000000",
  22441=>"000000001",
  22442=>"111111111",
  22443=>"000000000",
  22444=>"000000000",
  22445=>"001000100",
  22446=>"000111111",
  22447=>"000000000",
  22448=>"111111111",
  22449=>"110111001",
  22450=>"000000000",
  22451=>"000000000",
  22452=>"100111001",
  22453=>"000010111",
  22454=>"111111111",
  22455=>"111111110",
  22456=>"000000001",
  22457=>"000011011",
  22458=>"111011101",
  22459=>"111111111",
  22460=>"110110111",
  22461=>"111001100",
  22462=>"001001011",
  22463=>"000000000",
  22464=>"000111111",
  22465=>"000000000",
  22466=>"000000001",
  22467=>"000011011",
  22468=>"110110101",
  22469=>"000010011",
  22470=>"100000000",
  22471=>"000000011",
  22472=>"000010110",
  22473=>"111111110",
  22474=>"111101101",
  22475=>"111111111",
  22476=>"010100010",
  22477=>"000000001",
  22478=>"000000000",
  22479=>"000111011",
  22480=>"000000010",
  22481=>"000010011",
  22482=>"100110110",
  22483=>"000000000",
  22484=>"111111111",
  22485=>"000010100",
  22486=>"001000000",
  22487=>"000000000",
  22488=>"000000000",
  22489=>"111001000",
  22490=>"111000000",
  22491=>"110110000",
  22492=>"111111111",
  22493=>"001001001",
  22494=>"110110000",
  22495=>"000000000",
  22496=>"111110110",
  22497=>"000000111",
  22498=>"111110110",
  22499=>"111111111",
  22500=>"111110111",
  22501=>"011010000",
  22502=>"000000000",
  22503=>"000000000",
  22504=>"111111111",
  22505=>"111111111",
  22506=>"011000000",
  22507=>"000111111",
  22508=>"000000000",
  22509=>"000001001",
  22510=>"000000000",
  22511=>"001000000",
  22512=>"000000000",
  22513=>"011111000",
  22514=>"111111111",
  22515=>"011111000",
  22516=>"000100111",
  22517=>"111111011",
  22518=>"110110100",
  22519=>"000100100",
  22520=>"111111111",
  22521=>"000010110",
  22522=>"111100000",
  22523=>"110000000",
  22524=>"111111111",
  22525=>"111110011",
  22526=>"111111110",
  22527=>"111110110",
  22528=>"001011111",
  22529=>"111001001",
  22530=>"101101111",
  22531=>"111111111",
  22532=>"000000000",
  22533=>"000000000",
  22534=>"000111111",
  22535=>"111111111",
  22536=>"111001100",
  22537=>"000000000",
  22538=>"000000100",
  22539=>"000000101",
  22540=>"000000000",
  22541=>"010000000",
  22542=>"111110011",
  22543=>"000000011",
  22544=>"000000000",
  22545=>"000111011",
  22546=>"000110000",
  22547=>"001000001",
  22548=>"111111111",
  22549=>"000000000",
  22550=>"001000000",
  22551=>"001011000",
  22552=>"111111001",
  22553=>"011111110",
  22554=>"000000000",
  22555=>"000000000",
  22556=>"000000000",
  22557=>"101111110",
  22558=>"111111100",
  22559=>"111111111",
  22560=>"001101111",
  22561=>"110111101",
  22562=>"000000000",
  22563=>"111111110",
  22564=>"000000000",
  22565=>"001000000",
  22566=>"001000000",
  22567=>"111111111",
  22568=>"000000000",
  22569=>"000000000",
  22570=>"111111111",
  22571=>"111111111",
  22572=>"001001000",
  22573=>"111111111",
  22574=>"000000100",
  22575=>"001000000",
  22576=>"000110110",
  22577=>"010110000",
  22578=>"000110110",
  22579=>"111111001",
  22580=>"000001001",
  22581=>"100000100",
  22582=>"101100111",
  22583=>"100100111",
  22584=>"111011001",
  22585=>"101000001",
  22586=>"000000000",
  22587=>"000110111",
  22588=>"111111111",
  22589=>"111111111",
  22590=>"000001111",
  22591=>"000000011",
  22592=>"000001111",
  22593=>"111011000",
  22594=>"000010000",
  22595=>"111000000",
  22596=>"000001111",
  22597=>"000000000",
  22598=>"000000000",
  22599=>"000000100",
  22600=>"111111110",
  22601=>"100111111",
  22602=>"111111111",
  22603=>"001000111",
  22604=>"001111111",
  22605=>"000100111",
  22606=>"011000000",
  22607=>"000000000",
  22608=>"111111011",
  22609=>"000100100",
  22610=>"100000001",
  22611=>"000000000",
  22612=>"111111111",
  22613=>"000000000",
  22614=>"111111111",
  22615=>"101101000",
  22616=>"000000001",
  22617=>"000000000",
  22618=>"000000101",
  22619=>"110110111",
  22620=>"111101101",
  22621=>"111111111",
  22622=>"001111000",
  22623=>"111111111",
  22624=>"100000000",
  22625=>"111100101",
  22626=>"111111111",
  22627=>"000000100",
  22628=>"100000000",
  22629=>"111111111",
  22630=>"111111001",
  22631=>"000000000",
  22632=>"000000000",
  22633=>"111111110",
  22634=>"111111111",
  22635=>"110111001",
  22636=>"000010111",
  22637=>"111000000",
  22638=>"000000000",
  22639=>"000110000",
  22640=>"111101111",
  22641=>"001001111",
  22642=>"111110111",
  22643=>"000000000",
  22644=>"111111111",
  22645=>"111111111",
  22646=>"111111110",
  22647=>"000000000",
  22648=>"000000000",
  22649=>"000000000",
  22650=>"111110100",
  22651=>"111000000",
  22652=>"110110110",
  22653=>"111111000",
  22654=>"100000000",
  22655=>"000000000",
  22656=>"111000000",
  22657=>"011001000",
  22658=>"111111110",
  22659=>"000000000",
  22660=>"111111111",
  22661=>"111000000",
  22662=>"000000100",
  22663=>"100111111",
  22664=>"000011110",
  22665=>"000000000",
  22666=>"111111011",
  22667=>"000000000",
  22668=>"001100110",
  22669=>"100000000",
  22670=>"100100111",
  22671=>"011011001",
  22672=>"111111111",
  22673=>"101001001",
  22674=>"001000001",
  22675=>"100100100",
  22676=>"101001000",
  22677=>"000000000",
  22678=>"000000001",
  22679=>"111111011",
  22680=>"001001001",
  22681=>"111111100",
  22682=>"000000000",
  22683=>"111111111",
  22684=>"000001111",
  22685=>"011001111",
  22686=>"111111111",
  22687=>"111111111",
  22688=>"000100100",
  22689=>"000000000",
  22690=>"111111111",
  22691=>"000010110",
  22692=>"000000101",
  22693=>"000000000",
  22694=>"111111100",
  22695=>"000000011",
  22696=>"111101111",
  22697=>"000000010",
  22698=>"111111110",
  22699=>"000000000",
  22700=>"000000000",
  22701=>"000000000",
  22702=>"000000001",
  22703=>"111111111",
  22704=>"111110111",
  22705=>"110110010",
  22706=>"111111111",
  22707=>"100111100",
  22708=>"000000000",
  22709=>"000000000",
  22710=>"000000000",
  22711=>"111111111",
  22712=>"100100110",
  22713=>"000000100",
  22714=>"001000000",
  22715=>"111101111",
  22716=>"000000110",
  22717=>"111111110",
  22718=>"000000000",
  22719=>"111111111",
  22720=>"000000000",
  22721=>"111111111",
  22722=>"111111111",
  22723=>"111111111",
  22724=>"111111111",
  22725=>"111111111",
  22726=>"111111111",
  22727=>"101111111",
  22728=>"000000000",
  22729=>"000100001",
  22730=>"000110110",
  22731=>"000000000",
  22732=>"111111111",
  22733=>"000100000",
  22734=>"101111111",
  22735=>"000000000",
  22736=>"011111010",
  22737=>"000100111",
  22738=>"010000000",
  22739=>"000010111",
  22740=>"000000000",
  22741=>"110000000",
  22742=>"000001000",
  22743=>"011010000",
  22744=>"111111111",
  22745=>"111101100",
  22746=>"000000000",
  22747=>"000000000",
  22748=>"111111111",
  22749=>"100100101",
  22750=>"011001000",
  22751=>"100100000",
  22752=>"000000000",
  22753=>"010111111",
  22754=>"111111111",
  22755=>"111111111",
  22756=>"000000000",
  22757=>"111111100",
  22758=>"111111111",
  22759=>"001001000",
  22760=>"000000111",
  22761=>"000111111",
  22762=>"111111111",
  22763=>"000000000",
  22764=>"000000000",
  22765=>"000000000",
  22766=>"000000000",
  22767=>"000000000",
  22768=>"111100000",
  22769=>"111111111",
  22770=>"111111111",
  22771=>"000000100",
  22772=>"111011000",
  22773=>"111111111",
  22774=>"000000000",
  22775=>"000000000",
  22776=>"111111100",
  22777=>"101111111",
  22778=>"000000000",
  22779=>"001000000",
  22780=>"111111111",
  22781=>"001001000",
  22782=>"110111111",
  22783=>"110111111",
  22784=>"000000000",
  22785=>"111111111",
  22786=>"000000000",
  22787=>"011011001",
  22788=>"111111000",
  22789=>"111111000",
  22790=>"000000000",
  22791=>"101101111",
  22792=>"000001000",
  22793=>"000000000",
  22794=>"000000000",
  22795=>"000000000",
  22796=>"111101111",
  22797=>"000110111",
  22798=>"110100000",
  22799=>"000000000",
  22800=>"000000000",
  22801=>"101001000",
  22802=>"000000000",
  22803=>"000100101",
  22804=>"000000000",
  22805=>"101001111",
  22806=>"110110110",
  22807=>"000000000",
  22808=>"111111111",
  22809=>"111111111",
  22810=>"000000000",
  22811=>"000000000",
  22812=>"000001001",
  22813=>"000000000",
  22814=>"110111110",
  22815=>"111000111",
  22816=>"000000000",
  22817=>"000000101",
  22818=>"000000000",
  22819=>"000000000",
  22820=>"000110011",
  22821=>"111111111",
  22822=>"111000000",
  22823=>"001001111",
  22824=>"110000011",
  22825=>"000000000",
  22826=>"111111111",
  22827=>"111111111",
  22828=>"110111110",
  22829=>"111111000",
  22830=>"111111111",
  22831=>"000000000",
  22832=>"000000000",
  22833=>"001000000",
  22834=>"000000010",
  22835=>"111111000",
  22836=>"101000101",
  22837=>"111111111",
  22838=>"110101111",
  22839=>"111111110",
  22840=>"111111110",
  22841=>"111111000",
  22842=>"000111111",
  22843=>"000000110",
  22844=>"000000000",
  22845=>"000100111",
  22846=>"001111111",
  22847=>"011001000",
  22848=>"111111000",
  22849=>"101111101",
  22850=>"100111111",
  22851=>"100100100",
  22852=>"110111110",
  22853=>"110110010",
  22854=>"000000000",
  22855=>"000000000",
  22856=>"111111110",
  22857=>"000010000",
  22858=>"000000000",
  22859=>"101111111",
  22860=>"000000000",
  22861=>"011000000",
  22862=>"000000000",
  22863=>"100000000",
  22864=>"000111111",
  22865=>"000000000",
  22866=>"101000000",
  22867=>"000000001",
  22868=>"000111111",
  22869=>"011011011",
  22870=>"111111111",
  22871=>"110100100",
  22872=>"110111111",
  22873=>"000000000",
  22874=>"000000000",
  22875=>"111111001",
  22876=>"111111111",
  22877=>"111111011",
  22878=>"000000001",
  22879=>"100111100",
  22880=>"111111111",
  22881=>"111000000",
  22882=>"011000000",
  22883=>"111111111",
  22884=>"111111100",
  22885=>"001011011",
  22886=>"000000001",
  22887=>"000000000",
  22888=>"000000100",
  22889=>"111111111",
  22890=>"110110111",
  22891=>"000000101",
  22892=>"000000000",
  22893=>"111001000",
  22894=>"000000000",
  22895=>"110111111",
  22896=>"000000000",
  22897=>"000010000",
  22898=>"000000000",
  22899=>"000000000",
  22900=>"000110000",
  22901=>"111111111",
  22902=>"000000101",
  22903=>"000000111",
  22904=>"000000000",
  22905=>"000011111",
  22906=>"000000000",
  22907=>"001011011",
  22908=>"000110111",
  22909=>"111111111",
  22910=>"000000000",
  22911=>"000000000",
  22912=>"011001000",
  22913=>"000000011",
  22914=>"000000000",
  22915=>"111111111",
  22916=>"000110000",
  22917=>"111111000",
  22918=>"000101111",
  22919=>"000000000",
  22920=>"000000000",
  22921=>"111110100",
  22922=>"100100100",
  22923=>"111111111",
  22924=>"111101101",
  22925=>"111111111",
  22926=>"100001001",
  22927=>"110100000",
  22928=>"011111111",
  22929=>"000000000",
  22930=>"000001001",
  22931=>"000000000",
  22932=>"000000011",
  22933=>"000000000",
  22934=>"111111000",
  22935=>"000000001",
  22936=>"000000000",
  22937=>"111111110",
  22938=>"110000000",
  22939=>"111111111",
  22940=>"000000000",
  22941=>"001101111",
  22942=>"000000000",
  22943=>"000000000",
  22944=>"000110010",
  22945=>"000000111",
  22946=>"111100000",
  22947=>"111111111",
  22948=>"111111000",
  22949=>"000000000",
  22950=>"111111111",
  22951=>"000110111",
  22952=>"000110110",
  22953=>"111100100",
  22954=>"000000000",
  22955=>"111000000",
  22956=>"000000010",
  22957=>"111111110",
  22958=>"000100111",
  22959=>"000000011",
  22960=>"111100111",
  22961=>"111000000",
  22962=>"111111011",
  22963=>"000000000",
  22964=>"000000101",
  22965=>"111000000",
  22966=>"100111111",
  22967=>"000111111",
  22968=>"101001001",
  22969=>"001101111",
  22970=>"100110011",
  22971=>"110110001",
  22972=>"000000000",
  22973=>"111111001",
  22974=>"111111111",
  22975=>"111111011",
  22976=>"000000000",
  22977=>"000000000",
  22978=>"011001111",
  22979=>"000000000",
  22980=>"101001111",
  22981=>"000111100",
  22982=>"101001101",
  22983=>"111000000",
  22984=>"000000000",
  22985=>"100110000",
  22986=>"000000000",
  22987=>"010010000",
  22988=>"000000000",
  22989=>"111111111",
  22990=>"111101101",
  22991=>"111111111",
  22992=>"000010011",
  22993=>"110100111",
  22994=>"111111111",
  22995=>"110110000",
  22996=>"110110011",
  22997=>"101111111",
  22998=>"101111111",
  22999=>"100111001",
  23000=>"100000001",
  23001=>"000110111",
  23002=>"001001011",
  23003=>"111111111",
  23004=>"110111111",
  23005=>"111111111",
  23006=>"100110111",
  23007=>"011111011",
  23008=>"001001101",
  23009=>"000100000",
  23010=>"111111101",
  23011=>"111111111",
  23012=>"110111000",
  23013=>"111111111",
  23014=>"111000000",
  23015=>"111111111",
  23016=>"001000000",
  23017=>"101011000",
  23018=>"111000000",
  23019=>"111111100",
  23020=>"111011101",
  23021=>"000000000",
  23022=>"101101101",
  23023=>"000100001",
  23024=>"000000000",
  23025=>"001000100",
  23026=>"001001001",
  23027=>"111111111",
  23028=>"000100000",
  23029=>"000000000",
  23030=>"000000110",
  23031=>"001111000",
  23032=>"100100100",
  23033=>"001001001",
  23034=>"110111000",
  23035=>"111111111",
  23036=>"011000110",
  23037=>"111001111",
  23038=>"001011011",
  23039=>"000000000",
  23040=>"000000100",
  23041=>"000000000",
  23042=>"101101000",
  23043=>"000101111",
  23044=>"110111110",
  23045=>"000000001",
  23046=>"000000111",
  23047=>"101101100",
  23048=>"011001001",
  23049=>"000000111",
  23050=>"000000000",
  23051=>"000000011",
  23052=>"000000010",
  23053=>"001001111",
  23054=>"100111011",
  23055=>"111100111",
  23056=>"000000110",
  23057=>"011111111",
  23058=>"100110110",
  23059=>"000000000",
  23060=>"111111111",
  23061=>"000000000",
  23062=>"111111100",
  23063=>"110110111",
  23064=>"000000010",
  23065=>"000000111",
  23066=>"111000001",
  23067=>"111111010",
  23068=>"000111111",
  23069=>"111111110",
  23070=>"101000000",
  23071=>"000111111",
  23072=>"000100101",
  23073=>"110111111",
  23074=>"111110111",
  23075=>"110011000",
  23076=>"100000000",
  23077=>"001111011",
  23078=>"000000111",
  23079=>"000010000",
  23080=>"100000000",
  23081=>"101000000",
  23082=>"000101111",
  23083=>"111111000",
  23084=>"111000111",
  23085=>"100100000",
  23086=>"000110100",
  23087=>"111111111",
  23088=>"000001111",
  23089=>"000110111",
  23090=>"100000111",
  23091=>"111001111",
  23092=>"111111011",
  23093=>"110111111",
  23094=>"100100100",
  23095=>"000011111",
  23096=>"000000110",
  23097=>"110000000",
  23098=>"000000001",
  23099=>"111111111",
  23100=>"001011111",
  23101=>"111000000",
  23102=>"111111000",
  23103=>"111100000",
  23104=>"111111111",
  23105=>"011000000",
  23106=>"111111000",
  23107=>"111000000",
  23108=>"001001011",
  23109=>"100000000",
  23110=>"101001000",
  23111=>"111000000",
  23112=>"111100000",
  23113=>"000000100",
  23114=>"111110111",
  23115=>"000000011",
  23116=>"111111000",
  23117=>"000000000",
  23118=>"101001000",
  23119=>"000000011",
  23120=>"111000000",
  23121=>"000000110",
  23122=>"001001001",
  23123=>"110100100",
  23124=>"111111100",
  23125=>"111111000",
  23126=>"110110011",
  23127=>"000000000",
  23128=>"100000100",
  23129=>"100000000",
  23130=>"100100011",
  23131=>"011010000",
  23132=>"111111111",
  23133=>"000000000",
  23134=>"000001000",
  23135=>"100000000",
  23136=>"000000000",
  23137=>"000000111",
  23138=>"101100100",
  23139=>"111111001",
  23140=>"000000000",
  23141=>"000000110",
  23142=>"000000011",
  23143=>"000000100",
  23144=>"000000000",
  23145=>"000001001",
  23146=>"000000000",
  23147=>"000001111",
  23148=>"010111110",
  23149=>"000000000",
  23150=>"011000010",
  23151=>"111000101",
  23152=>"100110000",
  23153=>"111111111",
  23154=>"111000000",
  23155=>"000110111",
  23156=>"111100010",
  23157=>"110000000",
  23158=>"111111111",
  23159=>"100101010",
  23160=>"000111100",
  23161=>"111110110",
  23162=>"000000000",
  23163=>"110110110",
  23164=>"110110110",
  23165=>"110000000",
  23166=>"000000000",
  23167=>"100111111",
  23168=>"110111101",
  23169=>"000000000",
  23170=>"000100111",
  23171=>"111111111",
  23172=>"111111111",
  23173=>"001011111",
  23174=>"000100101",
  23175=>"001111110",
  23176=>"000011000",
  23177=>"101001000",
  23178=>"111111111",
  23179=>"111111111",
  23180=>"000000111",
  23181=>"111000000",
  23182=>"000001111",
  23183=>"111111010",
  23184=>"000001111",
  23185=>"000111000",
  23186=>"000000111",
  23187=>"001111011",
  23188=>"000000001",
  23189=>"110010000",
  23190=>"100100100",
  23191=>"001001001",
  23192=>"000000001",
  23193=>"000000000",
  23194=>"011000000",
  23195=>"000101100",
  23196=>"001000000",
  23197=>"101111111",
  23198=>"101110110",
  23199=>"000000000",
  23200=>"111111000",
  23201=>"000100111",
  23202=>"111101101",
  23203=>"001111111",
  23204=>"000000000",
  23205=>"111100000",
  23206=>"000000111",
  23207=>"001000111",
  23208=>"000000000",
  23209=>"111111111",
  23210=>"100111000",
  23211=>"000000110",
  23212=>"111111111",
  23213=>"111111000",
  23214=>"000000000",
  23215=>"110110111",
  23216=>"000000000",
  23217=>"000000110",
  23218=>"111111011",
  23219=>"111111000",
  23220=>"100100110",
  23221=>"000100111",
  23222=>"000000111",
  23223=>"111111000",
  23224=>"000000000",
  23225=>"001000000",
  23226=>"000000111",
  23227=>"111011000",
  23228=>"000000111",
  23229=>"111110111",
  23230=>"101000000",
  23231=>"000000000",
  23232=>"000000000",
  23233=>"000011001",
  23234=>"000000000",
  23235=>"001000001",
  23236=>"001100001",
  23237=>"111111111",
  23238=>"000001000",
  23239=>"000000111",
  23240=>"011001000",
  23241=>"111110000",
  23242=>"000000011",
  23243=>"000000011",
  23244=>"011000011",
  23245=>"000000001",
  23246=>"111000111",
  23247=>"000100000",
  23248=>"001000100",
  23249=>"000000100",
  23250=>"000110000",
  23251=>"111100000",
  23252=>"000000000",
  23253=>"111111110",
  23254=>"100010000",
  23255=>"000101100",
  23256=>"111111000",
  23257=>"000000111",
  23258=>"000000001",
  23259=>"000000000",
  23260=>"111010000",
  23261=>"000000000",
  23262=>"000111001",
  23263=>"100000000",
  23264=>"000000000",
  23265=>"111111000",
  23266=>"000100001",
  23267=>"110110110",
  23268=>"111111111",
  23269=>"110000001",
  23270=>"000000111",
  23271=>"000000111",
  23272=>"001000000",
  23273=>"000000000",
  23274=>"111110000",
  23275=>"000000000",
  23276=>"001000111",
  23277=>"011000000",
  23278=>"111101111",
  23279=>"000100110",
  23280=>"000000001",
  23281=>"110010000",
  23282=>"111101101",
  23283=>"000000000",
  23284=>"111111000",
  23285=>"111000000",
  23286=>"100111000",
  23287=>"011000000",
  23288=>"111111111",
  23289=>"000000111",
  23290=>"111101000",
  23291=>"111011001",
  23292=>"111010000",
  23293=>"111111111",
  23294=>"110000101",
  23295=>"000000000",
  23296=>"100000000",
  23297=>"011111000",
  23298=>"111111110",
  23299=>"101110000",
  23300=>"000000000",
  23301=>"111000000",
  23302=>"000000011",
  23303=>"110111111",
  23304=>"111111110",
  23305=>"000000011",
  23306=>"000000000",
  23307=>"111111000",
  23308=>"001001001",
  23309=>"100111011",
  23310=>"111111000",
  23311=>"000000111",
  23312=>"111100000",
  23313=>"000100111",
  23314=>"111000000",
  23315=>"000000000",
  23316=>"000000000",
  23317=>"111110110",
  23318=>"111111110",
  23319=>"111111111",
  23320=>"000001001",
  23321=>"000000000",
  23322=>"111111000",
  23323=>"000000000",
  23324=>"111011011",
  23325=>"001101111",
  23326=>"110000000",
  23327=>"000000000",
  23328=>"000101000",
  23329=>"000100111",
  23330=>"000000001",
  23331=>"111011101",
  23332=>"111000100",
  23333=>"111111111",
  23334=>"101000110",
  23335=>"111001110",
  23336=>"000000001",
  23337=>"111111000",
  23338=>"110000100",
  23339=>"000000000",
  23340=>"110000111",
  23341=>"011010111",
  23342=>"000000101",
  23343=>"001000000",
  23344=>"100111100",
  23345=>"110000000",
  23346=>"000110110",
  23347=>"000100111",
  23348=>"111000000",
  23349=>"111011000",
  23350=>"111000000",
  23351=>"000000111",
  23352=>"111001000",
  23353=>"111111111",
  23354=>"000000111",
  23355=>"100000000",
  23356=>"000000000",
  23357=>"000000001",
  23358=>"011111111",
  23359=>"111100100",
  23360=>"111100101",
  23361=>"111001010",
  23362=>"111110011",
  23363=>"000000000",
  23364=>"000000000",
  23365=>"111111111",
  23366=>"111110110",
  23367=>"011011011",
  23368=>"111111000",
  23369=>"000000000",
  23370=>"000000000",
  23371=>"111111111",
  23372=>"000000000",
  23373=>"111000000",
  23374=>"000010000",
  23375=>"111111000",
  23376=>"111001001",
  23377=>"001101111",
  23378=>"000000111",
  23379=>"000000000",
  23380=>"111000000",
  23381=>"011111001",
  23382=>"001000110",
  23383=>"111110111",
  23384=>"000011010",
  23385=>"000010000",
  23386=>"110000111",
  23387=>"110111110",
  23388=>"000101001",
  23389=>"111111111",
  23390=>"111100000",
  23391=>"000000000",
  23392=>"000000000",
  23393=>"000000111",
  23394=>"000001100",
  23395=>"001111111",
  23396=>"111111111",
  23397=>"010111110",
  23398=>"001001111",
  23399=>"000111111",
  23400=>"111111111",
  23401=>"011000000",
  23402=>"010000000",
  23403=>"111111001",
  23404=>"000100100",
  23405=>"000100111",
  23406=>"011000000",
  23407=>"000000111",
  23408=>"111000000",
  23409=>"001000111",
  23410=>"001111110",
  23411=>"011010111",
  23412=>"011111101",
  23413=>"100101110",
  23414=>"001101111",
  23415=>"101100100",
  23416=>"111000000",
  23417=>"111010111",
  23418=>"000000000",
  23419=>"110111111",
  23420=>"000101111",
  23421=>"100110000",
  23422=>"000000111",
  23423=>"111111111",
  23424=>"011111010",
  23425=>"111111110",
  23426=>"011110110",
  23427=>"000000000",
  23428=>"111011000",
  23429=>"000110000",
  23430=>"111000000",
  23431=>"110000000",
  23432=>"100000000",
  23433=>"111111110",
  23434=>"111111000",
  23435=>"000000000",
  23436=>"111111111",
  23437=>"001111111",
  23438=>"110111111",
  23439=>"111111101",
  23440=>"000101100",
  23441=>"100110111",
  23442=>"111010110",
  23443=>"010000000",
  23444=>"000000000",
  23445=>"000010000",
  23446=>"001001001",
  23447=>"110111111",
  23448=>"111111110",
  23449=>"110000101",
  23450=>"000000000",
  23451=>"101101101",
  23452=>"111111111",
  23453=>"110110110",
  23454=>"000000000",
  23455=>"010011001",
  23456=>"111111111",
  23457=>"011111101",
  23458=>"000000000",
  23459=>"000000001",
  23460=>"111110111",
  23461=>"000000111",
  23462=>"000000111",
  23463=>"111110000",
  23464=>"111111110",
  23465=>"111111100",
  23466=>"111111000",
  23467=>"000000111",
  23468=>"000000000",
  23469=>"111111000",
  23470=>"000001111",
  23471=>"000111111",
  23472=>"111111100",
  23473=>"110000000",
  23474=>"001000111",
  23475=>"111110000",
  23476=>"101000000",
  23477=>"001000111",
  23478=>"000000100",
  23479=>"000000111",
  23480=>"000000100",
  23481=>"000000000",
  23482=>"010000000",
  23483=>"110110100",
  23484=>"111111111",
  23485=>"111111000",
  23486=>"001001001",
  23487=>"011100100",
  23488=>"111001111",
  23489=>"111111111",
  23490=>"001000100",
  23491=>"111111000",
  23492=>"111111001",
  23493=>"001111111",
  23494=>"000000000",
  23495=>"000000001",
  23496=>"111000111",
  23497=>"111111000",
  23498=>"000000000",
  23499=>"011011011",
  23500=>"000000111",
  23501=>"000000111",
  23502=>"100000111",
  23503=>"000000000",
  23504=>"000000000",
  23505=>"111000000",
  23506=>"111111111",
  23507=>"010010111",
  23508=>"010010011",
  23509=>"110111000",
  23510=>"111111111",
  23511=>"111111111",
  23512=>"000000001",
  23513=>"101111110",
  23514=>"000100000",
  23515=>"111101101",
  23516=>"001111111",
  23517=>"111111111",
  23518=>"000111000",
  23519=>"001100100",
  23520=>"111111011",
  23521=>"000000000",
  23522=>"110111111",
  23523=>"100100101",
  23524=>"111111111",
  23525=>"010000000",
  23526=>"000000000",
  23527=>"000000000",
  23528=>"001111111",
  23529=>"000000000",
  23530=>"111110000",
  23531=>"000000001",
  23532=>"001111100",
  23533=>"011111111",
  23534=>"000011000",
  23535=>"111111000",
  23536=>"000000111",
  23537=>"000000110",
  23538=>"111001000",
  23539=>"000011001",
  23540=>"111010110",
  23541=>"000000000",
  23542=>"111110110",
  23543=>"111111101",
  23544=>"000011011",
  23545=>"111101001",
  23546=>"000000000",
  23547=>"111001001",
  23548=>"000100111",
  23549=>"000000100",
  23550=>"100000000",
  23551=>"000000111",
  23552=>"111110111",
  23553=>"001000000",
  23554=>"001101111",
  23555=>"111111111",
  23556=>"000000000",
  23557=>"101000001",
  23558=>"100100000",
  23559=>"000000000",
  23560=>"000000000",
  23561=>"001011000",
  23562=>"111100000",
  23563=>"000111111",
  23564=>"100100100",
  23565=>"111111111",
  23566=>"001000001",
  23567=>"110000000",
  23568=>"000000000",
  23569=>"110111011",
  23570=>"111111111",
  23571=>"110000000",
  23572=>"111100000",
  23573=>"111111111",
  23574=>"111111111",
  23575=>"111111111",
  23576=>"111101110",
  23577=>"111111000",
  23578=>"001000000",
  23579=>"110000100",
  23580=>"000100111",
  23581=>"111011111",
  23582=>"000000000",
  23583=>"001001111",
  23584=>"001000000",
  23585=>"110111111",
  23586=>"101000100",
  23587=>"111001111",
  23588=>"110110111",
  23589=>"000000000",
  23590=>"000011111",
  23591=>"011011001",
  23592=>"001000000",
  23593=>"000000000",
  23594=>"000000111",
  23595=>"111000000",
  23596=>"011001001",
  23597=>"111111110",
  23598=>"001001000",
  23599=>"111111000",
  23600=>"111111111",
  23601=>"111101000",
  23602=>"001001001",
  23603=>"100000110",
  23604=>"001111100",
  23605=>"101101110",
  23606=>"000000001",
  23607=>"100000000",
  23608=>"111110110",
  23609=>"100110111",
  23610=>"110111100",
  23611=>"111111001",
  23612=>"000000100",
  23613=>"111111010",
  23614=>"001000001",
  23615=>"111111111",
  23616=>"111100100",
  23617=>"001011111",
  23618=>"101000100",
  23619=>"101100110",
  23620=>"000000000",
  23621=>"110111010",
  23622=>"000000000",
  23623=>"100000000",
  23624=>"111110100",
  23625=>"011011111",
  23626=>"100000000",
  23627=>"111000000",
  23628=>"001000000",
  23629=>"111111111",
  23630=>"100100000",
  23631=>"000000000",
  23632=>"111111111",
  23633=>"111011011",
  23634=>"110000111",
  23635=>"001001001",
  23636=>"100100100",
  23637=>"000000101",
  23638=>"111000001",
  23639=>"101101000",
  23640=>"111111111",
  23641=>"000000000",
  23642=>"001001111",
  23643=>"101101111",
  23644=>"000000000",
  23645=>"111111111",
  23646=>"011111000",
  23647=>"000000111",
  23648=>"111101111",
  23649=>"010001001",
  23650=>"000000000",
  23651=>"000000000",
  23652=>"000000000",
  23653=>"110000000",
  23654=>"111100100",
  23655=>"000000000",
  23656=>"000000001",
  23657=>"100101111",
  23658=>"000001000",
  23659=>"111111111",
  23660=>"100000000",
  23661=>"111001000",
  23662=>"000000001",
  23663=>"010000000",
  23664=>"000000000",
  23665=>"100000000",
  23666=>"001001011",
  23667=>"111111111",
  23668=>"100000000",
  23669=>"111100000",
  23670=>"000000000",
  23671=>"111111111",
  23672=>"111101111",
  23673=>"000000000",
  23674=>"000000000",
  23675=>"000000000",
  23676=>"100100000",
  23677=>"110000001",
  23678=>"000000000",
  23679=>"000001000",
  23680=>"000111111",
  23681=>"110110000",
  23682=>"000000000",
  23683=>"111111111",
  23684=>"111111111",
  23685=>"111111111",
  23686=>"000000111",
  23687=>"110110111",
  23688=>"000000000",
  23689=>"010000000",
  23690=>"100011001",
  23691=>"111100000",
  23692=>"111111111",
  23693=>"000000000",
  23694=>"100000000",
  23695=>"111001000",
  23696=>"000000011",
  23697=>"111000000",
  23698=>"000100111",
  23699=>"100000000",
  23700=>"100111110",
  23701=>"101000000",
  23702=>"001000000",
  23703=>"011001111",
  23704=>"011111111",
  23705=>"111111111",
  23706=>"111111101",
  23707=>"000000000",
  23708=>"100000000",
  23709=>"000000100",
  23710=>"101000000",
  23711=>"110100100",
  23712=>"000001000",
  23713=>"000000000",
  23714=>"000110110",
  23715=>"000000000",
  23716=>"000000000",
  23717=>"010110011",
  23718=>"111001000",
  23719=>"010011110",
  23720=>"111101001",
  23721=>"000000000",
  23722=>"111111011",
  23723=>"111111111",
  23724=>"100111111",
  23725=>"001011111",
  23726=>"100000000",
  23727=>"000000111",
  23728=>"111111000",
  23729=>"111011011",
  23730=>"111111111",
  23731=>"000000100",
  23732=>"001001111",
  23733=>"110111111",
  23734=>"000111111",
  23735=>"111111100",
  23736=>"100001111",
  23737=>"101100100",
  23738=>"111111000",
  23739=>"111011111",
  23740=>"100100000",
  23741=>"111111101",
  23742=>"111000000",
  23743=>"111111111",
  23744=>"111111111",
  23745=>"100001011",
  23746=>"110100000",
  23747=>"000000000",
  23748=>"010000111",
  23749=>"000000100",
  23750=>"011110100",
  23751=>"110111011",
  23752=>"110111111",
  23753=>"110000000",
  23754=>"100100100",
  23755=>"000000000",
  23756=>"100111111",
  23757=>"110110001",
  23758=>"000000000",
  23759=>"000000011",
  23760=>"000000001",
  23761=>"000000101",
  23762=>"000000000",
  23763=>"111111100",
  23764=>"111001011",
  23765=>"110110110",
  23766=>"001111111",
  23767=>"111110100",
  23768=>"110111111",
  23769=>"010000000",
  23770=>"001000000",
  23771=>"000111111",
  23772=>"000100110",
  23773=>"001111111",
  23774=>"101001111",
  23775=>"100000000",
  23776=>"011000110",
  23777=>"000001001",
  23778=>"000000000",
  23779=>"111101111",
  23780=>"110110100",
  23781=>"000111001",
  23782=>"011011011",
  23783=>"110111001",
  23784=>"000000000",
  23785=>"010011111",
  23786=>"111000001",
  23787=>"000000000",
  23788=>"000011001",
  23789=>"000001011",
  23790=>"000000001",
  23791=>"111110111",
  23792=>"000000000",
  23793=>"000000011",
  23794=>"000000111",
  23795=>"110100011",
  23796=>"000000111",
  23797=>"000000100",
  23798=>"100101111",
  23799=>"001011111",
  23800=>"000000000",
  23801=>"000010010",
  23802=>"101001000",
  23803=>"001111111",
  23804=>"011011011",
  23805=>"111011011",
  23806=>"000000110",
  23807=>"110110110",
  23808=>"101001001",
  23809=>"100100111",
  23810=>"000010110",
  23811=>"000000000",
  23812=>"100000000",
  23813=>"000000001",
  23814=>"000000000",
  23815=>"111100101",
  23816=>"000000000",
  23817=>"111111111",
  23818=>"111111111",
  23819=>"111001000",
  23820=>"100100100",
  23821=>"111111001",
  23822=>"000000000",
  23823=>"000000000",
  23824=>"111111111",
  23825=>"000100100",
  23826=>"111111111",
  23827=>"111111111",
  23828=>"000000000",
  23829=>"111010111",
  23830=>"100001001",
  23831=>"111111111",
  23832=>"000011011",
  23833=>"111111111",
  23834=>"110101111",
  23835=>"111110000",
  23836=>"000000000",
  23837=>"111011111",
  23838=>"000010011",
  23839=>"111111111",
  23840=>"111111000",
  23841=>"000000000",
  23842=>"111010111",
  23843=>"111000111",
  23844=>"000110111",
  23845=>"000000111",
  23846=>"011111111",
  23847=>"111111111",
  23848=>"100110111",
  23849=>"101000000",
  23850=>"111110110",
  23851=>"111100000",
  23852=>"000000000",
  23853=>"111111011",
  23854=>"000000111",
  23855=>"101111011",
  23856=>"111011001",
  23857=>"110000000",
  23858=>"001001001",
  23859=>"000000000",
  23860=>"000000000",
  23861=>"111100100",
  23862=>"000000000",
  23863=>"000100100",
  23864=>"011001001",
  23865=>"000000000",
  23866=>"001100100",
  23867=>"000000000",
  23868=>"001001001",
  23869=>"100000000",
  23870=>"000000000",
  23871=>"101111000",
  23872=>"000000010",
  23873=>"111111111",
  23874=>"111111111",
  23875=>"111111011",
  23876=>"000000000",
  23877=>"111001000",
  23878=>"111111111",
  23879=>"000000001",
  23880=>"111111111",
  23881=>"000000100",
  23882=>"111000000",
  23883=>"111111111",
  23884=>"100000111",
  23885=>"000001111",
  23886=>"101011011",
  23887=>"111000000",
  23888=>"111111001",
  23889=>"011000001",
  23890=>"000000111",
  23891=>"001011111",
  23892=>"000000100",
  23893=>"011011011",
  23894=>"000001111",
  23895=>"000000001",
  23896=>"111111111",
  23897=>"111111111",
  23898=>"001111111",
  23899=>"001000011",
  23900=>"000000000",
  23901=>"111111111",
  23902=>"100100000",
  23903=>"111101101",
  23904=>"000000000",
  23905=>"000011111",
  23906=>"000001000",
  23907=>"000000000",
  23908=>"100000000",
  23909=>"100000000",
  23910=>"111111111",
  23911=>"111111111",
  23912=>"000100111",
  23913=>"000000000",
  23914=>"000000001",
  23915=>"111111011",
  23916=>"110000000",
  23917=>"011001101",
  23918=>"000000000",
  23919=>"000000000",
  23920=>"000000000",
  23921=>"111111110",
  23922=>"000000001",
  23923=>"111000111",
  23924=>"111101000",
  23925=>"000110110",
  23926=>"000000000",
  23927=>"000000110",
  23928=>"001000000",
  23929=>"000000001",
  23930=>"111111111",
  23931=>"000000000",
  23932=>"111010000",
  23933=>"000000000",
  23934=>"000000000",
  23935=>"000001111",
  23936=>"001001001",
  23937=>"000000000",
  23938=>"111111101",
  23939=>"111000000",
  23940=>"000000000",
  23941=>"000011011",
  23942=>"000000001",
  23943=>"000011011",
  23944=>"001001001",
  23945=>"011111111",
  23946=>"111111111",
  23947=>"000000011",
  23948=>"111111111",
  23949=>"100100000",
  23950=>"110111011",
  23951=>"000000000",
  23952=>"000000000",
  23953=>"000000000",
  23954=>"111111111",
  23955=>"000000000",
  23956=>"000000000",
  23957=>"000011011",
  23958=>"000000000",
  23959=>"111000000",
  23960=>"110000000",
  23961=>"000011110",
  23962=>"100000000",
  23963=>"111111111",
  23964=>"000000000",
  23965=>"001000000",
  23966=>"100100111",
  23967=>"000000000",
  23968=>"111011111",
  23969=>"011001000",
  23970=>"111000001",
  23971=>"011001111",
  23972=>"101111100",
  23973=>"111111111",
  23974=>"111111111",
  23975=>"001111111",
  23976=>"010010000",
  23977=>"100100110",
  23978=>"100110110",
  23979=>"111000001",
  23980=>"000101001",
  23981=>"000000101",
  23982=>"000000011",
  23983=>"111011001",
  23984=>"111111111",
  23985=>"000000110",
  23986=>"001001000",
  23987=>"110100000",
  23988=>"111011011",
  23989=>"101001000",
  23990=>"110111001",
  23991=>"000111111",
  23992=>"110011111",
  23993=>"111111111",
  23994=>"100000000",
  23995=>"000100101",
  23996=>"001011011",
  23997=>"000111111",
  23998=>"001000000",
  23999=>"101101001",
  24000=>"111001011",
  24001=>"011111111",
  24002=>"000011001",
  24003=>"000000000",
  24004=>"101000000",
  24005=>"011111110",
  24006=>"000001000",
  24007=>"001001101",
  24008=>"000000011",
  24009=>"110010111",
  24010=>"000000000",
  24011=>"000000000",
  24012=>"111111000",
  24013=>"000000000",
  24014=>"001111111",
  24015=>"111110110",
  24016=>"001001000",
  24017=>"111111111",
  24018=>"000000100",
  24019=>"000000000",
  24020=>"001001000",
  24021=>"100000000",
  24022=>"000000000",
  24023=>"011011011",
  24024=>"111110110",
  24025=>"000000011",
  24026=>"001000000",
  24027=>"000000000",
  24028=>"110110111",
  24029=>"100000000",
  24030=>"111111111",
  24031=>"101101010",
  24032=>"000000000",
  24033=>"111111111",
  24034=>"000000000",
  24035=>"000000000",
  24036=>"011000000",
  24037=>"111111111",
  24038=>"111111000",
  24039=>"111110111",
  24040=>"000000000",
  24041=>"100101000",
  24042=>"000111110",
  24043=>"111111111",
  24044=>"111101111",
  24045=>"110110110",
  24046=>"101101111",
  24047=>"110000000",
  24048=>"000000000",
  24049=>"000000000",
  24050=>"111111111",
  24051=>"001000001",
  24052=>"000000000",
  24053=>"000000000",
  24054=>"000000000",
  24055=>"100000000",
  24056=>"000110000",
  24057=>"100000001",
  24058=>"110000000",
  24059=>"111101111",
  24060=>"001000111",
  24061=>"111111111",
  24062=>"000000110",
  24063=>"111111111",
  24064=>"000000000",
  24065=>"100100000",
  24066=>"111111111",
  24067=>"000000010",
  24068=>"110010010",
  24069=>"110110110",
  24070=>"111000111",
  24071=>"111111000",
  24072=>"001000000",
  24073=>"010000010",
  24074=>"111111100",
  24075=>"011101111",
  24076=>"000000000",
  24077=>"111100110",
  24078=>"001101101",
  24079=>"111111111",
  24080=>"111111111",
  24081=>"011011111",
  24082=>"000000000",
  24083=>"000000000",
  24084=>"000000000",
  24085=>"000000000",
  24086=>"100000000",
  24087=>"000000000",
  24088=>"110000100",
  24089=>"011001000",
  24090=>"001000000",
  24091=>"110100111",
  24092=>"000000000",
  24093=>"001000110",
  24094=>"101000110",
  24095=>"111111111",
  24096=>"111001000",
  24097=>"111000110",
  24098=>"000000000",
  24099=>"011011011",
  24100=>"111111110",
  24101=>"111001000",
  24102=>"000000000",
  24103=>"111110110",
  24104=>"111111110",
  24105=>"000000000",
  24106=>"000010010",
  24107=>"111111111",
  24108=>"000000000",
  24109=>"110100110",
  24110=>"011010000",
  24111=>"100110000",
  24112=>"000000000",
  24113=>"000000000",
  24114=>"111111111",
  24115=>"110000000",
  24116=>"100100000",
  24117=>"100001000",
  24118=>"111111110",
  24119=>"011001000",
  24120=>"100000011",
  24121=>"111001011",
  24122=>"000000000",
  24123=>"100000100",
  24124=>"111101100",
  24125=>"110111111",
  24126=>"111111101",
  24127=>"000000000",
  24128=>"111101000",
  24129=>"111111111",
  24130=>"000000000",
  24131=>"111001111",
  24132=>"011001011",
  24133=>"011000000",
  24134=>"011001001",
  24135=>"001000000",
  24136=>"000000001",
  24137=>"001001001",
  24138=>"000000000",
  24139=>"111011001",
  24140=>"110111111",
  24141=>"111101101",
  24142=>"111100000",
  24143=>"111111111",
  24144=>"111000000",
  24145=>"111111111",
  24146=>"000000100",
  24147=>"000000000",
  24148=>"111111111",
  24149=>"001001001",
  24150=>"000000100",
  24151=>"000000000",
  24152=>"111111111",
  24153=>"000000100",
  24154=>"000000000",
  24155=>"110100100",
  24156=>"000000001",
  24157=>"111111111",
  24158=>"000000100",
  24159=>"111111111",
  24160=>"100110100",
  24161=>"111111010",
  24162=>"111111111",
  24163=>"011110110",
  24164=>"011111111",
  24165=>"100000000",
  24166=>"000101111",
  24167=>"111111111",
  24168=>"000100000",
  24169=>"111111111",
  24170=>"000000000",
  24171=>"111011000",
  24172=>"001111110",
  24173=>"001000000",
  24174=>"000111111",
  24175=>"011111001",
  24176=>"000000000",
  24177=>"000011111",
  24178=>"110110010",
  24179=>"111111111",
  24180=>"000000000",
  24181=>"111111110",
  24182=>"000101111",
  24183=>"111101110",
  24184=>"000000000",
  24185=>"000000000",
  24186=>"011000000",
  24187=>"111101111",
  24188=>"111110111",
  24189=>"000000000",
  24190=>"000000000",
  24191=>"010010000",
  24192=>"000000000",
  24193=>"101001000",
  24194=>"111111000",
  24195=>"000000000",
  24196=>"111111111",
  24197=>"111001011",
  24198=>"000000000",
  24199=>"111111111",
  24200=>"000000011",
  24201=>"000000100",
  24202=>"000001000",
  24203=>"010000001",
  24204=>"111111111",
  24205=>"111111111",
  24206=>"110011111",
  24207=>"000000000",
  24208=>"000000000",
  24209=>"000000000",
  24210=>"000000000",
  24211=>"000010000",
  24212=>"000000000",
  24213=>"111101100",
  24214=>"011111110",
  24215=>"001011111",
  24216=>"000000000",
  24217=>"101000111",
  24218=>"111000000",
  24219=>"111110000",
  24220=>"111111110",
  24221=>"111111111",
  24222=>"101101101",
  24223=>"000000001",
  24224=>"101000000",
  24225=>"000000000",
  24226=>"111111111",
  24227=>"000100100",
  24228=>"000000000",
  24229=>"001000100",
  24230=>"111111111",
  24231=>"111100000",
  24232=>"111111111",
  24233=>"000000000",
  24234=>"011001000",
  24235=>"111111111",
  24236=>"111011010",
  24237=>"111101111",
  24238=>"111111111",
  24239=>"111100001",
  24240=>"111111100",
  24241=>"101011111",
  24242=>"110110000",
  24243=>"111110000",
  24244=>"000111111",
  24245=>"101001000",
  24246=>"111111111",
  24247=>"111111000",
  24248=>"100000100",
  24249=>"111111000",
  24250=>"000000000",
  24251=>"110100100",
  24252=>"000000000",
  24253=>"111111111",
  24254=>"000000000",
  24255=>"111111111",
  24256=>"010010000",
  24257=>"111000000",
  24258=>"101111111",
  24259=>"111111111",
  24260=>"000000000",
  24261=>"011011001",
  24262=>"100000000",
  24263=>"111111111",
  24264=>"110110000",
  24265=>"111111111",
  24266=>"110000100",
  24267=>"111111011",
  24268=>"100100100",
  24269=>"011111111",
  24270=>"100110100",
  24271=>"000000000",
  24272=>"011011011",
  24273=>"111010000",
  24274=>"110100110",
  24275=>"100100101",
  24276=>"000000101",
  24277=>"000000000",
  24278=>"000000000",
  24279=>"110000000",
  24280=>"000000000",
  24281=>"000000111",
  24282=>"111100000",
  24283=>"000100111",
  24284=>"111111100",
  24285=>"000000100",
  24286=>"111111110",
  24287=>"101000011",
  24288=>"010111111",
  24289=>"111111111",
  24290=>"000000000",
  24291=>"111111111",
  24292=>"000000101",
  24293=>"000011011",
  24294=>"000000000",
  24295=>"001010110",
  24296=>"111111111",
  24297=>"111111111",
  24298=>"111111111",
  24299=>"101101001",
  24300=>"100111001",
  24301=>"000000000",
  24302=>"111011110",
  24303=>"111110110",
  24304=>"000000000",
  24305=>"000000000",
  24306=>"000110100",
  24307=>"000000000",
  24308=>"001000010",
  24309=>"111111111",
  24310=>"101110111",
  24311=>"000110111",
  24312=>"000000100",
  24313=>"111111111",
  24314=>"111101111",
  24315=>"000010101",
  24316=>"111111101",
  24317=>"100000001",
  24318=>"011000000",
  24319=>"100000100",
  24320=>"111111111",
  24321=>"001000000",
  24322=>"001001001",
  24323=>"000000000",
  24324=>"111110100",
  24325=>"000110110",
  24326=>"101101100",
  24327=>"111101111",
  24328=>"111110110",
  24329=>"000011111",
  24330=>"111111111",
  24331=>"000000110",
  24332=>"110110000",
  24333=>"111111111",
  24334=>"000000000",
  24335=>"000000000",
  24336=>"101101111",
  24337=>"100000000",
  24338=>"111111111",
  24339=>"010010110",
  24340=>"010000000",
  24341=>"000000000",
  24342=>"110110110",
  24343=>"100000000",
  24344=>"100000000",
  24345=>"111111111",
  24346=>"000110000",
  24347=>"111111101",
  24348=>"111100000",
  24349=>"111111111",
  24350=>"111111100",
  24351=>"110100100",
  24352=>"111101101",
  24353=>"000000000",
  24354=>"111111111",
  24355=>"011011111",
  24356=>"111000100",
  24357=>"000000000",
  24358=>"000000000",
  24359=>"111011011",
  24360=>"000110111",
  24361=>"100000000",
  24362=>"000000000",
  24363=>"001101101",
  24364=>"011111111",
  24365=>"011011111",
  24366=>"111111111",
  24367=>"111000000",
  24368=>"001011111",
  24369=>"000000000",
  24370=>"000000000",
  24371=>"000110000",
  24372=>"111101010",
  24373=>"001001011",
  24374=>"111101100",
  24375=>"000000000",
  24376=>"000000000",
  24377=>"000000111",
  24378=>"111111111",
  24379=>"100110111",
  24380=>"000000000",
  24381=>"101100111",
  24382=>"110111001",
  24383=>"000000100",
  24384=>"000000000",
  24385=>"000000000",
  24386=>"000100100",
  24387=>"000100000",
  24388=>"111111111",
  24389=>"000000000",
  24390=>"111111111",
  24391=>"111110111",
  24392=>"111111111",
  24393=>"000000000",
  24394=>"110110000",
  24395=>"110111010",
  24396=>"111011111",
  24397=>"000111111",
  24398=>"000000100",
  24399=>"110111111",
  24400=>"001001000",
  24401=>"111001011",
  24402=>"000000000",
  24403=>"000000000",
  24404=>"000000000",
  24405=>"011011001",
  24406=>"000000000",
  24407=>"000000000",
  24408=>"000000000",
  24409=>"000000000",
  24410=>"100101111",
  24411=>"000000000",
  24412=>"000000000",
  24413=>"111000000",
  24414=>"111111111",
  24415=>"111111111",
  24416=>"000001011",
  24417=>"000000000",
  24418=>"110110111",
  24419=>"000000001",
  24420=>"111001000",
  24421=>"000000000",
  24422=>"100100100",
  24423=>"111111111",
  24424=>"111000000",
  24425=>"011010000",
  24426=>"110000000",
  24427=>"000000000",
  24428=>"111101111",
  24429=>"011111111",
  24430=>"000000000",
  24431=>"110000000",
  24432=>"111000000",
  24433=>"001000000",
  24434=>"000001101",
  24435=>"000011110",
  24436=>"111111111",
  24437=>"000000000",
  24438=>"000000000",
  24439=>"000000000",
  24440=>"000000011",
  24441=>"000000000",
  24442=>"000100100",
  24443=>"111011001",
  24444=>"011001001",
  24445=>"111111111",
  24446=>"111001001",
  24447=>"011111111",
  24448=>"110000010",
  24449=>"111111111",
  24450=>"111111001",
  24451=>"111111111",
  24452=>"001001111",
  24453=>"111111111",
  24454=>"111101100",
  24455=>"100110000",
  24456=>"000111111",
  24457=>"001001011",
  24458=>"100100100",
  24459=>"011010010",
  24460=>"111111111",
  24461=>"100100100",
  24462=>"110110111",
  24463=>"000001001",
  24464=>"000000000",
  24465=>"111001001",
  24466=>"011111000",
  24467=>"000000000",
  24468=>"000000000",
  24469=>"000000000",
  24470=>"100100000",
  24471=>"111111111",
  24472=>"000000010",
  24473=>"111001011",
  24474=>"110001111",
  24475=>"000000111",
  24476=>"111100000",
  24477=>"101001111",
  24478=>"000000000",
  24479=>"111111111",
  24480=>"111111111",
  24481=>"001000001",
  24482=>"111000111",
  24483=>"111111111",
  24484=>"111011011",
  24485=>"111111111",
  24486=>"111100100",
  24487=>"000100111",
  24488=>"000010000",
  24489=>"000000010",
  24490=>"111010000",
  24491=>"000000000",
  24492=>"000000000",
  24493=>"001111111",
  24494=>"110111000",
  24495=>"111111111",
  24496=>"001000000",
  24497=>"011000000",
  24498=>"111000000",
  24499=>"111110000",
  24500=>"000000011",
  24501=>"100000000",
  24502=>"111000111",
  24503=>"000000000",
  24504=>"000000110",
  24505=>"000111111",
  24506=>"111000000",
  24507=>"101001011",
  24508=>"000000000",
  24509=>"111111111",
  24510=>"001000000",
  24511=>"100100100",
  24512=>"100111111",
  24513=>"000000000",
  24514=>"011111010",
  24515=>"000000000",
  24516=>"111111111",
  24517=>"111111111",
  24518=>"000000000",
  24519=>"000000000",
  24520=>"100000000",
  24521=>"100100000",
  24522=>"111000111",
  24523=>"000000111",
  24524=>"000100111",
  24525=>"000001000",
  24526=>"110111111",
  24527=>"011111011",
  24528=>"000000000",
  24529=>"000000000",
  24530=>"000000000",
  24531=>"111001001",
  24532=>"000000000",
  24533=>"011000110",
  24534=>"100000000",
  24535=>"000100100",
  24536=>"100000101",
  24537=>"111011001",
  24538=>"000000000",
  24539=>"111111111",
  24540=>"000000000",
  24541=>"011001000",
  24542=>"110110111",
  24543=>"111110000",
  24544=>"000010000",
  24545=>"111111111",
  24546=>"000000111",
  24547=>"111111111",
  24548=>"000010111",
  24549=>"101111111",
  24550=>"010111110",
  24551=>"000000000",
  24552=>"111111111",
  24553=>"110111111",
  24554=>"111111111",
  24555=>"000000110",
  24556=>"100110110",
  24557=>"000110110",
  24558=>"000111111",
  24559=>"111111111",
  24560=>"110110110",
  24561=>"000000100",
  24562=>"111111111",
  24563=>"000000000",
  24564=>"111111111",
  24565=>"111000011",
  24566=>"000000000",
  24567=>"000000000",
  24568=>"000010011",
  24569=>"000000000",
  24570=>"111111111",
  24571=>"111111111",
  24572=>"000000000",
  24573=>"111011011",
  24574=>"011000101",
  24575=>"000000000",
  24576=>"111001000",
  24577=>"111101000",
  24578=>"000000000",
  24579=>"111111111",
  24580=>"011000111",
  24581=>"111011111",
  24582=>"000000000",
  24583=>"001000111",
  24584=>"111110000",
  24585=>"000111111",
  24586=>"111010000",
  24587=>"000000000",
  24588=>"111111111",
  24589=>"001011000",
  24590=>"101100111",
  24591=>"111111111",
  24592=>"000100100",
  24593=>"000000000",
  24594=>"111001011",
  24595=>"111110111",
  24596=>"001001010",
  24597=>"000000111",
  24598=>"111011111",
  24599=>"011111111",
  24600=>"110110000",
  24601=>"000110100",
  24602=>"111111111",
  24603=>"001001000",
  24604=>"101000100",
  24605=>"100110111",
  24606=>"000010010",
  24607=>"000000101",
  24608=>"000000010",
  24609=>"000100110",
  24610=>"000100100",
  24611=>"000000000",
  24612=>"001001001",
  24613=>"011011011",
  24614=>"000000000",
  24615=>"111111111",
  24616=>"111111110",
  24617=>"000111111",
  24618=>"111011000",
  24619=>"001111111",
  24620=>"000000111",
  24621=>"111100100",
  24622=>"000011111",
  24623=>"000010000",
  24624=>"000000110",
  24625=>"111111111",
  24626=>"001000000",
  24627=>"011111011",
  24628=>"111011011",
  24629=>"000000100",
  24630=>"111011111",
  24631=>"000000000",
  24632=>"000000000",
  24633=>"011000001",
  24634=>"100000001",
  24635=>"111111000",
  24636=>"100100101",
  24637=>"011011000",
  24638=>"111100000",
  24639=>"111111111",
  24640=>"001011111",
  24641=>"000000000",
  24642=>"000111111",
  24643=>"110010110",
  24644=>"000000000",
  24645=>"010000001",
  24646=>"111111000",
  24647=>"111001011",
  24648=>"001001001",
  24649=>"101000000",
  24650=>"000000000",
  24651=>"000000110",
  24652=>"100000110",
  24653=>"000000111",
  24654=>"000111011",
  24655=>"000000100",
  24656=>"010111111",
  24657=>"111111001",
  24658=>"111010100",
  24659=>"100000000",
  24660=>"010000000",
  24661=>"111111111",
  24662=>"111111011",
  24663=>"111111111",
  24664=>"111110111",
  24665=>"111000000",
  24666=>"011001000",
  24667=>"001001000",
  24668=>"000000000",
  24669=>"001001000",
  24670=>"001010111",
  24671=>"110110000",
  24672=>"000110111",
  24673=>"110111111",
  24674=>"111001111",
  24675=>"111100111",
  24676=>"100111100",
  24677=>"101000000",
  24678=>"000011000",
  24679=>"001001011",
  24680=>"000000000",
  24681=>"111111111",
  24682=>"111111111",
  24683=>"000000000",
  24684=>"111101100",
  24685=>"000000011",
  24686=>"111110000",
  24687=>"001011111",
  24688=>"111111111",
  24689=>"010010001",
  24690=>"000001001",
  24691=>"000000110",
  24692=>"111111111",
  24693=>"011111111",
  24694=>"111110000",
  24695=>"000000000",
  24696=>"000000010",
  24697=>"111011001",
  24698=>"001011111",
  24699=>"000000001",
  24700=>"100100100",
  24701=>"011011111",
  24702=>"111011111",
  24703=>"000111010",
  24704=>"000000000",
  24705=>"000000111",
  24706=>"000000000",
  24707=>"000000000",
  24708=>"111111111",
  24709=>"111111111",
  24710=>"111111111",
  24711=>"111111110",
  24712=>"111111110",
  24713=>"011011001",
  24714=>"000000000",
  24715=>"001001111",
  24716=>"001000100",
  24717=>"100110000",
  24718=>"000000001",
  24719=>"011000110",
  24720=>"101101100",
  24721=>"000000000",
  24722=>"111000000",
  24723=>"011111101",
  24724=>"000001111",
  24725=>"111100000",
  24726=>"111111111",
  24727=>"111110000",
  24728=>"011001011",
  24729=>"001111111",
  24730=>"001001000",
  24731=>"001001111",
  24732=>"011001001",
  24733=>"111111110",
  24734=>"110001001",
  24735=>"000000000",
  24736=>"000000000",
  24737=>"101111011",
  24738=>"111110110",
  24739=>"111011000",
  24740=>"111011111",
  24741=>"000000000",
  24742=>"000111111",
  24743=>"000000001",
  24744=>"111111111",
  24745=>"000111111",
  24746=>"000000000",
  24747=>"110100101",
  24748=>"111011000",
  24749=>"111111011",
  24750=>"000000110",
  24751=>"111000100",
  24752=>"111111100",
  24753=>"000000001",
  24754=>"000000100",
  24755=>"000000111",
  24756=>"011011000",
  24757=>"001001001",
  24758=>"000111111",
  24759=>"011111111",
  24760=>"000010010",
  24761=>"011001011",
  24762=>"001000000",
  24763=>"111001111",
  24764=>"111111001",
  24765=>"000011111",
  24766=>"000000000",
  24767=>"011000000",
  24768=>"110110111",
  24769=>"000000110",
  24770=>"011011111",
  24771=>"111111011",
  24772=>"111100000",
  24773=>"111111111",
  24774=>"001001001",
  24775=>"111111111",
  24776=>"111111011",
  24777=>"111001101",
  24778=>"011001011",
  24779=>"000001000",
  24780=>"000001000",
  24781=>"111111100",
  24782=>"010000001",
  24783=>"111010000",
  24784=>"110000000",
  24785=>"010000000",
  24786=>"111000000",
  24787=>"000011111",
  24788=>"000100000",
  24789=>"110100101",
  24790=>"111111000",
  24791=>"000000000",
  24792=>"111111111",
  24793=>"000000110",
  24794=>"111000110",
  24795=>"011111101",
  24796=>"111111100",
  24797=>"000100110",
  24798=>"000100111",
  24799=>"000000000",
  24800=>"000001111",
  24801=>"111111111",
  24802=>"011000000",
  24803=>"100111111",
  24804=>"111111011",
  24805=>"100100001",
  24806=>"000000110",
  24807=>"000000000",
  24808=>"111111101",
  24809=>"111111111",
  24810=>"011111111",
  24811=>"000011111",
  24812=>"111100000",
  24813=>"111111111",
  24814=>"111111100",
  24815=>"111111111",
  24816=>"000000000",
  24817=>"001110100",
  24818=>"000000111",
  24819=>"011011111",
  24820=>"111111111",
  24821=>"111011000",
  24822=>"000111001",
  24823=>"111111111",
  24824=>"000111111",
  24825=>"000000000",
  24826=>"111000011",
  24827=>"000001000",
  24828=>"000000100",
  24829=>"111110111",
  24830=>"000011111",
  24831=>"011011111",
  24832=>"011011110",
  24833=>"110110100",
  24834=>"000000000",
  24835=>"111001101",
  24836=>"000000111",
  24837=>"110000011",
  24838=>"000000000",
  24839=>"010000011",
  24840=>"011111110",
  24841=>"000100111",
  24842=>"111000000",
  24843=>"000000000",
  24844=>"111111001",
  24845=>"000011010",
  24846=>"110111011",
  24847=>"101000000",
  24848=>"000000000",
  24849=>"000000000",
  24850=>"111111000",
  24851=>"111001000",
  24852=>"001001001",
  24853=>"100100101",
  24854=>"110110110",
  24855=>"000010010",
  24856=>"000100010",
  24857=>"010000000",
  24858=>"011000000",
  24859=>"000000111",
  24860=>"110110100",
  24861=>"000000010",
  24862=>"001111011",
  24863=>"111111010",
  24864=>"001000000",
  24865=>"000010011",
  24866=>"001000001",
  24867=>"111100110",
  24868=>"000000000",
  24869=>"111000110",
  24870=>"110100100",
  24871=>"000000110",
  24872=>"101000000",
  24873=>"000000011",
  24874=>"111111111",
  24875=>"000001011",
  24876=>"111011011",
  24877=>"000000110",
  24878=>"111111001",
  24879=>"000000000",
  24880=>"100100010",
  24881=>"111011111",
  24882=>"011000000",
  24883=>"011111111",
  24884=>"011111111",
  24885=>"111101111",
  24886=>"000111000",
  24887=>"111110111",
  24888=>"001111111",
  24889=>"000000000",
  24890=>"011111010",
  24891=>"111111111",
  24892=>"000000110",
  24893=>"000000011",
  24894=>"111111111",
  24895=>"000000000",
  24896=>"000101100",
  24897=>"000000000",
  24898=>"010111111",
  24899=>"100000000",
  24900=>"000000111",
  24901=>"000000111",
  24902=>"111111100",
  24903=>"111111000",
  24904=>"000111111",
  24905=>"011000000",
  24906=>"111011000",
  24907=>"000000100",
  24908=>"000000100",
  24909=>"000100111",
  24910=>"111111011",
  24911=>"001001101",
  24912=>"000100100",
  24913=>"010011111",
  24914=>"100000111",
  24915=>"000011000",
  24916=>"111111111",
  24917=>"110000001",
  24918=>"000011111",
  24919=>"111111111",
  24920=>"111111111",
  24921=>"000000000",
  24922=>"110111111",
  24923=>"001011111",
  24924=>"000000000",
  24925=>"111010111",
  24926=>"111111000",
  24927=>"000000000",
  24928=>"011111111",
  24929=>"000000000",
  24930=>"001110110",
  24931=>"000000000",
  24932=>"001010110",
  24933=>"100111000",
  24934=>"111111111",
  24935=>"110111000",
  24936=>"000000001",
  24937=>"001000000",
  24938=>"110110000",
  24939=>"111111110",
  24940=>"000000000",
  24941=>"010111111",
  24942=>"000011000",
  24943=>"100100110",
  24944=>"001011111",
  24945=>"000011111",
  24946=>"011011011",
  24947=>"110110110",
  24948=>"111111001",
  24949=>"011001100",
  24950=>"101000111",
  24951=>"000000000",
  24952=>"000000000",
  24953=>"000000100",
  24954=>"011001011",
  24955=>"000011001",
  24956=>"111100000",
  24957=>"011011111",
  24958=>"000000011",
  24959=>"101111111",
  24960=>"111001000",
  24961=>"001111111",
  24962=>"011111111",
  24963=>"111111111",
  24964=>"111111111",
  24965=>"001111111",
  24966=>"011111000",
  24967=>"111111111",
  24968=>"000000000",
  24969=>"000000000",
  24970=>"111011000",
  24971=>"111001000",
  24972=>"111001001",
  24973=>"000000000",
  24974=>"001000000",
  24975=>"111101111",
  24976=>"000111111",
  24977=>"100110111",
  24978=>"000000000",
  24979=>"000000001",
  24980=>"000000011",
  24981=>"010110000",
  24982=>"111011011",
  24983=>"111110110",
  24984=>"101100111",
  24985=>"111001001",
  24986=>"011111111",
  24987=>"111111111",
  24988=>"111111000",
  24989=>"111110110",
  24990=>"000001001",
  24991=>"111111111",
  24992=>"000111011",
  24993=>"100100100",
  24994=>"111000100",
  24995=>"011000100",
  24996=>"111111111",
  24997=>"111111111",
  24998=>"000111111",
  24999=>"011111111",
  25000=>"011010001",
  25001=>"011011000",
  25002=>"000001111",
  25003=>"010011000",
  25004=>"000100000",
  25005=>"000111111",
  25006=>"111111100",
  25007=>"110110111",
  25008=>"111000000",
  25009=>"110000000",
  25010=>"000000001",
  25011=>"000000000",
  25012=>"000000000",
  25013=>"000100110",
  25014=>"000000000",
  25015=>"000000001",
  25016=>"000000111",
  25017=>"111001111",
  25018=>"000000100",
  25019=>"001011011",
  25020=>"110111111",
  25021=>"111110110",
  25022=>"111111111",
  25023=>"011000111",
  25024=>"111111100",
  25025=>"000000000",
  25026=>"000000000",
  25027=>"111111111",
  25028=>"111011111",
  25029=>"011001100",
  25030=>"011111111",
  25031=>"001001011",
  25032=>"001000000",
  25033=>"001000000",
  25034=>"011010010",
  25035=>"111000000",
  25036=>"000010011",
  25037=>"111111111",
  25038=>"111111111",
  25039=>"110101101",
  25040=>"111111111",
  25041=>"000001000",
  25042=>"111111111",
  25043=>"111111101",
  25044=>"111111011",
  25045=>"111011000",
  25046=>"111111011",
  25047=>"111110000",
  25048=>"011111111",
  25049=>"010011111",
  25050=>"111111111",
  25051=>"000001000",
  25052=>"111111011",
  25053=>"111111111",
  25054=>"000000000",
  25055=>"000000011",
  25056=>"001011111",
  25057=>"000000010",
  25058=>"000000001",
  25059=>"111111000",
  25060=>"000111111",
  25061=>"001011010",
  25062=>"000000000",
  25063=>"000000100",
  25064=>"000001111",
  25065=>"100101101",
  25066=>"010111111",
  25067=>"000110010",
  25068=>"011000000",
  25069=>"110010000",
  25070=>"000000000",
  25071=>"000001001",
  25072=>"010000111",
  25073=>"100000000",
  25074=>"011011001",
  25075=>"011001001",
  25076=>"111111111",
  25077=>"110111111",
  25078=>"000000000",
  25079=>"111111111",
  25080=>"001001001",
  25081=>"100100100",
  25082=>"111111010",
  25083=>"111011011",
  25084=>"110000001",
  25085=>"000110111",
  25086=>"001000001",
  25087=>"000011111",
  25088=>"011011111",
  25089=>"111000000",
  25090=>"110000011",
  25091=>"000000011",
  25092=>"011011000",
  25093=>"000000011",
  25094=>"011000000",
  25095=>"111100111",
  25096=>"111111111",
  25097=>"111100000",
  25098=>"000111111",
  25099=>"000110111",
  25100=>"001011011",
  25101=>"111100000",
  25102=>"100000000",
  25103=>"111000000",
  25104=>"011000000",
  25105=>"111111001",
  25106=>"111011010",
  25107=>"000000001",
  25108=>"111000000",
  25109=>"000100110",
  25110=>"111111111",
  25111=>"111001000",
  25112=>"111000000",
  25113=>"000010000",
  25114=>"000000000",
  25115=>"101100000",
  25116=>"000000000",
  25117=>"001111000",
  25118=>"111110000",
  25119=>"111111000",
  25120=>"100100001",
  25121=>"000000000",
  25122=>"001001000",
  25123=>"111111111",
  25124=>"001000000",
  25125=>"001001000",
  25126=>"111000000",
  25127=>"111111111",
  25128=>"000000111",
  25129=>"111111110",
  25130=>"011000100",
  25131=>"100110100",
  25132=>"111111000",
  25133=>"111111000",
  25134=>"000000001",
  25135=>"011111111",
  25136=>"000000010",
  25137=>"000000000",
  25138=>"000000000",
  25139=>"111101000",
  25140=>"000001011",
  25141=>"001001000",
  25142=>"001000000",
  25143=>"000110111",
  25144=>"100111011",
  25145=>"000111111",
  25146=>"101101111",
  25147=>"111011001",
  25148=>"111111000",
  25149=>"111111100",
  25150=>"000000000",
  25151=>"001000100",
  25152=>"011111010",
  25153=>"000100110",
  25154=>"111111111",
  25155=>"111001000",
  25156=>"011000100",
  25157=>"001111101",
  25158=>"000000100",
  25159=>"001000000",
  25160=>"000100000",
  25161=>"111111111",
  25162=>"111111001",
  25163=>"111111000",
  25164=>"111111111",
  25165=>"111111000",
  25166=>"111000000",
  25167=>"111111111",
  25168=>"111111111",
  25169=>"000110111",
  25170=>"000000110",
  25171=>"111000000",
  25172=>"010010000",
  25173=>"000100000",
  25174=>"111111011",
  25175=>"011110110",
  25176=>"111111111",
  25177=>"111000100",
  25178=>"111000001",
  25179=>"100111111",
  25180=>"111100111",
  25181=>"111101000",
  25182=>"000000100",
  25183=>"111100000",
  25184=>"000101010",
  25185=>"111011000",
  25186=>"110110000",
  25187=>"000100000",
  25188=>"000000010",
  25189=>"000000000",
  25190=>"111111111",
  25191=>"111101100",
  25192=>"111100000",
  25193=>"000111111",
  25194=>"000100111",
  25195=>"111111111",
  25196=>"000110100",
  25197=>"100000000",
  25198=>"000001001",
  25199=>"110111101",
  25200=>"000111111",
  25201=>"000000111",
  25202=>"000111100",
  25203=>"110010000",
  25204=>"111111011",
  25205=>"001111111",
  25206=>"011010000",
  25207=>"000000000",
  25208=>"000000000",
  25209=>"100110010",
  25210=>"010010000",
  25211=>"000000101",
  25212=>"000000000",
  25213=>"000000101",
  25214=>"000000000",
  25215=>"000000000",
  25216=>"001000000",
  25217=>"110110110",
  25218=>"111101111",
  25219=>"111010000",
  25220=>"000101011",
  25221=>"111000000",
  25222=>"000111111",
  25223=>"000000011",
  25224=>"111111011",
  25225=>"111111000",
  25226=>"000101000",
  25227=>"111111000",
  25228=>"000001111",
  25229=>"000000000",
  25230=>"111111000",
  25231=>"111111100",
  25232=>"000000000",
  25233=>"000000000",
  25234=>"000000000",
  25235=>"000000000",
  25236=>"100111001",
  25237=>"000000000",
  25238=>"101100111",
  25239=>"111000011",
  25240=>"001000011",
  25241=>"000000000",
  25242=>"111000000",
  25243=>"000000000",
  25244=>"000000111",
  25245=>"000000100",
  25246=>"001000000",
  25247=>"111111111",
  25248=>"111000000",
  25249=>"100111111",
  25250=>"000000000",
  25251=>"000000110",
  25252=>"101001111",
  25253=>"101001001",
  25254=>"111110110",
  25255=>"000000110",
  25256=>"000000100",
  25257=>"000000110",
  25258=>"111111000",
  25259=>"000000111",
  25260=>"100001111",
  25261=>"001111000",
  25262=>"000000001",
  25263=>"111111000",
  25264=>"010111100",
  25265=>"100111000",
  25266=>"111111111",
  25267=>"111000111",
  25268=>"111111000",
  25269=>"000000111",
  25270=>"001000000",
  25271=>"111111100",
  25272=>"111111000",
  25273=>"010111111",
  25274=>"000000101",
  25275=>"001101111",
  25276=>"000000000",
  25277=>"001111111",
  25278=>"100001000",
  25279=>"001011011",
  25280=>"111111111",
  25281=>"111111111",
  25282=>"001111111",
  25283=>"111111010",
  25284=>"000111111",
  25285=>"000000111",
  25286=>"110000101",
  25287=>"000100110",
  25288=>"111111111",
  25289=>"111111111",
  25290=>"111001000",
  25291=>"111111111",
  25292=>"111111000",
  25293=>"111011001",
  25294=>"000000111",
  25295=>"001000000",
  25296=>"100100001",
  25297=>"111000000",
  25298=>"000001001",
  25299=>"101111111",
  25300=>"011001000",
  25301=>"000000000",
  25302=>"111110000",
  25303=>"111001001",
  25304=>"000110110",
  25305=>"001111000",
  25306=>"111111111",
  25307=>"111001000",
  25308=>"111000000",
  25309=>"000000000",
  25310=>"111111111",
  25311=>"001001001",
  25312=>"111111000",
  25313=>"110000000",
  25314=>"111110110",
  25315=>"000000000",
  25316=>"000000000",
  25317=>"001100100",
  25318=>"110100111",
  25319=>"110110000",
  25320=>"000000000",
  25321=>"000000000",
  25322=>"000111111",
  25323=>"111001000",
  25324=>"101111001",
  25325=>"111111111",
  25326=>"000000111",
  25327=>"000000000",
  25328=>"111111111",
  25329=>"100000000",
  25330=>"000000000",
  25331=>"111111111",
  25332=>"000101101",
  25333=>"111111011",
  25334=>"110000000",
  25335=>"000110001",
  25336=>"111111111",
  25337=>"011111000",
  25338=>"000000000",
  25339=>"000110000",
  25340=>"111111000",
  25341=>"110010010",
  25342=>"101000111",
  25343=>"001000000",
  25344=>"111000101",
  25345=>"001010000",
  25346=>"000000000",
  25347=>"010110000",
  25348=>"111000000",
  25349=>"000000111",
  25350=>"000001011",
  25351=>"000000000",
  25352=>"110111111",
  25353=>"000010111",
  25354=>"111010000",
  25355=>"111011001",
  25356=>"100110111",
  25357=>"001001001",
  25358=>"000000100",
  25359=>"111111000",
  25360=>"001000000",
  25361=>"000111111",
  25362=>"010011011",
  25363=>"000111111",
  25364=>"000111111",
  25365=>"000111000",
  25366=>"000100000",
  25367=>"000000000",
  25368=>"100101111",
  25369=>"011111000",
  25370=>"111111000",
  25371=>"111111111",
  25372=>"001001001",
  25373=>"111111000",
  25374=>"000000101",
  25375=>"111000000",
  25376=>"111000100",
  25377=>"111111000",
  25378=>"001101101",
  25379=>"000000000",
  25380=>"000000000",
  25381=>"111111001",
  25382=>"100100000",
  25383=>"100111111",
  25384=>"000000000",
  25385=>"000100111",
  25386=>"000111111",
  25387=>"000111111",
  25388=>"000000000",
  25389=>"001011111",
  25390=>"000100111",
  25391=>"000000110",
  25392=>"000000000",
  25393=>"010110110",
  25394=>"111111111",
  25395=>"000111111",
  25396=>"111100110",
  25397=>"111110010",
  25398=>"111110110",
  25399=>"000000111",
  25400=>"001111111",
  25401=>"111000000",
  25402=>"111100100",
  25403=>"111101000",
  25404=>"001000000",
  25405=>"100000000",
  25406=>"111110000",
  25407=>"111000100",
  25408=>"010111111",
  25409=>"100100000",
  25410=>"001000011",
  25411=>"000011000",
  25412=>"111111110",
  25413=>"111000011",
  25414=>"111111101",
  25415=>"000011000",
  25416=>"001011000",
  25417=>"111000000",
  25418=>"000110110",
  25419=>"110111001",
  25420=>"111111111",
  25421=>"110111111",
  25422=>"111111000",
  25423=>"111111100",
  25424=>"111110110",
  25425=>"000000000",
  25426=>"000111111",
  25427=>"001011111",
  25428=>"000000011",
  25429=>"011011011",
  25430=>"000000111",
  25431=>"100000000",
  25432=>"000111111",
  25433=>"100100100",
  25434=>"000011111",
  25435=>"000001111",
  25436=>"000000000",
  25437=>"001001101",
  25438=>"000000111",
  25439=>"111011000",
  25440=>"000111011",
  25441=>"000000000",
  25442=>"111111001",
  25443=>"111111011",
  25444=>"111111000",
  25445=>"000000000",
  25446=>"101101111",
  25447=>"000111111",
  25448=>"011011111",
  25449=>"110111100",
  25450=>"000000000",
  25451=>"000011001",
  25452=>"111111110",
  25453=>"111000111",
  25454=>"111111111",
  25455=>"100000000",
  25456=>"000010011",
  25457=>"000000110",
  25458=>"000000101",
  25459=>"000000000",
  25460=>"000111110",
  25461=>"000001001",
  25462=>"110111111",
  25463=>"000100100",
  25464=>"000000000",
  25465=>"111111000",
  25466=>"101000000",
  25467=>"111111111",
  25468=>"111111111",
  25469=>"001101111",
  25470=>"111111111",
  25471=>"111111000",
  25472=>"001011000",
  25473=>"011011110",
  25474=>"000000010",
  25475=>"000000000",
  25476=>"110010000",
  25477=>"111111111",
  25478=>"000110111",
  25479=>"111101000",
  25480=>"111111111",
  25481=>"101000110",
  25482=>"000000111",
  25483=>"111111111",
  25484=>"111000000",
  25485=>"111111000",
  25486=>"000000000",
  25487=>"110000000",
  25488=>"110000000",
  25489=>"001011000",
  25490=>"110111111",
  25491=>"000000000",
  25492=>"001001111",
  25493=>"111111111",
  25494=>"111111111",
  25495=>"100110000",
  25496=>"000011111",
  25497=>"000000000",
  25498=>"011000011",
  25499=>"000001111",
  25500=>"111110000",
  25501=>"011111111",
  25502=>"000101111",
  25503=>"111111111",
  25504=>"111111110",
  25505=>"110111011",
  25506=>"111111111",
  25507=>"000000111",
  25508=>"000110110",
  25509=>"111111111",
  25510=>"000000111",
  25511=>"111000000",
  25512=>"111111111",
  25513=>"011010000",
  25514=>"000000100",
  25515=>"000000000",
  25516=>"000000000",
  25517=>"000000100",
  25518=>"111000110",
  25519=>"111011000",
  25520=>"111010011",
  25521=>"110111110",
  25522=>"100000000",
  25523=>"100110111",
  25524=>"000100111",
  25525=>"000000100",
  25526=>"011111100",
  25527=>"000000111",
  25528=>"111111111",
  25529=>"001001111",
  25530=>"111111110",
  25531=>"000000000",
  25532=>"000011111",
  25533=>"000000000",
  25534=>"100101111",
  25535=>"000100110",
  25536=>"000000000",
  25537=>"111000000",
  25538=>"111111011",
  25539=>"111111000",
  25540=>"000111111",
  25541=>"000100000",
  25542=>"111111011",
  25543=>"010011111",
  25544=>"000111100",
  25545=>"111001000",
  25546=>"110110110",
  25547=>"001000000",
  25548=>"001001000",
  25549=>"111111011",
  25550=>"100000000",
  25551=>"000000000",
  25552=>"110111100",
  25553=>"100100110",
  25554=>"110101011",
  25555=>"000000000",
  25556=>"001000000",
  25557=>"111000000",
  25558=>"000011000",
  25559=>"100111111",
  25560=>"111001001",
  25561=>"111111010",
  25562=>"000000000",
  25563=>"000000111",
  25564=>"110000000",
  25565=>"001000000",
  25566=>"111111111",
  25567=>"000000000",
  25568=>"000110110",
  25569=>"011010000",
  25570=>"000000111",
  25571=>"111000000",
  25572=>"000000000",
  25573=>"111110000",
  25574=>"111101111",
  25575=>"110110100",
  25576=>"000000000",
  25577=>"100111111",
  25578=>"000000000",
  25579=>"000011000",
  25580=>"000111001",
  25581=>"101101001",
  25582=>"111111000",
  25583=>"111001111",
  25584=>"110000000",
  25585=>"000000001",
  25586=>"000001000",
  25587=>"000000000",
  25588=>"100000000",
  25589=>"000111111",
  25590=>"011000111",
  25591=>"000001001",
  25592=>"010111000",
  25593=>"001111111",
  25594=>"011011010",
  25595=>"111111111",
  25596=>"000000110",
  25597=>"111111100",
  25598=>"000111100",
  25599=>"011000000",
  25600=>"000000000",
  25601=>"111111111",
  25602=>"001000000",
  25603=>"111111111",
  25604=>"001101101",
  25605=>"111011001",
  25606=>"111111111",
  25607=>"111111100",
  25608=>"111100000",
  25609=>"111110110",
  25610=>"110100000",
  25611=>"111110011",
  25612=>"100100100",
  25613=>"010000000",
  25614=>"000011111",
  25615=>"000000000",
  25616=>"000000111",
  25617=>"000111011",
  25618=>"111111111",
  25619=>"011010000",
  25620=>"000000100",
  25621=>"111111000",
  25622=>"111111111",
  25623=>"000000000",
  25624=>"000000000",
  25625=>"011111010",
  25626=>"001000000",
  25627=>"111111110",
  25628=>"111111100",
  25629=>"000100111",
  25630=>"111011100",
  25631=>"100010111",
  25632=>"000001111",
  25633=>"000000000",
  25634=>"000000000",
  25635=>"100000000",
  25636=>"000000000",
  25637=>"000000000",
  25638=>"111111101",
  25639=>"111111111",
  25640=>"111111011",
  25641=>"000001001",
  25642=>"110111111",
  25643=>"111111111",
  25644=>"111111111",
  25645=>"010010000",
  25646=>"000000000",
  25647=>"111000101",
  25648=>"111111111",
  25649=>"110000101",
  25650=>"000010011",
  25651=>"000110110",
  25652=>"000100100",
  25653=>"000000000",
  25654=>"111111111",
  25655=>"111101000",
  25656=>"110110111",
  25657=>"101000000",
  25658=>"111111111",
  25659=>"000000000",
  25660=>"111111111",
  25661=>"001000000",
  25662=>"000010110",
  25663=>"000000000",
  25664=>"101111110",
  25665=>"111011000",
  25666=>"100000101",
  25667=>"000000100",
  25668=>"111110110",
  25669=>"000000000",
  25670=>"110110100",
  25671=>"111111111",
  25672=>"100011001",
  25673=>"000000001",
  25674=>"001011000",
  25675=>"100000111",
  25676=>"101111111",
  25677=>"001111000",
  25678=>"000000000",
  25679=>"000111111",
  25680=>"111100000",
  25681=>"000000000",
  25682=>"000000000",
  25683=>"001001101",
  25684=>"000001001",
  25685=>"100000000",
  25686=>"111111111",
  25687=>"000000000",
  25688=>"100000000",
  25689=>"000000000",
  25690=>"111111111",
  25691=>"010011000",
  25692=>"000111111",
  25693=>"111111110",
  25694=>"001011011",
  25695=>"110011111",
  25696=>"111111111",
  25697=>"000000000",
  25698=>"001000111",
  25699=>"111111111",
  25700=>"111100000",
  25701=>"100101111",
  25702=>"111111111",
  25703=>"000000000",
  25704=>"000000000",
  25705=>"001000000",
  25706=>"111000000",
  25707=>"010010010",
  25708=>"011111111",
  25709=>"111111111",
  25710=>"000000000",
  25711=>"011111111",
  25712=>"000000000",
  25713=>"000000000",
  25714=>"111001001",
  25715=>"000011111",
  25716=>"000000000",
  25717=>"010111111",
  25718=>"000000000",
  25719=>"100000101",
  25720=>"100000000",
  25721=>"000000000",
  25722=>"000000000",
  25723=>"000000000",
  25724=>"001111111",
  25725=>"000000000",
  25726=>"111111111",
  25727=>"111111001",
  25728=>"001101111",
  25729=>"010011111",
  25730=>"000000101",
  25731=>"110110100",
  25732=>"100100111",
  25733=>"000000000",
  25734=>"001000000",
  25735=>"000011111",
  25736=>"111110111",
  25737=>"111111111",
  25738=>"000000000",
  25739=>"110111111",
  25740=>"111111111",
  25741=>"000000000",
  25742=>"100100000",
  25743=>"111111111",
  25744=>"000000000",
  25745=>"111111111",
  25746=>"000000100",
  25747=>"101000000",
  25748=>"100100100",
  25749=>"011011111",
  25750=>"000000000",
  25751=>"000000000",
  25752=>"001001000",
  25753=>"000000000",
  25754=>"000100110",
  25755=>"000100010",
  25756=>"010111111",
  25757=>"000000000",
  25758=>"000000000",
  25759=>"000000000",
  25760=>"001000000",
  25761=>"111110100",
  25762=>"000000000",
  25763=>"111000000",
  25764=>"000000000",
  25765=>"111111110",
  25766=>"000000000",
  25767=>"000000000",
  25768=>"111111111",
  25769=>"011000000",
  25770=>"000000000",
  25771=>"111111111",
  25772=>"000000000",
  25773=>"000100100",
  25774=>"111100100",
  25775=>"001111111",
  25776=>"000000111",
  25777=>"111111011",
  25778=>"111111111",
  25779=>"100000101",
  25780=>"111000000",
  25781=>"011000110",
  25782=>"000000000",
  25783=>"111111001",
  25784=>"111101111",
  25785=>"000000011",
  25786=>"000000000",
  25787=>"111111111",
  25788=>"111111111",
  25789=>"110010000",
  25790=>"000111111",
  25791=>"100100100",
  25792=>"110000000",
  25793=>"000000000",
  25794=>"000000000",
  25795=>"000000000",
  25796=>"000000001",
  25797=>"000000000",
  25798=>"110110110",
  25799=>"000100000",
  25800=>"111111111",
  25801=>"000111111",
  25802=>"111111111",
  25803=>"000000001",
  25804=>"000000000",
  25805=>"111111000",
  25806=>"000000000",
  25807=>"000000000",
  25808=>"111111111",
  25809=>"000001111",
  25810=>"000001111",
  25811=>"000000000",
  25812=>"000111111",
  25813=>"111111111",
  25814=>"111001011",
  25815=>"111111111",
  25816=>"000000000",
  25817=>"100111111",
  25818=>"111111111",
  25819=>"111111111",
  25820=>"110001111",
  25821=>"100110101",
  25822=>"000000000",
  25823=>"111101000",
  25824=>"000000001",
  25825=>"111111000",
  25826=>"110000000",
  25827=>"000000000",
  25828=>"111011100",
  25829=>"100100111",
  25830=>"111111111",
  25831=>"001100110",
  25832=>"000000000",
  25833=>"000000000",
  25834=>"111011111",
  25835=>"110011000",
  25836=>"000000111",
  25837=>"000000000",
  25838=>"000001000",
  25839=>"101111111",
  25840=>"110100000",
  25841=>"000000000",
  25842=>"000000100",
  25843=>"000000000",
  25844=>"001000000",
  25845=>"000111110",
  25846=>"110110010",
  25847=>"000000011",
  25848=>"110100111",
  25849=>"000001001",
  25850=>"000111111",
  25851=>"111111111",
  25852=>"011011010",
  25853=>"001111111",
  25854=>"011110111",
  25855=>"111111111",
  25856=>"000110000",
  25857=>"111101001",
  25858=>"001000000",
  25859=>"111111111",
  25860=>"100100100",
  25861=>"111111110",
  25862=>"101101101",
  25863=>"000001101",
  25864=>"000000000",
  25865=>"000000000",
  25866=>"100100101",
  25867=>"110110110",
  25868=>"000000111",
  25869=>"010010000",
  25870=>"101000000",
  25871=>"100111111",
  25872=>"111111100",
  25873=>"111100000",
  25874=>"000011000",
  25875=>"101110111",
  25876=>"000000000",
  25877=>"000110110",
  25878=>"001000000",
  25879=>"100000000",
  25880=>"001001000",
  25881=>"000000001",
  25882=>"000000000",
  25883=>"111011000",
  25884=>"111100000",
  25885=>"111111111",
  25886=>"110111111",
  25887=>"010111111",
  25888=>"110111111",
  25889=>"000000000",
  25890=>"000011111",
  25891=>"111111111",
  25892=>"100100001",
  25893=>"000000000",
  25894=>"001001001",
  25895=>"111111111",
  25896=>"111101110",
  25897=>"000000000",
  25898=>"100110101",
  25899=>"000110000",
  25900=>"010011011",
  25901=>"000000000",
  25902=>"100111111",
  25903=>"000000000",
  25904=>"111001001",
  25905=>"000000000",
  25906=>"101111111",
  25907=>"111111111",
  25908=>"111111111",
  25909=>"000000110",
  25910=>"001111110",
  25911=>"110110000",
  25912=>"000000000",
  25913=>"000000000",
  25914=>"001011000",
  25915=>"101001001",
  25916=>"000000000",
  25917=>"000010000",
  25918=>"101111111",
  25919=>"100100111",
  25920=>"111111000",
  25921=>"000000000",
  25922=>"111110110",
  25923=>"111111111",
  25924=>"111111111",
  25925=>"111111111",
  25926=>"000000000",
  25927=>"111111111",
  25928=>"000000000",
  25929=>"111111111",
  25930=>"000000000",
  25931=>"100101111",
  25932=>"110111111",
  25933=>"000001000",
  25934=>"111000000",
  25935=>"110111100",
  25936=>"000111111",
  25937=>"000000110",
  25938=>"000000001",
  25939=>"111111001",
  25940=>"000000000",
  25941=>"011011001",
  25942=>"101000101",
  25943=>"000110110",
  25944=>"000000000",
  25945=>"111001001",
  25946=>"111111111",
  25947=>"111111110",
  25948=>"000001101",
  25949=>"000111111",
  25950=>"000000000",
  25951=>"000111111",
  25952=>"111111111",
  25953=>"000000000",
  25954=>"000000000",
  25955=>"111111111",
  25956=>"000101011",
  25957=>"001001001",
  25958=>"100001000",
  25959=>"000000100",
  25960=>"010111111",
  25961=>"011111111",
  25962=>"111111001",
  25963=>"000110010",
  25964=>"000001001",
  25965=>"000000000",
  25966=>"000000000",
  25967=>"111111111",
  25968=>"000000000",
  25969=>"000000111",
  25970=>"000000000",
  25971=>"011001001",
  25972=>"111111111",
  25973=>"100100000",
  25974=>"000110011",
  25975=>"000001010",
  25976=>"111111111",
  25977=>"111111111",
  25978=>"111111111",
  25979=>"000100100",
  25980=>"111011001",
  25981=>"111001000",
  25982=>"001001000",
  25983=>"101001011",
  25984=>"000000000",
  25985=>"101101000",
  25986=>"000000000",
  25987=>"000000000",
  25988=>"000110111",
  25989=>"000000000",
  25990=>"101000000",
  25991=>"100110100",
  25992=>"111000100",
  25993=>"111111111",
  25994=>"001111111",
  25995=>"111111111",
  25996=>"111101111",
  25997=>"000000010",
  25998=>"010000000",
  25999=>"011001000",
  26000=>"000000000",
  26001=>"111111111",
  26002=>"111001001",
  26003=>"000001011",
  26004=>"110110000",
  26005=>"000010010",
  26006=>"101111111",
  26007=>"100100100",
  26008=>"111100100",
  26009=>"011111111",
  26010=>"111111010",
  26011=>"000000100",
  26012=>"111111111",
  26013=>"111000000",
  26014=>"000000000",
  26015=>"000000000",
  26016=>"111111111",
  26017=>"111111011",
  26018=>"000000000",
  26019=>"000000100",
  26020=>"000000000",
  26021=>"000000000",
  26022=>"111101111",
  26023=>"000000000",
  26024=>"111111111",
  26025=>"000000000",
  26026=>"111111111",
  26027=>"000000110",
  26028=>"000000001",
  26029=>"000000000",
  26030=>"000000000",
  26031=>"111111111",
  26032=>"100100111",
  26033=>"010000000",
  26034=>"110100100",
  26035=>"101111010",
  26036=>"100000000",
  26037=>"000100111",
  26038=>"111111000",
  26039=>"111111111",
  26040=>"000010000",
  26041=>"001000000",
  26042=>"001001001",
  26043=>"111111100",
  26044=>"111111111",
  26045=>"111111101",
  26046=>"111000111",
  26047=>"001011000",
  26048=>"000000000",
  26049=>"111111111",
  26050=>"100000000",
  26051=>"010111000",
  26052=>"100100000",
  26053=>"000110110",
  26054=>"111111000",
  26055=>"111111111",
  26056=>"000000000",
  26057=>"010110000",
  26058=>"001111111",
  26059=>"000000011",
  26060=>"110000000",
  26061=>"111111111",
  26062=>"000000110",
  26063=>"001011001",
  26064=>"110100101",
  26065=>"000000000",
  26066=>"010011111",
  26067=>"000001001",
  26068=>"111111111",
  26069=>"001000000",
  26070=>"001011000",
  26071=>"011011011",
  26072=>"100111111",
  26073=>"000000000",
  26074=>"001000001",
  26075=>"000000000",
  26076=>"000011011",
  26077=>"000000010",
  26078=>"111110110",
  26079=>"000110000",
  26080=>"111111111",
  26081=>"000001000",
  26082=>"000000000",
  26083=>"100110111",
  26084=>"001111111",
  26085=>"001001011",
  26086=>"100111100",
  26087=>"001011111",
  26088=>"111100000",
  26089=>"111100100",
  26090=>"100111100",
  26091=>"110111011",
  26092=>"001000000",
  26093=>"000100000",
  26094=>"001001000",
  26095=>"000000000",
  26096=>"001111001",
  26097=>"111111111",
  26098=>"000000000",
  26099=>"111111111",
  26100=>"000000000",
  26101=>"000001111",
  26102=>"011111111",
  26103=>"011011000",
  26104=>"000000000",
  26105=>"000100101",
  26106=>"000000000",
  26107=>"111111110",
  26108=>"111111111",
  26109=>"111111111",
  26110=>"110111111",
  26111=>"001000100",
  26112=>"000000111",
  26113=>"111110000",
  26114=>"111111111",
  26115=>"111011000",
  26116=>"011001111",
  26117=>"100100000",
  26118=>"111111101",
  26119=>"111111111",
  26120=>"101111111",
  26121=>"000011111",
  26122=>"101000000",
  26123=>"000000011",
  26124=>"000000010",
  26125=>"110000111",
  26126=>"111110000",
  26127=>"111111111",
  26128=>"111111011",
  26129=>"000111111",
  26130=>"000000000",
  26131=>"100100111",
  26132=>"111111111",
  26133=>"010111111",
  26134=>"110000000",
  26135=>"111111111",
  26136=>"000000000",
  26137=>"000011100",
  26138=>"110110100",
  26139=>"111110010",
  26140=>"011111111",
  26141=>"000000000",
  26142=>"111010011",
  26143=>"000001101",
  26144=>"111111111",
  26145=>"111001001",
  26146=>"111111111",
  26147=>"000100000",
  26148=>"000000000",
  26149=>"011011011",
  26150=>"000000000",
  26151=>"111111111",
  26152=>"111111111",
  26153=>"010000000",
  26154=>"101101111",
  26155=>"100110011",
  26156=>"001001011",
  26157=>"000110110",
  26158=>"000111110",
  26159=>"000000000",
  26160=>"010110110",
  26161=>"101111110",
  26162=>"101101111",
  26163=>"000000000",
  26164=>"000000000",
  26165=>"000000000",
  26166=>"111111111",
  26167=>"001011111",
  26168=>"101001111",
  26169=>"000100111",
  26170=>"000000000",
  26171=>"100110111",
  26172=>"111110000",
  26173=>"000100111",
  26174=>"000000000",
  26175=>"110101001",
  26176=>"100100101",
  26177=>"001111111",
  26178=>"100111110",
  26179=>"011111111",
  26180=>"111111111",
  26181=>"000000011",
  26182=>"000111111",
  26183=>"001000000",
  26184=>"111111011",
  26185=>"000000001",
  26186=>"110000000",
  26187=>"000000111",
  26188=>"111111111",
  26189=>"000110111",
  26190=>"111111111",
  26191=>"100000011",
  26192=>"000000000",
  26193=>"000011011",
  26194=>"001011111",
  26195=>"000000100",
  26196=>"000011111",
  26197=>"011111011",
  26198=>"011111111",
  26199=>"111101111",
  26200=>"000000001",
  26201=>"000000000",
  26202=>"000111000",
  26203=>"000000110",
  26204=>"111011111",
  26205=>"111111001",
  26206=>"111111111",
  26207=>"000000000",
  26208=>"111000011",
  26209=>"111111111",
  26210=>"111111111",
  26211=>"000000111",
  26212=>"111111111",
  26213=>"111000111",
  26214=>"111000000",
  26215=>"000000000",
  26216=>"111110000",
  26217=>"000110010",
  26218=>"000100111",
  26219=>"001111111",
  26220=>"001001000",
  26221=>"110111110",
  26222=>"111111111",
  26223=>"000000000",
  26224=>"111110110",
  26225=>"011100111",
  26226=>"001100100",
  26227=>"100000000",
  26228=>"111011000",
  26229=>"000000000",
  26230=>"111101111",
  26231=>"000000000",
  26232=>"111110111",
  26233=>"111010000",
  26234=>"010011111",
  26235=>"111111111",
  26236=>"110010000",
  26237=>"011111000",
  26238=>"111111011",
  26239=>"111111111",
  26240=>"000011110",
  26241=>"111111111",
  26242=>"000000000",
  26243=>"000100111",
  26244=>"110000000",
  26245=>"111111111",
  26246=>"000000111",
  26247=>"111100111",
  26248=>"000000000",
  26249=>"000000000",
  26250=>"000000000",
  26251=>"111000000",
  26252=>"110100000",
  26253=>"000000111",
  26254=>"010110111",
  26255=>"001001000",
  26256=>"111111111",
  26257=>"000000001",
  26258=>"000001001",
  26259=>"000000000",
  26260=>"000000111",
  26261=>"000010000",
  26262=>"000000000",
  26263=>"001000001",
  26264=>"111111111",
  26265=>"111111111",
  26266=>"111111111",
  26267=>"001111111",
  26268=>"000000000",
  26269=>"111111101",
  26270=>"000000000",
  26271=>"111110000",
  26272=>"110101111",
  26273=>"011111000",
  26274=>"000010000",
  26275=>"000000100",
  26276=>"000100111",
  26277=>"000110110",
  26278=>"110110000",
  26279=>"000000001",
  26280=>"000001001",
  26281=>"111111111",
  26282=>"111111111",
  26283=>"011111010",
  26284=>"100101111",
  26285=>"000000000",
  26286=>"011010000",
  26287=>"111011010",
  26288=>"000001111",
  26289=>"001001001",
  26290=>"000011010",
  26291=>"111111111",
  26292=>"110000000",
  26293=>"111111100",
  26294=>"000010000",
  26295=>"000000110",
  26296=>"000000000",
  26297=>"000000000",
  26298=>"100111111",
  26299=>"110011111",
  26300=>"001111111",
  26301=>"000000000",
  26302=>"000100011",
  26303=>"111111111",
  26304=>"011111000",
  26305=>"001011111",
  26306=>"101001001",
  26307=>"111111111",
  26308=>"000000001",
  26309=>"111110110",
  26310=>"111000000",
  26311=>"000001000",
  26312=>"111101101",
  26313=>"001101111",
  26314=>"111111111",
  26315=>"111011001",
  26316=>"110111111",
  26317=>"000111111",
  26318=>"001000110",
  26319=>"000001001",
  26320=>"100100000",
  26321=>"111110111",
  26322=>"111111111",
  26323=>"000000000",
  26324=>"000000000",
  26325=>"110100100",
  26326=>"000010011",
  26327=>"000000000",
  26328=>"010110111",
  26329=>"000000000",
  26330=>"000000101",
  26331=>"101111111",
  26332=>"100000000",
  26333=>"000000011",
  26334=>"000000000",
  26335=>"111111111",
  26336=>"111111111",
  26337=>"111101100",
  26338=>"111111000",
  26339=>"000100111",
  26340=>"000000000",
  26341=>"000000000",
  26342=>"000000000",
  26343=>"111111111",
  26344=>"001001001",
  26345=>"100100111",
  26346=>"100000000",
  26347=>"111111111",
  26348=>"100000000",
  26349=>"011011000",
  26350=>"111111111",
  26351=>"111111111",
  26352=>"110000000",
  26353=>"100100111",
  26354=>"000000000",
  26355=>"110110110",
  26356=>"100111111",
  26357=>"000000000",
  26358=>"111111111",
  26359=>"000000000",
  26360=>"100000000",
  26361=>"110110110",
  26362=>"111111111",
  26363=>"000000000",
  26364=>"111000101",
  26365=>"111111000",
  26366=>"111111111",
  26367=>"111111111",
  26368=>"101011011",
  26369=>"011000001",
  26370=>"110111110",
  26371=>"111111111",
  26372=>"111111100",
  26373=>"000000000",
  26374=>"111111111",
  26375=>"111111111",
  26376=>"000000001",
  26377=>"011011110",
  26378=>"111100100",
  26379=>"100100000",
  26380=>"000000000",
  26381=>"111111110",
  26382=>"011111111",
  26383=>"000010000",
  26384=>"001001000",
  26385=>"111000010",
  26386=>"000000111",
  26387=>"000111001",
  26388=>"000001000",
  26389=>"000000010",
  26390=>"001001000",
  26391=>"000000000",
  26392=>"001001000",
  26393=>"111111000",
  26394=>"000000000",
  26395=>"111111101",
  26396=>"011011011",
  26397=>"111111111",
  26398=>"111100000",
  26399=>"100100000",
  26400=>"110110011",
  26401=>"111000111",
  26402=>"000110011",
  26403=>"111000100",
  26404=>"000000000",
  26405=>"100011011",
  26406=>"111111111",
  26407=>"000000111",
  26408=>"111111111",
  26409=>"101111110",
  26410=>"000010010",
  26411=>"101111111",
  26412=>"000000000",
  26413=>"111111111",
  26414=>"111101111",
  26415=>"111111111",
  26416=>"111011000",
  26417=>"000000111",
  26418=>"011010010",
  26419=>"111000000",
  26420=>"111111111",
  26421=>"000000111",
  26422=>"000000100",
  26423=>"011000101",
  26424=>"111110100",
  26425=>"111110111",
  26426=>"000001111",
  26427=>"111111111",
  26428=>"111111111",
  26429=>"000010000",
  26430=>"000000000",
  26431=>"111111111",
  26432=>"111111000",
  26433=>"000000000",
  26434=>"001101111",
  26435=>"100100111",
  26436=>"001100100",
  26437=>"001000111",
  26438=>"010000000",
  26439=>"110111110",
  26440=>"111111111",
  26441=>"111111111",
  26442=>"111011000",
  26443=>"111001001",
  26444=>"000000000",
  26445=>"110100000",
  26446=>"111111111",
  26447=>"111111011",
  26448=>"000100100",
  26449=>"100000000",
  26450=>"111111000",
  26451=>"111111111",
  26452=>"111111111",
  26453=>"001001001",
  26454=>"000110110",
  26455=>"000011111",
  26456=>"111111110",
  26457=>"110111100",
  26458=>"011000001",
  26459=>"110111000",
  26460=>"001111111",
  26461=>"011011011",
  26462=>"000000000",
  26463=>"000000000",
  26464=>"101111111",
  26465=>"111111111",
  26466=>"000011111",
  26467=>"100000111",
  26468=>"111001001",
  26469=>"011111111",
  26470=>"111111000",
  26471=>"001001000",
  26472=>"111100000",
  26473=>"010010000",
  26474=>"000000000",
  26475=>"000100000",
  26476=>"111001000",
  26477=>"110110111",
  26478=>"011000000",
  26479=>"000000000",
  26480=>"000000111",
  26481=>"111111111",
  26482=>"111000000",
  26483=>"101000000",
  26484=>"111111111",
  26485=>"111111111",
  26486=>"101101101",
  26487=>"111111111",
  26488=>"110111110",
  26489=>"111010111",
  26490=>"111111111",
  26491=>"000000000",
  26492=>"000111111",
  26493=>"000000000",
  26494=>"110111111",
  26495=>"000000000",
  26496=>"011111111",
  26497=>"110111111",
  26498=>"000000000",
  26499=>"111101101",
  26500=>"111111111",
  26501=>"111110101",
  26502=>"100000000",
  26503=>"000000010",
  26504=>"000000000",
  26505=>"000000000",
  26506=>"100000111",
  26507=>"000110111",
  26508=>"000000000",
  26509=>"000000000",
  26510=>"100111011",
  26511=>"000000001",
  26512=>"011011001",
  26513=>"111010000",
  26514=>"111111000",
  26515=>"111111111",
  26516=>"000000000",
  26517=>"000110000",
  26518=>"000001000",
  26519=>"000000000",
  26520=>"111111111",
  26521=>"010011100",
  26522=>"111111111",
  26523=>"001111111",
  26524=>"111111111",
  26525=>"111111111",
  26526=>"000000000",
  26527=>"000101111",
  26528=>"111111000",
  26529=>"110110111",
  26530=>"000000110",
  26531=>"111111000",
  26532=>"111110110",
  26533=>"111111011",
  26534=>"000000000",
  26535=>"000110111",
  26536=>"000000000",
  26537=>"101111111",
  26538=>"000000100",
  26539=>"000000000",
  26540=>"000000000",
  26541=>"110000111",
  26542=>"000111111",
  26543=>"111111011",
  26544=>"000000010",
  26545=>"100100000",
  26546=>"000001111",
  26547=>"000000010",
  26548=>"111000011",
  26549=>"011000100",
  26550=>"100101111",
  26551=>"000110111",
  26552=>"110111001",
  26553=>"111110111",
  26554=>"011000000",
  26555=>"011000111",
  26556=>"111001001",
  26557=>"111111111",
  26558=>"111111111",
  26559=>"000010011",
  26560=>"000000000",
  26561=>"111111011",
  26562=>"111111111",
  26563=>"100000111",
  26564=>"001111111",
  26565=>"001001111",
  26566=>"110111111",
  26567=>"000111111",
  26568=>"111111111",
  26569=>"110110111",
  26570=>"000110110",
  26571=>"011001000",
  26572=>"010010000",
  26573=>"111111000",
  26574=>"000010110",
  26575=>"000000101",
  26576=>"111000000",
  26577=>"000000000",
  26578=>"111111111",
  26579=>"111111111",
  26580=>"110110010",
  26581=>"000000111",
  26582=>"000001011",
  26583=>"000000010",
  26584=>"111111111",
  26585=>"000110110",
  26586=>"111100000",
  26587=>"000000111",
  26588=>"001101001",
  26589=>"111111111",
  26590=>"001100111",
  26591=>"101101101",
  26592=>"000110111",
  26593=>"011011111",
  26594=>"111111001",
  26595=>"100000000",
  26596=>"110111001",
  26597=>"000000111",
  26598=>"000000000",
  26599=>"000000000",
  26600=>"000000001",
  26601=>"101111111",
  26602=>"011000100",
  26603=>"000000001",
  26604=>"111111111",
  26605=>"000000000",
  26606=>"111111111",
  26607=>"110111111",
  26608=>"000000010",
  26609=>"000110110",
  26610=>"001000000",
  26611=>"111111111",
  26612=>"000000000",
  26613=>"000011111",
  26614=>"110000000",
  26615=>"111011111",
  26616=>"000000011",
  26617=>"100000000",
  26618=>"000111101",
  26619=>"110110000",
  26620=>"000000000",
  26621=>"000001111",
  26622=>"000100110",
  26623=>"110110110",
  26624=>"010110100",
  26625=>"011011011",
  26626=>"101101001",
  26627=>"111111111",
  26628=>"011001111",
  26629=>"010000000",
  26630=>"000000111",
  26631=>"111111111",
  26632=>"111101001",
  26633=>"111111100",
  26634=>"011011111",
  26635=>"000010011",
  26636=>"000000111",
  26637=>"111010010",
  26638=>"000000001",
  26639=>"001111010",
  26640=>"000000000",
  26641=>"111101111",
  26642=>"000010000",
  26643=>"001001111",
  26644=>"111000100",
  26645=>"111111111",
  26646=>"010010000",
  26647=>"111111110",
  26648=>"001001000",
  26649=>"111101101",
  26650=>"111111111",
  26651=>"101001111",
  26652=>"000110111",
  26653=>"111110111",
  26654=>"001011110",
  26655=>"001011111",
  26656=>"010111111",
  26657=>"000000000",
  26658=>"001001001",
  26659=>"111110110",
  26660=>"000000000",
  26661=>"111111111",
  26662=>"111111111",
  26663=>"011001000",
  26664=>"010000010",
  26665=>"111111101",
  26666=>"111111111",
  26667=>"000000000",
  26668=>"111011000",
  26669=>"000111111",
  26670=>"000000111",
  26671=>"011011111",
  26672=>"000010010",
  26673=>"011101111",
  26674=>"100100111",
  26675=>"000110010",
  26676=>"000111110",
  26677=>"001001011",
  26678=>"000000000",
  26679=>"111111111",
  26680=>"111111000",
  26681=>"010111000",
  26682=>"000010000",
  26683=>"000000000",
  26684=>"100100000",
  26685=>"000100100",
  26686=>"001011111",
  26687=>"000000000",
  26688=>"010010010",
  26689=>"100111001",
  26690=>"011000001",
  26691=>"011111110",
  26692=>"110000110",
  26693=>"001001111",
  26694=>"000000110",
  26695=>"111111101",
  26696=>"001111001",
  26697=>"000000000",
  26698=>"000000000",
  26699=>"010110110",
  26700=>"000000000",
  26701=>"001000000",
  26702=>"111101000",
  26703=>"000000000",
  26704=>"111000000",
  26705=>"000110100",
  26706=>"011011011",
  26707=>"101001101",
  26708=>"000000111",
  26709=>"111011011",
  26710=>"011001000",
  26711=>"000000100",
  26712=>"001001111",
  26713=>"000000000",
  26714=>"010111111",
  26715=>"110000111",
  26716=>"100001111",
  26717=>"111111111",
  26718=>"000000000",
  26719=>"110110100",
  26720=>"000000000",
  26721=>"000000000",
  26722=>"000000011",
  26723=>"000000000",
  26724=>"000000000",
  26725=>"000000000",
  26726=>"001000000",
  26727=>"111000000",
  26728=>"011000000",
  26729=>"000000000",
  26730=>"010010011",
  26731=>"111111111",
  26732=>"000001001",
  26733=>"111111111",
  26734=>"000000000",
  26735=>"101101000",
  26736=>"111000000",
  26737=>"000101011",
  26738=>"001001111",
  26739=>"100110111",
  26740=>"101101111",
  26741=>"000000000",
  26742=>"100111111",
  26743=>"000000010",
  26744=>"000000010",
  26745=>"001000000",
  26746=>"111111111",
  26747=>"011111111",
  26748=>"001000000",
  26749=>"111111011",
  26750=>"011011010",
  26751=>"111011000",
  26752=>"100100000",
  26753=>"111111111",
  26754=>"000000101",
  26755=>"100100001",
  26756=>"111010000",
  26757=>"101000000",
  26758=>"111111111",
  26759=>"000000000",
  26760=>"000010000",
  26761=>"110100000",
  26762=>"111001101",
  26763=>"000001000",
  26764=>"111100010",
  26765=>"111111111",
  26766=>"000111110",
  26767=>"001000101",
  26768=>"111111000",
  26769=>"111111111",
  26770=>"000000000",
  26771=>"000000010",
  26772=>"110110110",
  26773=>"010001001",
  26774=>"011000000",
  26775=>"111111111",
  26776=>"111110000",
  26777=>"111111110",
  26778=>"111001100",
  26779=>"100000000",
  26780=>"110110110",
  26781=>"010010010",
  26782=>"110110000",
  26783=>"111111101",
  26784=>"000000111",
  26785=>"111111111",
  26786=>"011110110",
  26787=>"111110000",
  26788=>"000000011",
  26789=>"101111111",
  26790=>"000000000",
  26791=>"010010010",
  26792=>"000000010",
  26793=>"000000000",
  26794=>"000000000",
  26795=>"111111111",
  26796=>"000110110",
  26797=>"011001011",
  26798=>"010010000",
  26799=>"000000000",
  26800=>"000111000",
  26801=>"011110111",
  26802=>"101100100",
  26803=>"000000100",
  26804=>"111111101",
  26805=>"000000000",
  26806=>"001001001",
  26807=>"000000000",
  26808=>"000111110",
  26809=>"000000000",
  26810=>"110000100",
  26811=>"000101101",
  26812=>"111111000",
  26813=>"000000000",
  26814=>"000000000",
  26815=>"111111111",
  26816=>"010000000",
  26817=>"111110110",
  26818=>"000001000",
  26819=>"000000011",
  26820=>"000000000",
  26821=>"011010111",
  26822=>"100000000",
  26823=>"000000010",
  26824=>"111111111",
  26825=>"000000000",
  26826=>"110110110",
  26827=>"111110111",
  26828=>"011111111",
  26829=>"110110111",
  26830=>"111110110",
  26831=>"000111111",
  26832=>"111111101",
  26833=>"101101111",
  26834=>"000010000",
  26835=>"000000101",
  26836=>"000000010",
  26837=>"111111111",
  26838=>"000000000",
  26839=>"111111110",
  26840=>"101111111",
  26841=>"111111000",
  26842=>"000110110",
  26843=>"000011011",
  26844=>"111111101",
  26845=>"100111001",
  26846=>"000000000",
  26847=>"000110000",
  26848=>"000100111",
  26849=>"100100101",
  26850=>"111111111",
  26851=>"100100110",
  26852=>"111010111",
  26853=>"000000000",
  26854=>"000000000",
  26855=>"000000110",
  26856=>"000011011",
  26857=>"110110110",
  26858=>"111111111",
  26859=>"000111111",
  26860=>"000000100",
  26861=>"111000000",
  26862=>"000011000",
  26863=>"110110000",
  26864=>"111011011",
  26865=>"000100100",
  26866=>"000000000",
  26867=>"111101001",
  26868=>"000000001",
  26869=>"000011011",
  26870=>"000110101",
  26871=>"111011010",
  26872=>"000000000",
  26873=>"111111111",
  26874=>"000110100",
  26875=>"111111111",
  26876=>"111111001",
  26877=>"000000010",
  26878=>"111110111",
  26879=>"000001111",
  26880=>"011011011",
  26881=>"000000011",
  26882=>"111001000",
  26883=>"000000000",
  26884=>"111111011",
  26885=>"110010000",
  26886=>"000000000",
  26887=>"111111000",
  26888=>"000100000",
  26889=>"111111111",
  26890=>"111100000",
  26891=>"001111111",
  26892=>"000000000",
  26893=>"000100101",
  26894=>"011111110",
  26895=>"000000000",
  26896=>"000000000",
  26897=>"100000000",
  26898=>"100101111",
  26899=>"000010011",
  26900=>"000000000",
  26901=>"000011111",
  26902=>"001001001",
  26903=>"000100111",
  26904=>"111111110",
  26905=>"000000000",
  26906=>"110110110",
  26907=>"000000000",
  26908=>"010100100",
  26909=>"111011000",
  26910=>"011111111",
  26911=>"000000000",
  26912=>"001010000",
  26913=>"111111111",
  26914=>"111111111",
  26915=>"011011111",
  26916=>"000100111",
  26917=>"110111111",
  26918=>"000000100",
  26919=>"111100001",
  26920=>"000000000",
  26921=>"001000100",
  26922=>"111111111",
  26923=>"111111111",
  26924=>"011111111",
  26925=>"000000000",
  26926=>"000111000",
  26927=>"000000000",
  26928=>"001101111",
  26929=>"000000000",
  26930=>"111111111",
  26931=>"111101111",
  26932=>"111000000",
  26933=>"000000000",
  26934=>"000000000",
  26935=>"000011111",
  26936=>"000000000",
  26937=>"000000111",
  26938=>"010000100",
  26939=>"000000000",
  26940=>"000110110",
  26941=>"011111010",
  26942=>"111000000",
  26943=>"000000000",
  26944=>"000111111",
  26945=>"110111111",
  26946=>"110111111",
  26947=>"111011000",
  26948=>"111111000",
  26949=>"011111000",
  26950=>"011111111",
  26951=>"111111111",
  26952=>"000000000",
  26953=>"111001011",
  26954=>"110110010",
  26955=>"110110000",
  26956=>"110110111",
  26957=>"101111111",
  26958=>"001001000",
  26959=>"001111110",
  26960=>"000000000",
  26961=>"111101000",
  26962=>"111110110",
  26963=>"111111011",
  26964=>"000000110",
  26965=>"000000001",
  26966=>"000001111",
  26967=>"111111111",
  26968=>"000111100",
  26969=>"111111111",
  26970=>"000000001",
  26971=>"000000010",
  26972=>"101111110",
  26973=>"111000100",
  26974=>"110111000",
  26975=>"111100111",
  26976=>"111111111",
  26977=>"111111111",
  26978=>"111111001",
  26979=>"000101111",
  26980=>"110010100",
  26981=>"010010000",
  26982=>"111111111",
  26983=>"111111111",
  26984=>"111111110",
  26985=>"000111111",
  26986=>"111111111",
  26987=>"010010000",
  26988=>"001001001",
  26989=>"110111111",
  26990=>"011111111",
  26991=>"100111000",
  26992=>"111111111",
  26993=>"111000000",
  26994=>"110111011",
  26995=>"111001000",
  26996=>"101111111",
  26997=>"011011001",
  26998=>"100110011",
  26999=>"000101111",
  27000=>"111001001",
  27001=>"111111111",
  27002=>"100100000",
  27003=>"011100110",
  27004=>"000001011",
  27005=>"000000000",
  27006=>"011011010",
  27007=>"111000000",
  27008=>"000110110",
  27009=>"011011110",
  27010=>"000000000",
  27011=>"001000001",
  27012=>"001000000",
  27013=>"000000111",
  27014=>"100000000",
  27015=>"001111111",
  27016=>"010000000",
  27017=>"000111111",
  27018=>"000100000",
  27019=>"100111111",
  27020=>"000000100",
  27021=>"001011011",
  27022=>"000110111",
  27023=>"100100111",
  27024=>"000000101",
  27025=>"011000000",
  27026=>"001000010",
  27027=>"011111110",
  27028=>"000000000",
  27029=>"000000000",
  27030=>"000001011",
  27031=>"000000001",
  27032=>"000111111",
  27033=>"000000110",
  27034=>"001001110",
  27035=>"000011000",
  27036=>"001000000",
  27037=>"011000000",
  27038=>"011000010",
  27039=>"111111100",
  27040=>"111001001",
  27041=>"100100100",
  27042=>"000101111",
  27043=>"100111111",
  27044=>"010000000",
  27045=>"000000100",
  27046=>"111000000",
  27047=>"000000000",
  27048=>"000000000",
  27049=>"000111111",
  27050=>"000000001",
  27051=>"111100010",
  27052=>"111111111",
  27053=>"000010011",
  27054=>"110110111",
  27055=>"011111111",
  27056=>"000000000",
  27057=>"010111010",
  27058=>"000000000",
  27059=>"000000000",
  27060=>"110000000",
  27061=>"111011000",
  27062=>"111001101",
  27063=>"111000111",
  27064=>"110010000",
  27065=>"000000000",
  27066=>"101101111",
  27067=>"010011011",
  27068=>"000000000",
  27069=>"000111111",
  27070=>"000001000",
  27071=>"000011011",
  27072=>"111110100",
  27073=>"110111110",
  27074=>"111111111",
  27075=>"000000000",
  27076=>"111111110",
  27077=>"000111111",
  27078=>"110111111",
  27079=>"000000000",
  27080=>"000111111",
  27081=>"000011011",
  27082=>"000000000",
  27083=>"000100100",
  27084=>"110111000",
  27085=>"000000000",
  27086=>"000110000",
  27087=>"000000000",
  27088=>"000000000",
  27089=>"011011111",
  27090=>"011111111",
  27091=>"111111111",
  27092=>"001000000",
  27093=>"010110100",
  27094=>"000011111",
  27095=>"000011001",
  27096=>"000111011",
  27097=>"111110100",
  27098=>"111111111",
  27099=>"000000100",
  27100=>"111011000",
  27101=>"001001011",
  27102=>"000000000",
  27103=>"011011001",
  27104=>"110100111",
  27105=>"111111111",
  27106=>"000011001",
  27107=>"000001001",
  27108=>"000100011",
  27109=>"000000100",
  27110=>"100000000",
  27111=>"101101101",
  27112=>"111111011",
  27113=>"110111011",
  27114=>"111110100",
  27115=>"000000000",
  27116=>"010011011",
  27117=>"000000100",
  27118=>"100011111",
  27119=>"000000000",
  27120=>"111111111",
  27121=>"111111101",
  27122=>"011011011",
  27123=>"111111100",
  27124=>"110100011",
  27125=>"001001111",
  27126=>"011111010",
  27127=>"001111111",
  27128=>"000000000",
  27129=>"010010000",
  27130=>"011111111",
  27131=>"100100000",
  27132=>"000000000",
  27133=>"001001111",
  27134=>"000000111",
  27135=>"000000001",
  27136=>"000110110",
  27137=>"111000000",
  27138=>"000000000",
  27139=>"000000000",
  27140=>"000111111",
  27141=>"111011000",
  27142=>"000000000",
  27143=>"000000000",
  27144=>"111101111",
  27145=>"011111111",
  27146=>"110000000",
  27147=>"111011111",
  27148=>"000000000",
  27149=>"111010000",
  27150=>"111111011",
  27151=>"000111111",
  27152=>"100000111",
  27153=>"110110111",
  27154=>"000000000",
  27155=>"111000000",
  27156=>"000000000",
  27157=>"100111111",
  27158=>"000010010",
  27159=>"110110100",
  27160=>"000100111",
  27161=>"110000000",
  27162=>"111010000",
  27163=>"111111000",
  27164=>"110110110",
  27165=>"000000011",
  27166=>"101101111",
  27167=>"000000011",
  27168=>"010011010",
  27169=>"111111111",
  27170=>"111100001",
  27171=>"011011010",
  27172=>"100000000",
  27173=>"111111101",
  27174=>"001001111",
  27175=>"111111111",
  27176=>"110110101",
  27177=>"000000000",
  27178=>"001000000",
  27179=>"000000011",
  27180=>"111111111",
  27181=>"101111111",
  27182=>"111100110",
  27183=>"111111111",
  27184=>"000110111",
  27185=>"000000000",
  27186=>"111111100",
  27187=>"111111111",
  27188=>"111111000",
  27189=>"100110110",
  27190=>"000111000",
  27191=>"011011000",
  27192=>"000010010",
  27193=>"011010111",
  27194=>"000000000",
  27195=>"111111100",
  27196=>"011001000",
  27197=>"001000000",
  27198=>"000000000",
  27199=>"111111111",
  27200=>"000011011",
  27201=>"000000000",
  27202=>"111111000",
  27203=>"001011000",
  27204=>"110100110",
  27205=>"111111111",
  27206=>"100100110",
  27207=>"111111111",
  27208=>"110111110",
  27209=>"111111100",
  27210=>"000000011",
  27211=>"010111111",
  27212=>"000000000",
  27213=>"111000111",
  27214=>"111100110",
  27215=>"000001001",
  27216=>"100001101",
  27217=>"111111000",
  27218=>"111111000",
  27219=>"110110000",
  27220=>"111111111",
  27221=>"100000000",
  27222=>"000110110",
  27223=>"111111001",
  27224=>"001000111",
  27225=>"000110110",
  27226=>"001000000",
  27227=>"110100110",
  27228=>"000001000",
  27229=>"110000101",
  27230=>"000000000",
  27231=>"000000100",
  27232=>"000000000",
  27233=>"101000000",
  27234=>"000000000",
  27235=>"111111000",
  27236=>"000101111",
  27237=>"010011100",
  27238=>"000111111",
  27239=>"111111111",
  27240=>"111000000",
  27241=>"011000110",
  27242=>"000000011",
  27243=>"111111101",
  27244=>"100101010",
  27245=>"111110111",
  27246=>"111111000",
  27247=>"111111100",
  27248=>"111111110",
  27249=>"111111111",
  27250=>"111000000",
  27251=>"011111111",
  27252=>"111111111",
  27253=>"100100110",
  27254=>"110000000",
  27255=>"111001000",
  27256=>"111110000",
  27257=>"111011010",
  27258=>"111111111",
  27259=>"110000000",
  27260=>"011111110",
  27261=>"111000111",
  27262=>"110000110",
  27263=>"110110110",
  27264=>"000000000",
  27265=>"110100000",
  27266=>"111111111",
  27267=>"111111111",
  27268=>"111111111",
  27269=>"111000011",
  27270=>"111011001",
  27271=>"010110110",
  27272=>"111111111",
  27273=>"110001001",
  27274=>"100100100",
  27275=>"100111101",
  27276=>"011101011",
  27277=>"000010000",
  27278=>"110010010",
  27279=>"011011011",
  27280=>"000000000",
  27281=>"111111111",
  27282=>"110000000",
  27283=>"000000000",
  27284=>"111111111",
  27285=>"000001101",
  27286=>"111111111",
  27287=>"000000000",
  27288=>"111111111",
  27289=>"101101101",
  27290=>"101000000",
  27291=>"000110011",
  27292=>"000000000",
  27293=>"111111110",
  27294=>"011001000",
  27295=>"000000000",
  27296=>"111110111",
  27297=>"100110011",
  27298=>"100000000",
  27299=>"111111001",
  27300=>"000110110",
  27301=>"111100000",
  27302=>"111111111",
  27303=>"111111011",
  27304=>"000000101",
  27305=>"101000000",
  27306=>"111111111",
  27307=>"100111111",
  27308=>"001000000",
  27309=>"001001001",
  27310=>"000000000",
  27311=>"111111110",
  27312=>"000010000",
  27313=>"100010110",
  27314=>"111111010",
  27315=>"111111000",
  27316=>"111111000",
  27317=>"111100100",
  27318=>"101000000",
  27319=>"000000001",
  27320=>"111111111",
  27321=>"111111111",
  27322=>"000000100",
  27323=>"011001101",
  27324=>"111111111",
  27325=>"011001001",
  27326=>"111111001",
  27327=>"000000000",
  27328=>"110001000",
  27329=>"111111011",
  27330=>"000010011",
  27331=>"000111111",
  27332=>"000000000",
  27333=>"111011000",
  27334=>"001111111",
  27335=>"111111111",
  27336=>"001010111",
  27337=>"000011011",
  27338=>"000010010",
  27339=>"011100000",
  27340=>"010000000",
  27341=>"000000100",
  27342=>"000001011",
  27343=>"000000111",
  27344=>"000110101",
  27345=>"001111111",
  27346=>"000000000",
  27347=>"100000100",
  27348=>"000001001",
  27349=>"111000000",
  27350=>"001111111",
  27351=>"001111000",
  27352=>"000110010",
  27353=>"011001000",
  27354=>"000000000",
  27355=>"000010010",
  27356=>"001000000",
  27357=>"000000000",
  27358=>"111111111",
  27359=>"110000000",
  27360=>"110000000",
  27361=>"110000111",
  27362=>"100000100",
  27363=>"000000001",
  27364=>"110111111",
  27365=>"111111110",
  27366=>"111110111",
  27367=>"001001111",
  27368=>"111111111",
  27369=>"000100000",
  27370=>"111011000",
  27371=>"111000111",
  27372=>"000000000",
  27373=>"000000101",
  27374=>"000100000",
  27375=>"000000111",
  27376=>"011111111",
  27377=>"111111111",
  27378=>"111111101",
  27379=>"000001111",
  27380=>"000000001",
  27381=>"110110110",
  27382=>"000000000",
  27383=>"111111111",
  27384=>"000000000",
  27385=>"111111111",
  27386=>"000000000",
  27387=>"010000000",
  27388=>"111001000",
  27389=>"100000111",
  27390=>"000000111",
  27391=>"000001000",
  27392=>"111111101",
  27393=>"000011011",
  27394=>"111111010",
  27395=>"011011011",
  27396=>"110110110",
  27397=>"000000010",
  27398=>"011001111",
  27399=>"110011000",
  27400=>"000111011",
  27401=>"111111110",
  27402=>"111111111",
  27403=>"000010111",
  27404=>"110110110",
  27405=>"111111101",
  27406=>"001111100",
  27407=>"000110000",
  27408=>"000110111",
  27409=>"000101100",
  27410=>"111000000",
  27411=>"100110010",
  27412=>"000000001",
  27413=>"100101111",
  27414=>"111111000",
  27415=>"111111111",
  27416=>"001111111",
  27417=>"000100111",
  27418=>"001000000",
  27419=>"111011111",
  27420=>"111011011",
  27421=>"011011110",
  27422=>"111111111",
  27423=>"000110111",
  27424=>"011111010",
  27425=>"010111111",
  27426=>"000000000",
  27427=>"111111001",
  27428=>"000001111",
  27429=>"111111111",
  27430=>"001101101",
  27431=>"000011001",
  27432=>"111010000",
  27433=>"000011111",
  27434=>"111011111",
  27435=>"000000110",
  27436=>"110001001",
  27437=>"011111011",
  27438=>"111111000",
  27439=>"000000000",
  27440=>"000000111",
  27441=>"000000000",
  27442=>"110111111",
  27443=>"000000111",
  27444=>"110000000",
  27445=>"100000000",
  27446=>"000100111",
  27447=>"111111111",
  27448=>"111111000",
  27449=>"001101111",
  27450=>"111111111",
  27451=>"011000000",
  27452=>"000000000",
  27453=>"111111010",
  27454=>"011110110",
  27455=>"111111000",
  27456=>"000000000",
  27457=>"110000000",
  27458=>"111111101",
  27459=>"001000000",
  27460=>"111011010",
  27461=>"111101111",
  27462=>"111111111",
  27463=>"000100000",
  27464=>"111000100",
  27465=>"111111111",
  27466=>"011000000",
  27467=>"110110110",
  27468=>"111111111",
  27469=>"001011010",
  27470=>"011111111",
  27471=>"111111110",
  27472=>"101100100",
  27473=>"000000101",
  27474=>"100000111",
  27475=>"000000000",
  27476=>"000010111",
  27477=>"100100111",
  27478=>"111000001",
  27479=>"000000000",
  27480=>"000000000",
  27481=>"001111111",
  27482=>"000100000",
  27483=>"000000000",
  27484=>"111111111",
  27485=>"111111100",
  27486=>"000000001",
  27487=>"001011111",
  27488=>"000110110",
  27489=>"111110110",
  27490=>"011010111",
  27491=>"000000001",
  27492=>"000000000",
  27493=>"000000011",
  27494=>"111000000",
  27495=>"111111111",
  27496=>"011010110",
  27497=>"111111110",
  27498=>"000000000",
  27499=>"100100100",
  27500=>"111011011",
  27501=>"000001111",
  27502=>"111010000",
  27503=>"000110010",
  27504=>"111111111",
  27505=>"000000000",
  27506=>"000000000",
  27507=>"000000000",
  27508=>"000000000",
  27509=>"010010111",
  27510=>"010111111",
  27511=>"111000001",
  27512=>"000000000",
  27513=>"111111111",
  27514=>"000000111",
  27515=>"010011011",
  27516=>"000111111",
  27517=>"111111111",
  27518=>"000000001",
  27519=>"111111111",
  27520=>"010000111",
  27521=>"111111111",
  27522=>"111111111",
  27523=>"000000000",
  27524=>"111111000",
  27525=>"111111111",
  27526=>"010000000",
  27527=>"100000011",
  27528=>"111111111",
  27529=>"111001000",
  27530=>"000000101",
  27531=>"000000000",
  27532=>"010000111",
  27533=>"000000000",
  27534=>"110111111",
  27535=>"000000000",
  27536=>"111111111",
  27537=>"000001001",
  27538=>"111111111",
  27539=>"000000000",
  27540=>"011000111",
  27541=>"111111000",
  27542=>"001111111",
  27543=>"100100100",
  27544=>"000000110",
  27545=>"000010110",
  27546=>"111111111",
  27547=>"111000111",
  27548=>"000000011",
  27549=>"110000000",
  27550=>"000001000",
  27551=>"010110000",
  27552=>"101100101",
  27553=>"100100100",
  27554=>"000000000",
  27555=>"000111111",
  27556=>"111111111",
  27557=>"111001001",
  27558=>"111110111",
  27559=>"111000000",
  27560=>"111101111",
  27561=>"000000000",
  27562=>"000100001",
  27563=>"111111111",
  27564=>"000000000",
  27565=>"000010010",
  27566=>"000000010",
  27567=>"000111011",
  27568=>"000011011",
  27569=>"110110010",
  27570=>"011000000",
  27571=>"000000000",
  27572=>"000000000",
  27573=>"010010111",
  27574=>"111111011",
  27575=>"000001111",
  27576=>"111111110",
  27577=>"000000000",
  27578=>"010011011",
  27579=>"001000000",
  27580=>"001101111",
  27581=>"010100111",
  27582=>"010111111",
  27583=>"011000000",
  27584=>"111111000",
  27585=>"010011011",
  27586=>"111111111",
  27587=>"000000000",
  27588=>"001001011",
  27589=>"000111110",
  27590=>"000000110",
  27591=>"000000000",
  27592=>"000111101",
  27593=>"111110011",
  27594=>"011011111",
  27595=>"000111100",
  27596=>"111111000",
  27597=>"000000111",
  27598=>"011000000",
  27599=>"000100000",
  27600=>"000000000",
  27601=>"100101111",
  27602=>"001111111",
  27603=>"001001101",
  27604=>"000000000",
  27605=>"000000110",
  27606=>"000000000",
  27607=>"011011011",
  27608=>"000011011",
  27609=>"111011001",
  27610=>"000110111",
  27611=>"111111011",
  27612=>"011111011",
  27613=>"000000000",
  27614=>"000100000",
  27615=>"000000001",
  27616=>"000000000",
  27617=>"111110010",
  27618=>"010110000",
  27619=>"111011011",
  27620=>"111111011",
  27621=>"101001111",
  27622=>"010111110",
  27623=>"000101111",
  27624=>"110111111",
  27625=>"000000010",
  27626=>"011010000",
  27627=>"010000000",
  27628=>"100000000",
  27629=>"101101101",
  27630=>"111111111",
  27631=>"110010000",
  27632=>"000000000",
  27633=>"000000001",
  27634=>"111001000",
  27635=>"000000000",
  27636=>"000000000",
  27637=>"111111111",
  27638=>"011111111",
  27639=>"001001001",
  27640=>"000010111",
  27641=>"100100100",
  27642=>"000000000",
  27643=>"110010000",
  27644=>"010110111",
  27645=>"111111111",
  27646=>"011001001",
  27647=>"110101100",
  27648=>"000000000",
  27649=>"000000001",
  27650=>"111001000",
  27651=>"111111111",
  27652=>"001001000",
  27653=>"001000001",
  27654=>"111110000",
  27655=>"111111111",
  27656=>"000000111",
  27657=>"110000000",
  27658=>"000001001",
  27659=>"001000000",
  27660=>"001010011",
  27661=>"110100100",
  27662=>"000000000",
  27663=>"110100000",
  27664=>"000000100",
  27665=>"000000000",
  27666=>"000000000",
  27667=>"111111111",
  27668=>"000111111",
  27669=>"000111111",
  27670=>"000000110",
  27671=>"001000000",
  27672=>"011001001",
  27673=>"000000000",
  27674=>"000000000",
  27675=>"011000000",
  27676=>"111011011",
  27677=>"001001001",
  27678=>"111001111",
  27679=>"111101111",
  27680=>"111111000",
  27681=>"110110110",
  27682=>"001111111",
  27683=>"011000000",
  27684=>"010100100",
  27685=>"000110010",
  27686=>"001111111",
  27687=>"001101000",
  27688=>"110100110",
  27689=>"010011111",
  27690=>"000000000",
  27691=>"111100000",
  27692=>"111111111",
  27693=>"100100100",
  27694=>"110000001",
  27695=>"111000000",
  27696=>"111111111",
  27697=>"100100000",
  27698=>"001011111",
  27699=>"000000000",
  27700=>"000000000",
  27701=>"111000000",
  27702=>"000000100",
  27703=>"111111111",
  27704=>"000000000",
  27705=>"011011111",
  27706=>"000010000",
  27707=>"000111111",
  27708=>"111111111",
  27709=>"000000001",
  27710=>"111111100",
  27711=>"000000000",
  27712=>"011001001",
  27713=>"111111111",
  27714=>"000000000",
  27715=>"111111111",
  27716=>"111111001",
  27717=>"011111111",
  27718=>"001001000",
  27719=>"001000111",
  27720=>"011001001",
  27721=>"000000000",
  27722=>"000000000",
  27723=>"111000000",
  27724=>"000000000",
  27725=>"000000111",
  27726=>"001000000",
  27727=>"111111010",
  27728=>"000010000",
  27729=>"111111111",
  27730=>"000000000",
  27731=>"111001000",
  27732=>"000000000",
  27733=>"000100110",
  27734=>"111111111",
  27735=>"000000000",
  27736=>"010010110",
  27737=>"000000001",
  27738=>"111111111",
  27739=>"001111111",
  27740=>"000000011",
  27741=>"111100111",
  27742=>"000111000",
  27743=>"011011011",
  27744=>"000000000",
  27745=>"100000000",
  27746=>"111000100",
  27747=>"111111111",
  27748=>"000110000",
  27749=>"000000000",
  27750=>"111111111",
  27751=>"000000000",
  27752=>"000000000",
  27753=>"000000000",
  27754=>"111000000",
  27755=>"111111111",
  27756=>"111011111",
  27757=>"000000000",
  27758=>"010000110",
  27759=>"001000000",
  27760=>"101111111",
  27761=>"000000110",
  27762=>"001000001",
  27763=>"000000011",
  27764=>"111110110",
  27765=>"111111111",
  27766=>"000000000",
  27767=>"111111111",
  27768=>"111111111",
  27769=>"011111111",
  27770=>"110100101",
  27771=>"000000000",
  27772=>"011011000",
  27773=>"111111111",
  27774=>"000001000",
  27775=>"111111111",
  27776=>"000010010",
  27777=>"000000000",
  27778=>"000000011",
  27779=>"000000000",
  27780=>"100110100",
  27781=>"000010110",
  27782=>"000000000",
  27783=>"000111111",
  27784=>"111111110",
  27785=>"000000000",
  27786=>"111111111",
  27787=>"111111111",
  27788=>"000000000",
  27789=>"111111111",
  27790=>"111111110",
  27791=>"111111111",
  27792=>"000000000",
  27793=>"101100111",
  27794=>"000010111",
  27795=>"000000010",
  27796=>"011000111",
  27797=>"000100101",
  27798=>"000011010",
  27799=>"111111111",
  27800=>"000000111",
  27801=>"011000000",
  27802=>"111110111",
  27803=>"000000000",
  27804=>"110111000",
  27805=>"000000000",
  27806=>"100100000",
  27807=>"011011010",
  27808=>"011000010",
  27809=>"001000000",
  27810=>"000000000",
  27811=>"000000000",
  27812=>"111011000",
  27813=>"011111100",
  27814=>"111111111",
  27815=>"100110000",
  27816=>"000000110",
  27817=>"111111000",
  27818=>"101000000",
  27819=>"000000001",
  27820=>"110111010",
  27821=>"111001011",
  27822=>"100100000",
  27823=>"000000111",
  27824=>"111111111",
  27825=>"000000011",
  27826=>"111111111",
  27827=>"111111111",
  27828=>"111111110",
  27829=>"100111101",
  27830=>"111110110",
  27831=>"111100110",
  27832=>"000000010",
  27833=>"000000000",
  27834=>"000000000",
  27835=>"111010111",
  27836=>"000000100",
  27837=>"110010110",
  27838=>"000100100",
  27839=>"000001111",
  27840=>"111111111",
  27841=>"111111110",
  27842=>"000000100",
  27843=>"111111111",
  27844=>"000000000",
  27845=>"000000000",
  27846=>"111101000",
  27847=>"100000011",
  27848=>"000000000",
  27849=>"111111111",
  27850=>"010000001",
  27851=>"000000111",
  27852=>"000000000",
  27853=>"000010000",
  27854=>"000000000",
  27855=>"111100100",
  27856=>"001001000",
  27857=>"000000001",
  27858=>"000110100",
  27859=>"111111111",
  27860=>"011010011",
  27861=>"001000000",
  27862=>"000000111",
  27863=>"111111000",
  27864=>"110001111",
  27865=>"000000000",
  27866=>"000000000",
  27867=>"000111111",
  27868=>"001111110",
  27869=>"100101111",
  27870=>"111111111",
  27871=>"000110000",
  27872=>"010010010",
  27873=>"000000000",
  27874=>"111111111",
  27875=>"011000000",
  27876=>"010010000",
  27877=>"000011110",
  27878=>"111110110",
  27879=>"000011011",
  27880=>"000000000",
  27881=>"111111111",
  27882=>"111111100",
  27883=>"001001000",
  27884=>"000000000",
  27885=>"111011011",
  27886=>"111111011",
  27887=>"111110111",
  27888=>"000000000",
  27889=>"011010010",
  27890=>"111111000",
  27891=>"100010111",
  27892=>"111110100",
  27893=>"000100100",
  27894=>"000000000",
  27895=>"111111111",
  27896=>"111111111",
  27897=>"000000000",
  27898=>"101111000",
  27899=>"001001111",
  27900=>"001111111",
  27901=>"111001111",
  27902=>"111111100",
  27903=>"000000000",
  27904=>"000000000",
  27905=>"101001001",
  27906=>"000000000",
  27907=>"000100111",
  27908=>"011111111",
  27909=>"110110010",
  27910=>"111111111",
  27911=>"000000000",
  27912=>"001011001",
  27913=>"000011111",
  27914=>"000000100",
  27915=>"000000000",
  27916=>"000000000",
  27917=>"001000000",
  27918=>"111111000",
  27919=>"010111111",
  27920=>"111111111",
  27921=>"110111111",
  27922=>"000000001",
  27923=>"001000000",
  27924=>"000000000",
  27925=>"110111111",
  27926=>"001001001",
  27927=>"011010000",
  27928=>"111111000",
  27929=>"000011111",
  27930=>"000000111",
  27931=>"011111111",
  27932=>"000001111",
  27933=>"000000011",
  27934=>"111111111",
  27935=>"001111111",
  27936=>"000011011",
  27937=>"011111111",
  27938=>"000000000",
  27939=>"000000000",
  27940=>"000000000",
  27941=>"111111111",
  27942=>"111110101",
  27943=>"000000111",
  27944=>"111111111",
  27945=>"010011111",
  27946=>"000111111",
  27947=>"111111111",
  27948=>"001110110",
  27949=>"000000111",
  27950=>"000000010",
  27951=>"000000110",
  27952=>"111000000",
  27953=>"010110100",
  27954=>"000111111",
  27955=>"111010110",
  27956=>"000000001",
  27957=>"000000111",
  27958=>"111111001",
  27959=>"000000001",
  27960=>"000000000",
  27961=>"000000000",
  27962=>"000000000",
  27963=>"000000000",
  27964=>"111111111",
  27965=>"000000101",
  27966=>"010000010",
  27967=>"000000110",
  27968=>"111000111",
  27969=>"111101111",
  27970=>"001000000",
  27971=>"111111111",
  27972=>"111111111",
  27973=>"111111111",
  27974=>"000000000",
  27975=>"111111110",
  27976=>"000000000",
  27977=>"000000011",
  27978=>"111111111",
  27979=>"000000110",
  27980=>"110111110",
  27981=>"000000111",
  27982=>"111111000",
  27983=>"111111110",
  27984=>"000000000",
  27985=>"001000110",
  27986=>"111111111",
  27987=>"111111011",
  27988=>"100000110",
  27989=>"111111011",
  27990=>"000000100",
  27991=>"010000000",
  27992=>"111011111",
  27993=>"111111111",
  27994=>"110000110",
  27995=>"000000000",
  27996=>"110010111",
  27997=>"000000000",
  27998=>"111000110",
  27999=>"110110111",
  28000=>"000100000",
  28001=>"000000011",
  28002=>"111111111",
  28003=>"000000000",
  28004=>"111110110",
  28005=>"111111111",
  28006=>"111111011",
  28007=>"111111111",
  28008=>"101100001",
  28009=>"000000101",
  28010=>"111111111",
  28011=>"000000000",
  28012=>"000000000",
  28013=>"110000000",
  28014=>"000000000",
  28015=>"100000000",
  28016=>"000000000",
  28017=>"111111011",
  28018=>"010000000",
  28019=>"101000000",
  28020=>"000000000",
  28021=>"000000001",
  28022=>"111111111",
  28023=>"000000100",
  28024=>"111011011",
  28025=>"000011111",
  28026=>"111111111",
  28027=>"000011111",
  28028=>"111111111",
  28029=>"101110110",
  28030=>"000001001",
  28031=>"111111111",
  28032=>"011010000",
  28033=>"111111111",
  28034=>"111110111",
  28035=>"111111111",
  28036=>"001001111",
  28037=>"000000000",
  28038=>"111111000",
  28039=>"010010000",
  28040=>"000000000",
  28041=>"001001000",
  28042=>"111011000",
  28043=>"000000000",
  28044=>"111111111",
  28045=>"100100000",
  28046=>"000010000",
  28047=>"111111111",
  28048=>"000000010",
  28049=>"000000000",
  28050=>"000000000",
  28051=>"111110110",
  28052=>"111101000",
  28053=>"000010000",
  28054=>"001000000",
  28055=>"001000001",
  28056=>"011001000",
  28057=>"111111000",
  28058=>"000000000",
  28059=>"111110100",
  28060=>"111111111",
  28061=>"100100111",
  28062=>"011001000",
  28063=>"000110100",
  28064=>"000000000",
  28065=>"001001011",
  28066=>"101011111",
  28067=>"000000101",
  28068=>"110000000",
  28069=>"111111111",
  28070=>"101000111",
  28071=>"000000000",
  28072=>"000001001",
  28073=>"111111111",
  28074=>"110100100",
  28075=>"111111111",
  28076=>"000000000",
  28077=>"001011001",
  28078=>"000110111",
  28079=>"101111111",
  28080=>"111111111",
  28081=>"000000001",
  28082=>"111001100",
  28083=>"111110100",
  28084=>"111111111",
  28085=>"011011000",
  28086=>"000000000",
  28087=>"111111111",
  28088=>"000000011",
  28089=>"111111111",
  28090=>"000000000",
  28091=>"100000001",
  28092=>"111100100",
  28093=>"000000000",
  28094=>"011000000",
  28095=>"100100000",
  28096=>"000000111",
  28097=>"000001111",
  28098=>"110110010",
  28099=>"111110111",
  28100=>"111111001",
  28101=>"111110010",
  28102=>"111111111",
  28103=>"101111011",
  28104=>"001000000",
  28105=>"000000000",
  28106=>"000000011",
  28107=>"000000000",
  28108=>"111110001",
  28109=>"011001011",
  28110=>"111111110",
  28111=>"111110110",
  28112=>"111000000",
  28113=>"001011111",
  28114=>"111111111",
  28115=>"000000000",
  28116=>"000000000",
  28117=>"000000000",
  28118=>"111000000",
  28119=>"000101001",
  28120=>"111111111",
  28121=>"000000000",
  28122=>"000000011",
  28123=>"000000111",
  28124=>"000111111",
  28125=>"111000000",
  28126=>"111101111",
  28127=>"101110111",
  28128=>"111000000",
  28129=>"011011000",
  28130=>"000110111",
  28131=>"000000000",
  28132=>"110000000",
  28133=>"000000111",
  28134=>"100101111",
  28135=>"000000000",
  28136=>"001011110",
  28137=>"011011111",
  28138=>"111111111",
  28139=>"101111111",
  28140=>"011111011",
  28141=>"110110100",
  28142=>"001001011",
  28143=>"111001000",
  28144=>"010000000",
  28145=>"000000000",
  28146=>"111100100",
  28147=>"111011111",
  28148=>"110011010",
  28149=>"000100111",
  28150=>"010000000",
  28151=>"000000000",
  28152=>"000000000",
  28153=>"000000000",
  28154=>"000001000",
  28155=>"000000000",
  28156=>"001001000",
  28157=>"011111111",
  28158=>"000000000",
  28159=>"111111010",
  28160=>"010010000",
  28161=>"111111001",
  28162=>"111111111",
  28163=>"110110111",
  28164=>"011001001",
  28165=>"000000101",
  28166=>"011000111",
  28167=>"111111111",
  28168=>"000000000",
  28169=>"001001000",
  28170=>"000000000",
  28171=>"000000000",
  28172=>"111011000",
  28173=>"111111111",
  28174=>"000110111",
  28175=>"111111111",
  28176=>"111000000",
  28177=>"110111111",
  28178=>"000000000",
  28179=>"110111110",
  28180=>"000001011",
  28181=>"111001000",
  28182=>"111111100",
  28183=>"001001001",
  28184=>"111111111",
  28185=>"100111011",
  28186=>"000000100",
  28187=>"110100100",
  28188=>"000000000",
  28189=>"000000000",
  28190=>"000011111",
  28191=>"000000000",
  28192=>"101000010",
  28193=>"011111111",
  28194=>"011011011",
  28195=>"000000001",
  28196=>"111111111",
  28197=>"111111111",
  28198=>"111111111",
  28199=>"000000000",
  28200=>"111111100",
  28201=>"010110010",
  28202=>"000000000",
  28203=>"010100111",
  28204=>"001001000",
  28205=>"111111111",
  28206=>"000000000",
  28207=>"110110110",
  28208=>"100110111",
  28209=>"111111000",
  28210=>"000000001",
  28211=>"000100000",
  28212=>"111111101",
  28213=>"011001001",
  28214=>"111001110",
  28215=>"111011011",
  28216=>"000000111",
  28217=>"001011000",
  28218=>"111111111",
  28219=>"110110111",
  28220=>"000000000",
  28221=>"111111101",
  28222=>"000000000",
  28223=>"111111111",
  28224=>"111111110",
  28225=>"111111111",
  28226=>"011000000",
  28227=>"000000000",
  28228=>"111011001",
  28229=>"000000000",
  28230=>"000010111",
  28231=>"111111111",
  28232=>"110110110",
  28233=>"000111111",
  28234=>"101100101",
  28235=>"011111111",
  28236=>"000000000",
  28237=>"111111111",
  28238=>"000101100",
  28239=>"001001111",
  28240=>"101001111",
  28241=>"111111111",
  28242=>"111011010",
  28243=>"001001001",
  28244=>"001010010",
  28245=>"111111111",
  28246=>"110111100",
  28247=>"111111111",
  28248=>"000000000",
  28249=>"100000100",
  28250=>"000000110",
  28251=>"111111111",
  28252=>"011010100",
  28253=>"000000000",
  28254=>"000000011",
  28255=>"111100000",
  28256=>"000001001",
  28257=>"001000000",
  28258=>"000000000",
  28259=>"001001000",
  28260=>"000111110",
  28261=>"000000000",
  28262=>"000000000",
  28263=>"001000000",
  28264=>"000000000",
  28265=>"000100000",
  28266=>"111111111",
  28267=>"110010011",
  28268=>"000000000",
  28269=>"000000010",
  28270=>"110110111",
  28271=>"000000000",
  28272=>"000001000",
  28273=>"000110100",
  28274=>"111111100",
  28275=>"010000000",
  28276=>"111111111",
  28277=>"111001001",
  28278=>"000100000",
  28279=>"011011011",
  28280=>"000000000",
  28281=>"110000101",
  28282=>"010000000",
  28283=>"000000100",
  28284=>"000000000",
  28285=>"011001101",
  28286=>"000000000",
  28287=>"111111111",
  28288=>"001000000",
  28289=>"110111111",
  28290=>"111111100",
  28291=>"000000000",
  28292=>"000000000",
  28293=>"111111111",
  28294=>"000000000",
  28295=>"100000000",
  28296=>"111111111",
  28297=>"101100000",
  28298=>"000000000",
  28299=>"000000010",
  28300=>"000010010",
  28301=>"111000000",
  28302=>"110111000",
  28303=>"111111111",
  28304=>"000000000",
  28305=>"111000001",
  28306=>"000000000",
  28307=>"110110110",
  28308=>"111111100",
  28309=>"011111110",
  28310=>"011111111",
  28311=>"111111111",
  28312=>"000000000",
  28313=>"111111111",
  28314=>"111011111",
  28315=>"011001001",
  28316=>"111000111",
  28317=>"011000000",
  28318=>"111111111",
  28319=>"111100111",
  28320=>"000000000",
  28321=>"111111001",
  28322=>"111111111",
  28323=>"000000111",
  28324=>"010011111",
  28325=>"110111111",
  28326=>"100111111",
  28327=>"010000000",
  28328=>"010111100",
  28329=>"000000000",
  28330=>"000010000",
  28331=>"001001111",
  28332=>"111111111",
  28333=>"111110100",
  28334=>"000000000",
  28335=>"111000011",
  28336=>"000011000",
  28337=>"111111111",
  28338=>"111111111",
  28339=>"111101111",
  28340=>"111111000",
  28341=>"100111111",
  28342=>"100111111",
  28343=>"000000000",
  28344=>"111111111",
  28345=>"000000000",
  28346=>"000111110",
  28347=>"000001001",
  28348=>"000110100",
  28349=>"001000000",
  28350=>"101100100",
  28351=>"111010000",
  28352=>"111001001",
  28353=>"001001111",
  28354=>"111111111",
  28355=>"000000000",
  28356=>"000001111",
  28357=>"111111111",
  28358=>"111111111",
  28359=>"000000000",
  28360=>"110110111",
  28361=>"000000000",
  28362=>"000000000",
  28363=>"111111111",
  28364=>"111111111",
  28365=>"111111111",
  28366=>"111111101",
  28367=>"111111111",
  28368=>"000000111",
  28369=>"110010000",
  28370=>"000000000",
  28371=>"111111111",
  28372=>"000000100",
  28373=>"000001111",
  28374=>"000000000",
  28375=>"111111111",
  28376=>"110000000",
  28377=>"111111111",
  28378=>"111101000",
  28379=>"000111000",
  28380=>"111001000",
  28381=>"111111111",
  28382=>"001000100",
  28383=>"001000101",
  28384=>"111000000",
  28385=>"000000000",
  28386=>"000000000",
  28387=>"000110110",
  28388=>"111111010",
  28389=>"110111111",
  28390=>"111111111",
  28391=>"111111110",
  28392=>"110111110",
  28393=>"000110000",
  28394=>"000000000",
  28395=>"111111111",
  28396=>"011011000",
  28397=>"000000010",
  28398=>"000111111",
  28399=>"000111111",
  28400=>"111101111",
  28401=>"000010000",
  28402=>"000000000",
  28403=>"000000010",
  28404=>"111111111",
  28405=>"111011000",
  28406=>"011011000",
  28407=>"111110110",
  28408=>"000000000",
  28409=>"000000000",
  28410=>"000000000",
  28411=>"000000010",
  28412=>"111110111",
  28413=>"100010000",
  28414=>"111111111",
  28415=>"111101101",
  28416=>"011000010",
  28417=>"010110100",
  28418=>"000000000",
  28419=>"000000000",
  28420=>"111111111",
  28421=>"111111111",
  28422=>"000111111",
  28423=>"000000101",
  28424=>"000000001",
  28425=>"000000000",
  28426=>"111000110",
  28427=>"111100101",
  28428=>"001000000",
  28429=>"000000001",
  28430=>"000000100",
  28431=>"100001011",
  28432=>"011111110",
  28433=>"000000000",
  28434=>"011000000",
  28435=>"111111001",
  28436=>"111110111",
  28437=>"000000000",
  28438=>"001000001",
  28439=>"011011111",
  28440=>"000000111",
  28441=>"000000110",
  28442=>"000000100",
  28443=>"101111111",
  28444=>"001011011",
  28445=>"000000000",
  28446=>"001001111",
  28447=>"001111111",
  28448=>"000000000",
  28449=>"000000000",
  28450=>"111111111",
  28451=>"111111011",
  28452=>"000001001",
  28453=>"000000000",
  28454=>"110100110",
  28455=>"001001000",
  28456=>"000000000",
  28457=>"110110110",
  28458=>"111111111",
  28459=>"111111000",
  28460=>"110110111",
  28461=>"000000000",
  28462=>"101111111",
  28463=>"000000000",
  28464=>"111111100",
  28465=>"111011111",
  28466=>"000001001",
  28467=>"111101111",
  28468=>"000000111",
  28469=>"000000000",
  28470=>"000010111",
  28471=>"000000000",
  28472=>"010000001",
  28473=>"111111111",
  28474=>"000111111",
  28475=>"111111011",
  28476=>"000000000",
  28477=>"100100000",
  28478=>"111011100",
  28479=>"001000100",
  28480=>"011010000",
  28481=>"111111111",
  28482=>"000000000",
  28483=>"001001001",
  28484=>"111110000",
  28485=>"000000000",
  28486=>"111111100",
  28487=>"010110000",
  28488=>"000000000",
  28489=>"011011011",
  28490=>"001000000",
  28491=>"110110111",
  28492=>"000000000",
  28493=>"111110000",
  28494=>"111111111",
  28495=>"111111011",
  28496=>"000000001",
  28497=>"111111110",
  28498=>"111111101",
  28499=>"011101111",
  28500=>"000000111",
  28501=>"000010001",
  28502=>"100100100",
  28503=>"111111111",
  28504=>"111110111",
  28505=>"000000100",
  28506=>"101000000",
  28507=>"111111111",
  28508=>"010110000",
  28509=>"000000000",
  28510=>"111111111",
  28511=>"011111111",
  28512=>"111000000",
  28513=>"001111111",
  28514=>"000000001",
  28515=>"110101100",
  28516=>"000000100",
  28517=>"000000000",
  28518=>"111111101",
  28519=>"101111111",
  28520=>"110110100",
  28521=>"111110000",
  28522=>"000111000",
  28523=>"111111000",
  28524=>"111111111",
  28525=>"001000000",
  28526=>"111011011",
  28527=>"000111111",
  28528=>"000000000",
  28529=>"111111111",
  28530=>"000111011",
  28531=>"100000110",
  28532=>"110010000",
  28533=>"000000000",
  28534=>"010011110",
  28535=>"011111111",
  28536=>"000111111",
  28537=>"111000000",
  28538=>"100000000",
  28539=>"111000100",
  28540=>"111111000",
  28541=>"111111111",
  28542=>"000000000",
  28543=>"111100101",
  28544=>"000000000",
  28545=>"111111111",
  28546=>"001000000",
  28547=>"000000000",
  28548=>"000010000",
  28549=>"111111111",
  28550=>"111111111",
  28551=>"111111111",
  28552=>"000000000",
  28553=>"110100000",
  28554=>"110100111",
  28555=>"111111111",
  28556=>"111111011",
  28557=>"101011000",
  28558=>"000111111",
  28559=>"111000100",
  28560=>"000110111",
  28561=>"111111110",
  28562=>"000000001",
  28563=>"000000010",
  28564=>"111111111",
  28565=>"000000101",
  28566=>"111111111",
  28567=>"000000000",
  28568=>"111001000",
  28569=>"000000110",
  28570=>"100100100",
  28571=>"000000000",
  28572=>"000111000",
  28573=>"000000111",
  28574=>"001101111",
  28575=>"000000000",
  28576=>"001000000",
  28577=>"011010100",
  28578=>"100111110",
  28579=>"111111111",
  28580=>"111011001",
  28581=>"111111111",
  28582=>"000000000",
  28583=>"000000000",
  28584=>"000000011",
  28585=>"110111111",
  28586=>"000110111",
  28587=>"000000000",
  28588=>"000000000",
  28589=>"111101000",
  28590=>"111010011",
  28591=>"000001000",
  28592=>"111001000",
  28593=>"111110110",
  28594=>"111111111",
  28595=>"111111111",
  28596=>"000000000",
  28597=>"010111111",
  28598=>"000000100",
  28599=>"000000111",
  28600=>"000000000",
  28601=>"000000000",
  28602=>"001010001",
  28603=>"111100111",
  28604=>"000000000",
  28605=>"111000000",
  28606=>"101100000",
  28607=>"111111110",
  28608=>"000110111",
  28609=>"111111110",
  28610=>"000111111",
  28611=>"000000000",
  28612=>"000000111",
  28613=>"000110010",
  28614=>"000000000",
  28615=>"111110100",
  28616=>"000000000",
  28617=>"000000111",
  28618=>"000100100",
  28619=>"000000000",
  28620=>"000000000",
  28621=>"000000000",
  28622=>"100100111",
  28623=>"000100100",
  28624=>"000000000",
  28625=>"111111111",
  28626=>"111111000",
  28627=>"000000000",
  28628=>"010010011",
  28629=>"100110000",
  28630=>"011001111",
  28631=>"100100000",
  28632=>"000000010",
  28633=>"111000000",
  28634=>"111011000",
  28635=>"000010111",
  28636=>"000100000",
  28637=>"000000011",
  28638=>"111011000",
  28639=>"100100110",
  28640=>"000000000",
  28641=>"111111111",
  28642=>"000001111",
  28643=>"000000000",
  28644=>"000000000",
  28645=>"111111111",
  28646=>"111111101",
  28647=>"000000000",
  28648=>"000000100",
  28649=>"111000000",
  28650=>"110100000",
  28651=>"000000000",
  28652=>"000000000",
  28653=>"000000001",
  28654=>"011111111",
  28655=>"000000110",
  28656=>"000000111",
  28657=>"000101100",
  28658=>"110010111",
  28659=>"111110111",
  28660=>"111111111",
  28661=>"000011111",
  28662=>"000000000",
  28663=>"000000000",
  28664=>"000111110",
  28665=>"010000111",
  28666=>"110000000",
  28667=>"100000000",
  28668=>"000111111",
  28669=>"100000000",
  28670=>"000000000",
  28671=>"111111111",
  28672=>"111000010",
  28673=>"000000011",
  28674=>"001111111",
  28675=>"000000000",
  28676=>"110111111",
  28677=>"111111111",
  28678=>"000000000",
  28679=>"000000000",
  28680=>"000000000",
  28681=>"001011111",
  28682=>"111111111",
  28683=>"000011111",
  28684=>"000000100",
  28685=>"111111000",
  28686=>"101001001",
  28687=>"000111011",
  28688=>"111101000",
  28689=>"000000100",
  28690=>"000000000",
  28691=>"110100100",
  28692=>"111111011",
  28693=>"000000110",
  28694=>"001000000",
  28695=>"110100111",
  28696=>"111111111",
  28697=>"001001011",
  28698=>"111011011",
  28699=>"000111101",
  28700=>"000000000",
  28701=>"011000000",
  28702=>"000000100",
  28703=>"000001011",
  28704=>"111111111",
  28705=>"000100110",
  28706=>"000000000",
  28707=>"111100100",
  28708=>"000000000",
  28709=>"000000000",
  28710=>"000000000",
  28711=>"011001111",
  28712=>"001111111",
  28713=>"111111111",
  28714=>"111111111",
  28715=>"001000000",
  28716=>"100111101",
  28717=>"000001001",
  28718=>"111010110",
  28719=>"101101100",
  28720=>"111111011",
  28721=>"111001000",
  28722=>"000000000",
  28723=>"111110100",
  28724=>"000010000",
  28725=>"000000000",
  28726=>"100000000",
  28727=>"011111110",
  28728=>"000000000",
  28729=>"111011000",
  28730=>"000010111",
  28731=>"011111110",
  28732=>"111111111",
  28733=>"000111111",
  28734=>"000101111",
  28735=>"000000111",
  28736=>"101111000",
  28737=>"011100110",
  28738=>"111111111",
  28739=>"111011111",
  28740=>"100111110",
  28741=>"000100110",
  28742=>"000000000",
  28743=>"111111111",
  28744=>"001011011",
  28745=>"111000000",
  28746=>"111111111",
  28747=>"001001001",
  28748=>"111111011",
  28749=>"010010000",
  28750=>"011011111",
  28751=>"000000000",
  28752=>"000000000",
  28753=>"000000100",
  28754=>"000011011",
  28755=>"111000000",
  28756=>"111111111",
  28757=>"011011111",
  28758=>"000000000",
  28759=>"110101101",
  28760=>"000000000",
  28761=>"111111111",
  28762=>"110101111",
  28763=>"000000000",
  28764=>"111111111",
  28765=>"000111111",
  28766=>"111101000",
  28767=>"011000000",
  28768=>"111111110",
  28769=>"111111111",
  28770=>"010111011",
  28771=>"111111101",
  28772=>"001001100",
  28773=>"111111001",
  28774=>"000000011",
  28775=>"111111011",
  28776=>"000000000",
  28777=>"111111111",
  28778=>"111000000",
  28779=>"000000000",
  28780=>"111110100",
  28781=>"000011001",
  28782=>"111011101",
  28783=>"000000000",
  28784=>"010000000",
  28785=>"111101101",
  28786=>"000000010",
  28787=>"001011011",
  28788=>"111111111",
  28789=>"011001011",
  28790=>"111111111",
  28791=>"011111111",
  28792=>"000000000",
  28793=>"111111111",
  28794=>"111100100",
  28795=>"111111111",
  28796=>"100100111",
  28797=>"011111111",
  28798=>"000000000",
  28799=>"111111111",
  28800=>"000000111",
  28801=>"000000111",
  28802=>"111100000",
  28803=>"000000000",
  28804=>"000001001",
  28805=>"011011111",
  28806=>"101100000",
  28807=>"111111011",
  28808=>"001111111",
  28809=>"000110100",
  28810=>"111111111",
  28811=>"000000000",
  28812=>"000000100",
  28813=>"000111111",
  28814=>"011000001",
  28815=>"110111000",
  28816=>"111011011",
  28817=>"011111111",
  28818=>"111111101",
  28819=>"110010111",
  28820=>"111011000",
  28821=>"100101111",
  28822=>"111111111",
  28823=>"110000000",
  28824=>"110100000",
  28825=>"101111111",
  28826=>"000110100",
  28827=>"111111111",
  28828=>"111111111",
  28829=>"001011000",
  28830=>"111111000",
  28831=>"111100100",
  28832=>"110111000",
  28833=>"001111111",
  28834=>"001000011",
  28835=>"100110111",
  28836=>"110000110",
  28837=>"000011111",
  28838=>"000000100",
  28839=>"000000000",
  28840=>"000000000",
  28841=>"000000011",
  28842=>"000000000",
  28843=>"011111010",
  28844=>"001001000",
  28845=>"100010000",
  28846=>"100100010",
  28847=>"110000000",
  28848=>"111111111",
  28849=>"000000001",
  28850=>"110010010",
  28851=>"111000000",
  28852=>"000000000",
  28853=>"111111000",
  28854=>"000000000",
  28855=>"111111000",
  28856=>"111000000",
  28857=>"111111100",
  28858=>"111111100",
  28859=>"111111000",
  28860=>"111111000",
  28861=>"100000100",
  28862=>"100100111",
  28863=>"000000110",
  28864=>"111111111",
  28865=>"110000000",
  28866=>"111111111",
  28867=>"111111011",
  28868=>"111000010",
  28869=>"111111111",
  28870=>"001000111",
  28871=>"011111111",
  28872=>"000010000",
  28873=>"000000000",
  28874=>"111011111",
  28875=>"011111111",
  28876=>"111101110",
  28877=>"100101111",
  28878=>"011111000",
  28879=>"111111011",
  28880=>"000111111",
  28881=>"000000111",
  28882=>"001000011",
  28883=>"111111111",
  28884=>"100000000",
  28885=>"000000001",
  28886=>"111111111",
  28887=>"111111111",
  28888=>"111111011",
  28889=>"000000110",
  28890=>"111111111",
  28891=>"001011111",
  28892=>"111111111",
  28893=>"110000111",
  28894=>"111111010",
  28895=>"101111011",
  28896=>"000000000",
  28897=>"111111000",
  28898=>"111111100",
  28899=>"000011011",
  28900=>"111111111",
  28901=>"000000000",
  28902=>"111111111",
  28903=>"000111111",
  28904=>"111111111",
  28905=>"011111111",
  28906=>"111111111",
  28907=>"110000110",
  28908=>"011010011",
  28909=>"000000000",
  28910=>"001111111",
  28911=>"111000000",
  28912=>"111111111",
  28913=>"101111111",
  28914=>"000001000",
  28915=>"000000000",
  28916=>"000000000",
  28917=>"100110000",
  28918=>"000111111",
  28919=>"111111111",
  28920=>"000000000",
  28921=>"000011001",
  28922=>"000100000",
  28923=>"000000000",
  28924=>"000000000",
  28925=>"000000110",
  28926=>"000000000",
  28927=>"000100100",
  28928=>"111111111",
  28929=>"000000000",
  28930=>"111111111",
  28931=>"111111111",
  28932=>"111111111",
  28933=>"010111111",
  28934=>"111111111",
  28935=>"011011001",
  28936=>"000000000",
  28937=>"101000011",
  28938=>"001001001",
  28939=>"110111111",
  28940=>"111111111",
  28941=>"011101110",
  28942=>"000001110",
  28943=>"101101101",
  28944=>"000000111",
  28945=>"011010010",
  28946=>"111111111",
  28947=>"101111111",
  28948=>"001011111",
  28949=>"000000000",
  28950=>"000100100",
  28951=>"111111111",
  28952=>"000000000",
  28953=>"111010000",
  28954=>"000000000",
  28955=>"000111111",
  28956=>"000000000",
  28957=>"000000000",
  28958=>"000000000",
  28959=>"000000000",
  28960=>"000000111",
  28961=>"011011011",
  28962=>"101111111",
  28963=>"111111111",
  28964=>"110000000",
  28965=>"111111001",
  28966=>"001110000",
  28967=>"111000100",
  28968=>"000011111",
  28969=>"000000000",
  28970=>"100000011",
  28971=>"111000111",
  28972=>"110000000",
  28973=>"110100000",
  28974=>"000000101",
  28975=>"100000101",
  28976=>"111001001",
  28977=>"000000000",
  28978=>"000000000",
  28979=>"111111111",
  28980=>"111001000",
  28981=>"111001001",
  28982=>"000000011",
  28983=>"111111011",
  28984=>"110110111",
  28985=>"000000101",
  28986=>"011010000",
  28987=>"000101111",
  28988=>"000000000",
  28989=>"001000111",
  28990=>"001001011",
  28991=>"110111100",
  28992=>"001010010",
  28993=>"000000000",
  28994=>"111111101",
  28995=>"111111111",
  28996=>"111111001",
  28997=>"000000111",
  28998=>"000111111",
  28999=>"001101101",
  29000=>"001011001",
  29001=>"000110111",
  29002=>"110010000",
  29003=>"100000000",
  29004=>"111111000",
  29005=>"000000000",
  29006=>"110000000",
  29007=>"100000000",
  29008=>"000000000",
  29009=>"110010100",
  29010=>"111000001",
  29011=>"000001001",
  29012=>"111111000",
  29013=>"011001011",
  29014=>"000110100",
  29015=>"001011001",
  29016=>"111111111",
  29017=>"000000111",
  29018=>"111111111",
  29019=>"111111111",
  29020=>"000110110",
  29021=>"000000000",
  29022=>"011011111",
  29023=>"100111111",
  29024=>"111111111",
  29025=>"111111011",
  29026=>"000000001",
  29027=>"111111011",
  29028=>"000000111",
  29029=>"011001111",
  29030=>"001001000",
  29031=>"111111000",
  29032=>"000000000",
  29033=>"111111111",
  29034=>"001111101",
  29035=>"000000001",
  29036=>"000001001",
  29037=>"000000000",
  29038=>"111111111",
  29039=>"000000000",
  29040=>"000110000",
  29041=>"111001001",
  29042=>"111111111",
  29043=>"011000001",
  29044=>"000000000",
  29045=>"000000000",
  29046=>"000000000",
  29047=>"111111111",
  29048=>"000000000",
  29049=>"001111000",
  29050=>"111111010",
  29051=>"000001001",
  29052=>"001111111",
  29053=>"000110010",
  29054=>"000000000",
  29055=>"111111111",
  29056=>"100000000",
  29057=>"111111111",
  29058=>"011011011",
  29059=>"111111111",
  29060=>"001111000",
  29061=>"111111111",
  29062=>"111000111",
  29063=>"110110111",
  29064=>"001011111",
  29065=>"111111011",
  29066=>"000001111",
  29067=>"111111111",
  29068=>"001101111",
  29069=>"011000110",
  29070=>"111101111",
  29071=>"111111111",
  29072=>"110111011",
  29073=>"000100100",
  29074=>"001000010",
  29075=>"000000000",
  29076=>"000000000",
  29077=>"111111111",
  29078=>"111111111",
  29079=>"011111110",
  29080=>"000001111",
  29081=>"111111111",
  29082=>"100101111",
  29083=>"111111100",
  29084=>"000101111",
  29085=>"000000000",
  29086=>"011000000",
  29087=>"111111111",
  29088=>"000000000",
  29089=>"011011111",
  29090=>"111101001",
  29091=>"111111001",
  29092=>"001001001",
  29093=>"111111000",
  29094=>"000000111",
  29095=>"000000000",
  29096=>"111011000",
  29097=>"110111001",
  29098=>"000000000",
  29099=>"111111110",
  29100=>"000010000",
  29101=>"111101001",
  29102=>"011111000",
  29103=>"000000000",
  29104=>"111110000",
  29105=>"111111111",
  29106=>"001111000",
  29107=>"111110111",
  29108=>"110001011",
  29109=>"111111100",
  29110=>"100100100",
  29111=>"110110000",
  29112=>"111111111",
  29113=>"000000000",
  29114=>"000111011",
  29115=>"100000000",
  29116=>"000000000",
  29117=>"101101111",
  29118=>"100000000",
  29119=>"111110110",
  29120=>"111111000",
  29121=>"011000000",
  29122=>"111110111",
  29123=>"000000000",
  29124=>"111111111",
  29125=>"000000011",
  29126=>"111111111",
  29127=>"000101111",
  29128=>"110110100",
  29129=>"111111000",
  29130=>"000000100",
  29131=>"011001111",
  29132=>"111100000",
  29133=>"101111101",
  29134=>"101101011",
  29135=>"111111111",
  29136=>"001000110",
  29137=>"010000000",
  29138=>"000000110",
  29139=>"001001001",
  29140=>"111001011",
  29141=>"000110111",
  29142=>"010001000",
  29143=>"000000011",
  29144=>"111111111",
  29145=>"111111001",
  29146=>"111011011",
  29147=>"011000000",
  29148=>"001000000",
  29149=>"000000000",
  29150=>"001000011",
  29151=>"000000000",
  29152=>"000000000",
  29153=>"000100100",
  29154=>"000000011",
  29155=>"110110110",
  29156=>"100111111",
  29157=>"111111000",
  29158=>"010000000",
  29159=>"000111111",
  29160=>"011011111",
  29161=>"000000001",
  29162=>"110111111",
  29163=>"111111111",
  29164=>"110000000",
  29165=>"001111001",
  29166=>"000000000",
  29167=>"100111111",
  29168=>"000000000",
  29169=>"110000000",
  29170=>"011111111",
  29171=>"000110111",
  29172=>"000110110",
  29173=>"000101111",
  29174=>"000000000",
  29175=>"000000100",
  29176=>"111111111",
  29177=>"000111011",
  29178=>"001111111",
  29179=>"111111111",
  29180=>"000000000",
  29181=>"111111011",
  29182=>"001011011",
  29183=>"111011101",
  29184=>"000000000",
  29185=>"000000000",
  29186=>"001001000",
  29187=>"111110111",
  29188=>"010110010",
  29189=>"110110110",
  29190=>"111001101",
  29191=>"001111100",
  29192=>"000110111",
  29193=>"101001101",
  29194=>"000000000",
  29195=>"111111111",
  29196=>"100001001",
  29197=>"000000000",
  29198=>"111111111",
  29199=>"100000101",
  29200=>"000001001",
  29201=>"011001000",
  29202=>"001001101",
  29203=>"001001001",
  29204=>"111110010",
  29205=>"110111111",
  29206=>"000000000",
  29207=>"011011011",
  29208=>"111110110",
  29209=>"100001101",
  29210=>"001000111",
  29211=>"000000000",
  29212=>"100001101",
  29213=>"001000101",
  29214=>"100100100",
  29215=>"111011011",
  29216=>"000000000",
  29217=>"001001001",
  29218=>"001001111",
  29219=>"000111011",
  29220=>"000000000",
  29221=>"000001011",
  29222=>"011000000",
  29223=>"000000000",
  29224=>"100111111",
  29225=>"000010000",
  29226=>"101101001",
  29227=>"110111000",
  29228=>"000001000",
  29229=>"011001000",
  29230=>"100101111",
  29231=>"010010000",
  29232=>"101101001",
  29233=>"101001101",
  29234=>"011011011",
  29235=>"011011011",
  29236=>"001000000",
  29237=>"111001001",
  29238=>"111001001",
  29239=>"111111111",
  29240=>"000000000",
  29241=>"100010000",
  29242=>"101101101",
  29243=>"011011000",
  29244=>"101101101",
  29245=>"110000000",
  29246=>"011000001",
  29247=>"100101111",
  29248=>"110110111",
  29249=>"000000000",
  29250=>"100000000",
  29251=>"000111010",
  29252=>"000000000",
  29253=>"101100100",
  29254=>"110010000",
  29255=>"101101101",
  29256=>"000000000",
  29257=>"111011111",
  29258=>"111111111",
  29259=>"100101000",
  29260=>"111111111",
  29261=>"111111110",
  29262=>"001001001",
  29263=>"101101111",
  29264=>"000000111",
  29265=>"000110111",
  29266=>"111111111",
  29267=>"111101100",
  29268=>"101101101",
  29269=>"110110110",
  29270=>"101001001",
  29271=>"101100100",
  29272=>"110111111",
  29273=>"101101010",
  29274=>"000011000",
  29275=>"010010000",
  29276=>"010010011",
  29277=>"111101101",
  29278=>"111011111",
  29279=>"000111011",
  29280=>"000000000",
  29281=>"001000001",
  29282=>"101001001",
  29283=>"111011001",
  29284=>"001001001",
  29285=>"100000000",
  29286=>"000000100",
  29287=>"000000010",
  29288=>"111111111",
  29289=>"000000101",
  29290=>"110010000",
  29291=>"000001111",
  29292=>"010110110",
  29293=>"100000000",
  29294=>"110111101",
  29295=>"111110110",
  29296=>"001000000",
  29297=>"011111000",
  29298=>"000001111",
  29299=>"111000000",
  29300=>"111001000",
  29301=>"000000011",
  29302=>"000000000",
  29303=>"011001111",
  29304=>"111111111",
  29305=>"111111111",
  29306=>"111000001",
  29307=>"000001000",
  29308=>"100100110",
  29309=>"000001101",
  29310=>"101001000",
  29311=>"010111010",
  29312=>"111111111",
  29313=>"110110010",
  29314=>"000010100",
  29315=>"001001001",
  29316=>"111101111",
  29317=>"011000001",
  29318=>"001011000",
  29319=>"000000000",
  29320=>"110000000",
  29321=>"000101111",
  29322=>"111111111",
  29323=>"000100100",
  29324=>"010010011",
  29325=>"000000101",
  29326=>"111111111",
  29327=>"101001100",
  29328=>"100101000",
  29329=>"011111000",
  29330=>"000000001",
  29331=>"010110110",
  29332=>"110110010",
  29333=>"100100000",
  29334=>"000011001",
  29335=>"001111011",
  29336=>"001001001",
  29337=>"100111111",
  29338=>"111111001",
  29339=>"000000000",
  29340=>"110000011",
  29341=>"000000110",
  29342=>"101000100",
  29343=>"111111011",
  29344=>"110000000",
  29345=>"111111011",
  29346=>"100110111",
  29347=>"010111111",
  29348=>"110111011",
  29349=>"110100100",
  29350=>"010111111",
  29351=>"000000100",
  29352=>"010000000",
  29353=>"111111101",
  29354=>"111111111",
  29355=>"000111111",
  29356=>"111111011",
  29357=>"100110100",
  29358=>"111111111",
  29359=>"010110111",
  29360=>"010011011",
  29361=>"000100101",
  29362=>"101001001",
  29363=>"000000000",
  29364=>"011011111",
  29365=>"010000001",
  29366=>"001001101",
  29367=>"000000000",
  29368=>"100111111",
  29369=>"101111111",
  29370=>"110010001",
  29371=>"010011001",
  29372=>"110110111",
  29373=>"011000000",
  29374=>"000000000",
  29375=>"110010101",
  29376=>"000001001",
  29377=>"000000000",
  29378=>"111100100",
  29379=>"111000000",
  29380=>"101101101",
  29381=>"011000111",
  29382=>"111111000",
  29383=>"110110110",
  29384=>"000111011",
  29385=>"000000000",
  29386=>"110111000",
  29387=>"000000101",
  29388=>"110111111",
  29389=>"000000000",
  29390=>"001001001",
  29391=>"000000001",
  29392=>"000010110",
  29393=>"001001000",
  29394=>"111111110",
  29395=>"000000010",
  29396=>"111111111",
  29397=>"100000110",
  29398=>"001001100",
  29399=>"110110010",
  29400=>"110010000",
  29401=>"100000101",
  29402=>"000000000",
  29403=>"111100101",
  29404=>"110010110",
  29405=>"101111111",
  29406=>"010110010",
  29407=>"111100100",
  29408=>"001100000",
  29409=>"000000000",
  29410=>"011000010",
  29411=>"111111101",
  29412=>"111110110",
  29413=>"011010010",
  29414=>"101001101",
  29415=>"100000000",
  29416=>"100000000",
  29417=>"101100001",
  29418=>"111111111",
  29419=>"111111111",
  29420=>"111101101",
  29421=>"111010000",
  29422=>"111111101",
  29423=>"001101000",
  29424=>"000000001",
  29425=>"111111111",
  29426=>"010010010",
  29427=>"011001111",
  29428=>"000000000",
  29429=>"000000110",
  29430=>"011011011",
  29431=>"100000000",
  29432=>"111010000",
  29433=>"000001001",
  29434=>"100101101",
  29435=>"000100100",
  29436=>"001001001",
  29437=>"000000100",
  29438=>"111110010",
  29439=>"101000000",
  29440=>"110111101",
  29441=>"100100100",
  29442=>"100100100",
  29443=>"110110110",
  29444=>"011010011",
  29445=>"000000110",
  29446=>"001101001",
  29447=>"000111010",
  29448=>"000000000",
  29449=>"001001101",
  29450=>"110111000",
  29451=>"001001111",
  29452=>"000000001",
  29453=>"111111011",
  29454=>"000000000",
  29455=>"000100000",
  29456=>"000000101",
  29457=>"110111000",
  29458=>"000000110",
  29459=>"011111111",
  29460=>"111111111",
  29461=>"100000000",
  29462=>"100100100",
  29463=>"110110110",
  29464=>"111111111",
  29465=>"100100111",
  29466=>"110010010",
  29467=>"000011000",
  29468=>"100000001",
  29469=>"010000000",
  29470=>"000100111",
  29471=>"000001000",
  29472=>"111111011",
  29473=>"000010010",
  29474=>"100000100",
  29475=>"001001011",
  29476=>"001011011",
  29477=>"000111111",
  29478=>"000000100",
  29479=>"110110111",
  29480=>"000000100",
  29481=>"111101111",
  29482=>"101100101",
  29483=>"101101101",
  29484=>"010000000",
  29485=>"001001000",
  29486=>"111111000",
  29487=>"101101101",
  29488=>"110100100",
  29489=>"110010010",
  29490=>"001011011",
  29491=>"110010010",
  29492=>"000010010",
  29493=>"000100000",
  29494=>"110111110",
  29495=>"000001011",
  29496=>"010010111",
  29497=>"000100100",
  29498=>"110000000",
  29499=>"001001101",
  29500=>"110111011",
  29501=>"110100101",
  29502=>"110110110",
  29503=>"110111010",
  29504=>"000000000",
  29505=>"001101111",
  29506=>"101001000",
  29507=>"101101101",
  29508=>"101001001",
  29509=>"000101101",
  29510=>"100001101",
  29511=>"101101101",
  29512=>"101100000",
  29513=>"111110010",
  29514=>"000000010",
  29515=>"000000000",
  29516=>"010010000",
  29517=>"111111111",
  29518=>"101101111",
  29519=>"000000100",
  29520=>"100000000",
  29521=>"010010010",
  29522=>"111111111",
  29523=>"000000010",
  29524=>"111101101",
  29525=>"001011001",
  29526=>"010110101",
  29527=>"111111111",
  29528=>"001001001",
  29529=>"011010000",
  29530=>"000100100",
  29531=>"000001001",
  29532=>"011011011",
  29533=>"110110110",
  29534=>"000000001",
  29535=>"000000011",
  29536=>"111111111",
  29537=>"100000001",
  29538=>"011011011",
  29539=>"001001000",
  29540=>"011001011",
  29541=>"000000010",
  29542=>"000000111",
  29543=>"110110110",
  29544=>"001001101",
  29545=>"000000000",
  29546=>"110110011",
  29547=>"000010000",
  29548=>"100110110",
  29549=>"111111011",
  29550=>"000000000",
  29551=>"110000000",
  29552=>"111101000",
  29553=>"110000100",
  29554=>"000000001",
  29555=>"111111111",
  29556=>"100000000",
  29557=>"101101101",
  29558=>"110110011",
  29559=>"000000000",
  29560=>"100000000",
  29561=>"011000000",
  29562=>"110110010",
  29563=>"110110110",
  29564=>"110110110",
  29565=>"111011111",
  29566=>"000000011",
  29567=>"101000000",
  29568=>"000000101",
  29569=>"100010001",
  29570=>"100100100",
  29571=>"010110010",
  29572=>"000000010",
  29573=>"010010000",
  29574=>"001011011",
  29575=>"000000011",
  29576=>"001000000",
  29577=>"111110111",
  29578=>"100100100",
  29579=>"011011000",
  29580=>"111111010",
  29581=>"000101101",
  29582=>"000011101",
  29583=>"001001001",
  29584=>"010011010",
  29585=>"000000001",
  29586=>"110110111",
  29587=>"111010110",
  29588=>"000000000",
  29589=>"000010010",
  29590=>"011110110",
  29591=>"100000100",
  29592=>"111111000",
  29593=>"000000110",
  29594=>"001001101",
  29595=>"111111111",
  29596=>"000010010",
  29597=>"111111000",
  29598=>"100100111",
  29599=>"100000000",
  29600=>"000000000",
  29601=>"001011111",
  29602=>"111001000",
  29603=>"000001000",
  29604=>"001000001",
  29605=>"011111101",
  29606=>"111101000",
  29607=>"000110000",
  29608=>"010010010",
  29609=>"101111111",
  29610=>"100001001",
  29611=>"010010000",
  29612=>"010110000",
  29613=>"110111111",
  29614=>"100000111",
  29615=>"110000010",
  29616=>"111100101",
  29617=>"000001001",
  29618=>"000000100",
  29619=>"100110110",
  29620=>"000010000",
  29621=>"000000111",
  29622=>"111111011",
  29623=>"000100100",
  29624=>"110110110",
  29625=>"010010110",
  29626=>"100100100",
  29627=>"100111111",
  29628=>"111111111",
  29629=>"110110110",
  29630=>"001011000",
  29631=>"100100100",
  29632=>"111111111",
  29633=>"001001000",
  29634=>"001101101",
  29635=>"111111000",
  29636=>"111111001",
  29637=>"101101001",
  29638=>"110110110",
  29639=>"001111100",
  29640=>"011011001",
  29641=>"001001101",
  29642=>"000000100",
  29643=>"111011000",
  29644=>"110110000",
  29645=>"000000000",
  29646=>"110110110",
  29647=>"010000000",
  29648=>"011011011",
  29649=>"111101101",
  29650=>"110110000",
  29651=>"111111111",
  29652=>"001000001",
  29653=>"010010010",
  29654=>"110110110",
  29655=>"001000101",
  29656=>"000001001",
  29657=>"110000100",
  29658=>"000011111",
  29659=>"111111111",
  29660=>"111001001",
  29661=>"111001000",
  29662=>"111111100",
  29663=>"110100110",
  29664=>"111011111",
  29665=>"110111111",
  29666=>"111000101",
  29667=>"000000000",
  29668=>"110010111",
  29669=>"010010010",
  29670=>"101000000",
  29671=>"000000010",
  29672=>"110110110",
  29673=>"111111111",
  29674=>"000110011",
  29675=>"011111111",
  29676=>"000010000",
  29677=>"110011011",
  29678=>"001101101",
  29679=>"011010010",
  29680=>"100000100",
  29681=>"110010110",
  29682=>"101101111",
  29683=>"000000000",
  29684=>"111111101",
  29685=>"000010110",
  29686=>"111111101",
  29687=>"101111111",
  29688=>"010010000",
  29689=>"010000001",
  29690=>"000000111",
  29691=>"101000000",
  29692=>"011111111",
  29693=>"010010011",
  29694=>"110100000",
  29695=>"101101111",
  29696=>"111111111",
  29697=>"111111111",
  29698=>"101111001",
  29699=>"001011001",
  29700=>"001111011",
  29701=>"000011111",
  29702=>"000011011",
  29703=>"111111111",
  29704=>"110010011",
  29705=>"000000110",
  29706=>"111111111",
  29707=>"111111111",
  29708=>"000000100",
  29709=>"000000000",
  29710=>"111111111",
  29711=>"000000000",
  29712=>"111111111",
  29713=>"001111111",
  29714=>"000000000",
  29715=>"111111111",
  29716=>"111111111",
  29717=>"000000101",
  29718=>"000000000",
  29719=>"001101111",
  29720=>"011111111",
  29721=>"000000100",
  29722=>"111111010",
  29723=>"000000100",
  29724=>"110110110",
  29725=>"111111101",
  29726=>"000000000",
  29727=>"110111111",
  29728=>"000001011",
  29729=>"100110111",
  29730=>"100100010",
  29731=>"111111111",
  29732=>"001101001",
  29733=>"100011000",
  29734=>"111111111",
  29735=>"000000000",
  29736=>"000001011",
  29737=>"111110000",
  29738=>"000000000",
  29739=>"111110111",
  29740=>"000110111",
  29741=>"111111111",
  29742=>"111111111",
  29743=>"111111100",
  29744=>"000011000",
  29745=>"000000000",
  29746=>"111111111",
  29747=>"000110000",
  29748=>"000000000",
  29749=>"011011111",
  29750=>"111011001",
  29751=>"000011010",
  29752=>"110111111",
  29753=>"000010011",
  29754=>"000000000",
  29755=>"000000011",
  29756=>"111111110",
  29757=>"000000000",
  29758=>"101000000",
  29759=>"111111111",
  29760=>"111011011",
  29761=>"111001111",
  29762=>"000000111",
  29763=>"000000010",
  29764=>"000100100",
  29765=>"110110110",
  29766=>"110000101",
  29767=>"001000010",
  29768=>"000010011",
  29769=>"000000100",
  29770=>"101110111",
  29771=>"100100000",
  29772=>"111111111",
  29773=>"011000110",
  29774=>"111000111",
  29775=>"000000000",
  29776=>"111111000",
  29777=>"000000000",
  29778=>"111011001",
  29779=>"111110010",
  29780=>"000001111",
  29781=>"000111011",
  29782=>"111111111",
  29783=>"110010000",
  29784=>"000000000",
  29785=>"110111111",
  29786=>"101000010",
  29787=>"100001000",
  29788=>"000110110",
  29789=>"000000010",
  29790=>"010010000",
  29791=>"111111110",
  29792=>"000000000",
  29793=>"111000000",
  29794=>"011111100",
  29795=>"000000010",
  29796=>"100110000",
  29797=>"111111111",
  29798=>"100100100",
  29799=>"000000000",
  29800=>"110111111",
  29801=>"111010000",
  29802=>"111000000",
  29803=>"111001000",
  29804=>"111111011",
  29805=>"111111011",
  29806=>"100100100",
  29807=>"111111111",
  29808=>"110010010",
  29809=>"000110010",
  29810=>"111111011",
  29811=>"000001001",
  29812=>"111111110",
  29813=>"001100100",
  29814=>"111000000",
  29815=>"111111010",
  29816=>"011011010",
  29817=>"000000100",
  29818=>"000000000",
  29819=>"111111111",
  29820=>"001000000",
  29821=>"111011111",
  29822=>"000000000",
  29823=>"011111000",
  29824=>"111001111",
  29825=>"111110111",
  29826=>"000000000",
  29827=>"100100000",
  29828=>"000000000",
  29829=>"111111111",
  29830=>"000000110",
  29831=>"101111111",
  29832=>"011111111",
  29833=>"001000000",
  29834=>"000000000",
  29835=>"000000000",
  29836=>"000001001",
  29837=>"000000000",
  29838=>"000001000",
  29839=>"000000000",
  29840=>"000000000",
  29841=>"111111011",
  29842=>"111111111",
  29843=>"110010111",
  29844=>"001000011",
  29845=>"000000111",
  29846=>"111111111",
  29847=>"111000000",
  29848=>"111111111",
  29849=>"001001100",
  29850=>"000000000",
  29851=>"111101111",
  29852=>"100000000",
  29853=>"000000000",
  29854=>"100000000",
  29855=>"011111111",
  29856=>"111010011",
  29857=>"000000000",
  29858=>"000111011",
  29859=>"000000000",
  29860=>"001001100",
  29861=>"000000000",
  29862=>"000011010",
  29863=>"000000001",
  29864=>"111010111",
  29865=>"000000110",
  29866=>"111111111",
  29867=>"110110111",
  29868=>"000000010",
  29869=>"100100100",
  29870=>"101010110",
  29871=>"101111111",
  29872=>"000000101",
  29873=>"000000000",
  29874=>"011011011",
  29875=>"111111000",
  29876=>"111011111",
  29877=>"111111000",
  29878=>"111111111",
  29879=>"110000101",
  29880=>"000000000",
  29881=>"001001011",
  29882=>"111111011",
  29883=>"100010111",
  29884=>"000000000",
  29885=>"000000000",
  29886=>"111111111",
  29887=>"001001001",
  29888=>"111111110",
  29889=>"110111111",
  29890=>"000111111",
  29891=>"111111111",
  29892=>"111110010",
  29893=>"110111111",
  29894=>"100100000",
  29895=>"100111111",
  29896=>"111001011",
  29897=>"000000000",
  29898=>"000000101",
  29899=>"111111011",
  29900=>"111111111",
  29901=>"010111001",
  29902=>"001000111",
  29903=>"011000000",
  29904=>"011111111",
  29905=>"011001011",
  29906=>"111111010",
  29907=>"001100111",
  29908=>"110111000",
  29909=>"000000010",
  29910=>"110111111",
  29911=>"001010111",
  29912=>"111111111",
  29913=>"100010001",
  29914=>"111111000",
  29915=>"111111111",
  29916=>"101101101",
  29917=>"111111100",
  29918=>"111111010",
  29919=>"100111111",
  29920=>"111111111",
  29921=>"111111111",
  29922=>"000000000",
  29923=>"111001000",
  29924=>"101000111",
  29925=>"000000100",
  29926=>"111111110",
  29927=>"111011001",
  29928=>"000000000",
  29929=>"100110000",
  29930=>"111111111",
  29931=>"111000111",
  29932=>"000011000",
  29933=>"001111111",
  29934=>"111111111",
  29935=>"111111000",
  29936=>"111111001",
  29937=>"110000000",
  29938=>"001000000",
  29939=>"000000000",
  29940=>"000000000",
  29941=>"111111000",
  29942=>"100110010",
  29943=>"010000001",
  29944=>"000000000",
  29945=>"111111111",
  29946=>"111111110",
  29947=>"000010111",
  29948=>"011001000",
  29949=>"111111111",
  29950=>"110000000",
  29951=>"001011111",
  29952=>"000000000",
  29953=>"111110110",
  29954=>"000000000",
  29955=>"000110111",
  29956=>"000000000",
  29957=>"111111111",
  29958=>"100000111",
  29959=>"111101111",
  29960=>"110110111",
  29961=>"001001111",
  29962=>"111111000",
  29963=>"110110100",
  29964=>"000000001",
  29965=>"111000000",
  29966=>"010011100",
  29967=>"111000101",
  29968=>"111001000",
  29969=>"111111111",
  29970=>"111111010",
  29971=>"010000000",
  29972=>"111101100",
  29973=>"111001100",
  29974=>"000100000",
  29975=>"010111111",
  29976=>"000010010",
  29977=>"111111111",
  29978=>"001011011",
  29979=>"111111111",
  29980=>"001011111",
  29981=>"000001000",
  29982=>"000111111",
  29983=>"111111111",
  29984=>"110110110",
  29985=>"001100100",
  29986=>"011000000",
  29987=>"000000000",
  29988=>"000000000",
  29989=>"101001001",
  29990=>"000011011",
  29991=>"111110000",
  29992=>"111111111",
  29993=>"000000000",
  29994=>"000010010",
  29995=>"111111101",
  29996=>"000000000",
  29997=>"000000000",
  29998=>"111111111",
  29999=>"000000000",
  30000=>"111111111",
  30001=>"111111111",
  30002=>"000000000",
  30003=>"000000011",
  30004=>"111111111",
  30005=>"000000000",
  30006=>"010010000",
  30007=>"110000000",
  30008=>"111111111",
  30009=>"000000000",
  30010=>"011011000",
  30011=>"111111111",
  30012=>"100000100",
  30013=>"111110110",
  30014=>"000100111",
  30015=>"111111010",
  30016=>"100100101",
  30017=>"000000010",
  30018=>"111111111",
  30019=>"111111111",
  30020=>"001011011",
  30021=>"000011111",
  30022=>"111111111",
  30023=>"001001011",
  30024=>"000000000",
  30025=>"111111111",
  30026=>"001001111",
  30027=>"011011011",
  30028=>"111111000",
  30029=>"011010010",
  30030=>"100000000",
  30031=>"010000000",
  30032=>"000001000",
  30033=>"111111111",
  30034=>"000000000",
  30035=>"110110000",
  30036=>"000000000",
  30037=>"000000000",
  30038=>"001111011",
  30039=>"111111110",
  30040=>"111111000",
  30041=>"000010010",
  30042=>"000000000",
  30043=>"111111111",
  30044=>"000000000",
  30045=>"000000000",
  30046=>"000000000",
  30047=>"100110110",
  30048=>"000100111",
  30049=>"001011011",
  30050=>"111000011",
  30051=>"111111111",
  30052=>"001111010",
  30053=>"000110010",
  30054=>"111111101",
  30055=>"100100100",
  30056=>"000111110",
  30057=>"111110010",
  30058=>"011000000",
  30059=>"111111111",
  30060=>"011000110",
  30061=>"000001000",
  30062=>"111110000",
  30063=>"111111011",
  30064=>"000000000",
  30065=>"111111111",
  30066=>"000000000",
  30067=>"100000000",
  30068=>"111111111",
  30069=>"001000000",
  30070=>"010000000",
  30071=>"101000001",
  30072=>"000001011",
  30073=>"000000000",
  30074=>"000000100",
  30075=>"000000000",
  30076=>"111111111",
  30077=>"111110000",
  30078=>"111000000",
  30079=>"111100100",
  30080=>"111111111",
  30081=>"000000001",
  30082=>"011011111",
  30083=>"000000000",
  30084=>"000110110",
  30085=>"000000000",
  30086=>"000001000",
  30087=>"111101111",
  30088=>"000000000",
  30089=>"100110110",
  30090=>"110110100",
  30091=>"001000000",
  30092=>"000000000",
  30093=>"110111111",
  30094=>"111111000",
  30095=>"111111111",
  30096=>"000000000",
  30097=>"111111111",
  30098=>"000000000",
  30099=>"000000000",
  30100=>"000000000",
  30101=>"110111111",
  30102=>"000000000",
  30103=>"001001111",
  30104=>"000000111",
  30105=>"111111001",
  30106=>"100111111",
  30107=>"000010010",
  30108=>"000000010",
  30109=>"011010010",
  30110=>"000001001",
  30111=>"011010110",
  30112=>"001000111",
  30113=>"000000000",
  30114=>"100111111",
  30115=>"111111000",
  30116=>"100010000",
  30117=>"111111000",
  30118=>"000000000",
  30119=>"000000111",
  30120=>"111111111",
  30121=>"111111000",
  30122=>"100000000",
  30123=>"000001001",
  30124=>"111111111",
  30125=>"111011111",
  30126=>"000000001",
  30127=>"111111110",
  30128=>"111111011",
  30129=>"111111111",
  30130=>"001000000",
  30131=>"100110110",
  30132=>"000000110",
  30133=>"101111111",
  30134=>"111111111",
  30135=>"111111101",
  30136=>"111111111",
  30137=>"111111111",
  30138=>"000000000",
  30139=>"000000001",
  30140=>"111111011",
  30141=>"101111110",
  30142=>"000000100",
  30143=>"100000000",
  30144=>"000000000",
  30145=>"110111111",
  30146=>"111111011",
  30147=>"111111110",
  30148=>"111111111",
  30149=>"111110100",
  30150=>"111110010",
  30151=>"001100110",
  30152=>"000000000",
  30153=>"111111000",
  30154=>"101111111",
  30155=>"111111111",
  30156=>"010011111",
  30157=>"000011000",
  30158=>"111111111",
  30159=>"111011000",
  30160=>"001000001",
  30161=>"000000000",
  30162=>"111111111",
  30163=>"111111111",
  30164=>"101101111",
  30165=>"111111010",
  30166=>"111111010",
  30167=>"000000000",
  30168=>"111111111",
  30169=>"111000000",
  30170=>"000000000",
  30171=>"110010000",
  30172=>"011111111",
  30173=>"001111111",
  30174=>"111111111",
  30175=>"110100000",
  30176=>"111100000",
  30177=>"000011111",
  30178=>"100100000",
  30179=>"111111010",
  30180=>"111111111",
  30181=>"001001111",
  30182=>"110111111",
  30183=>"000000000",
  30184=>"100110110",
  30185=>"101111110",
  30186=>"111111111",
  30187=>"000111111",
  30188=>"111111111",
  30189=>"100111111",
  30190=>"100111111",
  30191=>"001111110",
  30192=>"000011000",
  30193=>"111000101",
  30194=>"000010110",
  30195=>"111111111",
  30196=>"000110000",
  30197=>"001111001",
  30198=>"111000000",
  30199=>"000000000",
  30200=>"111111111",
  30201=>"000001011",
  30202=>"111110110",
  30203=>"100110110",
  30204=>"111111111",
  30205=>"111110001",
  30206=>"111111111",
  30207=>"101000111",
  30208=>"011111111",
  30209=>"000000011",
  30210=>"111000111",
  30211=>"110111111",
  30212=>"000000111",
  30213=>"111000000",
  30214=>"111111000",
  30215=>"111111111",
  30216=>"000000000",
  30217=>"110000000",
  30218=>"000000000",
  30219=>"000010010",
  30220=>"000011001",
  30221=>"111111010",
  30222=>"111111111",
  30223=>"001111111",
  30224=>"001000000",
  30225=>"111111110",
  30226=>"100000101",
  30227=>"000000001",
  30228=>"000000000",
  30229=>"000000000",
  30230=>"000001101",
  30231=>"011000000",
  30232=>"011111111",
  30233=>"100100111",
  30234=>"111000110",
  30235=>"001000000",
  30236=>"011111111",
  30237=>"000000000",
  30238=>"111111011",
  30239=>"111110000",
  30240=>"111101000",
  30241=>"111100000",
  30242=>"111111111",
  30243=>"111111111",
  30244=>"111100000",
  30245=>"100111111",
  30246=>"111111111",
  30247=>"100111111",
  30248=>"111111000",
  30249=>"000000000",
  30250=>"111111111",
  30251=>"111111000",
  30252=>"000000000",
  30253=>"111111111",
  30254=>"111001001",
  30255=>"111110111",
  30256=>"010111000",
  30257=>"111010000",
  30258=>"100000000",
  30259=>"011000011",
  30260=>"000101111",
  30261=>"000000000",
  30262=>"000000000",
  30263=>"110111001",
  30264=>"000000000",
  30265=>"011000000",
  30266=>"111001001",
  30267=>"111111000",
  30268=>"000000111",
  30269=>"110111001",
  30270=>"111111110",
  30271=>"000000001",
  30272=>"111111111",
  30273=>"000000000",
  30274=>"111000000",
  30275=>"111010111",
  30276=>"111111011",
  30277=>"000000111",
  30278=>"000000110",
  30279=>"111111110",
  30280=>"111111111",
  30281=>"000000100",
  30282=>"110101111",
  30283=>"000111111",
  30284=>"110110000",
  30285=>"011000000",
  30286=>"000000000",
  30287=>"111111000",
  30288=>"001000000",
  30289=>"101000000",
  30290=>"000000000",
  30291=>"000111000",
  30292=>"000000000",
  30293=>"000000000",
  30294=>"000011111",
  30295=>"000101111",
  30296=>"001000000",
  30297=>"101000111",
  30298=>"000000000",
  30299=>"111000000",
  30300=>"001000000",
  30301=>"000110000",
  30302=>"111111110",
  30303=>"111111000",
  30304=>"110110000",
  30305=>"000000000",
  30306=>"000000000",
  30307=>"000010111",
  30308=>"100000010",
  30309=>"001011110",
  30310=>"000111110",
  30311=>"111111111",
  30312=>"111000000",
  30313=>"101101001",
  30314=>"111000111",
  30315=>"000111011",
  30316=>"110111110",
  30317=>"111000000",
  30318=>"111111110",
  30319=>"000100110",
  30320=>"111000011",
  30321=>"001111111",
  30322=>"100000100",
  30323=>"111111001",
  30324=>"111101000",
  30325=>"001001001",
  30326=>"111100000",
  30327=>"110100000",
  30328=>"000101110",
  30329=>"111111011",
  30330=>"000000000",
  30331=>"000000000",
  30332=>"110110110",
  30333=>"000000111",
  30334=>"101000000",
  30335=>"111111111",
  30336=>"111000111",
  30337=>"000000000",
  30338=>"001001001",
  30339=>"000111000",
  30340=>"111000010",
  30341=>"101000111",
  30342=>"111110000",
  30343=>"001000000",
  30344=>"000000000",
  30345=>"000000101",
  30346=>"000010000",
  30347=>"111000111",
  30348=>"001101100",
  30349=>"000100100",
  30350=>"100000000",
  30351=>"111111111",
  30352=>"000000010",
  30353=>"111111000",
  30354=>"111000000",
  30355=>"111111000",
  30356=>"001111000",
  30357=>"000000111",
  30358=>"011111111",
  30359=>"111111111",
  30360=>"000000101",
  30361=>"000000000",
  30362=>"011001011",
  30363=>"111111000",
  30364=>"101111111",
  30365=>"000000000",
  30366=>"000010011",
  30367=>"000000001",
  30368=>"000000000",
  30369=>"001000000",
  30370=>"000000111",
  30371=>"000000000",
  30372=>"010010110",
  30373=>"000111111",
  30374=>"011111101",
  30375=>"111010001",
  30376=>"110111010",
  30377=>"000000000",
  30378=>"000010111",
  30379=>"000000110",
  30380=>"111111000",
  30381=>"111000000",
  30382=>"000000000",
  30383=>"000110000",
  30384=>"110111001",
  30385=>"111111011",
  30386=>"111111011",
  30387=>"110101111",
  30388=>"111111000",
  30389=>"101100100",
  30390=>"000000000",
  30391=>"000000111",
  30392=>"000000101",
  30393=>"111111111",
  30394=>"111011001",
  30395=>"010000000",
  30396=>"111111010",
  30397=>"111111111",
  30398=>"100000100",
  30399=>"001000000",
  30400=>"010111111",
  30401=>"001001111",
  30402=>"111111111",
  30403=>"000111111",
  30404=>"111111111",
  30405=>"000111111",
  30406=>"011111001",
  30407=>"000000000",
  30408=>"000000001",
  30409=>"110111110",
  30410=>"000000110",
  30411=>"111111000",
  30412=>"000000100",
  30413=>"111111111",
  30414=>"111111000",
  30415=>"111011100",
  30416=>"011000000",
  30417=>"000000000",
  30418=>"111100000",
  30419=>"000000000",
  30420=>"000000111",
  30421=>"110100100",
  30422=>"110010000",
  30423=>"101101000",
  30424=>"000000001",
  30425=>"111111100",
  30426=>"000000000",
  30427=>"010111100",
  30428=>"111100000",
  30429=>"100110111",
  30430=>"000000000",
  30431=>"000111111",
  30432=>"000000001",
  30433=>"111011000",
  30434=>"111000000",
  30435=>"001000000",
  30436=>"111000001",
  30437=>"111100001",
  30438=>"000001100",
  30439=>"000110000",
  30440=>"000000111",
  30441=>"101000111",
  30442=>"111000100",
  30443=>"111111000",
  30444=>"000000001",
  30445=>"000000000",
  30446=>"011011010",
  30447=>"000111111",
  30448=>"010100111",
  30449=>"000000111",
  30450=>"000000101",
  30451=>"000000111",
  30452=>"001100111",
  30453=>"111111000",
  30454=>"011011000",
  30455=>"010010000",
  30456=>"110110111",
  30457=>"111111000",
  30458=>"011111111",
  30459=>"001001000",
  30460=>"000100110",
  30461=>"000000111",
  30462=>"111000000",
  30463=>"111000000",
  30464=>"000000000",
  30465=>"000000011",
  30466=>"111111110",
  30467=>"111110000",
  30468=>"111111000",
  30469=>"000000000",
  30470=>"111111101",
  30471=>"111101111",
  30472=>"111000000",
  30473=>"000000000",
  30474=>"111111111",
  30475=>"111111010",
  30476=>"000000000",
  30477=>"000000111",
  30478=>"001111111",
  30479=>"000111011",
  30480=>"000000000",
  30481=>"000000000",
  30482=>"100000110",
  30483=>"000111111",
  30484=>"000000000",
  30485=>"000000111",
  30486=>"111110110",
  30487=>"101111000",
  30488=>"111111000",
  30489=>"000000000",
  30490=>"110000111",
  30491=>"000000101",
  30492=>"001011111",
  30493=>"000000000",
  30494=>"000111111",
  30495=>"111100100",
  30496=>"000111000",
  30497=>"000110000",
  30498=>"111111000",
  30499=>"111111110",
  30500=>"111111111",
  30501=>"000110000",
  30502=>"000000000",
  30503=>"000111000",
  30504=>"001001011",
  30505=>"001111111",
  30506=>"000000001",
  30507=>"000000010",
  30508=>"111000000",
  30509=>"111011010",
  30510=>"111111111",
  30511=>"000000001",
  30512=>"111111100",
  30513=>"000000111",
  30514=>"000000000",
  30515=>"111111000",
  30516=>"000111000",
  30517=>"011111111",
  30518=>"000000111",
  30519=>"111011000",
  30520=>"111111000",
  30521=>"111100111",
  30522=>"010111111",
  30523=>"001000000",
  30524=>"000000011",
  30525=>"000000000",
  30526=>"000111011",
  30527=>"101111110",
  30528=>"001000000",
  30529=>"000000000",
  30530=>"000111110",
  30531=>"011110110",
  30532=>"000000111",
  30533=>"000111111",
  30534=>"111001000",
  30535=>"111111000",
  30536=>"001001000",
  30537=>"000000000",
  30538=>"001000000",
  30539=>"111100000",
  30540=>"110111111",
  30541=>"001001111",
  30542=>"111111000",
  30543=>"000011111",
  30544=>"111000100",
  30545=>"011000000",
  30546=>"111100011",
  30547=>"011000000",
  30548=>"000000010",
  30549=>"011111000",
  30550=>"000000000",
  30551=>"111111111",
  30552=>"111111000",
  30553=>"000111111",
  30554=>"111111000",
  30555=>"000000000",
  30556=>"100110111",
  30557=>"000000111",
  30558=>"101000001",
  30559=>"110110111",
  30560=>"000100000",
  30561=>"111111000",
  30562=>"111111100",
  30563=>"000110111",
  30564=>"011111111",
  30565=>"000000000",
  30566=>"001000000",
  30567=>"111111000",
  30568=>"010111100",
  30569=>"111101000",
  30570=>"110110110",
  30571=>"110110110",
  30572=>"011011110",
  30573=>"111000111",
  30574=>"000101111",
  30575=>"000011111",
  30576=>"111111001",
  30577=>"001111111",
  30578=>"111111111",
  30579=>"111111111",
  30580=>"111111000",
  30581=>"101111111",
  30582=>"000000000",
  30583=>"000000000",
  30584=>"000111111",
  30585=>"000000000",
  30586=>"111111111",
  30587=>"010000001",
  30588=>"011111011",
  30589=>"111111000",
  30590=>"000000111",
  30591=>"000111111",
  30592=>"000000000",
  30593=>"001000000",
  30594=>"000000110",
  30595=>"100000000",
  30596=>"011000111",
  30597=>"001111111",
  30598=>"111111111",
  30599=>"110111000",
  30600=>"000000111",
  30601=>"000000111",
  30602=>"000001111",
  30603=>"111111000",
  30604=>"101111111",
  30605=>"000000000",
  30606=>"101100000",
  30607=>"000000000",
  30608=>"011011000",
  30609=>"001000011",
  30610=>"100100000",
  30611=>"000000100",
  30612=>"111111111",
  30613=>"000000000",
  30614=>"000000000",
  30615=>"110111000",
  30616=>"111001000",
  30617=>"110111011",
  30618=>"001000111",
  30619=>"000111001",
  30620=>"111010000",
  30621=>"111111000",
  30622=>"000000011",
  30623=>"000000111",
  30624=>"111111101",
  30625=>"110110000",
  30626=>"000111111",
  30627=>"110111000",
  30628=>"001000101",
  30629=>"000001011",
  30630=>"111111111",
  30631=>"111111100",
  30632=>"011011111",
  30633=>"000000000",
  30634=>"111000000",
  30635=>"000000000",
  30636=>"000001111",
  30637=>"001000001",
  30638=>"001111011",
  30639=>"111111000",
  30640=>"111000000",
  30641=>"101000000",
  30642=>"110010111",
  30643=>"111000000",
  30644=>"000000111",
  30645=>"111000000",
  30646=>"100111111",
  30647=>"000000000",
  30648=>"000000000",
  30649=>"111111111",
  30650=>"111111111",
  30651=>"000001101",
  30652=>"111000101",
  30653=>"111000100",
  30654=>"001000101",
  30655=>"000100000",
  30656=>"111111000",
  30657=>"000100111",
  30658=>"001111111",
  30659=>"000000000",
  30660=>"101110001",
  30661=>"000000000",
  30662=>"001001001",
  30663=>"000101101",
  30664=>"000110000",
  30665=>"111011000",
  30666=>"000000000",
  30667=>"111111111",
  30668=>"000100000",
  30669=>"111001000",
  30670=>"000000000",
  30671=>"000000100",
  30672=>"000000011",
  30673=>"000111011",
  30674=>"111111001",
  30675=>"001011111",
  30676=>"111111100",
  30677=>"000000111",
  30678=>"000000000",
  30679=>"100110111",
  30680=>"000000000",
  30681=>"001000111",
  30682=>"000011111",
  30683=>"111110111",
  30684=>"011010000",
  30685=>"100100111",
  30686=>"110100001",
  30687=>"010000111",
  30688=>"111111111",
  30689=>"111111111",
  30690=>"111111111",
  30691=>"000000000",
  30692=>"111011000",
  30693=>"000111111",
  30694=>"111101001",
  30695=>"000111111",
  30696=>"111111111",
  30697=>"111111111",
  30698=>"111010000",
  30699=>"000000000",
  30700=>"000000110",
  30701=>"111111000",
  30702=>"000000011",
  30703=>"111111111",
  30704=>"110011111",
  30705=>"000111111",
  30706=>"111111000",
  30707=>"110010000",
  30708=>"111000011",
  30709=>"110010111",
  30710=>"111111000",
  30711=>"111001000",
  30712=>"000000111",
  30713=>"010000001",
  30714=>"111111100",
  30715=>"111111110",
  30716=>"000000100",
  30717=>"011001000",
  30718=>"111011010",
  30719=>"100000000",
  30720=>"110000000",
  30721=>"111000000",
  30722=>"000000001",
  30723=>"111111000",
  30724=>"000000000",
  30725=>"000000111",
  30726=>"001000001",
  30727=>"000000000",
  30728=>"000000100",
  30729=>"000000000",
  30730=>"000111111",
  30731=>"111110100",
  30732=>"001100001",
  30733=>"111011000",
  30734=>"011100100",
  30735=>"101000001",
  30736=>"000000010",
  30737=>"000000111",
  30738=>"011001011",
  30739=>"111111111",
  30740=>"011000000",
  30741=>"111111111",
  30742=>"110111111",
  30743=>"100111000",
  30744=>"100111110",
  30745=>"111001000",
  30746=>"001000000",
  30747=>"111111100",
  30748=>"101000000",
  30749=>"000001000",
  30750=>"011000000",
  30751=>"001111000",
  30752=>"100010111",
  30753=>"000101111",
  30754=>"000111111",
  30755=>"000000000",
  30756=>"000010000",
  30757=>"000001101",
  30758=>"000000000",
  30759=>"111111101",
  30760=>"110110110",
  30761=>"000111111",
  30762=>"100111111",
  30763=>"000000000",
  30764=>"001111110",
  30765=>"000011111",
  30766=>"111011000",
  30767=>"111000000",
  30768=>"000111111",
  30769=>"110100000",
  30770=>"000111111",
  30771=>"111111011",
  30772=>"000000100",
  30773=>"001001001",
  30774=>"101111111",
  30775=>"111000000",
  30776=>"011111011",
  30777=>"111111111",
  30778=>"111111001",
  30779=>"110111111",
  30780=>"000000111",
  30781=>"100000000",
  30782=>"100100111",
  30783=>"111111111",
  30784=>"100000000",
  30785=>"000000100",
  30786=>"111110110",
  30787=>"000001100",
  30788=>"000110000",
  30789=>"111000000",
  30790=>"011000111",
  30791=>"000000000",
  30792=>"000111000",
  30793=>"011000000",
  30794=>"011111111",
  30795=>"100100111",
  30796=>"111000000",
  30797=>"111111000",
  30798=>"100100111",
  30799=>"000000111",
  30800=>"001000000",
  30801=>"000000111",
  30802=>"111000000",
  30803=>"000001011",
  30804=>"000000000",
  30805=>"111111100",
  30806=>"000000101",
  30807=>"000011001",
  30808=>"001110000",
  30809=>"001000000",
  30810=>"000000000",
  30811=>"000110111",
  30812=>"000000100",
  30813=>"111111111",
  30814=>"000000011",
  30815=>"011111000",
  30816=>"000000100",
  30817=>"111111111",
  30818=>"100100100",
  30819=>"000000000",
  30820=>"111111111",
  30821=>"000000101",
  30822=>"000000000",
  30823=>"000111111",
  30824=>"111100111",
  30825=>"001000001",
  30826=>"111001111",
  30827=>"111111111",
  30828=>"000111110",
  30829=>"100100111",
  30830=>"110110000",
  30831=>"010011110",
  30832=>"011011111",
  30833=>"000000000",
  30834=>"111000111",
  30835=>"000000000",
  30836=>"000000000",
  30837=>"111101111",
  30838=>"000100110",
  30839=>"000000011",
  30840=>"111111100",
  30841=>"111000000",
  30842=>"111110110",
  30843=>"010000000",
  30844=>"000110000",
  30845=>"000000000",
  30846=>"100110111",
  30847=>"111111001",
  30848=>"111111111",
  30849=>"111111011",
  30850=>"111111111",
  30851=>"010000000",
  30852=>"100110100",
  30853=>"100101111",
  30854=>"111111111",
  30855=>"000010000",
  30856=>"111111001",
  30857=>"000000000",
  30858=>"001000000",
  30859=>"000000000",
  30860=>"001000000",
  30861=>"000000111",
  30862=>"111111111",
  30863=>"000000000",
  30864=>"110000000",
  30865=>"000000001",
  30866=>"000000000",
  30867=>"000111111",
  30868=>"000001000",
  30869=>"000100111",
  30870=>"001001111",
  30871=>"000001001",
  30872=>"000000000",
  30873=>"111111101",
  30874=>"111111111",
  30875=>"111100000",
  30876=>"001000111",
  30877=>"111000000",
  30878=>"000111111",
  30879=>"011001111",
  30880=>"000000100",
  30881=>"011111111",
  30882=>"111111111",
  30883=>"100110110",
  30884=>"010000110",
  30885=>"111101111",
  30886=>"111111000",
  30887=>"011010011",
  30888=>"111000111",
  30889=>"111111011",
  30890=>"000000000",
  30891=>"000001000",
  30892=>"010000011",
  30893=>"000001111",
  30894=>"000000100",
  30895=>"111011000",
  30896=>"111111000",
  30897=>"010011001",
  30898=>"111111111",
  30899=>"111111111",
  30900=>"111010000",
  30901=>"011111111",
  30902=>"000111111",
  30903=>"111110111",
  30904=>"000000110",
  30905=>"011111111",
  30906=>"011011000",
  30907=>"101111011",
  30908=>"000110111",
  30909=>"111111001",
  30910=>"111110011",
  30911=>"101000000",
  30912=>"000100000",
  30913=>"111111111",
  30914=>"101000000",
  30915=>"111111000",
  30916=>"111111111",
  30917=>"000000001",
  30918=>"111000110",
  30919=>"111111111",
  30920=>"001111011",
  30921=>"111111110",
  30922=>"000100000",
  30923=>"101000111",
  30924=>"110000000",
  30925=>"000101001",
  30926=>"001000000",
  30927=>"001000000",
  30928=>"001001111",
  30929=>"111111111",
  30930=>"111000000",
  30931=>"001000000",
  30932=>"010110110",
  30933=>"110111110",
  30934=>"000000000",
  30935=>"010011000",
  30936=>"011011111",
  30937=>"100100111",
  30938=>"000000000",
  30939=>"000000000",
  30940=>"111011000",
  30941=>"000011000",
  30942=>"101111111",
  30943=>"001000000",
  30944=>"111000000",
  30945=>"000111111",
  30946=>"111011000",
  30947=>"000001101",
  30948=>"000111111",
  30949=>"000000110",
  30950=>"111000000",
  30951=>"000100101",
  30952=>"100111100",
  30953=>"111000000",
  30954=>"001000000",
  30955=>"100111000",
  30956=>"010010000",
  30957=>"111000000",
  30958=>"000000111",
  30959=>"000000111",
  30960=>"000000000",
  30961=>"000011111",
  30962=>"111110100",
  30963=>"000001001",
  30964=>"111000001",
  30965=>"000110110",
  30966=>"001000000",
  30967=>"000111001",
  30968=>"111111111",
  30969=>"111010000",
  30970=>"011111111",
  30971=>"100100000",
  30972=>"000000000",
  30973=>"000111110",
  30974=>"111111001",
  30975=>"111011011",
  30976=>"100000000",
  30977=>"000000000",
  30978=>"010000111",
  30979=>"111111111",
  30980=>"111000000",
  30981=>"000000111",
  30982=>"000111111",
  30983=>"111111101",
  30984=>"111110111",
  30985=>"111000000",
  30986=>"010111111",
  30987=>"100101001",
  30988=>"000000000",
  30989=>"000000111",
  30990=>"011111111",
  30991=>"000000000",
  30992=>"010111011",
  30993=>"111110000",
  30994=>"011000000",
  30995=>"000111111",
  30996=>"000000000",
  30997=>"000000000",
  30998=>"111111111",
  30999=>"110110000",
  31000=>"111111110",
  31001=>"001000011",
  31002=>"000000000",
  31003=>"001011111",
  31004=>"011111111",
  31005=>"011000000",
  31006=>"111001001",
  31007=>"111100100",
  31008=>"000111010",
  31009=>"111110000",
  31010=>"011111000",
  31011=>"000111111",
  31012=>"000000110",
  31013=>"110000111",
  31014=>"000000000",
  31015=>"111111000",
  31016=>"000110110",
  31017=>"000010111",
  31018=>"101000000",
  31019=>"000000000",
  31020=>"100010001",
  31021=>"000011000",
  31022=>"001111111",
  31023=>"100000000",
  31024=>"000000100",
  31025=>"000000000",
  31026=>"011010110",
  31027=>"000000000",
  31028=>"111100000",
  31029=>"000000000",
  31030=>"000000000",
  31031=>"101100111",
  31032=>"000000000",
  31033=>"001000000",
  31034=>"000000000",
  31035=>"110000000",
  31036=>"011001000",
  31037=>"001111100",
  31038=>"000100000",
  31039=>"111111000",
  31040=>"000000011",
  31041=>"111000000",
  31042=>"000000100",
  31043=>"001111111",
  31044=>"000000100",
  31045=>"000000000",
  31046=>"111011010",
  31047=>"001000111",
  31048=>"000010010",
  31049=>"111000000",
  31050=>"011000000",
  31051=>"111000100",
  31052=>"110111111",
  31053=>"001000000",
  31054=>"000111111",
  31055=>"100110000",
  31056=>"011111111",
  31057=>"101100000",
  31058=>"010111110",
  31059=>"000000100",
  31060=>"000000000",
  31061=>"000001001",
  31062=>"000000011",
  31063=>"111000000",
  31064=>"111011000",
  31065=>"111000111",
  31066=>"011000000",
  31067=>"110000000",
  31068=>"110111101",
  31069=>"010010000",
  31070=>"111000111",
  31071=>"001000000",
  31072=>"111000101",
  31073=>"001000000",
  31074=>"101101111",
  31075=>"111000111",
  31076=>"001111111",
  31077=>"000000000",
  31078=>"000000000",
  31079=>"000000000",
  31080=>"000000000",
  31081=>"101000000",
  31082=>"000000000",
  31083=>"100111000",
  31084=>"000111110",
  31085=>"110000000",
  31086=>"111111111",
  31087=>"000000000",
  31088=>"000000101",
  31089=>"000101000",
  31090=>"111001001",
  31091=>"100100100",
  31092=>"000110000",
  31093=>"100000000",
  31094=>"111111111",
  31095=>"100000000",
  31096=>"111000000",
  31097=>"111111111",
  31098=>"000000110",
  31099=>"110111000",
  31100=>"011011010",
  31101=>"000111111",
  31102=>"000000000",
  31103=>"101000000",
  31104=>"000100001",
  31105=>"111111111",
  31106=>"111100100",
  31107=>"000000000",
  31108=>"111011011",
  31109=>"000111011",
  31110=>"110000001",
  31111=>"000000000",
  31112=>"000001111",
  31113=>"111111111",
  31114=>"000000000",
  31115=>"100001000",
  31116=>"111001000",
  31117=>"111000000",
  31118=>"000111111",
  31119=>"000111111",
  31120=>"000000011",
  31121=>"111111111",
  31122=>"011000001",
  31123=>"100000000",
  31124=>"000111111",
  31125=>"000011000",
  31126=>"000000000",
  31127=>"000000000",
  31128=>"111000000",
  31129=>"000000010",
  31130=>"111011000",
  31131=>"100110011",
  31132=>"110111000",
  31133=>"101111111",
  31134=>"110110000",
  31135=>"000000000",
  31136=>"111111111",
  31137=>"111111111",
  31138=>"111110101",
  31139=>"001000000",
  31140=>"011000001",
  31141=>"111111111",
  31142=>"111000000",
  31143=>"000110111",
  31144=>"110110100",
  31145=>"000100111",
  31146=>"100110110",
  31147=>"000000000",
  31148=>"000000000",
  31149=>"111001000",
  31150=>"111010000",
  31151=>"000111100",
  31152=>"111000000",
  31153=>"000000001",
  31154=>"111111111",
  31155=>"000110110",
  31156=>"010111111",
  31157=>"000000000",
  31158=>"110000000",
  31159=>"111011110",
  31160=>"000000110",
  31161=>"100111110",
  31162=>"000000000",
  31163=>"111111011",
  31164=>"101000010",
  31165=>"111111111",
  31166=>"000000101",
  31167=>"000011111",
  31168=>"000111110",
  31169=>"111111111",
  31170=>"000000000",
  31171=>"011000000",
  31172=>"000011111",
  31173=>"111000000",
  31174=>"110000001",
  31175=>"110100000",
  31176=>"110010000",
  31177=>"000000000",
  31178=>"000000001",
  31179=>"111111000",
  31180=>"000000000",
  31181=>"000000000",
  31182=>"000010111",
  31183=>"000010111",
  31184=>"111000000",
  31185=>"000110111",
  31186=>"000000000",
  31187=>"000000000",
  31188=>"000000000",
  31189=>"001010011",
  31190=>"010000111",
  31191=>"110110000",
  31192=>"111111111",
  31193=>"000111011",
  31194=>"000000000",
  31195=>"000000000",
  31196=>"111110111",
  31197=>"101001101",
  31198=>"111000000",
  31199=>"000100100",
  31200=>"000000000",
  31201=>"011011111",
  31202=>"000000010",
  31203=>"111111011",
  31204=>"010111111",
  31205=>"100101000",
  31206=>"111111000",
  31207=>"011000000",
  31208=>"000111011",
  31209=>"111111011",
  31210=>"110110000",
  31211=>"000111110",
  31212=>"000000100",
  31213=>"000000000",
  31214=>"000110111",
  31215=>"101001111",
  31216=>"000100000",
  31217=>"100110111",
  31218=>"000111111",
  31219=>"111001111",
  31220=>"111111111",
  31221=>"011011111",
  31222=>"010111111",
  31223=>"000001011",
  31224=>"000000000",
  31225=>"000000000",
  31226=>"000000110",
  31227=>"010000000",
  31228=>"000111101",
  31229=>"101111111",
  31230=>"010000000",
  31231=>"111000110",
  31232=>"010000011",
  31233=>"111000000",
  31234=>"111001111",
  31235=>"101111111",
  31236=>"001001111",
  31237=>"000110110",
  31238=>"111111111",
  31239=>"111111111",
  31240=>"100000000",
  31241=>"111111000",
  31242=>"000001111",
  31243=>"000011000",
  31244=>"111111111",
  31245=>"111101111",
  31246=>"011011001",
  31247=>"111101101",
  31248=>"111111001",
  31249=>"011110100",
  31250=>"000000000",
  31251=>"111111111",
  31252=>"000000000",
  31253=>"001111111",
  31254=>"111111001",
  31255=>"011011000",
  31256=>"001000101",
  31257=>"100111111",
  31258=>"111011001",
  31259=>"000000110",
  31260=>"011111111",
  31261=>"000000000",
  31262=>"110000111",
  31263=>"100100100",
  31264=>"111001000",
  31265=>"111111110",
  31266=>"000000100",
  31267=>"001010111",
  31268=>"111111111",
  31269=>"000000000",
  31270=>"000000000",
  31271=>"010000000",
  31272=>"011011111",
  31273=>"000000000",
  31274=>"011011011",
  31275=>"011111111",
  31276=>"111111111",
  31277=>"110111111",
  31278=>"000000011",
  31279=>"000000100",
  31280=>"111001000",
  31281=>"111111000",
  31282=>"110100100",
  31283=>"100000000",
  31284=>"111000000",
  31285=>"011001111",
  31286=>"000000101",
  31287=>"010000000",
  31288=>"100000001",
  31289=>"111011011",
  31290=>"000000000",
  31291=>"101101011",
  31292=>"110110100",
  31293=>"111101111",
  31294=>"110111100",
  31295=>"111111111",
  31296=>"100000000",
  31297=>"111111001",
  31298=>"111111111",
  31299=>"111001001",
  31300=>"000000000",
  31301=>"011111011",
  31302=>"001001000",
  31303=>"000000000",
  31304=>"111111111",
  31305=>"111010111",
  31306=>"000000000",
  31307=>"000000000",
  31308=>"111111111",
  31309=>"110110000",
  31310=>"111111111",
  31311=>"000000001",
  31312=>"000000000",
  31313=>"001001001",
  31314=>"011000000",
  31315=>"010110000",
  31316=>"111101000",
  31317=>"000000000",
  31318=>"101100001",
  31319=>"000000000",
  31320=>"111111111",
  31321=>"000000111",
  31322=>"000000011",
  31323=>"111110111",
  31324=>"011111101",
  31325=>"111111111",
  31326=>"100000001",
  31327=>"000000000",
  31328=>"110000010",
  31329=>"111011011",
  31330=>"011111111",
  31331=>"111111111",
  31332=>"110100000",
  31333=>"011000101",
  31334=>"100100111",
  31335=>"011111111",
  31336=>"111011000",
  31337=>"111111111",
  31338=>"111111111",
  31339=>"000000000",
  31340=>"111111111",
  31341=>"000000011",
  31342=>"101101111",
  31343=>"111111111",
  31344=>"111000001",
  31345=>"010000000",
  31346=>"110000011",
  31347=>"001011001",
  31348=>"000000000",
  31349=>"111111111",
  31350=>"111111111",
  31351=>"000000000",
  31352=>"000000011",
  31353=>"011011011",
  31354=>"011000000",
  31355=>"001001001",
  31356=>"110100000",
  31357=>"111111101",
  31358=>"001011001",
  31359=>"111000000",
  31360=>"111000000",
  31361=>"111011000",
  31362=>"111111100",
  31363=>"110111011",
  31364=>"111111011",
  31365=>"000000000",
  31366=>"000000011",
  31367=>"111111111",
  31368=>"111111111",
  31369=>"000111111",
  31370=>"000001001",
  31371=>"000001011",
  31372=>"111000110",
  31373=>"100111111",
  31374=>"111101011",
  31375=>"111111111",
  31376=>"101000100",
  31377=>"111111111",
  31378=>"010000000",
  31379=>"111110100",
  31380=>"000000000",
  31381=>"111111111",
  31382=>"111111111",
  31383=>"000000000",
  31384=>"101001101",
  31385=>"111111111",
  31386=>"101111111",
  31387=>"001001000",
  31388=>"000000000",
  31389=>"011001000",
  31390=>"100000010",
  31391=>"110111111",
  31392=>"100000000",
  31393=>"011011111",
  31394=>"111111111",
  31395=>"111111111",
  31396=>"111111111",
  31397=>"100101111",
  31398=>"111111000",
  31399=>"000000011",
  31400=>"000000000",
  31401=>"111000000",
  31402=>"000000111",
  31403=>"010010001",
  31404=>"111111111",
  31405=>"011000000",
  31406=>"000000000",
  31407=>"000000000",
  31408=>"111111111",
  31409=>"111111101",
  31410=>"011111011",
  31411=>"111111111",
  31412=>"111111111",
  31413=>"000000000",
  31414=>"111111111",
  31415=>"000000111",
  31416=>"001011011",
  31417=>"000010010",
  31418=>"000000000",
  31419=>"111111101",
  31420=>"000000010",
  31421=>"100100000",
  31422=>"000100111",
  31423=>"000000000",
  31424=>"100100100",
  31425=>"001000000",
  31426=>"111111111",
  31427=>"000110000",
  31428=>"111111111",
  31429=>"010010011",
  31430=>"000000111",
  31431=>"000010011",
  31432=>"000001001",
  31433=>"000000100",
  31434=>"010000000",
  31435=>"000000100",
  31436=>"100111000",
  31437=>"001001010",
  31438=>"111111110",
  31439=>"101100111",
  31440=>"111001111",
  31441=>"001001000",
  31442=>"111100100",
  31443=>"011000000",
  31444=>"100100101",
  31445=>"110100000",
  31446=>"110011000",
  31447=>"000000001",
  31448=>"110111111",
  31449=>"101101101",
  31450=>"000000000",
  31451=>"000000000",
  31452=>"000000100",
  31453=>"111101101",
  31454=>"000000000",
  31455=>"111111111",
  31456=>"000000000",
  31457=>"000000000",
  31458=>"001001111",
  31459=>"000000001",
  31460=>"101101100",
  31461=>"101111111",
  31462=>"111111110",
  31463=>"100111111",
  31464=>"111111111",
  31465=>"111111110",
  31466=>"000000000",
  31467=>"011101111",
  31468=>"111101001",
  31469=>"000100000",
  31470=>"000100110",
  31471=>"011111001",
  31472=>"001011000",
  31473=>"011000011",
  31474=>"111100100",
  31475=>"000000000",
  31476=>"000000000",
  31477=>"111100000",
  31478=>"101111111",
  31479=>"000000011",
  31480=>"000011111",
  31481=>"011111000",
  31482=>"110111100",
  31483=>"111111111",
  31484=>"110110111",
  31485=>"111000011",
  31486=>"001101101",
  31487=>"101111111",
  31488=>"000000000",
  31489=>"111000001",
  31490=>"011001001",
  31491=>"000000011",
  31492=>"111111111",
  31493=>"001000111",
  31494=>"000000000",
  31495=>"100000111",
  31496=>"000110010",
  31497=>"001000011",
  31498=>"001000101",
  31499=>"111111100",
  31500=>"000000000",
  31501=>"000000000",
  31502=>"000000001",
  31503=>"001001001",
  31504=>"110000001",
  31505=>"001001101",
  31506=>"000000111",
  31507=>"000111111",
  31508=>"000000000",
  31509=>"011000000",
  31510=>"111111110",
  31511=>"110100000",
  31512=>"011001000",
  31513=>"111111111",
  31514=>"111111111",
  31515=>"111111111",
  31516=>"011011001",
  31517=>"000000010",
  31518=>"111100111",
  31519=>"010110111",
  31520=>"001001000",
  31521=>"111111000",
  31522=>"000000000",
  31523=>"000000000",
  31524=>"000000100",
  31525=>"000000000",
  31526=>"110110111",
  31527=>"000000000",
  31528=>"000000111",
  31529=>"000000000",
  31530=>"111111110",
  31531=>"000001000",
  31532=>"110010000",
  31533=>"010110110",
  31534=>"111001000",
  31535=>"000000000",
  31536=>"111111110",
  31537=>"111111111",
  31538=>"010111110",
  31539=>"000000000",
  31540=>"011001000",
  31541=>"111011001",
  31542=>"000000001",
  31543=>"101100100",
  31544=>"111111111",
  31545=>"001000011",
  31546=>"111101100",
  31547=>"101000001",
  31548=>"100000011",
  31549=>"110111001",
  31550=>"111111111",
  31551=>"000000100",
  31552=>"100110000",
  31553=>"000000000",
  31554=>"111111111",
  31555=>"000011111",
  31556=>"011001000",
  31557=>"000000011",
  31558=>"111000000",
  31559=>"001000100",
  31560=>"111001000",
  31561=>"111000000",
  31562=>"010000011",
  31563=>"001011111",
  31564=>"011000001",
  31565=>"000000000",
  31566=>"000000000",
  31567=>"111111110",
  31568=>"111111111",
  31569=>"000000000",
  31570=>"000000000",
  31571=>"000000000",
  31572=>"001000000",
  31573=>"011011011",
  31574=>"111111111",
  31575=>"100101101",
  31576=>"111111100",
  31577=>"111111000",
  31578=>"001000000",
  31579=>"000000111",
  31580=>"011001000",
  31581=>"111111111",
  31582=>"011111111",
  31583=>"000000001",
  31584=>"111011011",
  31585=>"000000000",
  31586=>"111000000",
  31587=>"000000001",
  31588=>"000011111",
  31589=>"111111011",
  31590=>"000000111",
  31591=>"000000000",
  31592=>"110110110",
  31593=>"111000000",
  31594=>"111110010",
  31595=>"111111101",
  31596=>"111111100",
  31597=>"000000000",
  31598=>"000000000",
  31599=>"111001111",
  31600=>"111111111",
  31601=>"000000000",
  31602=>"011011000",
  31603=>"000000000",
  31604=>"111111111",
  31605=>"111111111",
  31606=>"111101001",
  31607=>"001111000",
  31608=>"111111110",
  31609=>"001000111",
  31610=>"000000100",
  31611=>"111001111",
  31612=>"111000000",
  31613=>"111111111",
  31614=>"111001001",
  31615=>"000100100",
  31616=>"111011111",
  31617=>"011000000",
  31618=>"100110110",
  31619=>"000000000",
  31620=>"011001110",
  31621=>"111111111",
  31622=>"111111111",
  31623=>"110000011",
  31624=>"000000000",
  31625=>"111111111",
  31626=>"001000000",
  31627=>"111111011",
  31628=>"000011111",
  31629=>"100100101",
  31630=>"000000000",
  31631=>"000000000",
  31632=>"011000000",
  31633=>"000100101",
  31634=>"111111111",
  31635=>"010110111",
  31636=>"000001111",
  31637=>"110110000",
  31638=>"100110110",
  31639=>"011111110",
  31640=>"111001001",
  31641=>"100000000",
  31642=>"111111111",
  31643=>"111111011",
  31644=>"000000000",
  31645=>"111111111",
  31646=>"100000000",
  31647=>"110111000",
  31648=>"110110100",
  31649=>"111000000",
  31650=>"111100000",
  31651=>"000001011",
  31652=>"011011001",
  31653=>"000000000",
  31654=>"000000000",
  31655=>"000000110",
  31656=>"000000000",
  31657=>"010000000",
  31658=>"000000000",
  31659=>"011000000",
  31660=>"001000000",
  31661=>"000001111",
  31662=>"000100000",
  31663=>"101101111",
  31664=>"001111111",
  31665=>"000000000",
  31666=>"111111111",
  31667=>"100111111",
  31668=>"000000001",
  31669=>"110110110",
  31670=>"111000000",
  31671=>"111111111",
  31672=>"111111111",
  31673=>"101101000",
  31674=>"110100011",
  31675=>"011001000",
  31676=>"100000011",
  31677=>"111111000",
  31678=>"011010010",
  31679=>"001001001",
  31680=>"000000000",
  31681=>"111111000",
  31682=>"010000000",
  31683=>"111111111",
  31684=>"001011111",
  31685=>"111010100",
  31686=>"111111011",
  31687=>"111101101",
  31688=>"111101111",
  31689=>"100110100",
  31690=>"111000000",
  31691=>"011001111",
  31692=>"111011000",
  31693=>"110100111",
  31694=>"000000000",
  31695=>"100000000",
  31696=>"111000000",
  31697=>"000000000",
  31698=>"000000000",
  31699=>"111111111",
  31700=>"000111111",
  31701=>"100100110",
  31702=>"111110000",
  31703=>"110110010",
  31704=>"000001111",
  31705=>"000000000",
  31706=>"111001010",
  31707=>"000000111",
  31708=>"111111111",
  31709=>"111011011",
  31710=>"111111000",
  31711=>"111101111",
  31712=>"111011000",
  31713=>"111111111",
  31714=>"010011000",
  31715=>"111111111",
  31716=>"000000000",
  31717=>"001011011",
  31718=>"000000000",
  31719=>"000011111",
  31720=>"001011011",
  31721=>"100100101",
  31722=>"111000000",
  31723=>"111111111",
  31724=>"000000000",
  31725=>"000110010",
  31726=>"000000111",
  31727=>"000000011",
  31728=>"000100000",
  31729=>"000000000",
  31730=>"110111111",
  31731=>"011011111",
  31732=>"000111111",
  31733=>"111111111",
  31734=>"000101000",
  31735=>"000100000",
  31736=>"111000000",
  31737=>"000000000",
  31738=>"001000000",
  31739=>"000100110",
  31740=>"000000001",
  31741=>"001000000",
  31742=>"000000100",
  31743=>"100110110",
  31744=>"101111111",
  31745=>"101111111",
  31746=>"111101001",
  31747=>"111111110",
  31748=>"111101111",
  31749=>"000000011",
  31750=>"000000000",
  31751=>"111111111",
  31752=>"000000000",
  31753=>"111111101",
  31754=>"000000000",
  31755=>"100110110",
  31756=>"000000000",
  31757=>"000110111",
  31758=>"000000001",
  31759=>"000000000",
  31760=>"011000110",
  31761=>"000000100",
  31762=>"111110000",
  31763=>"000000000",
  31764=>"000000101",
  31765=>"000001000",
  31766=>"011000100",
  31767=>"100001000",
  31768=>"001000000",
  31769=>"100001011",
  31770=>"000000111",
  31771=>"001011001",
  31772=>"111111111",
  31773=>"000111111",
  31774=>"000001001",
  31775=>"011111110",
  31776=>"111111111",
  31777=>"000000100",
  31778=>"011110110",
  31779=>"001011011",
  31780=>"111111111",
  31781=>"000000001",
  31782=>"111111111",
  31783=>"000000111",
  31784=>"001000000",
  31785=>"000000000",
  31786=>"111111111",
  31787=>"000000000",
  31788=>"000000111",
  31789=>"111111111",
  31790=>"111000000",
  31791=>"000000000",
  31792=>"011111110",
  31793=>"000000000",
  31794=>"000000100",
  31795=>"100110010",
  31796=>"111001001",
  31797=>"101111111",
  31798=>"000001000",
  31799=>"010011001",
  31800=>"110110111",
  31801=>"000000111",
  31802=>"000000000",
  31803=>"001001000",
  31804=>"000000111",
  31805=>"001110100",
  31806=>"111111111",
  31807=>"000000000",
  31808=>"000000000",
  31809=>"111111000",
  31810=>"000000111",
  31811=>"111111111",
  31812=>"000000000",
  31813=>"111111111",
  31814=>"000000111",
  31815=>"111111100",
  31816=>"000000000",
  31817=>"111101111",
  31818=>"110100000",
  31819=>"111111111",
  31820=>"111011001",
  31821=>"110110000",
  31822=>"100111111",
  31823=>"111000001",
  31824=>"011011000",
  31825=>"000000000",
  31826=>"000000110",
  31827=>"001001111",
  31828=>"000000000",
  31829=>"000010110",
  31830=>"000000000",
  31831=>"110111110",
  31832=>"001000000",
  31833=>"111101101",
  31834=>"010000000",
  31835=>"110110110",
  31836=>"000110111",
  31837=>"110111110",
  31838=>"110000000",
  31839=>"000111111",
  31840=>"000000000",
  31841=>"001001111",
  31842=>"001000000",
  31843=>"000000000",
  31844=>"001001000",
  31845=>"000000000",
  31846=>"000011000",
  31847=>"000000000",
  31848=>"111111111",
  31849=>"111000000",
  31850=>"111000000",
  31851=>"000000010",
  31852=>"111111000",
  31853=>"111101111",
  31854=>"101000001",
  31855=>"010110110",
  31856=>"110110111",
  31857=>"000000000",
  31858=>"011001001",
  31859=>"001011111",
  31860=>"000000000",
  31861=>"111111111",
  31862=>"111011011",
  31863=>"000000000",
  31864=>"111111111",
  31865=>"000000111",
  31866=>"111001011",
  31867=>"100000001",
  31868=>"110111111",
  31869=>"000000000",
  31870=>"000000000",
  31871=>"000011011",
  31872=>"100100110",
  31873=>"111000000",
  31874=>"000000000",
  31875=>"111110011",
  31876=>"010111111",
  31877=>"000001001",
  31878=>"111110000",
  31879=>"001001110",
  31880=>"111111000",
  31881=>"111101101",
  31882=>"111111111",
  31883=>"111111111",
  31884=>"111000000",
  31885=>"000000000",
  31886=>"110000000",
  31887=>"000000000",
  31888=>"001001111",
  31889=>"000000101",
  31890=>"000000001",
  31891=>"000110110",
  31892=>"000000000",
  31893=>"000000001",
  31894=>"000100110",
  31895=>"111000111",
  31896=>"111111111",
  31897=>"111111111",
  31898=>"011011111",
  31899=>"010011111",
  31900=>"111111101",
  31901=>"110110110",
  31902=>"000001011",
  31903=>"000000111",
  31904=>"011000001",
  31905=>"000000001",
  31906=>"000111110",
  31907=>"000000000",
  31908=>"111000000",
  31909=>"110000110",
  31910=>"101101111",
  31911=>"011001101",
  31912=>"111000000",
  31913=>"000000111",
  31914=>"000000100",
  31915=>"000000000",
  31916=>"000000010",
  31917=>"010110010",
  31918=>"001100000",
  31919=>"000000000",
  31920=>"111010010",
  31921=>"100000110",
  31922=>"111111111",
  31923=>"000101111",
  31924=>"111111111",
  31925=>"111111110",
  31926=>"000110010",
  31927=>"111111000",
  31928=>"111111111",
  31929=>"111111101",
  31930=>"111001000",
  31931=>"111111100",
  31932=>"000110100",
  31933=>"100000111",
  31934=>"111111111",
  31935=>"000100111",
  31936=>"111111111",
  31937=>"000000000",
  31938=>"000000101",
  31939=>"110111110",
  31940=>"100111110",
  31941=>"110111000",
  31942=>"000001001",
  31943=>"111111000",
  31944=>"110111111",
  31945=>"110000111",
  31946=>"111111011",
  31947=>"000000101",
  31948=>"100011011",
  31949=>"000111111",
  31950=>"011111110",
  31951=>"101001001",
  31952=>"100000000",
  31953=>"111111110",
  31954=>"100111000",
  31955=>"000000000",
  31956=>"010010010",
  31957=>"111110111",
  31958=>"000000111",
  31959=>"111011111",
  31960=>"011111100",
  31961=>"000000001",
  31962=>"111001001",
  31963=>"000000110",
  31964=>"000001001",
  31965=>"000111111",
  31966=>"110100000",
  31967=>"011011000",
  31968=>"101000001",
  31969=>"011010111",
  31970=>"011111010",
  31971=>"111111111",
  31972=>"111111111",
  31973=>"111111001",
  31974=>"000100110",
  31975=>"111111111",
  31976=>"111000000",
  31977=>"111011011",
  31978=>"100100101",
  31979=>"001011101",
  31980=>"111111111",
  31981=>"000000000",
  31982=>"110010111",
  31983=>"111111111",
  31984=>"000000001",
  31985=>"110110111",
  31986=>"111101001",
  31987=>"011000001",
  31988=>"000000000",
  31989=>"000111111",
  31990=>"011011000",
  31991=>"000000110",
  31992=>"000000000",
  31993=>"000000000",
  31994=>"111010010",
  31995=>"001110100",
  31996=>"100111001",
  31997=>"101111111",
  31998=>"000000001",
  31999=>"110001110",
  32000=>"111100000",
  32001=>"001000000",
  32002=>"000110111",
  32003=>"001000111",
  32004=>"011100000",
  32005=>"000111110",
  32006=>"111101111",
  32007=>"111111000",
  32008=>"000000000",
  32009=>"000000111",
  32010=>"111111111",
  32011=>"100100101",
  32012=>"111101101",
  32013=>"110010011",
  32014=>"000100000",
  32015=>"110111000",
  32016=>"110000001",
  32017=>"110111111",
  32018=>"111111111",
  32019=>"110111110",
  32020=>"000000111",
  32021=>"010111111",
  32022=>"001000100",
  32023=>"110111110",
  32024=>"001011011",
  32025=>"111111111",
  32026=>"000000000",
  32027=>"111111100",
  32028=>"100101001",
  32029=>"111111111",
  32030=>"110110110",
  32031=>"000000000",
  32032=>"000000000",
  32033=>"100000000",
  32034=>"111000000",
  32035=>"111111111",
  32036=>"001000000",
  32037=>"111111111",
  32038=>"000000100",
  32039=>"110110100",
  32040=>"000101111",
  32041=>"000000000",
  32042=>"000000010",
  32043=>"111111000",
  32044=>"001001111",
  32045=>"000000001",
  32046=>"111111011",
  32047=>"110100110",
  32048=>"000000100",
  32049=>"000000110",
  32050=>"001001101",
  32051=>"011001011",
  32052=>"001100000",
  32053=>"101000110",
  32054=>"010000000",
  32055=>"001111111",
  32056=>"000100000",
  32057=>"100101101",
  32058=>"000000000",
  32059=>"000000000",
  32060=>"000000010",
  32061=>"111111111",
  32062=>"000000000",
  32063=>"000000011",
  32064=>"000000100",
  32065=>"000000001",
  32066=>"111111111",
  32067=>"000000001",
  32068=>"111010000",
  32069=>"000001011",
  32070=>"000001111",
  32071=>"001000110",
  32072=>"001000001",
  32073=>"010010000",
  32074=>"000110111",
  32075=>"000000001",
  32076=>"111111111",
  32077=>"111111111",
  32078=>"001000001",
  32079=>"110110110",
  32080=>"001101111",
  32081=>"000000111",
  32082=>"111111000",
  32083=>"000110110",
  32084=>"000000111",
  32085=>"011011001",
  32086=>"111111111",
  32087=>"000111111",
  32088=>"111111111",
  32089=>"011111011",
  32090=>"001000110",
  32091=>"111110110",
  32092=>"111111111",
  32093=>"000000000",
  32094=>"100000001",
  32095=>"111011111",
  32096=>"000000100",
  32097=>"111111111",
  32098=>"000000101",
  32099=>"000000010",
  32100=>"000000000",
  32101=>"000000101",
  32102=>"111000000",
  32103=>"000110111",
  32104=>"011111100",
  32105=>"000011000",
  32106=>"110111111",
  32107=>"000000100",
  32108=>"000000000",
  32109=>"011000011",
  32110=>"000110110",
  32111=>"000000110",
  32112=>"001000000",
  32113=>"110110111",
  32114=>"000000001",
  32115=>"111111111",
  32116=>"000000000",
  32117=>"001001001",
  32118=>"000000001",
  32119=>"110000011",
  32120=>"111000000",
  32121=>"010111111",
  32122=>"000001001",
  32123=>"000000000",
  32124=>"000000000",
  32125=>"001010000",
  32126=>"110010000",
  32127=>"000101111",
  32128=>"110111110",
  32129=>"010111000",
  32130=>"111111110",
  32131=>"001000000",
  32132=>"000011010",
  32133=>"000000000",
  32134=>"000001001",
  32135=>"000000110",
  32136=>"001001001",
  32137=>"101001001",
  32138=>"111111111",
  32139=>"111110010",
  32140=>"111111110",
  32141=>"110100000",
  32142=>"110110000",
  32143=>"000000000",
  32144=>"001001000",
  32145=>"111100000",
  32146=>"110111000",
  32147=>"000000100",
  32148=>"111111000",
  32149=>"010000010",
  32150=>"111111001",
  32151=>"101111101",
  32152=>"000111110",
  32153=>"000111111",
  32154=>"111111000",
  32155=>"101000001",
  32156=>"101000000",
  32157=>"111111000",
  32158=>"111111011",
  32159=>"101011000",
  32160=>"110111111",
  32161=>"111111111",
  32162=>"111110110",
  32163=>"111110000",
  32164=>"000000000",
  32165=>"111111111",
  32166=>"111001000",
  32167=>"111011011",
  32168=>"000000000",
  32169=>"111111011",
  32170=>"010010110",
  32171=>"001000000",
  32172=>"000110110",
  32173=>"000000000",
  32174=>"000000100",
  32175=>"000000000",
  32176=>"001001001",
  32177=>"111111111",
  32178=>"010000000",
  32179=>"000000000",
  32180=>"000000000",
  32181=>"001000000",
  32182=>"111111011",
  32183=>"000000000",
  32184=>"000011111",
  32185=>"111110000",
  32186=>"111110110",
  32187=>"000000000",
  32188=>"101101100",
  32189=>"000000000",
  32190=>"000000111",
  32191=>"001000000",
  32192=>"000001011",
  32193=>"111111111",
  32194=>"001001111",
  32195=>"000000000",
  32196=>"000001001",
  32197=>"001110110",
  32198=>"101011111",
  32199=>"000000111",
  32200=>"001100100",
  32201=>"000000100",
  32202=>"110000010",
  32203=>"011111111",
  32204=>"111010000",
  32205=>"110111111",
  32206=>"110011000",
  32207=>"000011111",
  32208=>"100101001",
  32209=>"111111001",
  32210=>"111111110",
  32211=>"111111111",
  32212=>"111000100",
  32213=>"111111000",
  32214=>"100000000",
  32215=>"011000000",
  32216=>"001000100",
  32217=>"110000000",
  32218=>"000000000",
  32219=>"111101000",
  32220=>"110010011",
  32221=>"111111111",
  32222=>"100001011",
  32223=>"000100000",
  32224=>"111111111",
  32225=>"111111111",
  32226=>"001111111",
  32227=>"000000110",
  32228=>"111111111",
  32229=>"111111000",
  32230=>"111110111",
  32231=>"000100110",
  32232=>"100110110",
  32233=>"011111111",
  32234=>"000000110",
  32235=>"110111111",
  32236=>"100000000",
  32237=>"101101101",
  32238=>"101001000",
  32239=>"111101111",
  32240=>"000000100",
  32241=>"000010010",
  32242=>"110100000",
  32243=>"111111000",
  32244=>"000000000",
  32245=>"010111111",
  32246=>"011001011",
  32247=>"000111111",
  32248=>"000000100",
  32249=>"001001001",
  32250=>"110110110",
  32251=>"111111001",
  32252=>"011001010",
  32253=>"001111100",
  32254=>"010000000",
  32255=>"001000000",
  32256=>"111111111",
  32257=>"111111000",
  32258=>"000111111",
  32259=>"011100101",
  32260=>"000011111",
  32261=>"001001000",
  32262=>"001111101",
  32263=>"000000100",
  32264=>"111111111",
  32265=>"000000111",
  32266=>"111111111",
  32267=>"100100000",
  32268=>"000001111",
  32269=>"000000000",
  32270=>"000000111",
  32271=>"001011110",
  32272=>"110110111",
  32273=>"000000000",
  32274=>"110000000",
  32275=>"111111111",
  32276=>"111010000",
  32277=>"110010111",
  32278=>"011110110",
  32279=>"111110110",
  32280=>"000000001",
  32281=>"001100100",
  32282=>"111111111",
  32283=>"111111100",
  32284=>"000000000",
  32285=>"100000000",
  32286=>"011011001",
  32287=>"000000011",
  32288=>"000000000",
  32289=>"101001000",
  32290=>"110000000",
  32291=>"100100111",
  32292=>"111111000",
  32293=>"111100000",
  32294=>"101111111",
  32295=>"111110000",
  32296=>"111011001",
  32297=>"111111111",
  32298=>"110101000",
  32299=>"000000000",
  32300=>"111000000",
  32301=>"100100111",
  32302=>"000100100",
  32303=>"111111111",
  32304=>"000100000",
  32305=>"000000000",
  32306=>"101110110",
  32307=>"011111111",
  32308=>"111111000",
  32309=>"000111011",
  32310=>"000000111",
  32311=>"011010000",
  32312=>"000000000",
  32313=>"101000001",
  32314=>"000000000",
  32315=>"111111110",
  32316=>"111100100",
  32317=>"111110110",
  32318=>"001111111",
  32319=>"111011111",
  32320=>"000000101",
  32321=>"000000000",
  32322=>"000000000",
  32323=>"111000011",
  32324=>"001000000",
  32325=>"111111111",
  32326=>"100001111",
  32327=>"000001111",
  32328=>"111011010",
  32329=>"001000000",
  32330=>"000000000",
  32331=>"111111111",
  32332=>"000000000",
  32333=>"111101101",
  32334=>"000000000",
  32335=>"000010100",
  32336=>"111111111",
  32337=>"000000000",
  32338=>"000000000",
  32339=>"011000000",
  32340=>"000000000",
  32341=>"000111111",
  32342=>"000000000",
  32343=>"000000000",
  32344=>"001001000",
  32345=>"000000101",
  32346=>"000111111",
  32347=>"100100000",
  32348=>"000000000",
  32349=>"000000000",
  32350=>"011000110",
  32351=>"100000000",
  32352=>"000000000",
  32353=>"000000000",
  32354=>"111111111",
  32355=>"000000000",
  32356=>"000000000",
  32357=>"000001001",
  32358=>"000000000",
  32359=>"000000000",
  32360=>"111000000",
  32361=>"000000110",
  32362=>"011010000",
  32363=>"100111111",
  32364=>"111111111",
  32365=>"000100100",
  32366=>"110110111",
  32367=>"011111111",
  32368=>"000000000",
  32369=>"000000000",
  32370=>"100000000",
  32371=>"001001000",
  32372=>"111101000",
  32373=>"000001001",
  32374=>"000000000",
  32375=>"110100100",
  32376=>"000000000",
  32377=>"000100000",
  32378=>"000001101",
  32379=>"110000000",
  32380=>"110110110",
  32381=>"110111110",
  32382=>"111111000",
  32383=>"111111111",
  32384=>"000000000",
  32385=>"001000000",
  32386=>"111111111",
  32387=>"000110000",
  32388=>"110110111",
  32389=>"000000000",
  32390=>"000000000",
  32391=>"000111111",
  32392=>"111111111",
  32393=>"011010000",
  32394=>"111111000",
  32395=>"000000000",
  32396=>"111110100",
  32397=>"010011011",
  32398=>"111111111",
  32399=>"100111111",
  32400=>"110110110",
  32401=>"111111100",
  32402=>"000000000",
  32403=>"000000011",
  32404=>"111111010",
  32405=>"111111011",
  32406=>"011000000",
  32407=>"011011111",
  32408=>"000100000",
  32409=>"111111111",
  32410=>"100000000",
  32411=>"000100110",
  32412=>"111110110",
  32413=>"001100000",
  32414=>"111110000",
  32415=>"000000000",
  32416=>"011000001",
  32417=>"000000110",
  32418=>"011000000",
  32419=>"111111111",
  32420=>"011001101",
  32421=>"011000110",
  32422=>"111111110",
  32423=>"110110011",
  32424=>"000100111",
  32425=>"000000111",
  32426=>"111111111",
  32427=>"111111111",
  32428=>"000000000",
  32429=>"111111011",
  32430=>"001000000",
  32431=>"000000000",
  32432=>"111111110",
  32433=>"000001011",
  32434=>"111111111",
  32435=>"111111111",
  32436=>"111111101",
  32437=>"010100101",
  32438=>"111111111",
  32439=>"111000111",
  32440=>"111111111",
  32441=>"111111111",
  32442=>"000000000",
  32443=>"000000000",
  32444=>"110100100",
  32445=>"111100100",
  32446=>"000000110",
  32447=>"111100111",
  32448=>"100111111",
  32449=>"111001001",
  32450=>"000000000",
  32451=>"000000111",
  32452=>"011000000",
  32453=>"111111110",
  32454=>"001011111",
  32455=>"101101001",
  32456=>"000000000",
  32457=>"000000010",
  32458=>"110111000",
  32459=>"011001000",
  32460=>"001000000",
  32461=>"000111111",
  32462=>"000000110",
  32463=>"000001101",
  32464=>"000000101",
  32465=>"000000000",
  32466=>"111111000",
  32467=>"000000001",
  32468=>"001110110",
  32469=>"101111111",
  32470=>"010011111",
  32471=>"111110000",
  32472=>"001101111",
  32473=>"111111000",
  32474=>"000000010",
  32475=>"000000000",
  32476=>"111010000",
  32477=>"000000000",
  32478=>"110111111",
  32479=>"001001000",
  32480=>"000000110",
  32481=>"000000000",
  32482=>"000000000",
  32483=>"000000010",
  32484=>"000101000",
  32485=>"001001001",
  32486=>"111011011",
  32487=>"111000001",
  32488=>"111111111",
  32489=>"000000111",
  32490=>"111111101",
  32491=>"111110000",
  32492=>"000000111",
  32493=>"111111111",
  32494=>"000000000",
  32495=>"000001000",
  32496=>"111111111",
  32497=>"111111111",
  32498=>"011011000",
  32499=>"000101001",
  32500=>"111111111",
  32501=>"000000001",
  32502=>"111111111",
  32503=>"000000000",
  32504=>"000000000",
  32505=>"000100100",
  32506=>"000000000",
  32507=>"010100100",
  32508=>"110110110",
  32509=>"110000000",
  32510=>"001111111",
  32511=>"110100100",
  32512=>"110110110",
  32513=>"011111111",
  32514=>"001001100",
  32515=>"000000001",
  32516=>"111101000",
  32517=>"010011111",
  32518=>"111110110",
  32519=>"000001011",
  32520=>"111111111",
  32521=>"000000000",
  32522=>"011001100",
  32523=>"000000000",
  32524=>"111111101",
  32525=>"110111110",
  32526=>"000101000",
  32527=>"000000000",
  32528=>"111101101",
  32529=>"100010010",
  32530=>"100100000",
  32531=>"000101101",
  32532=>"000000000",
  32533=>"111011000",
  32534=>"111011010",
  32535=>"000000000",
  32536=>"000000000",
  32537=>"111111101",
  32538=>"111111111",
  32539=>"111010000",
  32540=>"100111111",
  32541=>"000000111",
  32542=>"111111111",
  32543=>"000010000",
  32544=>"100100000",
  32545=>"000001111",
  32546=>"111000000",
  32547=>"111011000",
  32548=>"000001001",
  32549=>"111111111",
  32550=>"011011111",
  32551=>"110110100",
  32552=>"000000000",
  32553=>"000000000",
  32554=>"100110110",
  32555=>"000111111",
  32556=>"000000000",
  32557=>"001001000",
  32558=>"111000000",
  32559=>"000000000",
  32560=>"111111100",
  32561=>"111111110",
  32562=>"111011111",
  32563=>"111111110",
  32564=>"000000000",
  32565=>"001111111",
  32566=>"000000000",
  32567=>"111111111",
  32568=>"111111001",
  32569=>"000000000",
  32570=>"111100111",
  32571=>"000000000",
  32572=>"001000000",
  32573=>"100100000",
  32574=>"001000000",
  32575=>"000000000",
  32576=>"000000000",
  32577=>"000110111",
  32578=>"110111111",
  32579=>"101111111",
  32580=>"111110110",
  32581=>"110010000",
  32582=>"001000000",
  32583=>"011111011",
  32584=>"110000000",
  32585=>"111111111",
  32586=>"101100000",
  32587=>"111101000",
  32588=>"111111000",
  32589=>"010000000",
  32590=>"101100100",
  32591=>"000001001",
  32592=>"011111000",
  32593=>"000100111",
  32594=>"000000000",
  32595=>"111111111",
  32596=>"000000000",
  32597=>"011000000",
  32598=>"011001000",
  32599=>"000000000",
  32600=>"111111111",
  32601=>"111111111",
  32602=>"011111011",
  32603=>"001001001",
  32604=>"110111111",
  32605=>"011111111",
  32606=>"100000000",
  32607=>"100000000",
  32608=>"101101111",
  32609=>"111111000",
  32610=>"100100110",
  32611=>"110100110",
  32612=>"100100110",
  32613=>"111111000",
  32614=>"111011000",
  32615=>"111111001",
  32616=>"111111011",
  32617=>"111001101",
  32618=>"100100111",
  32619=>"000011111",
  32620=>"111001001",
  32621=>"000000001",
  32622=>"000011000",
  32623=>"111000000",
  32624=>"000000111",
  32625=>"000010010",
  32626=>"000111111",
  32627=>"111110010",
  32628=>"111000000",
  32629=>"110000111",
  32630=>"111110111",
  32631=>"000000000",
  32632=>"000000000",
  32633=>"110110000",
  32634=>"000000011",
  32635=>"000000000",
  32636=>"000000111",
  32637=>"001000000",
  32638=>"000000001",
  32639=>"000000000",
  32640=>"110000100",
  32641=>"001000000",
  32642=>"111111111",
  32643=>"000000000",
  32644=>"000000000",
  32645=>"111111101",
  32646=>"011111111",
  32647=>"000000010",
  32648=>"000010111",
  32649=>"111001111",
  32650=>"111111111",
  32651=>"000000000",
  32652=>"111111111",
  32653=>"001001001",
  32654=>"111111000",
  32655=>"111111000",
  32656=>"010000100",
  32657=>"111110111",
  32658=>"111111111",
  32659=>"100110010",
  32660=>"000101001",
  32661=>"000000000",
  32662=>"100101000",
  32663=>"000000011",
  32664=>"000000000",
  32665=>"000001111",
  32666=>"000100111",
  32667=>"110110110",
  32668=>"011001001",
  32669=>"111111000",
  32670=>"011011001",
  32671=>"000000000",
  32672=>"000000000",
  32673=>"011111111",
  32674=>"000000010",
  32675=>"000000000",
  32676=>"001000100",
  32677=>"111100000",
  32678=>"000011111",
  32679=>"000001000",
  32680=>"000000101",
  32681=>"110000000",
  32682=>"110110110",
  32683=>"111111000",
  32684=>"000000000",
  32685=>"010000000",
  32686=>"001011011",
  32687=>"111111000",
  32688=>"001010111",
  32689=>"111111111",
  32690=>"011011011",
  32691=>"111000000",
  32692=>"111111111",
  32693=>"001000000",
  32694=>"111111111",
  32695=>"110111111",
  32696=>"011000000",
  32697=>"011011000",
  32698=>"000000000",
  32699=>"111111111",
  32700=>"100100111",
  32701=>"111111111",
  32702=>"000000000",
  32703=>"110110100",
  32704=>"110110000",
  32705=>"010010110",
  32706=>"111111111",
  32707=>"000100111",
  32708=>"000000001",
  32709=>"011111110",
  32710=>"001000000",
  32711=>"111111111",
  32712=>"000100000",
  32713=>"001101100",
  32714=>"000000010",
  32715=>"100111111",
  32716=>"000000000",
  32717=>"000000000",
  32718=>"000000000",
  32719=>"001000000",
  32720=>"110110000",
  32721=>"111111111",
  32722=>"011001000",
  32723=>"111100111",
  32724=>"111100100",
  32725=>"000001000",
  32726=>"111011000",
  32727=>"000010000",
  32728=>"110111111",
  32729=>"000000011",
  32730=>"111111111",
  32731=>"000000000",
  32732=>"110110100",
  32733=>"011111111",
  32734=>"100000000",
  32735=>"111111011",
  32736=>"000000111",
  32737=>"111111111",
  32738=>"000000000",
  32739=>"111011011",
  32740=>"111111111",
  32741=>"000100111",
  32742=>"000111000",
  32743=>"111111111",
  32744=>"000000000",
  32745=>"001100100",
  32746=>"111000000",
  32747=>"011111000",
  32748=>"000000000",
  32749=>"001111100",
  32750=>"010000000",
  32751=>"000000011",
  32752=>"000000011",
  32753=>"000000000",
  32754=>"111011000",
  32755=>"000001011",
  32756=>"001000000",
  32757=>"111011000",
  32758=>"111111111",
  32759=>"110011001",
  32760=>"000101111",
  32761=>"011011011",
  32762=>"011011011",
  32763=>"000000110",
  32764=>"111111111",
  32765=>"001000000",
  32766=>"000000000",
  32767=>"111111111",
  32768=>"000000100",
  32769=>"000000000",
  32770=>"110000000",
  32771=>"000000000",
  32772=>"000011000",
  32773=>"000000000",
  32774=>"000000000",
  32775=>"101000000",
  32776=>"000000101",
  32777=>"111011001",
  32778=>"110100010",
  32779=>"000000111",
  32780=>"101111110",
  32781=>"111111111",
  32782=>"000000000",
  32783=>"111111000",
  32784=>"000000000",
  32785=>"111111111",
  32786=>"000110111",
  32787=>"111111111",
  32788=>"111111111",
  32789=>"100100000",
  32790=>"111111001",
  32791=>"000001000",
  32792=>"110110110",
  32793=>"000000111",
  32794=>"000000000",
  32795=>"011111111",
  32796=>"111111111",
  32797=>"110111111",
  32798=>"011010000",
  32799=>"000101111",
  32800=>"001000111",
  32801=>"111001000",
  32802=>"100100000",
  32803=>"110000000",
  32804=>"000001011",
  32805=>"000000111",
  32806=>"101001000",
  32807=>"111100000",
  32808=>"111111011",
  32809=>"111111111",
  32810=>"000000000",
  32811=>"111111110",
  32812=>"000000101",
  32813=>"111111000",
  32814=>"000010111",
  32815=>"100000000",
  32816=>"111111111",
  32817=>"110001001",
  32818=>"111111001",
  32819=>"000000010",
  32820=>"100100111",
  32821=>"000101111",
  32822=>"100000000",
  32823=>"000000000",
  32824=>"010011110",
  32825=>"000101111",
  32826=>"010111111",
  32827=>"110110111",
  32828=>"101111111",
  32829=>"110110111",
  32830=>"000001000",
  32831=>"111101001",
  32832=>"000000000",
  32833=>"100100000",
  32834=>"111111111",
  32835=>"111111111",
  32836=>"100110100",
  32837=>"001011100",
  32838=>"111011110",
  32839=>"111111100",
  32840=>"111111000",
  32841=>"000000010",
  32842=>"010110110",
  32843=>"000000001",
  32844=>"000000000",
  32845=>"111000000",
  32846=>"000011000",
  32847=>"000000011",
  32848=>"111111000",
  32849=>"111111111",
  32850=>"000000000",
  32851=>"110110100",
  32852=>"111111010",
  32853=>"111111111",
  32854=>"110100000",
  32855=>"111111000",
  32856=>"000000001",
  32857=>"001100101",
  32858=>"000111111",
  32859=>"010001001",
  32860=>"111111111",
  32861=>"101111001",
  32862=>"000000000",
  32863=>"111111000",
  32864=>"111101100",
  32865=>"000000000",
  32866=>"111000000",
  32867=>"000001001",
  32868=>"110110111",
  32869=>"111111101",
  32870=>"000111101",
  32871=>"111111111",
  32872=>"000000000",
  32873=>"010111111",
  32874=>"000110110",
  32875=>"001111100",
  32876=>"000000001",
  32877=>"000000000",
  32878=>"101101111",
  32879=>"000110010",
  32880=>"111000000",
  32881=>"100101111",
  32882=>"100100000",
  32883=>"000000111",
  32884=>"000000110",
  32885=>"000000000",
  32886=>"111111111",
  32887=>"111111111",
  32888=>"000000111",
  32889=>"111111111",
  32890=>"000000000",
  32891=>"000000000",
  32892=>"110100100",
  32893=>"000000101",
  32894=>"111111110",
  32895=>"000000000",
  32896=>"111111000",
  32897=>"110110110",
  32898=>"111111111",
  32899=>"111111111",
  32900=>"000000001",
  32901=>"000010111",
  32902=>"111101111",
  32903=>"000000000",
  32904=>"000000110",
  32905=>"000111111",
  32906=>"000000111",
  32907=>"001001001",
  32908=>"100110111",
  32909=>"111111111",
  32910=>"001111111",
  32911=>"111111000",
  32912=>"000000111",
  32913=>"000000000",
  32914=>"111111111",
  32915=>"110100111",
  32916=>"001001000",
  32917=>"010000000",
  32918=>"000000100",
  32919=>"110100000",
  32920=>"000000000",
  32921=>"100000100",
  32922=>"111011011",
  32923=>"111111100",
  32924=>"100000000",
  32925=>"011000001",
  32926=>"111001111",
  32927=>"111111111",
  32928=>"111111111",
  32929=>"000110111",
  32930=>"111110000",
  32931=>"011010000",
  32932=>"000000000",
  32933=>"110101111",
  32934=>"101101001",
  32935=>"000000000",
  32936=>"000000100",
  32937=>"100000000",
  32938=>"000000101",
  32939=>"111111111",
  32940=>"111111111",
  32941=>"000110111",
  32942=>"000000101",
  32943=>"110011011",
  32944=>"010111000",
  32945=>"001011011",
  32946=>"111111111",
  32947=>"011001000",
  32948=>"111111111",
  32949=>"000010000",
  32950=>"100010000",
  32951=>"111111100",
  32952=>"111001111",
  32953=>"111111111",
  32954=>"000000000",
  32955=>"111110111",
  32956=>"110000001",
  32957=>"111111111",
  32958=>"000000001",
  32959=>"101111010",
  32960=>"111000000",
  32961=>"111111101",
  32962=>"000000000",
  32963=>"111111101",
  32964=>"111111111",
  32965=>"101101011",
  32966=>"011111111",
  32967=>"000000111",
  32968=>"111111001",
  32969=>"000000001",
  32970=>"000000000",
  32971=>"000000000",
  32972=>"111110000",
  32973=>"001001000",
  32974=>"100100100",
  32975=>"000000011",
  32976=>"100000000",
  32977=>"111111011",
  32978=>"100001011",
  32979=>"111111111",
  32980=>"011011100",
  32981=>"000000000",
  32982=>"001000000",
  32983=>"000000001",
  32984=>"000010111",
  32985=>"110110110",
  32986=>"000000000",
  32987=>"111001101",
  32988=>"000100100",
  32989=>"000000000",
  32990=>"000000001",
  32991=>"000000100",
  32992=>"000000111",
  32993=>"000110110",
  32994=>"111111111",
  32995=>"000000000",
  32996=>"011011010",
  32997=>"111100000",
  32998=>"101001111",
  32999=>"111111111",
  33000=>"000000111",
  33001=>"111111101",
  33002=>"110111111",
  33003=>"110111101",
  33004=>"000101111",
  33005=>"100111111",
  33006=>"101000100",
  33007=>"000100111",
  33008=>"111111111",
  33009=>"111111011",
  33010=>"000000000",
  33011=>"001000000",
  33012=>"111111111",
  33013=>"010100000",
  33014=>"100101100",
  33015=>"010111111",
  33016=>"111111110",
  33017=>"000000000",
  33018=>"000000000",
  33019=>"110100000",
  33020=>"000000000",
  33021=>"000000000",
  33022=>"111111111",
  33023=>"110100101",
  33024=>"100100100",
  33025=>"111111100",
  33026=>"000001111",
  33027=>"100000000",
  33028=>"111000111",
  33029=>"100111111",
  33030=>"001001111",
  33031=>"111111000",
  33032=>"110010000",
  33033=>"000000000",
  33034=>"111101111",
  33035=>"001000010",
  33036=>"001001111",
  33037=>"000000000",
  33038=>"010110110",
  33039=>"111111111",
  33040=>"000000000",
  33041=>"000000000",
  33042=>"101111110",
  33043=>"110110110",
  33044=>"000011111",
  33045=>"110110001",
  33046=>"111111110",
  33047=>"111111111",
  33048=>"111111110",
  33049=>"101110010",
  33050=>"010100000",
  33051=>"110110010",
  33052=>"100000000",
  33053=>"110100011",
  33054=>"000000111",
  33055=>"000000101",
  33056=>"001000000",
  33057=>"111111010",
  33058=>"111111011",
  33059=>"100000010",
  33060=>"111111001",
  33061=>"000000000",
  33062=>"000000000",
  33063=>"000010111",
  33064=>"000000111",
  33065=>"000000000",
  33066=>"111010010",
  33067=>"001101111",
  33068=>"111111000",
  33069=>"000000000",
  33070=>"111111010",
  33071=>"000000000",
  33072=>"111111111",
  33073=>"000010000",
  33074=>"111111111",
  33075=>"000000011",
  33076=>"000000000",
  33077=>"111111111",
  33078=>"000010111",
  33079=>"100111011",
  33080=>"000000100",
  33081=>"100000000",
  33082=>"111111101",
  33083=>"111111111",
  33084=>"100100100",
  33085=>"110111111",
  33086=>"011111100",
  33087=>"111111111",
  33088=>"111001111",
  33089=>"110110000",
  33090=>"000000111",
  33091=>"111111111",
  33092=>"110110000",
  33093=>"000000000",
  33094=>"011011000",
  33095=>"000111111",
  33096=>"001000111",
  33097=>"010000000",
  33098=>"111111111",
  33099=>"001000001",
  33100=>"111010000",
  33101=>"110111111",
  33102=>"111111111",
  33103=>"000000000",
  33104=>"000000000",
  33105=>"111111111",
  33106=>"111111111",
  33107=>"000110111",
  33108=>"000000000",
  33109=>"001011001",
  33110=>"111000000",
  33111=>"111111111",
  33112=>"111111000",
  33113=>"111111111",
  33114=>"111111000",
  33115=>"000000000",
  33116=>"111111011",
  33117=>"111111010",
  33118=>"110000000",
  33119=>"110110100",
  33120=>"100011000",
  33121=>"111111100",
  33122=>"111100001",
  33123=>"111000000",
  33124=>"101001001",
  33125=>"001000000",
  33126=>"000000010",
  33127=>"000000000",
  33128=>"110110100",
  33129=>"111111110",
  33130=>"000000000",
  33131=>"111000000",
  33132=>"110100100",
  33133=>"100111111",
  33134=>"111000001",
  33135=>"000111111",
  33136=>"111111111",
  33137=>"100110111",
  33138=>"000000000",
  33139=>"111001000",
  33140=>"010000000",
  33141=>"100111101",
  33142=>"001000111",
  33143=>"111111000",
  33144=>"111100000",
  33145=>"000101001",
  33146=>"111111111",
  33147=>"110111111",
  33148=>"000000000",
  33149=>"000000101",
  33150=>"001000000",
  33151=>"000000100",
  33152=>"111001000",
  33153=>"100000000",
  33154=>"111110110",
  33155=>"000000000",
  33156=>"111011111",
  33157=>"010000000",
  33158=>"000000100",
  33159=>"000000111",
  33160=>"000100100",
  33161=>"111111111",
  33162=>"000000100",
  33163=>"100111110",
  33164=>"111111111",
  33165=>"111111000",
  33166=>"000000000",
  33167=>"111111111",
  33168=>"001001000",
  33169=>"000000000",
  33170=>"111011011",
  33171=>"001001000",
  33172=>"111111111",
  33173=>"011000000",
  33174=>"001001111",
  33175=>"000000011",
  33176=>"000000000",
  33177=>"111110000",
  33178=>"111110100",
  33179=>"000000000",
  33180=>"111111010",
  33181=>"111111111",
  33182=>"111011001",
  33183=>"000000101",
  33184=>"000000000",
  33185=>"110110000",
  33186=>"000000000",
  33187=>"000000000",
  33188=>"111001101",
  33189=>"010111110",
  33190=>"111111001",
  33191=>"010010000",
  33192=>"111010000",
  33193=>"000000000",
  33194=>"111111111",
  33195=>"011001001",
  33196=>"000000000",
  33197=>"000000000",
  33198=>"111111111",
  33199=>"000000000",
  33200=>"000000000",
  33201=>"100111111",
  33202=>"000000010",
  33203=>"011111111",
  33204=>"111011011",
  33205=>"000000000",
  33206=>"111101100",
  33207=>"000000111",
  33208=>"111111111",
  33209=>"000000000",
  33210=>"000110010",
  33211=>"101000000",
  33212=>"000000000",
  33213=>"001001001",
  33214=>"100100100",
  33215=>"111100000",
  33216=>"110010110",
  33217=>"111111111",
  33218=>"000001001",
  33219=>"001001101",
  33220=>"110110111",
  33221=>"001001011",
  33222=>"111111111",
  33223=>"111111111",
  33224=>"000000000",
  33225=>"110111000",
  33226=>"000000100",
  33227=>"000000000",
  33228=>"111111010",
  33229=>"111111011",
  33230=>"000000010",
  33231=>"000111111",
  33232=>"000111111",
  33233=>"000101011",
  33234=>"000000110",
  33235=>"011111111",
  33236=>"001001001",
  33237=>"111110111",
  33238=>"000000111",
  33239=>"001001000",
  33240=>"000000000",
  33241=>"010001011",
  33242=>"000000000",
  33243=>"111111111",
  33244=>"000000000",
  33245=>"001000000",
  33246=>"000001000",
  33247=>"111000100",
  33248=>"100000000",
  33249=>"000000000",
  33250=>"000000000",
  33251=>"000000100",
  33252=>"001000000",
  33253=>"111100001",
  33254=>"010000000",
  33255=>"111010000",
  33256=>"000010111",
  33257=>"000000000",
  33258=>"101000101",
  33259=>"000000000",
  33260=>"100100011",
  33261=>"000000000",
  33262=>"111111111",
  33263=>"001001011",
  33264=>"011011001",
  33265=>"111111100",
  33266=>"010011011",
  33267=>"111101100",
  33268=>"000011111",
  33269=>"111000000",
  33270=>"111000000",
  33271=>"100110111",
  33272=>"100110000",
  33273=>"111111111",
  33274=>"000000000",
  33275=>"100111111",
  33276=>"010000000",
  33277=>"111111110",
  33278=>"001111111",
  33279=>"111011011",
  33280=>"110000110",
  33281=>"000000110",
  33282=>"111111111",
  33283=>"000000001",
  33284=>"111111111",
  33285=>"101100110",
  33286=>"101000000",
  33287=>"001000000",
  33288=>"001000000",
  33289=>"010011011",
  33290=>"101001000",
  33291=>"000000000",
  33292=>"111111111",
  33293=>"111010100",
  33294=>"000000001",
  33295=>"111111111",
  33296=>"100110110",
  33297=>"000001111",
  33298=>"000001001",
  33299=>"011111011",
  33300=>"101101101",
  33301=>"001000111",
  33302=>"000000001",
  33303=>"100100001",
  33304=>"111000111",
  33305=>"011000000",
  33306=>"000000010",
  33307=>"111111111",
  33308=>"000000000",
  33309=>"011000101",
  33310=>"110000000",
  33311=>"001001000",
  33312=>"111111001",
  33313=>"110010010",
  33314=>"111110001",
  33315=>"000000000",
  33316=>"111110000",
  33317=>"111111100",
  33318=>"111010000",
  33319=>"010111111",
  33320=>"111011111",
  33321=>"000000000",
  33322=>"000000000",
  33323=>"000011111",
  33324=>"000000000",
  33325=>"000000000",
  33326=>"101111111",
  33327=>"100111111",
  33328=>"000000100",
  33329=>"000001001",
  33330=>"000000000",
  33331=>"011001101",
  33332=>"000000000",
  33333=>"110110111",
  33334=>"000000100",
  33335=>"111111111",
  33336=>"011011001",
  33337=>"111111110",
  33338=>"100000100",
  33339=>"000000110",
  33340=>"111100111",
  33341=>"111111111",
  33342=>"000011011",
  33343=>"000000000",
  33344=>"011001000",
  33345=>"000111111",
  33346=>"101100000",
  33347=>"000111011",
  33348=>"100100110",
  33349=>"111111000",
  33350=>"000001001",
  33351=>"000000000",
  33352=>"010000000",
  33353=>"111101111",
  33354=>"111011111",
  33355=>"011111010",
  33356=>"000010111",
  33357=>"111111000",
  33358=>"101000000",
  33359=>"000111111",
  33360=>"000000000",
  33361=>"000001100",
  33362=>"111111111",
  33363=>"100110100",
  33364=>"001001011",
  33365=>"011000000",
  33366=>"110110010",
  33367=>"110111111",
  33368=>"000010000",
  33369=>"111100100",
  33370=>"011011000",
  33371=>"111011011",
  33372=>"111111111",
  33373=>"111011000",
  33374=>"000000001",
  33375=>"001000100",
  33376=>"100111110",
  33377=>"100000000",
  33378=>"000000000",
  33379=>"000000100",
  33380=>"000000001",
  33381=>"011111000",
  33382=>"100110111",
  33383=>"101001111",
  33384=>"000000000",
  33385=>"000000111",
  33386=>"001000000",
  33387=>"000000011",
  33388=>"000000110",
  33389=>"111111111",
  33390=>"001111111",
  33391=>"111111110",
  33392=>"110000110",
  33393=>"000000111",
  33394=>"011001001",
  33395=>"101100111",
  33396=>"000000000",
  33397=>"111111101",
  33398=>"001000000",
  33399=>"111111111",
  33400=>"111111111",
  33401=>"111111001",
  33402=>"001001000",
  33403=>"111111111",
  33404=>"110100110",
  33405=>"111101001",
  33406=>"001110000",
  33407=>"010110110",
  33408=>"000111111",
  33409=>"001001111",
  33410=>"000000000",
  33411=>"001001000",
  33412=>"000000100",
  33413=>"111100100",
  33414=>"110100000",
  33415=>"000110110",
  33416=>"110111111",
  33417=>"000000000",
  33418=>"111000000",
  33419=>"111111100",
  33420=>"000000000",
  33421=>"111111110",
  33422=>"111000000",
  33423=>"001001011",
  33424=>"111111000",
  33425=>"111111111",
  33426=>"111111000",
  33427=>"111111010",
  33428=>"111111011",
  33429=>"110000000",
  33430=>"001001000",
  33431=>"110010000",
  33432=>"011011001",
  33433=>"010110000",
  33434=>"111110111",
  33435=>"000000000",
  33436=>"111011111",
  33437=>"100110111",
  33438=>"000000011",
  33439=>"101101000",
  33440=>"111111111",
  33441=>"111100110",
  33442=>"000000000",
  33443=>"111111111",
  33444=>"000100110",
  33445=>"111111111",
  33446=>"100000000",
  33447=>"111111111",
  33448=>"010010000",
  33449=>"000000000",
  33450=>"001001000",
  33451=>"011010110",
  33452=>"000001010",
  33453=>"000000000",
  33454=>"011011111",
  33455=>"000000111",
  33456=>"000111111",
  33457=>"001001011",
  33458=>"000101000",
  33459=>"000000000",
  33460=>"111100110",
  33461=>"010000000",
  33462=>"010000000",
  33463=>"000000000",
  33464=>"000101111",
  33465=>"000111111",
  33466=>"001111111",
  33467=>"010010110",
  33468=>"111111111",
  33469=>"000001111",
  33470=>"111111000",
  33471=>"111100100",
  33472=>"100000000",
  33473=>"111011001",
  33474=>"000000011",
  33475=>"000000000",
  33476=>"111111111",
  33477=>"011010000",
  33478=>"010010000",
  33479=>"000010000",
  33480=>"000000000",
  33481=>"100100100",
  33482=>"111111100",
  33483=>"001000000",
  33484=>"111111111",
  33485=>"001111100",
  33486=>"000000000",
  33487=>"000000000",
  33488=>"011011111",
  33489=>"111111110",
  33490=>"111111110",
  33491=>"111101101",
  33492=>"000100111",
  33493=>"111111111",
  33494=>"110000010",
  33495=>"111111010",
  33496=>"111111111",
  33497=>"111111001",
  33498=>"111111111",
  33499=>"111011111",
  33500=>"110110111",
  33501=>"000000001",
  33502=>"111100101",
  33503=>"000010010",
  33504=>"000000000",
  33505=>"001111111",
  33506=>"101101010",
  33507=>"111000000",
  33508=>"111011001",
  33509=>"011011110",
  33510=>"010110000",
  33511=>"000000000",
  33512=>"000000000",
  33513=>"000001011",
  33514=>"001000001",
  33515=>"001000000",
  33516=>"110000000",
  33517=>"111111111",
  33518=>"101100100",
  33519=>"000000000",
  33520=>"011011111",
  33521=>"111011111",
  33522=>"101000000",
  33523=>"110110111",
  33524=>"000001000",
  33525=>"111111101",
  33526=>"011111111",
  33527=>"000000000",
  33528=>"111111111",
  33529=>"110110110",
  33530=>"111110000",
  33531=>"010010000",
  33532=>"111011001",
  33533=>"110100100",
  33534=>"011000110",
  33535=>"101001000",
  33536=>"100111111",
  33537=>"010010000",
  33538=>"111111111",
  33539=>"000100100",
  33540=>"111111111",
  33541=>"001001111",
  33542=>"000000000",
  33543=>"111100000",
  33544=>"000000000",
  33545=>"000100100",
  33546=>"111000000",
  33547=>"111000001",
  33548=>"000000000",
  33549=>"000000000",
  33550=>"111111000",
  33551=>"000000001",
  33552=>"000000000",
  33553=>"111011111",
  33554=>"001000000",
  33555=>"100111111",
  33556=>"000000000",
  33557=>"100100100",
  33558=>"000000100",
  33559=>"111111001",
  33560=>"010010010",
  33561=>"000010111",
  33562=>"111111111",
  33563=>"111011000",
  33564=>"000000000",
  33565=>"000000000",
  33566=>"101101101",
  33567=>"111001111",
  33568=>"011111111",
  33569=>"000000000",
  33570=>"100101111",
  33571=>"001001111",
  33572=>"000000100",
  33573=>"100100100",
  33574=>"000001001",
  33575=>"100000001",
  33576=>"000000100",
  33577=>"001001001",
  33578=>"100000110",
  33579=>"001011000",
  33580=>"001011011",
  33581=>"000011011",
  33582=>"000000000",
  33583=>"000000000",
  33584=>"111011111",
  33585=>"000000000",
  33586=>"000000011",
  33587=>"111111111",
  33588=>"111111111",
  33589=>"101111101",
  33590=>"011011001",
  33591=>"110100000",
  33592=>"000000000",
  33593=>"000000000",
  33594=>"111001011",
  33595=>"000000000",
  33596=>"000000000",
  33597=>"010010000",
  33598=>"111000000",
  33599=>"001001001",
  33600=>"111111110",
  33601=>"000000000",
  33602=>"110110110",
  33603=>"111111111",
  33604=>"010000000",
  33605=>"111011000",
  33606=>"111000000",
  33607=>"000000000",
  33608=>"010010000",
  33609=>"000000000",
  33610=>"100000110",
  33611=>"000000000",
  33612=>"110000001",
  33613=>"111111011",
  33614=>"000000000",
  33615=>"010011111",
  33616=>"111110110",
  33617=>"111101000",
  33618=>"000000000",
  33619=>"111111111",
  33620=>"111111111",
  33621=>"001000001",
  33622=>"111111001",
  33623=>"001000000",
  33624=>"000000100",
  33625=>"111000000",
  33626=>"000000000",
  33627=>"000000111",
  33628=>"000000000",
  33629=>"011011001",
  33630=>"111111111",
  33631=>"111111011",
  33632=>"111011110",
  33633=>"000000000",
  33634=>"000010000",
  33635=>"000011011",
  33636=>"001000000",
  33637=>"000100111",
  33638=>"000111111",
  33639=>"001011011",
  33640=>"011001000",
  33641=>"000011000",
  33642=>"000111111",
  33643=>"000111110",
  33644=>"001000011",
  33645=>"000001011",
  33646=>"111111111",
  33647=>"000010000",
  33648=>"111111111",
  33649=>"111111010",
  33650=>"001000101",
  33651=>"001001000",
  33652=>"011011010",
  33653=>"000010110",
  33654=>"000000000",
  33655=>"011111111",
  33656=>"111000000",
  33657=>"110001001",
  33658=>"111111111",
  33659=>"111111111",
  33660=>"110111100",
  33661=>"111111111",
  33662=>"011011000",
  33663=>"111111111",
  33664=>"110100110",
  33665=>"000000000",
  33666=>"111111111",
  33667=>"111111101",
  33668=>"111101111",
  33669=>"100100110",
  33670=>"000000000",
  33671=>"100000001",
  33672=>"111111011",
  33673=>"111111111",
  33674=>"111111111",
  33675=>"111101101",
  33676=>"000001111",
  33677=>"011011110",
  33678=>"000000100",
  33679=>"000000000",
  33680=>"000000100",
  33681=>"010100111",
  33682=>"111111111",
  33683=>"111110000",
  33684=>"111111111",
  33685=>"000000000",
  33686=>"100110111",
  33687=>"000000000",
  33688=>"111111111",
  33689=>"000000000",
  33690=>"001000001",
  33691=>"111111001",
  33692=>"100000000",
  33693=>"010000111",
  33694=>"111111010",
  33695=>"001111101",
  33696=>"111000000",
  33697=>"111001001",
  33698=>"100000100",
  33699=>"111111111",
  33700=>"000000000",
  33701=>"000000000",
  33702=>"111111111",
  33703=>"111111111",
  33704=>"000001101",
  33705=>"001111111",
  33706=>"000000000",
  33707=>"000111111",
  33708=>"110000000",
  33709=>"101000100",
  33710=>"011000000",
  33711=>"000000000",
  33712=>"000000000",
  33713=>"010111110",
  33714=>"111111111",
  33715=>"011111111",
  33716=>"000000000",
  33717=>"111111101",
  33718=>"111001011",
  33719=>"000000000",
  33720=>"110110110",
  33721=>"000000000",
  33722=>"100100101",
  33723=>"111111010",
  33724=>"000000000",
  33725=>"000000000",
  33726=>"000000000",
  33727=>"000000000",
  33728=>"111111111",
  33729=>"000000000",
  33730=>"000000000",
  33731=>"111000000",
  33732=>"111111110",
  33733=>"111011000",
  33734=>"000000110",
  33735=>"011011000",
  33736=>"011111111",
  33737=>"000000000",
  33738=>"001000000",
  33739=>"000000000",
  33740=>"000000100",
  33741=>"110111110",
  33742=>"100110111",
  33743=>"111100110",
  33744=>"000000000",
  33745=>"001111000",
  33746=>"111111111",
  33747=>"000000111",
  33748=>"000001001",
  33749=>"111111111",
  33750=>"111111001",
  33751=>"111111111",
  33752=>"111101111",
  33753=>"101001000",
  33754=>"000000000",
  33755=>"000000000",
  33756=>"111111111",
  33757=>"000000001",
  33758=>"011111000",
  33759=>"111111101",
  33760=>"000010000",
  33761=>"100101000",
  33762=>"111111111",
  33763=>"001111111",
  33764=>"110111100",
  33765=>"000000000",
  33766=>"111111111",
  33767=>"111111111",
  33768=>"110010010",
  33769=>"000000110",
  33770=>"000100100",
  33771=>"000000000",
  33772=>"000110111",
  33773=>"001000000",
  33774=>"111111111",
  33775=>"000000000",
  33776=>"000000000",
  33777=>"100101111",
  33778=>"111111111",
  33779=>"111111100",
  33780=>"111111111",
  33781=>"000000111",
  33782=>"000000000",
  33783=>"000000110",
  33784=>"100000000",
  33785=>"000010000",
  33786=>"101100110",
  33787=>"011011000",
  33788=>"010110100",
  33789=>"100110100",
  33790=>"011111111",
  33791=>"110110110",
  33792=>"000000001",
  33793=>"000000000",
  33794=>"111000001",
  33795=>"110111111",
  33796=>"111111111",
  33797=>"011000011",
  33798=>"011111111",
  33799=>"000001111",
  33800=>"111000000",
  33801=>"010011011",
  33802=>"100000001",
  33803=>"011011001",
  33804=>"110111111",
  33805=>"111111000",
  33806=>"000000001",
  33807=>"111000111",
  33808=>"000000001",
  33809=>"010110100",
  33810=>"110111000",
  33811=>"000000111",
  33812=>"000000011",
  33813=>"011001000",
  33814=>"000000111",
  33815=>"100100110",
  33816=>"100000110",
  33817=>"000000011",
  33818=>"000111100",
  33819=>"000000000",
  33820=>"111111011",
  33821=>"110011000",
  33822=>"011011101",
  33823=>"011000000",
  33824=>"000000000",
  33825=>"001000001",
  33826=>"111011000",
  33827=>"000000101",
  33828=>"011000000",
  33829=>"001000000",
  33830=>"110111111",
  33831=>"000000101",
  33832=>"100111110",
  33833=>"100000000",
  33834=>"000000101",
  33835=>"001011000",
  33836=>"000111111",
  33837=>"000111000",
  33838=>"011011000",
  33839=>"000000000",
  33840=>"100100000",
  33841=>"000000000",
  33842=>"110111111",
  33843=>"110000000",
  33844=>"000000000",
  33845=>"000000110",
  33846=>"111011000",
  33847=>"111001101",
  33848=>"111111111",
  33849=>"000001101",
  33850=>"010000000",
  33851=>"001111111",
  33852=>"101100000",
  33853=>"000000000",
  33854=>"000000000",
  33855=>"000001111",
  33856=>"100000000",
  33857=>"000111111",
  33858=>"000000111",
  33859=>"001001001",
  33860=>"000001001",
  33861=>"001111111",
  33862=>"010110110",
  33863=>"001101000",
  33864=>"000000100",
  33865=>"000010000",
  33866=>"000000000",
  33867=>"000000000",
  33868=>"110111011",
  33869=>"101101000",
  33870=>"001001000",
  33871=>"011111111",
  33872=>"100000010",
  33873=>"100111111",
  33874=>"000000000",
  33875=>"111111111",
  33876=>"000111111",
  33877=>"110110100",
  33878=>"111111000",
  33879=>"111111000",
  33880=>"111111000",
  33881=>"000100100",
  33882=>"000110111",
  33883=>"100000100",
  33884=>"000000111",
  33885=>"100000111",
  33886=>"011011111",
  33887=>"111111111",
  33888=>"111111011",
  33889=>"111111001",
  33890=>"000000000",
  33891=>"111111010",
  33892=>"000000000",
  33893=>"000111111",
  33894=>"010011111",
  33895=>"010000000",
  33896=>"000000000",
  33897=>"001000000",
  33898=>"000000110",
  33899=>"000000000",
  33900=>"000000000",
  33901=>"000000111",
  33902=>"111111111",
  33903=>"111101100",
  33904=>"111111111",
  33905=>"000100111",
  33906=>"101110100",
  33907=>"111111011",
  33908=>"000000000",
  33909=>"000001001",
  33910=>"010111111",
  33911=>"000111011",
  33912=>"000000000",
  33913=>"000001011",
  33914=>"110111111",
  33915=>"000000000",
  33916=>"011001111",
  33917=>"000000000",
  33918=>"010111111",
  33919=>"000000000",
  33920=>"011011000",
  33921=>"000001001",
  33922=>"111111110",
  33923=>"111111000",
  33924=>"100111011",
  33925=>"001000000",
  33926=>"000001001",
  33927=>"111100100",
  33928=>"111111000",
  33929=>"100100111",
  33930=>"000000000",
  33931=>"111111000",
  33932=>"000010000",
  33933=>"001011001",
  33934=>"111111011",
  33935=>"111111111",
  33936=>"001000111",
  33937=>"111010000",
  33938=>"000000110",
  33939=>"111111000",
  33940=>"000111001",
  33941=>"111100000",
  33942=>"001000000",
  33943=>"000000000",
  33944=>"000000100",
  33945=>"011001000",
  33946=>"000000100",
  33947=>"100000000",
  33948=>"111111111",
  33949=>"110100111",
  33950=>"111001011",
  33951=>"011001011",
  33952=>"111111110",
  33953=>"000011011",
  33954=>"111111111",
  33955=>"111110111",
  33956=>"010010011",
  33957=>"001000011",
  33958=>"000000000",
  33959=>"111001111",
  33960=>"000111111",
  33961=>"000000000",
  33962=>"111000001",
  33963=>"010111000",
  33964=>"100001111",
  33965=>"000000000",
  33966=>"100001000",
  33967=>"000100100",
  33968=>"011111111",
  33969=>"011000000",
  33970=>"101101000",
  33971=>"100000000",
  33972=>"000010011",
  33973=>"000001100",
  33974=>"111111000",
  33975=>"111000000",
  33976=>"000011010",
  33977=>"000110110",
  33978=>"111100111",
  33979=>"111001111",
  33980=>"111111111",
  33981=>"001000000",
  33982=>"010000001",
  33983=>"111000000",
  33984=>"100000000",
  33985=>"110011000",
  33986=>"111000001",
  33987=>"111001000",
  33988=>"001000000",
  33989=>"110000000",
  33990=>"110110111",
  33991=>"111111011",
  33992=>"100111001",
  33993=>"111111111",
  33994=>"000111011",
  33995=>"000000001",
  33996=>"100000000",
  33997=>"111100100",
  33998=>"000000111",
  33999=>"110000111",
  34000=>"111111000",
  34001=>"001000000",
  34002=>"011011010",
  34003=>"111010000",
  34004=>"000000111",
  34005=>"111101100",
  34006=>"000000000",
  34007=>"000110110",
  34008=>"000011000",
  34009=>"000000011",
  34010=>"111000000",
  34011=>"111111111",
  34012=>"100000111",
  34013=>"000110010",
  34014=>"111111111",
  34015=>"111001111",
  34016=>"000000111",
  34017=>"000001011",
  34018=>"000110111",
  34019=>"000000000",
  34020=>"000111101",
  34021=>"111110110",
  34022=>"001000000",
  34023=>"000000000",
  34024=>"000001111",
  34025=>"001001111",
  34026=>"000000000",
  34027=>"111000001",
  34028=>"000110000",
  34029=>"101100100",
  34030=>"111011011",
  34031=>"111000000",
  34032=>"011000000",
  34033=>"111000000",
  34034=>"111111000",
  34035=>"100000001",
  34036=>"001000111",
  34037=>"000111110",
  34038=>"100111001",
  34039=>"111011001",
  34040=>"000000110",
  34041=>"100000000",
  34042=>"000000010",
  34043=>"011011001",
  34044=>"000011010",
  34045=>"001011001",
  34046=>"101000101",
  34047=>"010110111",
  34048=>"000000000",
  34049=>"100110110",
  34050=>"100011001",
  34051=>"100000111",
  34052=>"000000111",
  34053=>"000111000",
  34054=>"011001111",
  34055=>"001111111",
  34056=>"001000100",
  34057=>"000000000",
  34058=>"111110111",
  34059=>"111111011",
  34060=>"000000000",
  34061=>"111111111",
  34062=>"111111010",
  34063=>"111100000",
  34064=>"111011100",
  34065=>"111100000",
  34066=>"000000000",
  34067=>"111110000",
  34068=>"010110111",
  34069=>"000111000",
  34070=>"111111111",
  34071=>"000010010",
  34072=>"100111111",
  34073=>"111000000",
  34074=>"001000000",
  34075=>"000000001",
  34076=>"101101001",
  34077=>"110100000",
  34078=>"000000000",
  34079=>"111110010",
  34080=>"000000000",
  34081=>"000000001",
  34082=>"111111000",
  34083=>"100100100",
  34084=>"011111111",
  34085=>"100000001",
  34086=>"111100000",
  34087=>"000000001",
  34088=>"000000011",
  34089=>"000000000",
  34090=>"000100000",
  34091=>"000000111",
  34092=>"101101100",
  34093=>"011011000",
  34094=>"000000000",
  34095=>"000000010",
  34096=>"000100011",
  34097=>"111111100",
  34098=>"100100001",
  34099=>"100111000",
  34100=>"000000000",
  34101=>"000000000",
  34102=>"111001000",
  34103=>"111111111",
  34104=>"000111111",
  34105=>"000000001",
  34106=>"000000000",
  34107=>"111111111",
  34108=>"111111111",
  34109=>"000000000",
  34110=>"000000001",
  34111=>"000000000",
  34112=>"111101100",
  34113=>"100001111",
  34114=>"111001111",
  34115=>"000010000",
  34116=>"101011000",
  34117=>"110111111",
  34118=>"000000011",
  34119=>"000100000",
  34120=>"111111111",
  34121=>"010000000",
  34122=>"100111000",
  34123=>"000000000",
  34124=>"111101001",
  34125=>"000000111",
  34126=>"111000111",
  34127=>"000101111",
  34128=>"111100101",
  34129=>"000111111",
  34130=>"000000000",
  34131=>"100000011",
  34132=>"000010000",
  34133=>"001000010",
  34134=>"000000000",
  34135=>"101010111",
  34136=>"000111110",
  34137=>"100000000",
  34138=>"100111011",
  34139=>"000000000",
  34140=>"110000110",
  34141=>"000000111",
  34142=>"000000000",
  34143=>"101111111",
  34144=>"001001000",
  34145=>"111111111",
  34146=>"110111111",
  34147=>"000100000",
  34148=>"101110000",
  34149=>"111000000",
  34150=>"111111111",
  34151=>"111111111",
  34152=>"100000000",
  34153=>"011000000",
  34154=>"000100001",
  34155=>"111110100",
  34156=>"110001000",
  34157=>"111000111",
  34158=>"000000000",
  34159=>"111111111",
  34160=>"111000000",
  34161=>"111111111",
  34162=>"111001011",
  34163=>"011011000",
  34164=>"111001101",
  34165=>"000000000",
  34166=>"111111100",
  34167=>"111000000",
  34168=>"111111111",
  34169=>"111111111",
  34170=>"000000000",
  34171=>"111000100",
  34172=>"011011010",
  34173=>"110000000",
  34174=>"001000001",
  34175=>"001101111",
  34176=>"110111100",
  34177=>"111110100",
  34178=>"001011001",
  34179=>"000000000",
  34180=>"000000111",
  34181=>"000000001",
  34182=>"110110101",
  34183=>"000110111",
  34184=>"000000000",
  34185=>"110000100",
  34186=>"111111010",
  34187=>"000010000",
  34188=>"000000110",
  34189=>"111010000",
  34190=>"111111000",
  34191=>"000111000",
  34192=>"000000110",
  34193=>"110001001",
  34194=>"000000000",
  34195=>"111001111",
  34196=>"001011111",
  34197=>"011001001",
  34198=>"111111011",
  34199=>"111011111",
  34200=>"001111111",
  34201=>"110111111",
  34202=>"000111111",
  34203=>"001010000",
  34204=>"101001010",
  34205=>"111111001",
  34206=>"111001000",
  34207=>"111100000",
  34208=>"000000111",
  34209=>"100100110",
  34210=>"001011111",
  34211=>"001001001",
  34212=>"000111111",
  34213=>"111101111",
  34214=>"000111100",
  34215=>"111000001",
  34216=>"111111000",
  34217=>"100111011",
  34218=>"111111010",
  34219=>"111000000",
  34220=>"000000000",
  34221=>"101000000",
  34222=>"101001111",
  34223=>"111011111",
  34224=>"000000000",
  34225=>"000111101",
  34226=>"111111011",
  34227=>"000111111",
  34228=>"111111000",
  34229=>"000000001",
  34230=>"110111000",
  34231=>"111111000",
  34232=>"000001000",
  34233=>"100111111",
  34234=>"000111111",
  34235=>"000100110",
  34236=>"011111000",
  34237=>"110111111",
  34238=>"111011000",
  34239=>"100001110",
  34240=>"100100000",
  34241=>"000000000",
  34242=>"111001111",
  34243=>"001101101",
  34244=>"001000110",
  34245=>"001011111",
  34246=>"000001101",
  34247=>"000000010",
  34248=>"111111110",
  34249=>"000000111",
  34250=>"001111010",
  34251=>"111111111",
  34252=>"000000000",
  34253=>"000000001",
  34254=>"100011000",
  34255=>"001111000",
  34256=>"111110000",
  34257=>"000000111",
  34258=>"000000111",
  34259=>"101100111",
  34260=>"011011101",
  34261=>"100000101",
  34262=>"001000011",
  34263=>"011110010",
  34264=>"111110110",
  34265=>"000011111",
  34266=>"110110111",
  34267=>"111111000",
  34268=>"111111101",
  34269=>"001111100",
  34270=>"000000010",
  34271=>"011011010",
  34272=>"101111110",
  34273=>"011111111",
  34274=>"111111111",
  34275=>"001011001",
  34276=>"100111111",
  34277=>"000010101",
  34278=>"000011101",
  34279=>"111000110",
  34280=>"000000000",
  34281=>"111111111",
  34282=>"111000100",
  34283=>"001011001",
  34284=>"000000110",
  34285=>"011011011",
  34286=>"111101101",
  34287=>"000000000",
  34288=>"000000010",
  34289=>"110000000",
  34290=>"011111111",
  34291=>"000100100",
  34292=>"111011000",
  34293=>"111100000",
  34294=>"111111111",
  34295=>"001011000",
  34296=>"111000001",
  34297=>"010110110",
  34298=>"111111111",
  34299=>"000001000",
  34300=>"110100101",
  34301=>"100000011",
  34302=>"101111111",
  34303=>"000000000",
  34304=>"000000001",
  34305=>"110110100",
  34306=>"111101111",
  34307=>"001000001",
  34308=>"111111001",
  34309=>"100100101",
  34310=>"011111101",
  34311=>"111111111",
  34312=>"101001001",
  34313=>"000011111",
  34314=>"000000000",
  34315=>"111111111",
  34316=>"100111110",
  34317=>"111101100",
  34318=>"101111011",
  34319=>"010001011",
  34320=>"111111100",
  34321=>"000111111",
  34322=>"000000000",
  34323=>"000100000",
  34324=>"000000111",
  34325=>"111100000",
  34326=>"110110111",
  34327=>"111110110",
  34328=>"111111110",
  34329=>"101111111",
  34330=>"111111111",
  34331=>"011111111",
  34332=>"100000000",
  34333=>"000100100",
  34334=>"000001001",
  34335=>"101111011",
  34336=>"000000100",
  34337=>"110111111",
  34338=>"111110000",
  34339=>"111111110",
  34340=>"011000000",
  34341=>"000001001",
  34342=>"000000000",
  34343=>"000000011",
  34344=>"001011111",
  34345=>"000000000",
  34346=>"011111111",
  34347=>"000000111",
  34348=>"111111110",
  34349=>"111111000",
  34350=>"000001001",
  34351=>"111111111",
  34352=>"000100111",
  34353=>"000000001",
  34354=>"000100000",
  34355=>"010000000",
  34356=>"000000000",
  34357=>"000000000",
  34358=>"001000000",
  34359=>"000000100",
  34360=>"101001001",
  34361=>"110100100",
  34362=>"000111111",
  34363=>"111100111",
  34364=>"000000000",
  34365=>"111110100",
  34366=>"001000010",
  34367=>"111111000",
  34368=>"011000000",
  34369=>"000000000",
  34370=>"111111001",
  34371=>"111111111",
  34372=>"111001000",
  34373=>"001011011",
  34374=>"000000110",
  34375=>"000000000",
  34376=>"101111100",
  34377=>"111111111",
  34378=>"101110000",
  34379=>"110000000",
  34380=>"000000000",
  34381=>"111111111",
  34382=>"101000111",
  34383=>"000000000",
  34384=>"000000110",
  34385=>"000000000",
  34386=>"000000000",
  34387=>"111111011",
  34388=>"101111101",
  34389=>"000001111",
  34390=>"110000000",
  34391=>"111111100",
  34392=>"000000000",
  34393=>"100000111",
  34394=>"111001000",
  34395=>"110100101",
  34396=>"100110110",
  34397=>"111111111",
  34398=>"011111110",
  34399=>"001001001",
  34400=>"000000000",
  34401=>"000100110",
  34402=>"000101001",
  34403=>"100101000",
  34404=>"001001010",
  34405=>"000000001",
  34406=>"111111111",
  34407=>"011001111",
  34408=>"011111000",
  34409=>"111110000",
  34410=>"001000110",
  34411=>"000000000",
  34412=>"001000000",
  34413=>"001000000",
  34414=>"111111111",
  34415=>"001111111",
  34416=>"000000000",
  34417=>"111011000",
  34418=>"101001001",
  34419=>"000000011",
  34420=>"000000000",
  34421=>"011111111",
  34422=>"111000111",
  34423=>"111111110",
  34424=>"000111001",
  34425=>"000000000",
  34426=>"000000000",
  34427=>"101000000",
  34428=>"111110110",
  34429=>"011101000",
  34430=>"111111110",
  34431=>"000001000",
  34432=>"000000101",
  34433=>"000000110",
  34434=>"000000001",
  34435=>"100000111",
  34436=>"100000000",
  34437=>"100000111",
  34438=>"011010000",
  34439=>"000101111",
  34440=>"000111111",
  34441=>"111101110",
  34442=>"111111111",
  34443=>"001001001",
  34444=>"111111111",
  34445=>"111111000",
  34446=>"100000000",
  34447=>"011111000",
  34448=>"100100111",
  34449=>"000000001",
  34450=>"000100100",
  34451=>"000000000",
  34452=>"101001111",
  34453=>"110111111",
  34454=>"000000111",
  34455=>"100100100",
  34456=>"000000001",
  34457=>"100110111",
  34458=>"111000000",
  34459=>"111111011",
  34460=>"111000001",
  34461=>"100000000",
  34462=>"111111000",
  34463=>"000000000",
  34464=>"000100000",
  34465=>"000000110",
  34466=>"111111000",
  34467=>"111111111",
  34468=>"000111001",
  34469=>"110111111",
  34470=>"111111101",
  34471=>"000100000",
  34472=>"000000000",
  34473=>"100000000",
  34474=>"001001101",
  34475=>"100100111",
  34476=>"000111111",
  34477=>"100110111",
  34478=>"111100100",
  34479=>"001101110",
  34480=>"111110111",
  34481=>"001111111",
  34482=>"110111110",
  34483=>"000111000",
  34484=>"000010011",
  34485=>"111100100",
  34486=>"111101000",
  34487=>"111111111",
  34488=>"100100111",
  34489=>"100100111",
  34490=>"000000000",
  34491=>"100101001",
  34492=>"001001000",
  34493=>"101001101",
  34494=>"111111111",
  34495=>"000001000",
  34496=>"000000000",
  34497=>"111011010",
  34498=>"000111111",
  34499=>"111111111",
  34500=>"111111110",
  34501=>"000000110",
  34502=>"000000000",
  34503=>"100100000",
  34504=>"011011111",
  34505=>"000100000",
  34506=>"111111100",
  34507=>"000001000",
  34508=>"100100110",
  34509=>"100111111",
  34510=>"100000100",
  34511=>"010011111",
  34512=>"000000111",
  34513=>"000011111",
  34514=>"111101100",
  34515=>"111111001",
  34516=>"111111111",
  34517=>"100110000",
  34518=>"110000000",
  34519=>"111111111",
  34520=>"000000000",
  34521=>"111110110",
  34522=>"111000000",
  34523=>"100101111",
  34524=>"101111011",
  34525=>"000000000",
  34526=>"000000110",
  34527=>"000000100",
  34528=>"000000000",
  34529=>"000011011",
  34530=>"000110000",
  34531=>"111101100",
  34532=>"111111111",
  34533=>"000110000",
  34534=>"000000101",
  34535=>"111111111",
  34536=>"000000011",
  34537=>"111111111",
  34538=>"001000100",
  34539=>"110100000",
  34540=>"001001000",
  34541=>"001001111",
  34542=>"100000000",
  34543=>"000000000",
  34544=>"000000000",
  34545=>"000000000",
  34546=>"111110000",
  34547=>"000000000",
  34548=>"111111110",
  34549=>"111110111",
  34550=>"110111100",
  34551=>"110110111",
  34552=>"000000111",
  34553=>"100111111",
  34554=>"101101111",
  34555=>"111000000",
  34556=>"010011010",
  34557=>"000000001",
  34558=>"111110100",
  34559=>"111000000",
  34560=>"000000111",
  34561=>"100100100",
  34562=>"000000001",
  34563=>"001111000",
  34564=>"000000000",
  34565=>"000100000",
  34566=>"101100111",
  34567=>"011001111",
  34568=>"111100100",
  34569=>"000000000",
  34570=>"000000111",
  34571=>"111111111",
  34572=>"000000000",
  34573=>"000000101",
  34574=>"010111111",
  34575=>"010000111",
  34576=>"110100000",
  34577=>"001001111",
  34578=>"001001111",
  34579=>"100111111",
  34580=>"011111110",
  34581=>"011011011",
  34582=>"111111100",
  34583=>"000101100",
  34584=>"110111111",
  34585=>"011100011",
  34586=>"011011000",
  34587=>"111000000",
  34588=>"110110110",
  34589=>"011001000",
  34590=>"000000000",
  34591=>"000100101",
  34592=>"111111100",
  34593=>"100100000",
  34594=>"110100000",
  34595=>"101111111",
  34596=>"111111011",
  34597=>"000000101",
  34598=>"111111010",
  34599=>"001001011",
  34600=>"000111101",
  34601=>"000000000",
  34602=>"110100100",
  34603=>"000000100",
  34604=>"001011111",
  34605=>"000000000",
  34606=>"111110000",
  34607=>"111101110",
  34608=>"001001001",
  34609=>"010011111",
  34610=>"111111111",
  34611=>"110111111",
  34612=>"110100110",
  34613=>"000000000",
  34614=>"011111100",
  34615=>"111111100",
  34616=>"000000000",
  34617=>"111100111",
  34618=>"100001001",
  34619=>"111010110",
  34620=>"000000101",
  34621=>"001000000",
  34622=>"000000011",
  34623=>"000000101",
  34624=>"101100000",
  34625=>"111111000",
  34626=>"110111010",
  34627=>"000000000",
  34628=>"100001100",
  34629=>"111110000",
  34630=>"010011001",
  34631=>"001001001",
  34632=>"000000000",
  34633=>"000111111",
  34634=>"111111011",
  34635=>"000110000",
  34636=>"000000101",
  34637=>"111111000",
  34638=>"100000000",
  34639=>"000110110",
  34640=>"001111111",
  34641=>"110011111",
  34642=>"111111111",
  34643=>"111111111",
  34644=>"000001001",
  34645=>"011011011",
  34646=>"111111111",
  34647=>"111101110",
  34648=>"101000000",
  34649=>"110111000",
  34650=>"100101010",
  34651=>"000000000",
  34652=>"111100100",
  34653=>"000001010",
  34654=>"111011010",
  34655=>"000000100",
  34656=>"000000001",
  34657=>"101001000",
  34658=>"100100100",
  34659=>"100100111",
  34660=>"101111001",
  34661=>"111111101",
  34662=>"001001111",
  34663=>"100000101",
  34664=>"100100100",
  34665=>"101000100",
  34666=>"000000000",
  34667=>"111011000",
  34668=>"101001101",
  34669=>"000000000",
  34670=>"000001000",
  34671=>"111111111",
  34672=>"111111111",
  34673=>"111111111",
  34674=>"100000000",
  34675=>"000011000",
  34676=>"011111011",
  34677=>"001000000",
  34678=>"010000110",
  34679=>"011111000",
  34680=>"111101001",
  34681=>"111111011",
  34682=>"000000000",
  34683=>"110111110",
  34684=>"000011010",
  34685=>"100100100",
  34686=>"000111000",
  34687=>"000001111",
  34688=>"100000100",
  34689=>"100000000",
  34690=>"000001011",
  34691=>"111000000",
  34692=>"001011111",
  34693=>"000000000",
  34694=>"111111011",
  34695=>"100000000",
  34696=>"001000111",
  34697=>"000111001",
  34698=>"100000101",
  34699=>"110100000",
  34700=>"000001101",
  34701=>"110111100",
  34702=>"100100111",
  34703=>"000000000",
  34704=>"000001001",
  34705=>"001000111",
  34706=>"001001011",
  34707=>"000000000",
  34708=>"111000000",
  34709=>"000001011",
  34710=>"111111111",
  34711=>"001101001",
  34712=>"111111111",
  34713=>"000100111",
  34714=>"101100101",
  34715=>"000000100",
  34716=>"111001001",
  34717=>"100000000",
  34718=>"111000000",
  34719=>"111111111",
  34720=>"011010111",
  34721=>"000101101",
  34722=>"100000000",
  34723=>"001001001",
  34724=>"001000000",
  34725=>"001001000",
  34726=>"000000000",
  34727=>"100001000",
  34728=>"000000000",
  34729=>"111111010",
  34730=>"111101101",
  34731=>"001000000",
  34732=>"011001011",
  34733=>"111100101",
  34734=>"010011111",
  34735=>"111111100",
  34736=>"111111111",
  34737=>"000000000",
  34738=>"000000001",
  34739=>"001001111",
  34740=>"100110000",
  34741=>"000000000",
  34742=>"100000000",
  34743=>"000111111",
  34744=>"000000010",
  34745=>"000000000",
  34746=>"011011011",
  34747=>"000000000",
  34748=>"000000100",
  34749=>"111111111",
  34750=>"100100000",
  34751=>"100101101",
  34752=>"111111000",
  34753=>"111110000",
  34754=>"111111111",
  34755=>"000001001",
  34756=>"111100111",
  34757=>"110110110",
  34758=>"100100101",
  34759=>"000000100",
  34760=>"100000000",
  34761=>"100110000",
  34762=>"101001011",
  34763=>"000000000",
  34764=>"101000000",
  34765=>"100100000",
  34766=>"110100100",
  34767=>"111111111",
  34768=>"100111110",
  34769=>"010111010",
  34770=>"001001101",
  34771=>"000001001",
  34772=>"000001011",
  34773=>"111111111",
  34774=>"110111011",
  34775=>"000000000",
  34776=>"100100111",
  34777=>"100101000",
  34778=>"111011000",
  34779=>"001001111",
  34780=>"011111101",
  34781=>"000000000",
  34782=>"111111000",
  34783=>"110100101",
  34784=>"111111000",
  34785=>"000100000",
  34786=>"110111110",
  34787=>"001001111",
  34788=>"111111111",
  34789=>"011111111",
  34790=>"000000111",
  34791=>"111011011",
  34792=>"111111111",
  34793=>"001001000",
  34794=>"000000000",
  34795=>"111111001",
  34796=>"011101000",
  34797=>"000000000",
  34798=>"000000010",
  34799=>"000000111",
  34800=>"000000000",
  34801=>"010111111",
  34802=>"011101000",
  34803=>"100000000",
  34804=>"001000100",
  34805=>"011001011",
  34806=>"011111000",
  34807=>"100100110",
  34808=>"000111111",
  34809=>"000000000",
  34810=>"111001001",
  34811=>"100100111",
  34812=>"101001111",
  34813=>"000000111",
  34814=>"100100100",
  34815=>"111101111",
  34816=>"000001111",
  34817=>"011000011",
  34818=>"111101111",
  34819=>"111111110",
  34820=>"101111111",
  34821=>"000000111",
  34822=>"000000000",
  34823=>"111111111",
  34824=>"011000000",
  34825=>"111000000",
  34826=>"000100000",
  34827=>"100100001",
  34828=>"100100000",
  34829=>"111111111",
  34830=>"100110111",
  34831=>"000000000",
  34832=>"111001000",
  34833=>"111111000",
  34834=>"000001111",
  34835=>"000000101",
  34836=>"111111000",
  34837=>"000000000",
  34838=>"110000001",
  34839=>"111100100",
  34840=>"001000000",
  34841=>"100111111",
  34842=>"111001011",
  34843=>"111000100",
  34844=>"000000000",
  34845=>"101100101",
  34846=>"000011101",
  34847=>"111111010",
  34848=>"000000000",
  34849=>"111111000",
  34850=>"000000001",
  34851=>"111000100",
  34852=>"000000000",
  34853=>"111000000",
  34854=>"110100000",
  34855=>"000000000",
  34856=>"000100101",
  34857=>"000000000",
  34858=>"100000100",
  34859=>"100100010",
  34860=>"111011011",
  34861=>"000011111",
  34862=>"111011101",
  34863=>"000000000",
  34864=>"000000000",
  34865=>"111011000",
  34866=>"011000000",
  34867=>"110111011",
  34868=>"101101000",
  34869=>"111101000",
  34870=>"100100100",
  34871=>"111110100",
  34872=>"000000011",
  34873=>"000111011",
  34874=>"000000101",
  34875=>"111111111",
  34876=>"011001000",
  34877=>"000000000",
  34878=>"000110111",
  34879=>"000000000",
  34880=>"100011111",
  34881=>"000110100",
  34882=>"000011001",
  34883=>"111111011",
  34884=>"000001001",
  34885=>"111110100",
  34886=>"000111111",
  34887=>"111111100",
  34888=>"001011000",
  34889=>"000000111",
  34890=>"111111000",
  34891=>"000001000",
  34892=>"100000000",
  34893=>"110000000",
  34894=>"111101111",
  34895=>"011111111",
  34896=>"100000000",
  34897=>"000000111",
  34898=>"000000000",
  34899=>"111111111",
  34900=>"000000101",
  34901=>"111110000",
  34902=>"100101100",
  34903=>"111111000",
  34904=>"111111111",
  34905=>"001001101",
  34906=>"000000001",
  34907=>"110010011",
  34908=>"011010010",
  34909=>"011000000",
  34910=>"001111111",
  34911=>"111111111",
  34912=>"000111111",
  34913=>"000000000",
  34914=>"000000100",
  34915=>"111111111",
  34916=>"111011111",
  34917=>"000000000",
  34918=>"001000000",
  34919=>"000110100",
  34920=>"110111111",
  34921=>"111011111",
  34922=>"000000001",
  34923=>"000000000",
  34924=>"010111111",
  34925=>"110111111",
  34926=>"111101101",
  34927=>"111111111",
  34928=>"001000000",
  34929=>"100100100",
  34930=>"011011111",
  34931=>"000011111",
  34932=>"000000000",
  34933=>"000000110",
  34934=>"000000000",
  34935=>"111000000",
  34936=>"010111111",
  34937=>"000000000",
  34938=>"000000010",
  34939=>"000000000",
  34940=>"110111110",
  34941=>"111110000",
  34942=>"000100100",
  34943=>"111000000",
  34944=>"111111110",
  34945=>"000000000",
  34946=>"011111000",
  34947=>"001000000",
  34948=>"000011111",
  34949=>"000000000",
  34950=>"001011111",
  34951=>"000000000",
  34952=>"111111111",
  34953=>"111111111",
  34954=>"000000000",
  34955=>"000000011",
  34956=>"000111101",
  34957=>"000000001",
  34958=>"000111100",
  34959=>"000000000",
  34960=>"000000101",
  34961=>"111111111",
  34962=>"111110000",
  34963=>"000000100",
  34964=>"000110111",
  34965=>"111111101",
  34966=>"001111111",
  34967=>"101001111",
  34968=>"000100101",
  34969=>"000000111",
  34970=>"111001101",
  34971=>"000000111",
  34972=>"111110000",
  34973=>"100000000",
  34974=>"100101111",
  34975=>"111000000",
  34976=>"100000100",
  34977=>"000111111",
  34978=>"000000000",
  34979=>"000000000",
  34980=>"111000100",
  34981=>"000000111",
  34982=>"011010000",
  34983=>"111111000",
  34984=>"000011011",
  34985=>"000000101",
  34986=>"011000100",
  34987=>"001001001",
  34988=>"011111111",
  34989=>"001111111",
  34990=>"000001000",
  34991=>"011001111",
  34992=>"000000000",
  34993=>"001000000",
  34994=>"110110111",
  34995=>"000100100",
  34996=>"111111111",
  34997=>"000000000",
  34998=>"000000000",
  34999=>"000000000",
  35000=>"001111101",
  35001=>"000111111",
  35002=>"001001101",
  35003=>"010111101",
  35004=>"110000000",
  35005=>"000000010",
  35006=>"000000110",
  35007=>"000000000",
  35008=>"111111111",
  35009=>"000000000",
  35010=>"000100000",
  35011=>"000000000",
  35012=>"110010111",
  35013=>"000000001",
  35014=>"000111001",
  35015=>"111111001",
  35016=>"011011011",
  35017=>"111111111",
  35018=>"111000000",
  35019=>"111111110",
  35020=>"000100100",
  35021=>"001111111",
  35022=>"111000000",
  35023=>"000000001",
  35024=>"011000000",
  35025=>"010000001",
  35026=>"111111111",
  35027=>"111100110",
  35028=>"000000000",
  35029=>"111111111",
  35030=>"111110000",
  35031=>"001111111",
  35032=>"000000110",
  35033=>"101111000",
  35034=>"000000000",
  35035=>"100110110",
  35036=>"111111111",
  35037=>"110000000",
  35038=>"111000111",
  35039=>"000100111",
  35040=>"000111111",
  35041=>"000011011",
  35042=>"111001001",
  35043=>"000111001",
  35044=>"111111000",
  35045=>"111111110",
  35046=>"111111000",
  35047=>"110111100",
  35048=>"101111111",
  35049=>"100001000",
  35050=>"111111111",
  35051=>"101011000",
  35052=>"110110111",
  35053=>"111000000",
  35054=>"111000111",
  35055=>"011000111",
  35056=>"000101111",
  35057=>"001000100",
  35058=>"000000111",
  35059=>"100100111",
  35060=>"000000000",
  35061=>"111111111",
  35062=>"111111010",
  35063=>"000000110",
  35064=>"000000001",
  35065=>"110100000",
  35066=>"000000000",
  35067=>"111000000",
  35068=>"111100100",
  35069=>"110001001",
  35070=>"010000000",
  35071=>"001111110",
  35072=>"000100000",
  35073=>"001001000",
  35074=>"000000000",
  35075=>"000000000",
  35076=>"001111111",
  35077=>"001000000",
  35078=>"000000111",
  35079=>"000101111",
  35080=>"111100100",
  35081=>"000000000",
  35082=>"010111111",
  35083=>"000111111",
  35084=>"111110000",
  35085=>"000100111",
  35086=>"111111111",
  35087=>"000101111",
  35088=>"100000000",
  35089=>"111101111",
  35090=>"011001111",
  35091=>"000111111",
  35092=>"000000111",
  35093=>"000000000",
  35094=>"111100000",
  35095=>"000000111",
  35096=>"111101111",
  35097=>"000010000",
  35098=>"101000000",
  35099=>"111010000",
  35100=>"110100000",
  35101=>"111111000",
  35102=>"110000000",
  35103=>"000000101",
  35104=>"111100111",
  35105=>"000000000",
  35106=>"100000000",
  35107=>"110111111",
  35108=>"111000000",
  35109=>"111111110",
  35110=>"000000000",
  35111=>"100110111",
  35112=>"110111111",
  35113=>"111000000",
  35114=>"000100000",
  35115=>"000000000",
  35116=>"000111100",
  35117=>"100011011",
  35118=>"000000111",
  35119=>"000111111",
  35120=>"011011111",
  35121=>"111100100",
  35122=>"111111111",
  35123=>"111011000",
  35124=>"111100000",
  35125=>"111101100",
  35126=>"111100101",
  35127=>"000000000",
  35128=>"000000000",
  35129=>"111101101",
  35130=>"111010001",
  35131=>"111110100",
  35132=>"111101000",
  35133=>"100000000",
  35134=>"111001000",
  35135=>"001000000",
  35136=>"000000000",
  35137=>"000000000",
  35138=>"111111001",
  35139=>"000001111",
  35140=>"001011111",
  35141=>"111111111",
  35142=>"111111010",
  35143=>"001111111",
  35144=>"111110010",
  35145=>"111000000",
  35146=>"001011001",
  35147=>"010111111",
  35148=>"111110111",
  35149=>"101011111",
  35150=>"111100111",
  35151=>"100100000",
  35152=>"111111110",
  35153=>"000000100",
  35154=>"111111111",
  35155=>"111111110",
  35156=>"000000110",
  35157=>"001011001",
  35158=>"110000001",
  35159=>"111000000",
  35160=>"000000111",
  35161=>"000000000",
  35162=>"001000110",
  35163=>"000100101",
  35164=>"000000000",
  35165=>"011000111",
  35166=>"110001000",
  35167=>"000111100",
  35168=>"000000110",
  35169=>"111111011",
  35170=>"000111101",
  35171=>"011000001",
  35172=>"111001000",
  35173=>"111100100",
  35174=>"001000000",
  35175=>"101001001",
  35176=>"010010111",
  35177=>"000000000",
  35178=>"000000000",
  35179=>"000111111",
  35180=>"010011111",
  35181=>"111000000",
  35182=>"000000000",
  35183=>"111110001",
  35184=>"000100110",
  35185=>"011011000",
  35186=>"111000000",
  35187=>"011000001",
  35188=>"011000000",
  35189=>"001000000",
  35190=>"011111000",
  35191=>"011011110",
  35192=>"111011000",
  35193=>"111010000",
  35194=>"001000100",
  35195=>"010110100",
  35196=>"000000100",
  35197=>"011001000",
  35198=>"111111111",
  35199=>"010000100",
  35200=>"110111111",
  35201=>"000111111",
  35202=>"111111000",
  35203=>"000000111",
  35204=>"111110111",
  35205=>"111111111",
  35206=>"001111000",
  35207=>"011111111",
  35208=>"101001000",
  35209=>"000001000",
  35210=>"000000000",
  35211=>"011011011",
  35212=>"000111111",
  35213=>"110111000",
  35214=>"110111111",
  35215=>"000000000",
  35216=>"111010000",
  35217=>"100000011",
  35218=>"000100101",
  35219=>"111111000",
  35220=>"111100111",
  35221=>"000000000",
  35222=>"000000111",
  35223=>"001011011",
  35224=>"100110110",
  35225=>"000010111",
  35226=>"111000000",
  35227=>"100101111",
  35228=>"000111000",
  35229=>"000000000",
  35230=>"011001011",
  35231=>"111111000",
  35232=>"000000010",
  35233=>"111010100",
  35234=>"000010001",
  35235=>"111000000",
  35236=>"000000000",
  35237=>"000111111",
  35238=>"000000000",
  35239=>"111111111",
  35240=>"011111111",
  35241=>"111101111",
  35242=>"111111111",
  35243=>"100001100",
  35244=>"000000000",
  35245=>"000000111",
  35246=>"000111110",
  35247=>"000000001",
  35248=>"110111000",
  35249=>"000000000",
  35250=>"111000001",
  35251=>"111100100",
  35252=>"111000000",
  35253=>"111111111",
  35254=>"001001111",
  35255=>"111111111",
  35256=>"000000000",
  35257=>"010000000",
  35258=>"111111010",
  35259=>"101101011",
  35260=>"000000000",
  35261=>"011111111",
  35262=>"000000111",
  35263=>"111101001",
  35264=>"111111111",
  35265=>"111001000",
  35266=>"111111111",
  35267=>"000000000",
  35268=>"001111111",
  35269=>"000000000",
  35270=>"001000001",
  35271=>"111111001",
  35272=>"101111111",
  35273=>"010000000",
  35274=>"110100000",
  35275=>"111111111",
  35276=>"000000000",
  35277=>"111111111",
  35278=>"110111111",
  35279=>"000000000",
  35280=>"011000000",
  35281=>"000001111",
  35282=>"111111100",
  35283=>"111111111",
  35284=>"110110000",
  35285=>"110100101",
  35286=>"000000111",
  35287=>"001111100",
  35288=>"110000000",
  35289=>"000000000",
  35290=>"000000000",
  35291=>"110100000",
  35292=>"000000111",
  35293=>"110111111",
  35294=>"000000111",
  35295=>"000000000",
  35296=>"101000000",
  35297=>"111011110",
  35298=>"001111111",
  35299=>"000010111",
  35300=>"011011111",
  35301=>"000000100",
  35302=>"111111111",
  35303=>"111111111",
  35304=>"000100000",
  35305=>"111111111",
  35306=>"000000111",
  35307=>"100000111",
  35308=>"001001101",
  35309=>"110110111",
  35310=>"000001000",
  35311=>"010111111",
  35312=>"000000000",
  35313=>"000000000",
  35314=>"011101000",
  35315=>"010010011",
  35316=>"110000000",
  35317=>"000000111",
  35318=>"001000000",
  35319=>"101001001",
  35320=>"000000000",
  35321=>"110100000",
  35322=>"110000000",
  35323=>"000000000",
  35324=>"000100000",
  35325=>"011011011",
  35326=>"000100100",
  35327=>"000000111",
  35328=>"001000111",
  35329=>"000000000",
  35330=>"111001000",
  35331=>"000000111",
  35332=>"000000100",
  35333=>"001000110",
  35334=>"111111111",
  35335=>"101111111",
  35336=>"000000000",
  35337=>"110110111",
  35338=>"000000011",
  35339=>"111111100",
  35340=>"001101111",
  35341=>"110111111",
  35342=>"110110000",
  35343=>"000000001",
  35344=>"101100101",
  35345=>"001000111",
  35346=>"000000000",
  35347=>"111001101",
  35348=>"111100111",
  35349=>"111111111",
  35350=>"111111011",
  35351=>"100101100",
  35352=>"111001111",
  35353=>"111111011",
  35354=>"000000100",
  35355=>"100000000",
  35356=>"000000001",
  35357=>"100100000",
  35358=>"110110010",
  35359=>"111111111",
  35360=>"111111111",
  35361=>"110110000",
  35362=>"101001001",
  35363=>"110111111",
  35364=>"111000000",
  35365=>"111110111",
  35366=>"111111011",
  35367=>"111101010",
  35368=>"000001111",
  35369=>"111111000",
  35370=>"000000010",
  35371=>"110111001",
  35372=>"100100111",
  35373=>"000000000",
  35374=>"000000000",
  35375=>"111111111",
  35376=>"111011010",
  35377=>"000000000",
  35378=>"100000000",
  35379=>"000000011",
  35380=>"000000000",
  35381=>"111111000",
  35382=>"101000000",
  35383=>"110111011",
  35384=>"000001011",
  35385=>"111010101",
  35386=>"000000111",
  35387=>"000001000",
  35388=>"111101111",
  35389=>"111111000",
  35390=>"111111111",
  35391=>"000000000",
  35392=>"000000001",
  35393=>"001000001",
  35394=>"111000101",
  35395=>"100100111",
  35396=>"101001111",
  35397=>"010010000",
  35398=>"000000111",
  35399=>"111111111",
  35400=>"011111101",
  35401=>"111101000",
  35402=>"111011110",
  35403=>"000010010",
  35404=>"000001111",
  35405=>"111111000",
  35406=>"011000000",
  35407=>"110000110",
  35408=>"111111111",
  35409=>"101000000",
  35410=>"100000110",
  35411=>"001110110",
  35412=>"111101000",
  35413=>"111111011",
  35414=>"000000000",
  35415=>"001000000",
  35416=>"101101111",
  35417=>"111100000",
  35418=>"000000111",
  35419=>"111100100",
  35420=>"011011111",
  35421=>"000000000",
  35422=>"001000000",
  35423=>"000001000",
  35424=>"111000000",
  35425=>"111000000",
  35426=>"010010000",
  35427=>"000001001",
  35428=>"101101111",
  35429=>"011010000",
  35430=>"000000100",
  35431=>"000000000",
  35432=>"111001000",
  35433=>"111000000",
  35434=>"111000001",
  35435=>"000000111",
  35436=>"111111110",
  35437=>"000000000",
  35438=>"100100111",
  35439=>"111111111",
  35440=>"001001010",
  35441=>"110111111",
  35442=>"010010000",
  35443=>"110010001",
  35444=>"011000010",
  35445=>"000000101",
  35446=>"000000000",
  35447=>"000101101",
  35448=>"000000000",
  35449=>"011111011",
  35450=>"000000000",
  35451=>"000000000",
  35452=>"100110110",
  35453=>"011111111",
  35454=>"000000000",
  35455=>"000001000",
  35456=>"100111111",
  35457=>"101011110",
  35458=>"010000001",
  35459=>"111000001",
  35460=>"000000000",
  35461=>"101000100",
  35462=>"111111000",
  35463=>"111111111",
  35464=>"110111111",
  35465=>"001000111",
  35466=>"110000000",
  35467=>"000000000",
  35468=>"000000111",
  35469=>"111111110",
  35470=>"110110110",
  35471=>"000000000",
  35472=>"000110110",
  35473=>"011000001",
  35474=>"000000000",
  35475=>"110110111",
  35476=>"111100111",
  35477=>"101100100",
  35478=>"000110111",
  35479=>"000000111",
  35480=>"001000000",
  35481=>"111111000",
  35482=>"100111111",
  35483=>"000000111",
  35484=>"111100100",
  35485=>"111011101",
  35486=>"111111001",
  35487=>"000000111",
  35488=>"100000000",
  35489=>"100111111",
  35490=>"100111111",
  35491=>"000000000",
  35492=>"000001001",
  35493=>"101100111",
  35494=>"000000111",
  35495=>"010010110",
  35496=>"000000011",
  35497=>"011011011",
  35498=>"000000000",
  35499=>"111001101",
  35500=>"000000011",
  35501=>"000001000",
  35502=>"000000000",
  35503=>"111111111",
  35504=>"110111111",
  35505=>"111111111",
  35506=>"111111111",
  35507=>"110111111",
  35508=>"111111111",
  35509=>"000010000",
  35510=>"111111011",
  35511=>"111110100",
  35512=>"000000000",
  35513=>"000111111",
  35514=>"000000011",
  35515=>"111000000",
  35516=>"111000000",
  35517=>"110111100",
  35518=>"100000000",
  35519=>"000110111",
  35520=>"100100100",
  35521=>"000000000",
  35522=>"100000000",
  35523=>"111110000",
  35524=>"111111111",
  35525=>"000000001",
  35526=>"011011111",
  35527=>"111111111",
  35528=>"000010111",
  35529=>"111111000",
  35530=>"000000111",
  35531=>"000001000",
  35532=>"100100000",
  35533=>"100111111",
  35534=>"111101101",
  35535=>"011011001",
  35536=>"001011011",
  35537=>"000000000",
  35538=>"001000000",
  35539=>"000000011",
  35540=>"000100100",
  35541=>"111111111",
  35542=>"000000000",
  35543=>"000111111",
  35544=>"010110000",
  35545=>"001100000",
  35546=>"111111111",
  35547=>"101101100",
  35548=>"111111111",
  35549=>"111111000",
  35550=>"000000000",
  35551=>"001000000",
  35552=>"000000111",
  35553=>"111111010",
  35554=>"000000111",
  35555=>"100000000",
  35556=>"000000000",
  35557=>"100100000",
  35558=>"111100000",
  35559=>"100000110",
  35560=>"111111000",
  35561=>"000000000",
  35562=>"111000001",
  35563=>"001000001",
  35564=>"111011111",
  35565=>"000000000",
  35566=>"000001111",
  35567=>"011011001",
  35568=>"111100101",
  35569=>"011111011",
  35570=>"000111111",
  35571=>"000111111",
  35572=>"010111111",
  35573=>"000000000",
  35574=>"100001001",
  35575=>"000100111",
  35576=>"000000000",
  35577=>"001000000",
  35578=>"111111001",
  35579=>"111111111",
  35580=>"100100001",
  35581=>"101111111",
  35582=>"110001111",
  35583=>"101100100",
  35584=>"111111111",
  35585=>"001101111",
  35586=>"111011011",
  35587=>"110111111",
  35588=>"110100100",
  35589=>"000000111",
  35590=>"000000000",
  35591=>"000000011",
  35592=>"111110000",
  35593=>"000000111",
  35594=>"100000000",
  35595=>"000000000",
  35596=>"001001001",
  35597=>"000000000",
  35598=>"100111100",
  35599=>"100111101",
  35600=>"000100110",
  35601=>"000000111",
  35602=>"100100101",
  35603=>"000000001",
  35604=>"111111111",
  35605=>"000000000",
  35606=>"000110111",
  35607=>"011000011",
  35608=>"000000000",
  35609=>"111001000",
  35610=>"111100101",
  35611=>"111111111",
  35612=>"000000100",
  35613=>"110000000",
  35614=>"000000000",
  35615=>"000110110",
  35616=>"000000000",
  35617=>"000000110",
  35618=>"001011000",
  35619=>"000000000",
  35620=>"100110110",
  35621=>"111111111",
  35622=>"011111111",
  35623=>"000010010",
  35624=>"000000000",
  35625=>"111111000",
  35626=>"000000000",
  35627=>"000000000",
  35628=>"111011110",
  35629=>"000000011",
  35630=>"111000111",
  35631=>"111000000",
  35632=>"111000100",
  35633=>"110100000",
  35634=>"011111000",
  35635=>"000010000",
  35636=>"001001000",
  35637=>"011011011",
  35638=>"000000000",
  35639=>"000111111",
  35640=>"000000000",
  35641=>"000000000",
  35642=>"000000000",
  35643=>"101111111",
  35644=>"110001001",
  35645=>"111111111",
  35646=>"000000000",
  35647=>"111001000",
  35648=>"011101000",
  35649=>"111111011",
  35650=>"111111111",
  35651=>"000000000",
  35652=>"011000000",
  35653=>"010000111",
  35654=>"111111000",
  35655=>"001000101",
  35656=>"000000000",
  35657=>"011000000",
  35658=>"001000000",
  35659=>"011111111",
  35660=>"010011011",
  35661=>"100000000",
  35662=>"101000000",
  35663=>"111111011",
  35664=>"001001001",
  35665=>"000000111",
  35666=>"111011000",
  35667=>"000000100",
  35668=>"111111100",
  35669=>"011011000",
  35670=>"111111111",
  35671=>"000000000",
  35672=>"000000000",
  35673=>"111111000",
  35674=>"111101011",
  35675=>"111111000",
  35676=>"111101101",
  35677=>"111100111",
  35678=>"010000100",
  35679=>"011110100",
  35680=>"001111000",
  35681=>"011000000",
  35682=>"000000000",
  35683=>"101111111",
  35684=>"000011111",
  35685=>"000000000",
  35686=>"001111111",
  35687=>"000000000",
  35688=>"111110100",
  35689=>"110111011",
  35690=>"000000000",
  35691=>"111111000",
  35692=>"001000000",
  35693=>"000100111",
  35694=>"000001111",
  35695=>"000000000",
  35696=>"000000000",
  35697=>"010010000",
  35698=>"111111011",
  35699=>"000110110",
  35700=>"111011000",
  35701=>"000100011",
  35702=>"100000010",
  35703=>"010111111",
  35704=>"000000000",
  35705=>"011000000",
  35706=>"001111111",
  35707=>"110110110",
  35708=>"110110010",
  35709=>"001000000",
  35710=>"000000000",
  35711=>"111101111",
  35712=>"111111111",
  35713=>"000000000",
  35714=>"011110110",
  35715=>"001000000",
  35716=>"111000110",
  35717=>"111011111",
  35718=>"011011011",
  35719=>"111111111",
  35720=>"111111111",
  35721=>"010000100",
  35722=>"000000000",
  35723=>"000010000",
  35724=>"101000001",
  35725=>"100111011",
  35726=>"111111000",
  35727=>"001000011",
  35728=>"000000000",
  35729=>"111001000",
  35730=>"000000000",
  35731=>"001000100",
  35732=>"110111011",
  35733=>"000000000",
  35734=>"100100100",
  35735=>"011011001",
  35736=>"000000000",
  35737=>"111111111",
  35738=>"000000000",
  35739=>"000000000",
  35740=>"000000000",
  35741=>"000000011",
  35742=>"001000000",
  35743=>"111110110",
  35744=>"111110000",
  35745=>"000000001",
  35746=>"111111111",
  35747=>"100100000",
  35748=>"100000000",
  35749=>"000000000",
  35750=>"001000001",
  35751=>"111111101",
  35752=>"000000001",
  35753=>"011000000",
  35754=>"111001111",
  35755=>"001110111",
  35756=>"001001000",
  35757=>"111000000",
  35758=>"010010010",
  35759=>"111001000",
  35760=>"000000111",
  35761=>"001001111",
  35762=>"000001001",
  35763=>"000000000",
  35764=>"000100110",
  35765=>"111111111",
  35766=>"000000111",
  35767=>"111111001",
  35768=>"111001111",
  35769=>"101111010",
  35770=>"111000000",
  35771=>"011001011",
  35772=>"000000000",
  35773=>"111111010",
  35774=>"000000000",
  35775=>"000000000",
  35776=>"110110110",
  35777=>"111111111",
  35778=>"000001000",
  35779=>"000011011",
  35780=>"000011111",
  35781=>"010011100",
  35782=>"111111110",
  35783=>"000100100",
  35784=>"000111111",
  35785=>"000000000",
  35786=>"111110000",
  35787=>"111000111",
  35788=>"000000000",
  35789=>"100100100",
  35790=>"010010110",
  35791=>"001111111",
  35792=>"000011000",
  35793=>"001001111",
  35794=>"000000100",
  35795=>"000000111",
  35796=>"111111011",
  35797=>"111111111",
  35798=>"000001111",
  35799=>"111111100",
  35800=>"100100111",
  35801=>"000000000",
  35802=>"000000000",
  35803=>"000000000",
  35804=>"000000010",
  35805=>"100000000",
  35806=>"111000100",
  35807=>"000000000",
  35808=>"101110100",
  35809=>"000000011",
  35810=>"000111110",
  35811=>"111111111",
  35812=>"111111011",
  35813=>"101000000",
  35814=>"111011111",
  35815=>"111000000",
  35816=>"111111111",
  35817=>"111111111",
  35818=>"000000000",
  35819=>"100111111",
  35820=>"111110100",
  35821=>"001101000",
  35822=>"000100100",
  35823=>"001111111",
  35824=>"000101111",
  35825=>"011111111",
  35826=>"101000000",
  35827=>"001111111",
  35828=>"111001111",
  35829=>"111111111",
  35830=>"110110111",
  35831=>"000010000",
  35832=>"011000010",
  35833=>"001001001",
  35834=>"001101000",
  35835=>"000100111",
  35836=>"101111001",
  35837=>"111111111",
  35838=>"011111111",
  35839=>"101000000",
  35840=>"111110000",
  35841=>"000000000",
  35842=>"000100101",
  35843=>"111111000",
  35844=>"111111100",
  35845=>"111111001",
  35846=>"101000001",
  35847=>"100000000",
  35848=>"111111100",
  35849=>"110000001",
  35850=>"001000001",
  35851=>"111111111",
  35852=>"000001011",
  35853=>"000100000",
  35854=>"000000000",
  35855=>"101000111",
  35856=>"001111111",
  35857=>"010110101",
  35858=>"011000000",
  35859=>"111111011",
  35860=>"111111000",
  35861=>"111000010",
  35862=>"111111111",
  35863=>"100101111",
  35864=>"010010111",
  35865=>"111111000",
  35866=>"001000001",
  35867=>"000000000",
  35868=>"000011111",
  35869=>"111111000",
  35870=>"000000000",
  35871=>"111111000",
  35872=>"100111111",
  35873=>"111011000",
  35874=>"000000111",
  35875=>"111111110",
  35876=>"000000000",
  35877=>"000000101",
  35878=>"111011111",
  35879=>"000001111",
  35880=>"111000110",
  35881=>"101000000",
  35882=>"111010000",
  35883=>"111011100",
  35884=>"111101000",
  35885=>"111111101",
  35886=>"000011000",
  35887=>"111110000",
  35888=>"000100000",
  35889=>"000001111",
  35890=>"000101111",
  35891=>"111111000",
  35892=>"000000111",
  35893=>"000110111",
  35894=>"000000000",
  35895=>"111000000",
  35896=>"111111111",
  35897=>"111110111",
  35898=>"001000000",
  35899=>"100000000",
  35900=>"000000110",
  35901=>"111111110",
  35902=>"000010001",
  35903=>"101111001",
  35904=>"000000110",
  35905=>"000000110",
  35906=>"110111110",
  35907=>"100000000",
  35908=>"100001111",
  35909=>"100100000",
  35910=>"111100110",
  35911=>"000111111",
  35912=>"000011011",
  35913=>"000000000",
  35914=>"111111110",
  35915=>"000000100",
  35916=>"111111111",
  35917=>"000000111",
  35918=>"000000000",
  35919=>"110110010",
  35920=>"001000001",
  35921=>"000000000",
  35922=>"111111010",
  35923=>"001111111",
  35924=>"001001101",
  35925=>"011000111",
  35926=>"111011111",
  35927=>"110111111",
  35928=>"111111111",
  35929=>"100111111",
  35930=>"000000000",
  35931=>"111111000",
  35932=>"000111111",
  35933=>"111101000",
  35934=>"110111000",
  35935=>"111111000",
  35936=>"111100111",
  35937=>"111001111",
  35938=>"111000000",
  35939=>"000000111",
  35940=>"001001000",
  35941=>"111111000",
  35942=>"111111000",
  35943=>"001001000",
  35944=>"001000101",
  35945=>"111111111",
  35946=>"000000111",
  35947=>"000000000",
  35948=>"000110110",
  35949=>"000000000",
  35950=>"111111101",
  35951=>"000000000",
  35952=>"000000000",
  35953=>"111111000",
  35954=>"101111111",
  35955=>"000000111",
  35956=>"000000111",
  35957=>"001111011",
  35958=>"001001111",
  35959=>"000111111",
  35960=>"111111111",
  35961=>"000000100",
  35962=>"000111111",
  35963=>"111000111",
  35964=>"110111110",
  35965=>"011111111",
  35966=>"111111111",
  35967=>"111111110",
  35968=>"000000010",
  35969=>"110010001",
  35970=>"111000001",
  35971=>"010111111",
  35972=>"111110110",
  35973=>"111000100",
  35974=>"110110111",
  35975=>"100111100",
  35976=>"010110111",
  35977=>"111111000",
  35978=>"111111111",
  35979=>"000000100",
  35980=>"111000000",
  35981=>"101000111",
  35982=>"001000100",
  35983=>"000000110",
  35984=>"111111111",
  35985=>"000000000",
  35986=>"000000000",
  35987=>"000010111",
  35988=>"100110000",
  35989=>"000000000",
  35990=>"101001111",
  35991=>"101100111",
  35992=>"000000111",
  35993=>"000000111",
  35994=>"111000000",
  35995=>"000011010",
  35996=>"001000000",
  35997=>"100111000",
  35998=>"111101000",
  35999=>"110111100",
  36000=>"100000000",
  36001=>"000000000",
  36002=>"111000010",
  36003=>"000000101",
  36004=>"100111111",
  36005=>"011000000",
  36006=>"111001111",
  36007=>"000111111",
  36008=>"011011111",
  36009=>"111111101",
  36010=>"111010000",
  36011=>"011000011",
  36012=>"111001000",
  36013=>"110000000",
  36014=>"111111111",
  36015=>"111111000",
  36016=>"111111001",
  36017=>"111110000",
  36018=>"111111011",
  36019=>"111111111",
  36020=>"110110110",
  36021=>"011000111",
  36022=>"000000001",
  36023=>"000000111",
  36024=>"000000011",
  36025=>"111111111",
  36026=>"000111101",
  36027=>"111101111",
  36028=>"111111001",
  36029=>"111111111",
  36030=>"110000000",
  36031=>"000000111",
  36032=>"101000000",
  36033=>"011011111",
  36034=>"000000101",
  36035=>"101110111",
  36036=>"111110111",
  36037=>"111001111",
  36038=>"011111000",
  36039=>"000101111",
  36040=>"111100100",
  36041=>"000000000",
  36042=>"000000001",
  36043=>"111111111",
  36044=>"000000111",
  36045=>"010111111",
  36046=>"000110111",
  36047=>"000100110",
  36048=>"110010000",
  36049=>"100001000",
  36050=>"000000000",
  36051=>"110110000",
  36052=>"011011011",
  36053=>"111111111",
  36054=>"111111111",
  36055=>"001001101",
  36056=>"000100111",
  36057=>"111111111",
  36058=>"111000100",
  36059=>"111111111",
  36060=>"100100101",
  36061=>"110010000",
  36062=>"011011000",
  36063=>"101000001",
  36064=>"000000000",
  36065=>"111111111",
  36066=>"000000010",
  36067=>"100100111",
  36068=>"000111111",
  36069=>"111111000",
  36070=>"111111111",
  36071=>"000000000",
  36072=>"111000111",
  36073=>"111111001",
  36074=>"100111111",
  36075=>"111111111",
  36076=>"010111111",
  36077=>"000001111",
  36078=>"111000000",
  36079=>"000000000",
  36080=>"011111011",
  36081=>"010000001",
  36082=>"000111111",
  36083=>"111111000",
  36084=>"111111000",
  36085=>"111111111",
  36086=>"000000111",
  36087=>"000000111",
  36088=>"110010000",
  36089=>"101001111",
  36090=>"111001111",
  36091=>"010000000",
  36092=>"111111100",
  36093=>"000000011",
  36094=>"111000100",
  36095=>"111000000",
  36096=>"000000000",
  36097=>"000000000",
  36098=>"000000111",
  36099=>"111001111",
  36100=>"111000000",
  36101=>"101000000",
  36102=>"100101000",
  36103=>"111111111",
  36104=>"100111110",
  36105=>"000000110",
  36106=>"111111001",
  36107=>"111111111",
  36108=>"000000111",
  36109=>"111111111",
  36110=>"111111010",
  36111=>"000000000",
  36112=>"111000000",
  36113=>"111111110",
  36114=>"001000111",
  36115=>"111001001",
  36116=>"000000000",
  36117=>"000000000",
  36118=>"111111011",
  36119=>"000000111",
  36120=>"100110111",
  36121=>"111111000",
  36122=>"000000000",
  36123=>"100000001",
  36124=>"001011011",
  36125=>"000100111",
  36126=>"111111111",
  36127=>"110101000",
  36128=>"001101110",
  36129=>"000000110",
  36130=>"110110111",
  36131=>"000000000",
  36132=>"111000000",
  36133=>"111010000",
  36134=>"010110110",
  36135=>"000000001",
  36136=>"111111000",
  36137=>"111111000",
  36138=>"111011011",
  36139=>"011001011",
  36140=>"000011111",
  36141=>"000000111",
  36142=>"111111111",
  36143=>"000001001",
  36144=>"001001111",
  36145=>"011011011",
  36146=>"111110110",
  36147=>"111111010",
  36148=>"000000000",
  36149=>"011000000",
  36150=>"111100001",
  36151=>"101000111",
  36152=>"000000100",
  36153=>"000000100",
  36154=>"101000001",
  36155=>"000011111",
  36156=>"000000000",
  36157=>"000000111",
  36158=>"001011111",
  36159=>"011001000",
  36160=>"111100100",
  36161=>"111110000",
  36162=>"111011011",
  36163=>"000011011",
  36164=>"000000000",
  36165=>"100111000",
  36166=>"110111111",
  36167=>"000000111",
  36168=>"111001000",
  36169=>"110100110",
  36170=>"111111110",
  36171=>"110110010",
  36172=>"000000001",
  36173=>"111000011",
  36174=>"110111110",
  36175=>"000000010",
  36176=>"111100101",
  36177=>"000000111",
  36178=>"111111111",
  36179=>"000011111",
  36180=>"000000111",
  36181=>"011111111",
  36182=>"111111111",
  36183=>"101001001",
  36184=>"010010000",
  36185=>"111111111",
  36186=>"000000000",
  36187=>"110111110",
  36188=>"111111000",
  36189=>"000000000",
  36190=>"110000101",
  36191=>"011001111",
  36192=>"101111111",
  36193=>"111111111",
  36194=>"110100000",
  36195=>"111010000",
  36196=>"111110110",
  36197=>"001000000",
  36198=>"000000000",
  36199=>"001001101",
  36200=>"110000000",
  36201=>"111111001",
  36202=>"011111000",
  36203=>"100000000",
  36204=>"010111111",
  36205=>"010111111",
  36206=>"001111111",
  36207=>"111000110",
  36208=>"011000000",
  36209=>"111111101",
  36210=>"000000010",
  36211=>"011111111",
  36212=>"011111111",
  36213=>"000000000",
  36214=>"100000111",
  36215=>"111111111",
  36216=>"101000000",
  36217=>"111111000",
  36218=>"111010000",
  36219=>"111111100",
  36220=>"100000100",
  36221=>"111011111",
  36222=>"111110110",
  36223=>"111111000",
  36224=>"100110000",
  36225=>"111100111",
  36226=>"011011000",
  36227=>"111111100",
  36228=>"010000000",
  36229=>"000000011",
  36230=>"111110111",
  36231=>"111100000",
  36232=>"111111111",
  36233=>"100000011",
  36234=>"111111101",
  36235=>"000110111",
  36236=>"111000001",
  36237=>"000011111",
  36238=>"001000001",
  36239=>"111110000",
  36240=>"111111100",
  36241=>"000000110",
  36242=>"100100111",
  36243=>"000000001",
  36244=>"000000111",
  36245=>"000000110",
  36246=>"110000000",
  36247=>"000000111",
  36248=>"101001011",
  36249=>"110000000",
  36250=>"000100111",
  36251=>"111111000",
  36252=>"000000000",
  36253=>"110111001",
  36254=>"000000111",
  36255=>"111110111",
  36256=>"000000111",
  36257=>"100100100",
  36258=>"101001111",
  36259=>"111111010",
  36260=>"100000001",
  36261=>"111111111",
  36262=>"111111111",
  36263=>"111111111",
  36264=>"000000110",
  36265=>"000000000",
  36266=>"100000000",
  36267=>"111111111",
  36268=>"000000000",
  36269=>"101110110",
  36270=>"000000000",
  36271=>"001011000",
  36272=>"100100000",
  36273=>"000111111",
  36274=>"000000111",
  36275=>"001000001",
  36276=>"000000000",
  36277=>"111101111",
  36278=>"111111101",
  36279=>"011011011",
  36280=>"011111111",
  36281=>"000000011",
  36282=>"111100000",
  36283=>"111111010",
  36284=>"111111111",
  36285=>"110001111",
  36286=>"000111111",
  36287=>"011011011",
  36288=>"111111111",
  36289=>"111111111",
  36290=>"111000000",
  36291=>"111111000",
  36292=>"000000100",
  36293=>"111100000",
  36294=>"000000111",
  36295=>"000000111",
  36296=>"101100111",
  36297=>"010011111",
  36298=>"111000101",
  36299=>"001111011",
  36300=>"110000000",
  36301=>"111010110",
  36302=>"001000000",
  36303=>"111111011",
  36304=>"000100110",
  36305=>"111111000",
  36306=>"000001111",
  36307=>"011010011",
  36308=>"000000001",
  36309=>"111111110",
  36310=>"101001001",
  36311=>"000000110",
  36312=>"111111000",
  36313=>"000000000",
  36314=>"111111000",
  36315=>"111011111",
  36316=>"001000110",
  36317=>"111000000",
  36318=>"000100111",
  36319=>"000010111",
  36320=>"111110111",
  36321=>"111111000",
  36322=>"000000111",
  36323=>"111000110",
  36324=>"000000000",
  36325=>"111111001",
  36326=>"111111001",
  36327=>"000000111",
  36328=>"001000111",
  36329=>"111011000",
  36330=>"000000000",
  36331=>"011111111",
  36332=>"101111000",
  36333=>"110000100",
  36334=>"000001001",
  36335=>"110110111",
  36336=>"000001111",
  36337=>"111000000",
  36338=>"000000111",
  36339=>"111101011",
  36340=>"110111111",
  36341=>"000000000",
  36342=>"000000110",
  36343=>"000000100",
  36344=>"001111111",
  36345=>"000000100",
  36346=>"000000000",
  36347=>"110001001",
  36348=>"000000000",
  36349=>"111000000",
  36350=>"000100010",
  36351=>"000000111",
  36352=>"001001000",
  36353=>"111001000",
  36354=>"111000111",
  36355=>"000000111",
  36356=>"010110111",
  36357=>"001111111",
  36358=>"111000000",
  36359=>"111000000",
  36360=>"000001000",
  36361=>"111110111",
  36362=>"001000001",
  36363=>"001011111",
  36364=>"111000000",
  36365=>"000000100",
  36366=>"000000011",
  36367=>"111111111",
  36368=>"010111111",
  36369=>"000000111",
  36370=>"000111010",
  36371=>"000000000",
  36372=>"001011001",
  36373=>"011011011",
  36374=>"000000110",
  36375=>"000100110",
  36376=>"100110100",
  36377=>"011110100",
  36378=>"000100111",
  36379=>"111111011",
  36380=>"111000000",
  36381=>"001001111",
  36382=>"100110000",
  36383=>"111111000",
  36384=>"111111000",
  36385=>"000000101",
  36386=>"000001111",
  36387=>"000000000",
  36388=>"100000000",
  36389=>"000111111",
  36390=>"000000001",
  36391=>"000111111",
  36392=>"000000111",
  36393=>"000110000",
  36394=>"111000000",
  36395=>"111000000",
  36396=>"111111010",
  36397=>"001001111",
  36398=>"110100011",
  36399=>"000000100",
  36400=>"010111000",
  36401=>"000000000",
  36402=>"000000011",
  36403=>"100111111",
  36404=>"001101111",
  36405=>"011011001",
  36406=>"000001001",
  36407=>"100100111",
  36408=>"000000011",
  36409=>"000000111",
  36410=>"111100111",
  36411=>"110000001",
  36412=>"000000000",
  36413=>"001000000",
  36414=>"001000000",
  36415=>"110100000",
  36416=>"011110110",
  36417=>"100111110",
  36418=>"111111111",
  36419=>"000000001",
  36420=>"000111000",
  36421=>"111110100",
  36422=>"111010111",
  36423=>"001000010",
  36424=>"111011000",
  36425=>"111010000",
  36426=>"000000001",
  36427=>"111111011",
  36428=>"111111111",
  36429=>"111111000",
  36430=>"100000111",
  36431=>"000000001",
  36432=>"111111111",
  36433=>"111000001",
  36434=>"000000100",
  36435=>"101100000",
  36436=>"111000000",
  36437=>"100111111",
  36438=>"011000100",
  36439=>"111111110",
  36440=>"001000000",
  36441=>"111111111",
  36442=>"111011000",
  36443=>"000111100",
  36444=>"111011111",
  36445=>"000111110",
  36446=>"111101000",
  36447=>"011111111",
  36448=>"000001000",
  36449=>"000000000",
  36450=>"000010000",
  36451=>"000000000",
  36452=>"111000110",
  36453=>"111000111",
  36454=>"111001100",
  36455=>"000000101",
  36456=>"111111011",
  36457=>"110100000",
  36458=>"000101111",
  36459=>"000000000",
  36460=>"000000000",
  36461=>"010110000",
  36462=>"111111001",
  36463=>"010000111",
  36464=>"111111000",
  36465=>"000001111",
  36466=>"111011001",
  36467=>"011011000",
  36468=>"010000000",
  36469=>"000100101",
  36470=>"000000000",
  36471=>"000011111",
  36472=>"000000000",
  36473=>"111000111",
  36474=>"000000000",
  36475=>"111000000",
  36476=>"000001110",
  36477=>"111111111",
  36478=>"000000000",
  36479=>"111011000",
  36480=>"000111010",
  36481=>"110100011",
  36482=>"010010111",
  36483=>"111011101",
  36484=>"110000000",
  36485=>"111111001",
  36486=>"110111111",
  36487=>"111000100",
  36488=>"111111111",
  36489=>"111110110",
  36490=>"000111000",
  36491=>"001000000",
  36492=>"001000000",
  36493=>"111111111",
  36494=>"011010110",
  36495=>"000000000",
  36496=>"000000101",
  36497=>"111011000",
  36498=>"000110000",
  36499=>"000100111",
  36500=>"111000000",
  36501=>"011001001",
  36502=>"000011111",
  36503=>"111000001",
  36504=>"100000000",
  36505=>"000000000",
  36506=>"000111111",
  36507=>"000101000",
  36508=>"111111111",
  36509=>"000100100",
  36510=>"101101111",
  36511=>"001000001",
  36512=>"100110000",
  36513=>"000000000",
  36514=>"000000000",
  36515=>"000111111",
  36516=>"011001111",
  36517=>"111100000",
  36518=>"101111001",
  36519=>"101101101",
  36520=>"000100111",
  36521=>"000000011",
  36522=>"011000000",
  36523=>"000111111",
  36524=>"000000011",
  36525=>"011010011",
  36526=>"111111111",
  36527=>"000111011",
  36528=>"111101000",
  36529=>"110010010",
  36530=>"010111111",
  36531=>"011101000",
  36532=>"100111111",
  36533=>"000111111",
  36534=>"011111000",
  36535=>"101111101",
  36536=>"111111111",
  36537=>"111111111",
  36538=>"111000000",
  36539=>"001101000",
  36540=>"000000000",
  36541=>"111111101",
  36542=>"000000100",
  36543=>"000000000",
  36544=>"111100110",
  36545=>"001000111",
  36546=>"111000100",
  36547=>"000000000",
  36548=>"111100111",
  36549=>"001000001",
  36550=>"100000100",
  36551=>"000000000",
  36552=>"000110111",
  36553=>"110000000",
  36554=>"000000100",
  36555=>"111111000",
  36556=>"111101101",
  36557=>"001111001",
  36558=>"101111111",
  36559=>"111111111",
  36560=>"000010000",
  36561=>"000000010",
  36562=>"000000100",
  36563=>"111111111",
  36564=>"000000001",
  36565=>"011001011",
  36566=>"000000000",
  36567=>"100110000",
  36568=>"100000111",
  36569=>"101100100",
  36570=>"111001111",
  36571=>"111101000",
  36572=>"000101111",
  36573=>"111000011",
  36574=>"000000000",
  36575=>"111000000",
  36576=>"001111111",
  36577=>"111111000",
  36578=>"000110000",
  36579=>"001111010",
  36580=>"000000001",
  36581=>"001111011",
  36582=>"111000111",
  36583=>"001000011",
  36584=>"111111000",
  36585=>"000000000",
  36586=>"111111011",
  36587=>"111111000",
  36588=>"000000000",
  36589=>"001001111",
  36590=>"000111111",
  36591=>"111111111",
  36592=>"110111111",
  36593=>"011111011",
  36594=>"000001111",
  36595=>"000000101",
  36596=>"000111110",
  36597=>"110111111",
  36598=>"000000000",
  36599=>"111000000",
  36600=>"100000101",
  36601=>"000000000",
  36602=>"000000000",
  36603=>"000000010",
  36604=>"001101000",
  36605=>"000100111",
  36606=>"000000001",
  36607=>"111000000",
  36608=>"101000100",
  36609=>"000110011",
  36610=>"100000000",
  36611=>"000100111",
  36612=>"111011111",
  36613=>"111000110",
  36614=>"000000111",
  36615=>"110111110",
  36616=>"000000000",
  36617=>"111111000",
  36618=>"111111010",
  36619=>"111111100",
  36620=>"000000000",
  36621=>"101001000",
  36622=>"000000001",
  36623=>"111111110",
  36624=>"100100100",
  36625=>"000000111",
  36626=>"111000111",
  36627=>"000001111",
  36628=>"000000110",
  36629=>"111011001",
  36630=>"001001101",
  36631=>"000000000",
  36632=>"000001101",
  36633=>"111001111",
  36634=>"110100111",
  36635=>"101111111",
  36636=>"011011000",
  36637=>"111100000",
  36638=>"111000000",
  36639=>"000000000",
  36640=>"000000100",
  36641=>"111011000",
  36642=>"111111000",
  36643=>"000110000",
  36644=>"110111000",
  36645=>"111000000",
  36646=>"101000110",
  36647=>"110111000",
  36648=>"000000111",
  36649=>"000100010",
  36650=>"000000111",
  36651=>"000111101",
  36652=>"111111000",
  36653=>"000000001",
  36654=>"000000111",
  36655=>"010111111",
  36656=>"111000001",
  36657=>"000000000",
  36658=>"111000000",
  36659=>"000000111",
  36660=>"011111011",
  36661=>"101111111",
  36662=>"000000000",
  36663=>"111000101",
  36664=>"000111001",
  36665=>"011011001",
  36666=>"000000000",
  36667=>"111111011",
  36668=>"000000000",
  36669=>"000111111",
  36670=>"000000000",
  36671=>"001001111",
  36672=>"011011000",
  36673=>"111111110",
  36674=>"111000000",
  36675=>"111111111",
  36676=>"000000010",
  36677=>"111111111",
  36678=>"000000000",
  36679=>"000000110",
  36680=>"000000000",
  36681=>"000000000",
  36682=>"000000000",
  36683=>"101111111",
  36684=>"000100111",
  36685=>"000110000",
  36686=>"100100000",
  36687=>"111110000",
  36688=>"000111111",
  36689=>"001001111",
  36690=>"111111000",
  36691=>"001001000",
  36692=>"010001111",
  36693=>"000111011",
  36694=>"000110111",
  36695=>"110111111",
  36696=>"111111111",
  36697=>"001111001",
  36698=>"111111110",
  36699=>"001000110",
  36700=>"011101000",
  36701=>"100110111",
  36702=>"101101101",
  36703=>"011000101",
  36704=>"000111111",
  36705=>"000000111",
  36706=>"001001100",
  36707=>"111110000",
  36708=>"001001001",
  36709=>"000000000",
  36710=>"000110000",
  36711=>"000000000",
  36712=>"011001101",
  36713=>"111111111",
  36714=>"111111000",
  36715=>"000110000",
  36716=>"111111100",
  36717=>"000000111",
  36718=>"101111111",
  36719=>"000000000",
  36720=>"000111110",
  36721=>"110110111",
  36722=>"011001000",
  36723=>"000111011",
  36724=>"000000000",
  36725=>"010110111",
  36726=>"000000000",
  36727=>"110010000",
  36728=>"000111010",
  36729=>"001000000",
  36730=>"111011111",
  36731=>"001000000",
  36732=>"111111110",
  36733=>"000000000",
  36734=>"000000000",
  36735=>"111111110",
  36736=>"100000100",
  36737=>"111101010",
  36738=>"110111001",
  36739=>"000000000",
  36740=>"111111111",
  36741=>"111111111",
  36742=>"000110110",
  36743=>"111101000",
  36744=>"111000111",
  36745=>"000000000",
  36746=>"000000110",
  36747=>"000010111",
  36748=>"011111111",
  36749=>"111110110",
  36750=>"111001001",
  36751=>"111000101",
  36752=>"000000000",
  36753=>"110111111",
  36754=>"111111111",
  36755=>"111100111",
  36756=>"100111000",
  36757=>"001111111",
  36758=>"111010010",
  36759=>"000000011",
  36760=>"001011111",
  36761=>"110010000",
  36762=>"000000000",
  36763=>"111111111",
  36764=>"111111110",
  36765=>"001000000",
  36766=>"110000000",
  36767=>"111111001",
  36768=>"000000000",
  36769=>"001111110",
  36770=>"111110000",
  36771=>"011011000",
  36772=>"111111110",
  36773=>"111111111",
  36774=>"011000111",
  36775=>"001011001",
  36776=>"111111111",
  36777=>"000000000",
  36778=>"001000110",
  36779=>"001001100",
  36780=>"000000000",
  36781=>"000000000",
  36782=>"111010011",
  36783=>"011010000",
  36784=>"111010000",
  36785=>"010111000",
  36786=>"000000100",
  36787=>"111111111",
  36788=>"100001011",
  36789=>"000000001",
  36790=>"010111111",
  36791=>"110111111",
  36792=>"000000000",
  36793=>"111111001",
  36794=>"111100001",
  36795=>"110111111",
  36796=>"001111111",
  36797=>"000000000",
  36798=>"000000111",
  36799=>"000101000",
  36800=>"000100111",
  36801=>"000001000",
  36802=>"011001000",
  36803=>"000111111",
  36804=>"101000111",
  36805=>"100100110",
  36806=>"001001011",
  36807=>"000000011",
  36808=>"111111111",
  36809=>"000011000",
  36810=>"001000010",
  36811=>"111111111",
  36812=>"111111111",
  36813=>"000000111",
  36814=>"111000000",
  36815=>"000000100",
  36816=>"000000000",
  36817=>"011111011",
  36818=>"111011111",
  36819=>"011111111",
  36820=>"000000010",
  36821=>"111000000",
  36822=>"000000000",
  36823=>"111100000",
  36824=>"101000011",
  36825=>"111111000",
  36826=>"111111100",
  36827=>"111011101",
  36828=>"110000110",
  36829=>"000000000",
  36830=>"001000111",
  36831=>"000001001",
  36832=>"000000011",
  36833=>"001111111",
  36834=>"011000100",
  36835=>"111000100",
  36836=>"000000000",
  36837=>"101000000",
  36838=>"110110100",
  36839=>"000001000",
  36840=>"001000000",
  36841=>"001001111",
  36842=>"001001111",
  36843=>"000100111",
  36844=>"111000000",
  36845=>"000000110",
  36846=>"011001000",
  36847=>"000111111",
  36848=>"000000000",
  36849=>"111111111",
  36850=>"000100111",
  36851=>"111111000",
  36852=>"000101111",
  36853=>"001000000",
  36854=>"011000000",
  36855=>"011010000",
  36856=>"000111111",
  36857=>"011011010",
  36858=>"000000000",
  36859=>"001011111",
  36860=>"000100111",
  36861=>"111111110",
  36862=>"111111111",
  36863=>"000000000",
  36864=>"000000000",
  36865=>"000000000",
  36866=>"000000000",
  36867=>"000110111",
  36868=>"000000000",
  36869=>"111110100",
  36870=>"000000000",
  36871=>"000000000",
  36872=>"111111111",
  36873=>"000000111",
  36874=>"110111111",
  36875=>"001111111",
  36876=>"001001001",
  36877=>"111111101",
  36878=>"100100001",
  36879=>"000100110",
  36880=>"001100001",
  36881=>"111111111",
  36882=>"000000000",
  36883=>"111111110",
  36884=>"000000001",
  36885=>"000000001",
  36886=>"110100100",
  36887=>"000000110",
  36888=>"011111011",
  36889=>"000000000",
  36890=>"111001000",
  36891=>"000111111",
  36892=>"111111111",
  36893=>"000010010",
  36894=>"011011011",
  36895=>"110011011",
  36896=>"111111111",
  36897=>"001001001",
  36898=>"000000010",
  36899=>"111111111",
  36900=>"000100100",
  36901=>"000011010",
  36902=>"000000000",
  36903=>"111111111",
  36904=>"011010010",
  36905=>"001001111",
  36906=>"111111111",
  36907=>"111111111",
  36908=>"111111111",
  36909=>"111111111",
  36910=>"111000000",
  36911=>"111111111",
  36912=>"000000000",
  36913=>"111111111",
  36914=>"001001011",
  36915=>"000000000",
  36916=>"111111100",
  36917=>"000000000",
  36918=>"001111100",
  36919=>"100111111",
  36920=>"000000000",
  36921=>"000000011",
  36922=>"000000000",
  36923=>"000000000",
  36924=>"000000111",
  36925=>"111111111",
  36926=>"111111111",
  36927=>"111111010",
  36928=>"000000000",
  36929=>"101000000",
  36930=>"000000000",
  36931=>"000000100",
  36932=>"100001001",
  36933=>"100110111",
  36934=>"000000000",
  36935=>"000000000",
  36936=>"111111001",
  36937=>"000000111",
  36938=>"111110000",
  36939=>"101101111",
  36940=>"000000100",
  36941=>"111111111",
  36942=>"001000000",
  36943=>"111111111",
  36944=>"111001000",
  36945=>"011111100",
  36946=>"000001001",
  36947=>"001011001",
  36948=>"000000000",
  36949=>"111110010",
  36950=>"001000100",
  36951=>"111111111",
  36952=>"011011111",
  36953=>"000010000",
  36954=>"000010111",
  36955=>"111111100",
  36956=>"111111101",
  36957=>"000000000",
  36958=>"000000000",
  36959=>"100000000",
  36960=>"000000100",
  36961=>"111011011",
  36962=>"000000011",
  36963=>"001000111",
  36964=>"000000000",
  36965=>"000000001",
  36966=>"111111111",
  36967=>"000000000",
  36968=>"110111111",
  36969=>"111111011",
  36970=>"111010000",
  36971=>"101101111",
  36972=>"111001011",
  36973=>"111111111",
  36974=>"111111111",
  36975=>"011000000",
  36976=>"100100100",
  36977=>"000000000",
  36978=>"001101111",
  36979=>"000000100",
  36980=>"111111111",
  36981=>"001001000",
  36982=>"011111111",
  36983=>"000000000",
  36984=>"000001111",
  36985=>"111000000",
  36986=>"000000111",
  36987=>"000000000",
  36988=>"000100100",
  36989=>"000000000",
  36990=>"111011001",
  36991=>"111100000",
  36992=>"000001000",
  36993=>"010000111",
  36994=>"111111101",
  36995=>"000100000",
  36996=>"110000000",
  36997=>"000000000",
  36998=>"111111110",
  36999=>"111111111",
  37000=>"000000000",
  37001=>"000000000",
  37002=>"000000000",
  37003=>"000001101",
  37004=>"101101000",
  37005=>"000111011",
  37006=>"110100110",
  37007=>"111111111",
  37008=>"000000000",
  37009=>"011001101",
  37010=>"000001001",
  37011=>"000000000",
  37012=>"011000000",
  37013=>"011011001",
  37014=>"000000000",
  37015=>"110111111",
  37016=>"000000001",
  37017=>"000000100",
  37018=>"111111111",
  37019=>"111110111",
  37020=>"111111100",
  37021=>"000101000",
  37022=>"111000000",
  37023=>"100000000",
  37024=>"011111111",
  37025=>"111000000",
  37026=>"010000000",
  37027=>"010000000",
  37028=>"011111111",
  37029=>"101111111",
  37030=>"000000001",
  37031=>"101100000",
  37032=>"000111111",
  37033=>"000111111",
  37034=>"110110110",
  37035=>"101000000",
  37036=>"000000000",
  37037=>"100000000",
  37038=>"000000000",
  37039=>"111111000",
  37040=>"111110000",
  37041=>"100100100",
  37042=>"000111111",
  37043=>"001000111",
  37044=>"110100000",
  37045=>"011111001",
  37046=>"001000100",
  37047=>"000000000",
  37048=>"000101011",
  37049=>"011111000",
  37050=>"000100100",
  37051=>"110110000",
  37052=>"011011000",
  37053=>"000001000",
  37054=>"111001001",
  37055=>"101000101",
  37056=>"111111111",
  37057=>"101101000",
  37058=>"000000000",
  37059=>"111111111",
  37060=>"110110110",
  37061=>"000000000",
  37062=>"001100100",
  37063=>"000000000",
  37064=>"000000000",
  37065=>"111100000",
  37066=>"011100100",
  37067=>"000001101",
  37068=>"000000000",
  37069=>"000010011",
  37070=>"100011110",
  37071=>"110111111",
  37072=>"011100110",
  37073=>"110011011",
  37074=>"011111111",
  37075=>"000000000",
  37076=>"001000000",
  37077=>"000000001",
  37078=>"111111111",
  37079=>"100111111",
  37080=>"000001011",
  37081=>"000111111",
  37082=>"000000000",
  37083=>"000000000",
  37084=>"111100111",
  37085=>"111111111",
  37086=>"111001001",
  37087=>"100000000",
  37088=>"000000000",
  37089=>"000000000",
  37090=>"000000000",
  37091=>"000000000",
  37092=>"001000000",
  37093=>"110110000",
  37094=>"111011010",
  37095=>"000000000",
  37096=>"111111111",
  37097=>"000000000",
  37098=>"110111000",
  37099=>"111111111",
  37100=>"000000000",
  37101=>"010111111",
  37102=>"111111111",
  37103=>"111111001",
  37104=>"000000000",
  37105=>"000000000",
  37106=>"111110111",
  37107=>"000000000",
  37108=>"111111111",
  37109=>"111111001",
  37110=>"111001011",
  37111=>"000000000",
  37112=>"110111111",
  37113=>"000000000",
  37114=>"000000000",
  37115=>"000000000",
  37116=>"011011000",
  37117=>"111011001",
  37118=>"100000111",
  37119=>"000000000",
  37120=>"000000000",
  37121=>"101101001",
  37122=>"111111010",
  37123=>"000000000",
  37124=>"110001111",
  37125=>"111000000",
  37126=>"100111111",
  37127=>"000001111",
  37128=>"000111111",
  37129=>"000000000",
  37130=>"111111111",
  37131=>"100100000",
  37132=>"001111111",
  37133=>"011001000",
  37134=>"111111111",
  37135=>"000100111",
  37136=>"000000001",
  37137=>"100110100",
  37138=>"001000000",
  37139=>"011111000",
  37140=>"001011000",
  37141=>"001001001",
  37142=>"001001001",
  37143=>"111111111",
  37144=>"000000100",
  37145=>"011011000",
  37146=>"111000000",
  37147=>"111111111",
  37148=>"111111111",
  37149=>"001011000",
  37150=>"000000000",
  37151=>"001001000",
  37152=>"000000000",
  37153=>"111100101",
  37154=>"000000000",
  37155=>"000100110",
  37156=>"000000100",
  37157=>"000000000",
  37158=>"110110110",
  37159=>"001101111",
  37160=>"111111000",
  37161=>"000000000",
  37162=>"000000110",
  37163=>"000000011",
  37164=>"000101111",
  37165=>"111101110",
  37166=>"000000000",
  37167=>"000000001",
  37168=>"111111111",
  37169=>"000001001",
  37170=>"000000000",
  37171=>"000000000",
  37172=>"000000001",
  37173=>"001000100",
  37174=>"110100001",
  37175=>"100100000",
  37176=>"000000000",
  37177=>"100000001",
  37178=>"110110111",
  37179=>"111111100",
  37180=>"111111111",
  37181=>"000000000",
  37182=>"000000000",
  37183=>"111100100",
  37184=>"000000000",
  37185=>"010111111",
  37186=>"000010000",
  37187=>"000000100",
  37188=>"111111001",
  37189=>"001001000",
  37190=>"101011111",
  37191=>"000000000",
  37192=>"111010010",
  37193=>"111111111",
  37194=>"000000000",
  37195=>"000000000",
  37196=>"111111111",
  37197=>"000000000",
  37198=>"111000000",
  37199=>"011110000",
  37200=>"100111111",
  37201=>"110111111",
  37202=>"111111111",
  37203=>"111111111",
  37204=>"001000000",
  37205=>"001011000",
  37206=>"111111111",
  37207=>"111111111",
  37208=>"000000000",
  37209=>"111111111",
  37210=>"100000000",
  37211=>"111110100",
  37212=>"000000000",
  37213=>"111111111",
  37214=>"000000000",
  37215=>"000110110",
  37216=>"001000000",
  37217=>"001000001",
  37218=>"000000000",
  37219=>"111111111",
  37220=>"100110110",
  37221=>"000000000",
  37222=>"000000000",
  37223=>"111111111",
  37224=>"111110111",
  37225=>"000000000",
  37226=>"111111111",
  37227=>"101100101",
  37228=>"111111111",
  37229=>"000000000",
  37230=>"111011000",
  37231=>"100100101",
  37232=>"000000001",
  37233=>"111111111",
  37234=>"000000000",
  37235=>"111011000",
  37236=>"111111111",
  37237=>"100001001",
  37238=>"000000001",
  37239=>"100111001",
  37240=>"111111111",
  37241=>"011111111",
  37242=>"111111111",
  37243=>"000011011",
  37244=>"111101101",
  37245=>"001001000",
  37246=>"111111111",
  37247=>"000000000",
  37248=>"111110001",
  37249=>"001000111",
  37250=>"001000000",
  37251=>"001000010",
  37252=>"111111000",
  37253=>"000111111",
  37254=>"101111110",
  37255=>"011011110",
  37256=>"000000000",
  37257=>"111111111",
  37258=>"100101001",
  37259=>"000000000",
  37260=>"111111111",
  37261=>"001001001",
  37262=>"100000000",
  37263=>"110110111",
  37264=>"011011001",
  37265=>"111111011",
  37266=>"011011000",
  37267=>"111011011",
  37268=>"000000000",
  37269=>"000010000",
  37270=>"000000000",
  37271=>"100100100",
  37272=>"101111110",
  37273=>"111001011",
  37274=>"110111111",
  37275=>"000100000",
  37276=>"111111111",
  37277=>"000111111",
  37278=>"010000000",
  37279=>"000111111",
  37280=>"000011001",
  37281=>"001001000",
  37282=>"110010000",
  37283=>"000111111",
  37284=>"000000000",
  37285=>"000011001",
  37286=>"000000000",
  37287=>"111100110",
  37288=>"111111000",
  37289=>"110110100",
  37290=>"010000000",
  37291=>"111011000",
  37292=>"000001111",
  37293=>"000000000",
  37294=>"111111111",
  37295=>"001001011",
  37296=>"000000110",
  37297=>"000011000",
  37298=>"100111011",
  37299=>"000001011",
  37300=>"111100101",
  37301=>"000000000",
  37302=>"111111111",
  37303=>"111111111",
  37304=>"111001000",
  37305=>"101111000",
  37306=>"111111101",
  37307=>"011011000",
  37308=>"111111110",
  37309=>"111111111",
  37310=>"000000100",
  37311=>"101111111",
  37312=>"000000000",
  37313=>"111111111",
  37314=>"000000101",
  37315=>"111111111",
  37316=>"001011000",
  37317=>"000000000",
  37318=>"111111111",
  37319=>"011011111",
  37320=>"000000000",
  37321=>"000000000",
  37322=>"100100100",
  37323=>"000000001",
  37324=>"101111101",
  37325=>"001000000",
  37326=>"000000000",
  37327=>"000000000",
  37328=>"111000000",
  37329=>"110111111",
  37330=>"111111111",
  37331=>"000001001",
  37332=>"111000000",
  37333=>"011101000",
  37334=>"111000111",
  37335=>"110110111",
  37336=>"100100000",
  37337=>"111110000",
  37338=>"111111110",
  37339=>"000100101",
  37340=>"101000011",
  37341=>"000111011",
  37342=>"000001011",
  37343=>"111100001",
  37344=>"111111110",
  37345=>"111111100",
  37346=>"000000000",
  37347=>"111111000",
  37348=>"010011000",
  37349=>"011001001",
  37350=>"111100111",
  37351=>"110010000",
  37352=>"000000100",
  37353=>"000001101",
  37354=>"000000000",
  37355=>"000000000",
  37356=>"000000000",
  37357=>"000110110",
  37358=>"000011011",
  37359=>"000000000",
  37360=>"111111111",
  37361=>"001001111",
  37362=>"111110100",
  37363=>"000000000",
  37364=>"111110100",
  37365=>"011101100",
  37366=>"111111111",
  37367=>"101111111",
  37368=>"001001111",
  37369=>"100100000",
  37370=>"111011001",
  37371=>"001000000",
  37372=>"111111000",
  37373=>"000000000",
  37374=>"001000000",
  37375=>"101001111",
  37376=>"101011011",
  37377=>"111111110",
  37378=>"000000001",
  37379=>"100000000",
  37380=>"001000000",
  37381=>"001000000",
  37382=>"111001001",
  37383=>"000000101",
  37384=>"111111111",
  37385=>"111000000",
  37386=>"011011001",
  37387=>"000100100",
  37388=>"000000000",
  37389=>"000001011",
  37390=>"100000011",
  37391=>"111111110",
  37392=>"000001011",
  37393=>"010011001",
  37394=>"000000000",
  37395=>"111000000",
  37396=>"001000101",
  37397=>"000000000",
  37398=>"000000000",
  37399=>"000000111",
  37400=>"001000110",
  37401=>"000100000",
  37402=>"100000000",
  37403=>"000110010",
  37404=>"111001001",
  37405=>"010010010",
  37406=>"000001101",
  37407=>"000000001",
  37408=>"110110010",
  37409=>"100110110",
  37410=>"110110100",
  37411=>"101111101",
  37412=>"110110000",
  37413=>"111111000",
  37414=>"000000000",
  37415=>"000000000",
  37416=>"100100110",
  37417=>"000000000",
  37418=>"111100111",
  37419=>"111110000",
  37420=>"000000111",
  37421=>"110001000",
  37422=>"111111001",
  37423=>"010001000",
  37424=>"101000110",
  37425=>"011010000",
  37426=>"100000100",
  37427=>"000100010",
  37428=>"000100110",
  37429=>"110110010",
  37430=>"000000000",
  37431=>"001000100",
  37432=>"000100111",
  37433=>"000000110",
  37434=>"001101111",
  37435=>"000101100",
  37436=>"010001000",
  37437=>"000000000",
  37438=>"111111111",
  37439=>"011000000",
  37440=>"111111000",
  37441=>"001001111",
  37442=>"000000000",
  37443=>"000000101",
  37444=>"000100100",
  37445=>"000000100",
  37446=>"000001000",
  37447=>"111111111",
  37448=>"110110000",
  37449=>"111001111",
  37450=>"000000110",
  37451=>"000001111",
  37452=>"110110111",
  37453=>"001011111",
  37454=>"111000000",
  37455=>"000000000",
  37456=>"001111111",
  37457=>"001001000",
  37458=>"111111011",
  37459=>"110100110",
  37460=>"111111001",
  37461=>"111111000",
  37462=>"000001111",
  37463=>"001000000",
  37464=>"100100000",
  37465=>"101001111",
  37466=>"111111111",
  37467=>"110111110",
  37468=>"100100000",
  37469=>"110110111",
  37470=>"111110110",
  37471=>"110010110",
  37472=>"000111110",
  37473=>"110110000",
  37474=>"000000111",
  37475=>"011011111",
  37476=>"000000110",
  37477=>"010011000",
  37478=>"001001111",
  37479=>"000000001",
  37480=>"111111111",
  37481=>"000000001",
  37482=>"001000001",
  37483=>"111111110",
  37484=>"111111111",
  37485=>"000000000",
  37486=>"111011111",
  37487=>"011111011",
  37488=>"110000000",
  37489=>"110110000",
  37490=>"101010000",
  37491=>"000110111",
  37492=>"101111111",
  37493=>"111111111",
  37494=>"001000000",
  37495=>"001001111",
  37496=>"000001110",
  37497=>"000101000",
  37498=>"000000000",
  37499=>"000000000",
  37500=>"100110111",
  37501=>"000001001",
  37502=>"100000000",
  37503=>"001000000",
  37504=>"111100100",
  37505=>"100111111",
  37506=>"101000111",
  37507=>"001110110",
  37508=>"000001000",
  37509=>"001111111",
  37510=>"010010000",
  37511=>"000000001",
  37512=>"000000101",
  37513=>"110110110",
  37514=>"001000001",
  37515=>"000010011",
  37516=>"000000111",
  37517=>"010110110",
  37518=>"110110010",
  37519=>"000000000",
  37520=>"001000111",
  37521=>"000111011",
  37522=>"001011000",
  37523=>"001100111",
  37524=>"000001101",
  37525=>"001001001",
  37526=>"100111111",
  37527=>"100100111",
  37528=>"001000000",
  37529=>"001001001",
  37530=>"111111011",
  37531=>"001000001",
  37532=>"111100000",
  37533=>"001000001",
  37534=>"001000101",
  37535=>"000001011",
  37536=>"110000000",
  37537=>"010110000",
  37538=>"001001000",
  37539=>"001011011",
  37540=>"100000000",
  37541=>"110010000",
  37542=>"110110111",
  37543=>"000000000",
  37544=>"000000111",
  37545=>"000000000",
  37546=>"111111111",
  37547=>"101000111",
  37548=>"110000000",
  37549=>"110110110",
  37550=>"111110110",
  37551=>"000000100",
  37552=>"000000010",
  37553=>"111110000",
  37554=>"110110010",
  37555=>"101000000",
  37556=>"010011001",
  37557=>"001000001",
  37558=>"110110010",
  37559=>"001001001",
  37560=>"111111111",
  37561=>"111111111",
  37562=>"000000000",
  37563=>"011000000",
  37564=>"000000101",
  37565=>"111111111",
  37566=>"001101000",
  37567=>"101111111",
  37568=>"111111100",
  37569=>"000100111",
  37570=>"000000000",
  37571=>"110110010",
  37572=>"111111011",
  37573=>"000000000",
  37574=>"000000000",
  37575=>"000001111",
  37576=>"000000111",
  37577=>"001001001",
  37578=>"101101001",
  37579=>"100111110",
  37580=>"000000110",
  37581=>"000010111",
  37582=>"001000110",
  37583=>"110111000",
  37584=>"111111001",
  37585=>"001100110",
  37586=>"111110110",
  37587=>"000000001",
  37588=>"000000111",
  37589=>"110000110",
  37590=>"000000000",
  37591=>"011001001",
  37592=>"111111001",
  37593=>"011001111",
  37594=>"101111111",
  37595=>"110111111",
  37596=>"010000000",
  37597=>"000001001",
  37598=>"100110110",
  37599=>"001111110",
  37600=>"111111111",
  37601=>"010010001",
  37602=>"101000101",
  37603=>"001001001",
  37604=>"111111001",
  37605=>"110110111",
  37606=>"111111110",
  37607=>"100000000",
  37608=>"110111111",
  37609=>"000000001",
  37610=>"000100111",
  37611=>"000000000",
  37612=>"000000000",
  37613=>"101000000",
  37614=>"111111111",
  37615=>"000000101",
  37616=>"111101111",
  37617=>"101111111",
  37618=>"000000000",
  37619=>"000000100",
  37620=>"111010000",
  37621=>"011110010",
  37622=>"000111001",
  37623=>"111001000",
  37624=>"011000000",
  37625=>"111111111",
  37626=>"110111110",
  37627=>"000000000",
  37628=>"100100100",
  37629=>"011111111",
  37630=>"010001001",
  37631=>"110111000",
  37632=>"011111111",
  37633=>"001011011",
  37634=>"000000000",
  37635=>"110100111",
  37636=>"000110101",
  37637=>"111111110",
  37638=>"101101111",
  37639=>"000000111",
  37640=>"000000111",
  37641=>"000110001",
  37642=>"000000000",
  37643=>"000000111",
  37644=>"100000010",
  37645=>"000000000",
  37646=>"110111111",
  37647=>"111111000",
  37648=>"010001001",
  37649=>"111111001",
  37650=>"111111111",
  37651=>"111001001",
  37652=>"000000000",
  37653=>"001001001",
  37654=>"011110100",
  37655=>"000000000",
  37656=>"110110110",
  37657=>"001001000",
  37658=>"001000000",
  37659=>"110110110",
  37660=>"011000000",
  37661=>"111111000",
  37662=>"111111111",
  37663=>"000000000",
  37664=>"000000000",
  37665=>"001011111",
  37666=>"110111110",
  37667=>"000100110",
  37668=>"101111111",
  37669=>"110111111",
  37670=>"111111010",
  37671=>"110110110",
  37672=>"000000011",
  37673=>"110110110",
  37674=>"000110010",
  37675=>"111000000",
  37676=>"000000000",
  37677=>"011011000",
  37678=>"111010010",
  37679=>"100000110",
  37680=>"110110011",
  37681=>"100110111",
  37682=>"111111110",
  37683=>"111001000",
  37684=>"000101000",
  37685=>"000000000",
  37686=>"010010000",
  37687=>"111000000",
  37688=>"000110110",
  37689=>"100000101",
  37690=>"001001101",
  37691=>"110111100",
  37692=>"011111111",
  37693=>"011011000",
  37694=>"000010000",
  37695=>"110110010",
  37696=>"111000000",
  37697=>"100110111",
  37698=>"000000111",
  37699=>"101001111",
  37700=>"110110000",
  37701=>"000010011",
  37702=>"001001011",
  37703=>"010110110",
  37704=>"010010010",
  37705=>"000000111",
  37706=>"001000100",
  37707=>"100100100",
  37708=>"000000000",
  37709=>"111000000",
  37710=>"000000000",
  37711=>"001001000",
  37712=>"000000100",
  37713=>"000001100",
  37714=>"001001001",
  37715=>"111011111",
  37716=>"000000000",
  37717=>"011011000",
  37718=>"111111110",
  37719=>"001000000",
  37720=>"111111111",
  37721=>"110000000",
  37722=>"110110010",
  37723=>"111111111",
  37724=>"101101001",
  37725=>"111111000",
  37726=>"110110110",
  37727=>"100100100",
  37728=>"001001101",
  37729=>"111111111",
  37730=>"000100000",
  37731=>"100000000",
  37732=>"001101111",
  37733=>"010001000",
  37734=>"000000000",
  37735=>"001001111",
  37736=>"011011011",
  37737=>"010000100",
  37738=>"111011011",
  37739=>"111001001",
  37740=>"110110111",
  37741=>"110011111",
  37742=>"111111111",
  37743=>"011000000",
  37744=>"001111111",
  37745=>"111111111",
  37746=>"110110100",
  37747=>"111111111",
  37748=>"001111000",
  37749=>"001001101",
  37750=>"001101111",
  37751=>"100110000",
  37752=>"000000000",
  37753=>"001011011",
  37754=>"000000100",
  37755=>"011001011",
  37756=>"111111111",
  37757=>"110110110",
  37758=>"000000011",
  37759=>"110110111",
  37760=>"110111111",
  37761=>"111001001",
  37762=>"000001011",
  37763=>"011011011",
  37764=>"000100111",
  37765=>"111011111",
  37766=>"000000111",
  37767=>"111110010",
  37768=>"000000110",
  37769=>"010000110",
  37770=>"110110000",
  37771=>"101100111",
  37772=>"111001111",
  37773=>"010011011",
  37774=>"111111111",
  37775=>"111111110",
  37776=>"001000010",
  37777=>"000000101",
  37778=>"000111111",
  37779=>"101101111",
  37780=>"000000000",
  37781=>"000000001",
  37782=>"111100000",
  37783=>"001000000",
  37784=>"111011001",
  37785=>"111111111",
  37786=>"100000001",
  37787=>"111110000",
  37788=>"000100110",
  37789=>"000000000",
  37790=>"001000000",
  37791=>"000100111",
  37792=>"010111111",
  37793=>"001011111",
  37794=>"110111111",
  37795=>"000000000",
  37796=>"110000000",
  37797=>"000111111",
  37798=>"110100111",
  37799=>"000111110",
  37800=>"111111101",
  37801=>"000000111",
  37802=>"110010000",
  37803=>"001000000",
  37804=>"000001111",
  37805=>"110110000",
  37806=>"011011010",
  37807=>"000000011",
  37808=>"000000100",
  37809=>"110110111",
  37810=>"111111111",
  37811=>"000000000",
  37812=>"111100000",
  37813=>"111000111",
  37814=>"111111111",
  37815=>"000111001",
  37816=>"000111111",
  37817=>"000100110",
  37818=>"000000000",
  37819=>"101100110",
  37820=>"000000000",
  37821=>"000000001",
  37822=>"111111010",
  37823=>"000010111",
  37824=>"000000110",
  37825=>"101000000",
  37826=>"111111001",
  37827=>"110111111",
  37828=>"111110110",
  37829=>"000001001",
  37830=>"000000010",
  37831=>"001001011",
  37832=>"000000000",
  37833=>"111111000",
  37834=>"001000000",
  37835=>"000000001",
  37836=>"110010000",
  37837=>"111111111",
  37838=>"000010111",
  37839=>"110111011",
  37840=>"001001001",
  37841=>"000111110",
  37842=>"000111111",
  37843=>"000000000",
  37844=>"110000000",
  37845=>"000000010",
  37846=>"010110010",
  37847=>"001000000",
  37848=>"111111010",
  37849=>"011111111",
  37850=>"011111000",
  37851=>"000000000",
  37852=>"111011001",
  37853=>"110110110",
  37854=>"111010000",
  37855=>"000001011",
  37856=>"001001000",
  37857=>"000001001",
  37858=>"000000000",
  37859=>"111011111",
  37860=>"011001001",
  37861=>"001111101",
  37862=>"110110110",
  37863=>"111101001",
  37864=>"101111111",
  37865=>"111111101",
  37866=>"000010010",
  37867=>"111111111",
  37868=>"111000111",
  37869=>"111110000",
  37870=>"001000000",
  37871=>"001000110",
  37872=>"000000000",
  37873=>"010110110",
  37874=>"000100110",
  37875=>"100101011",
  37876=>"000001000",
  37877=>"101001000",
  37878=>"011000000",
  37879=>"000101011",
  37880=>"000000111",
  37881=>"111100100",
  37882=>"000000000",
  37883=>"101011111",
  37884=>"000001010",
  37885=>"010110110",
  37886=>"011111111",
  37887=>"001001000",
  37888=>"110000101",
  37889=>"000110111",
  37890=>"010010011",
  37891=>"100000011",
  37892=>"000000110",
  37893=>"001000011",
  37894=>"110110100",
  37895=>"111000000",
  37896=>"111000001",
  37897=>"000101100",
  37898=>"000000111",
  37899=>"110101101",
  37900=>"000000000",
  37901=>"110110000",
  37902=>"001111010",
  37903=>"111111010",
  37904=>"000000000",
  37905=>"111111110",
  37906=>"111111010",
  37907=>"111111111",
  37908=>"000000111",
  37909=>"000111011",
  37910=>"010011011",
  37911=>"001001000",
  37912=>"000001001",
  37913=>"001111111",
  37914=>"001000000",
  37915=>"001111111",
  37916=>"011111111",
  37917=>"010010011",
  37918=>"011000000",
  37919=>"111101100",
  37920=>"111001001",
  37921=>"011010000",
  37922=>"000000010",
  37923=>"111111111",
  37924=>"110111000",
  37925=>"111110100",
  37926=>"110100000",
  37927=>"000110111",
  37928=>"111111001",
  37929=>"000000100",
  37930=>"111001111",
  37931=>"000000001",
  37932=>"111111101",
  37933=>"101101111",
  37934=>"111000000",
  37935=>"010000000",
  37936=>"000000111",
  37937=>"111111100",
  37938=>"000001111",
  37939=>"000000001",
  37940=>"000110111",
  37941=>"111101000",
  37942=>"100000000",
  37943=>"100000000",
  37944=>"100000011",
  37945=>"000000011",
  37946=>"000000010",
  37947=>"111000000",
  37948=>"001000000",
  37949=>"000000011",
  37950=>"101001110",
  37951=>"011000000",
  37952=>"000100111",
  37953=>"000110111",
  37954=>"000010111",
  37955=>"000000000",
  37956=>"011111010",
  37957=>"111110000",
  37958=>"111011000",
  37959=>"000110110",
  37960=>"000000000",
  37961=>"000111111",
  37962=>"110110111",
  37963=>"111111110",
  37964=>"001111111",
  37965=>"110100100",
  37966=>"111000000",
  37967=>"100111111",
  37968=>"110100000",
  37969=>"000000010",
  37970=>"111001001",
  37971=>"111011111",
  37972=>"000000011",
  37973=>"000000000",
  37974=>"000000100",
  37975=>"001111000",
  37976=>"000010000",
  37977=>"001011111",
  37978=>"001000000",
  37979=>"000000000",
  37980=>"111111000",
  37981=>"000001011",
  37982=>"011000111",
  37983=>"011001001",
  37984=>"000000000",
  37985=>"000000000",
  37986=>"110000111",
  37987=>"111000001",
  37988=>"001000000",
  37989=>"000000000",
  37990=>"010111100",
  37991=>"110111110",
  37992=>"000100111",
  37993=>"000011111",
  37994=>"111111000",
  37995=>"111111100",
  37996=>"001000001",
  37997=>"110000000",
  37998=>"000000000",
  37999=>"111111111",
  38000=>"011000011",
  38001=>"111010110",
  38002=>"001000000",
  38003=>"111101100",
  38004=>"111000000",
  38005=>"110110100",
  38006=>"000000000",
  38007=>"110101000",
  38008=>"110111111",
  38009=>"010110000",
  38010=>"100000000",
  38011=>"111010000",
  38012=>"000001000",
  38013=>"111111100",
  38014=>"110000000",
  38015=>"110110100",
  38016=>"001111111",
  38017=>"011110111",
  38018=>"111111111",
  38019=>"000100000",
  38020=>"000000000",
  38021=>"111000001",
  38022=>"000000111",
  38023=>"000011111",
  38024=>"111010111",
  38025=>"011000100",
  38026=>"011111111",
  38027=>"011000000",
  38028=>"111111111",
  38029=>"011111111",
  38030=>"111011001",
  38031=>"111110000",
  38032=>"000000000",
  38033=>"101000000",
  38034=>"000000011",
  38035=>"110111111",
  38036=>"000111111",
  38037=>"111111111",
  38038=>"001111111",
  38039=>"000000000",
  38040=>"000001101",
  38041=>"110110000",
  38042=>"111100100",
  38043=>"110000000",
  38044=>"010111111",
  38045=>"111100000",
  38046=>"111101000",
  38047=>"111111111",
  38048=>"111111000",
  38049=>"000000000",
  38050=>"000011001",
  38051=>"111111111",
  38052=>"000100110",
  38053=>"111111110",
  38054=>"001011000",
  38055=>"111011000",
  38056=>"001000101",
  38057=>"111111111",
  38058=>"110111111",
  38059=>"011010000",
  38060=>"000001101",
  38061=>"011011000",
  38062=>"011111111",
  38063=>"001111111",
  38064=>"000111011",
  38065=>"111111110",
  38066=>"111111000",
  38067=>"111111010",
  38068=>"000000100",
  38069=>"000001111",
  38070=>"111000000",
  38071=>"110110110",
  38072=>"001000011",
  38073=>"000111111",
  38074=>"000000000",
  38075=>"000000001",
  38076=>"011011111",
  38077=>"111111100",
  38078=>"111111111",
  38079=>"100100111",
  38080=>"001000000",
  38081=>"011110110",
  38082=>"111101101",
  38083=>"000000110",
  38084=>"111111110",
  38085=>"011111000",
  38086=>"001111111",
  38087=>"001111111",
  38088=>"000000000",
  38089=>"000000111",
  38090=>"000011111",
  38091=>"111111000",
  38092=>"011111001",
  38093=>"111111111",
  38094=>"110110111",
  38095=>"111100000",
  38096=>"000000000",
  38097=>"000000111",
  38098=>"111001011",
  38099=>"000000000",
  38100=>"000000000",
  38101=>"010011011",
  38102=>"000000010",
  38103=>"000000100",
  38104=>"111000000",
  38105=>"111111111",
  38106=>"000000000",
  38107=>"110000001",
  38108=>"101000100",
  38109=>"000000000",
  38110=>"111111010",
  38111=>"010110000",
  38112=>"000000001",
  38113=>"000000110",
  38114=>"111111000",
  38115=>"011000000",
  38116=>"110110100",
  38117=>"111001111",
  38118=>"111110000",
  38119=>"111111000",
  38120=>"000001111",
  38121=>"111101000",
  38122=>"110100000",
  38123=>"000000001",
  38124=>"101111111",
  38125=>"000000111",
  38126=>"000111111",
  38127=>"000000111",
  38128=>"100000000",
  38129=>"000000000",
  38130=>"111111111",
  38131=>"000101101",
  38132=>"111111111",
  38133=>"000111111",
  38134=>"111111000",
  38135=>"111110000",
  38136=>"111111110",
  38137=>"111111111",
  38138=>"101111000",
  38139=>"000001001",
  38140=>"111101101",
  38141=>"100000111",
  38142=>"110000000",
  38143=>"110000000",
  38144=>"000000000",
  38145=>"000000010",
  38146=>"000000000",
  38147=>"000000011",
  38148=>"111000001",
  38149=>"000000000",
  38150=>"000000001",
  38151=>"000000111",
  38152=>"100110111",
  38153=>"000000101",
  38154=>"111111111",
  38155=>"000000000",
  38156=>"101101001",
  38157=>"111111010",
  38158=>"111111110",
  38159=>"000000000",
  38160=>"100001000",
  38161=>"000000000",
  38162=>"001000001",
  38163=>"001111100",
  38164=>"110110110",
  38165=>"111001111",
  38166=>"001000001",
  38167=>"001111111",
  38168=>"111111000",
  38169=>"100000100",
  38170=>"111111000",
  38171=>"111010001",
  38172=>"000100000",
  38173=>"000001111",
  38174=>"111111111",
  38175=>"111011111",
  38176=>"100001000",
  38177=>"001111111",
  38178=>"010010011",
  38179=>"000111111",
  38180=>"000111111",
  38181=>"000000000",
  38182=>"111011011",
  38183=>"000000000",
  38184=>"111111111",
  38185=>"110110111",
  38186=>"000000011",
  38187=>"001001011",
  38188=>"111111000",
  38189=>"011001001",
  38190=>"111010111",
  38191=>"000000000",
  38192=>"111111100",
  38193=>"111110000",
  38194=>"110110111",
  38195=>"111111111",
  38196=>"111001011",
  38197=>"110110011",
  38198=>"100000000",
  38199=>"001111011",
  38200=>"000001000",
  38201=>"001001111",
  38202=>"000000110",
  38203=>"000000011",
  38204=>"011011000",
  38205=>"011101000",
  38206=>"100000000",
  38207=>"111000000",
  38208=>"000000110",
  38209=>"001000000",
  38210=>"000000000",
  38211=>"000000000",
  38212=>"011011011",
  38213=>"000001011",
  38214=>"100000000",
  38215=>"000000000",
  38216=>"111111000",
  38217=>"000000111",
  38218=>"100100111",
  38219=>"001111111",
  38220=>"110110111",
  38221=>"111111010",
  38222=>"000100110",
  38223=>"111001001",
  38224=>"111011001",
  38225=>"000100100",
  38226=>"010110010",
  38227=>"111101001",
  38228=>"000000000",
  38229=>"110100000",
  38230=>"000000011",
  38231=>"111111100",
  38232=>"111111111",
  38233=>"000111001",
  38234=>"011110110",
  38235=>"001001100",
  38236=>"000111111",
  38237=>"111111111",
  38238=>"111011000",
  38239=>"010110100",
  38240=>"110110100",
  38241=>"000000000",
  38242=>"101100000",
  38243=>"010010111",
  38244=>"111111110",
  38245=>"000011111",
  38246=>"011000110",
  38247=>"000001001",
  38248=>"000011111",
  38249=>"001000000",
  38250=>"000000111",
  38251=>"000000100",
  38252=>"111111010",
  38253=>"000011001",
  38254=>"000011001",
  38255=>"000000000",
  38256=>"000010111",
  38257=>"111000000",
  38258=>"001011111",
  38259=>"111111001",
  38260=>"110100100",
  38261=>"111101111",
  38262=>"001001000",
  38263=>"001111000",
  38264=>"111000000",
  38265=>"111000111",
  38266=>"000000110",
  38267=>"011011001",
  38268=>"100100110",
  38269=>"000000000",
  38270=>"111111111",
  38271=>"100111111",
  38272=>"000000100",
  38273=>"000000000",
  38274=>"111101111",
  38275=>"000000110",
  38276=>"111111011",
  38277=>"000010000",
  38278=>"111100100",
  38279=>"000101111",
  38280=>"000000001",
  38281=>"111100000",
  38282=>"111001111",
  38283=>"011111010",
  38284=>"001111111",
  38285=>"001011000",
  38286=>"011010000",
  38287=>"111111111",
  38288=>"000000100",
  38289=>"000000101",
  38290=>"011111010",
  38291=>"011110000",
  38292=>"111011000",
  38293=>"000000000",
  38294=>"110110000",
  38295=>"000001110",
  38296=>"111110111",
  38297=>"000000001",
  38298=>"000000011",
  38299=>"001001000",
  38300=>"000100000",
  38301=>"100000011",
  38302=>"000000000",
  38303=>"000000000",
  38304=>"100100000",
  38305=>"011111000",
  38306=>"000000000",
  38307=>"110100101",
  38308=>"111100000",
  38309=>"110000010",
  38310=>"000000001",
  38311=>"000011111",
  38312=>"111101111",
  38313=>"001100100",
  38314=>"000011011",
  38315=>"001001000",
  38316=>"111100000",
  38317=>"111011000",
  38318=>"100111111",
  38319=>"001001111",
  38320=>"000000111",
  38321=>"000000000",
  38322=>"000000000",
  38323=>"111100011",
  38324=>"000010000",
  38325=>"000000100",
  38326=>"111111111",
  38327=>"100001111",
  38328=>"010010111",
  38329=>"011011111",
  38330=>"111100110",
  38331=>"111001011",
  38332=>"001001001",
  38333=>"111010111",
  38334=>"011000001",
  38335=>"000000000",
  38336=>"000011001",
  38337=>"001001111",
  38338=>"111111111",
  38339=>"000001011",
  38340=>"010010111",
  38341=>"001000001",
  38342=>"000011010",
  38343=>"000001111",
  38344=>"000100000",
  38345=>"000000000",
  38346=>"100100111",
  38347=>"000111111",
  38348=>"111010000",
  38349=>"111011000",
  38350=>"011011011",
  38351=>"111110111",
  38352=>"000000000",
  38353=>"011011011",
  38354=>"111111111",
  38355=>"011000010",
  38356=>"100111111",
  38357=>"100100100",
  38358=>"111111111",
  38359=>"001101111",
  38360=>"000111000",
  38361=>"111000100",
  38362=>"001001111",
  38363=>"111001000",
  38364=>"110111111",
  38365=>"111111111",
  38366=>"111111000",
  38367=>"000000000",
  38368=>"001000011",
  38369=>"111111011",
  38370=>"101001000",
  38371=>"000000100",
  38372=>"111111111",
  38373=>"111110000",
  38374=>"111111001",
  38375=>"111100100",
  38376=>"001000000",
  38377=>"011001000",
  38378=>"011001000",
  38379=>"111110000",
  38380=>"111111110",
  38381=>"101111111",
  38382=>"000001001",
  38383=>"001011111",
  38384=>"000000000",
  38385=>"001011011",
  38386=>"000000000",
  38387=>"000010111",
  38388=>"000000101",
  38389=>"111111110",
  38390=>"011111111",
  38391=>"010011111",
  38392=>"011001010",
  38393=>"001001101",
  38394=>"110001011",
  38395=>"000001011",
  38396=>"000001111",
  38397=>"000000011",
  38398=>"011111110",
  38399=>"111111111",
  38400=>"111111111",
  38401=>"001001001",
  38402=>"000000000",
  38403=>"111111011",
  38404=>"000000000",
  38405=>"000000000",
  38406=>"110110110",
  38407=>"011111111",
  38408=>"000000000",
  38409=>"111110111",
  38410=>"011111111",
  38411=>"111100101",
  38412=>"011011001",
  38413=>"111111111",
  38414=>"100000001",
  38415=>"111111111",
  38416=>"000000100",
  38417=>"111111100",
  38418=>"100111111",
  38419=>"000111111",
  38420=>"111100011",
  38421=>"001001100",
  38422=>"111111111",
  38423=>"111100000",
  38424=>"000010011",
  38425=>"110111011",
  38426=>"000000111",
  38427=>"100100111",
  38428=>"000000000",
  38429=>"010000000",
  38430=>"001111111",
  38431=>"011011000",
  38432=>"000000100",
  38433=>"000111111",
  38434=>"111111111",
  38435=>"000000000",
  38436=>"001001000",
  38437=>"111111111",
  38438=>"111001111",
  38439=>"111111100",
  38440=>"101111110",
  38441=>"000000100",
  38442=>"000000000",
  38443=>"100100110",
  38444=>"111111110",
  38445=>"000000000",
  38446=>"001001111",
  38447=>"111111100",
  38448=>"100110111",
  38449=>"110000000",
  38450=>"110111011",
  38451=>"110000000",
  38452=>"011001000",
  38453=>"111011001",
  38454=>"001100100",
  38455=>"000000000",
  38456=>"101001101",
  38457=>"100000110",
  38458=>"111111011",
  38459=>"010111111",
  38460=>"000000000",
  38461=>"000000111",
  38462=>"000001001",
  38463=>"000001001",
  38464=>"000000000",
  38465=>"111111100",
  38466=>"101000000",
  38467=>"100100111",
  38468=>"001001011",
  38469=>"011111110",
  38470=>"000100000",
  38471=>"111111111",
  38472=>"111000000",
  38473=>"110001001",
  38474=>"111111111",
  38475=>"101100100",
  38476=>"111111111",
  38477=>"111000000",
  38478=>"110000000",
  38479=>"000000000",
  38480=>"001101000",
  38481=>"000000000",
  38482=>"000000111",
  38483=>"000110111",
  38484=>"110111111",
  38485=>"110100000",
  38486=>"101101000",
  38487=>"100000110",
  38488=>"000000000",
  38489=>"011000011",
  38490=>"011010000",
  38491=>"111100000",
  38492=>"111111111",
  38493=>"111111111",
  38494=>"000000000",
  38495=>"111111011",
  38496=>"000000000",
  38497=>"100100001",
  38498=>"111111101",
  38499=>"000000000",
  38500=>"000110100",
  38501=>"001001000",
  38502=>"111111011",
  38503=>"000110111",
  38504=>"011001000",
  38505=>"000111111",
  38506=>"111110100",
  38507=>"011011000",
  38508=>"101100100",
  38509=>"000000000",
  38510=>"000000000",
  38511=>"111111110",
  38512=>"111111101",
  38513=>"101001011",
  38514=>"111111110",
  38515=>"000000000",
  38516=>"000000100",
  38517=>"011011111",
  38518=>"101111111",
  38519=>"000001011",
  38520=>"000000000",
  38521=>"111111111",
  38522=>"000001111",
  38523=>"100111111",
  38524=>"001001101",
  38525=>"111110101",
  38526=>"000000111",
  38527=>"000000101",
  38528=>"000000001",
  38529=>"100000000",
  38530=>"111000000",
  38531=>"111001001",
  38532=>"000100000",
  38533=>"010010110",
  38534=>"100111100",
  38535=>"000111011",
  38536=>"111001001",
  38537=>"000000000",
  38538=>"000000111",
  38539=>"000100111",
  38540=>"000000000",
  38541=>"000000000",
  38542=>"101000011",
  38543=>"000000010",
  38544=>"111111111",
  38545=>"010000110",
  38546=>"111111000",
  38547=>"000101111",
  38548=>"110000010",
  38549=>"110110000",
  38550=>"111111000",
  38551=>"000000000",
  38552=>"000000000",
  38553=>"000110111",
  38554=>"111111111",
  38555=>"110111011",
  38556=>"011000000",
  38557=>"001000000",
  38558=>"100100111",
  38559=>"111000100",
  38560=>"111111111",
  38561=>"111100000",
  38562=>"100111011",
  38563=>"110111111",
  38564=>"011111111",
  38565=>"011111000",
  38566=>"110110111",
  38567=>"100100000",
  38568=>"000100111",
  38569=>"000000000",
  38570=>"000000000",
  38571=>"101111001",
  38572=>"001111101",
  38573=>"111001001",
  38574=>"000000000",
  38575=>"100111001",
  38576=>"000111000",
  38577=>"001001011",
  38578=>"111111100",
  38579=>"111101101",
  38580=>"111111000",
  38581=>"000000000",
  38582=>"000001111",
  38583=>"000000000",
  38584=>"000000000",
  38585=>"111000000",
  38586=>"000000100",
  38587=>"011111110",
  38588=>"111111111",
  38589=>"000000000",
  38590=>"101111000",
  38591=>"000110111",
  38592=>"111111111",
  38593=>"100100100",
  38594=>"111111111",
  38595=>"000000000",
  38596=>"111111001",
  38597=>"111111111",
  38598=>"000100000",
  38599=>"111111101",
  38600=>"011111110",
  38601=>"101001111",
  38602=>"100000011",
  38603=>"111111111",
  38604=>"111100111",
  38605=>"000110111",
  38606=>"000111111",
  38607=>"000000000",
  38608=>"000000000",
  38609=>"010001000",
  38610=>"000000000",
  38611=>"000000000",
  38612=>"101111000",
  38613=>"000011111",
  38614=>"011011111",
  38615=>"100000000",
  38616=>"000000111",
  38617=>"100000000",
  38618=>"111111111",
  38619=>"110000000",
  38620=>"000110100",
  38621=>"101001000",
  38622=>"000000000",
  38623=>"001000000",
  38624=>"000000000",
  38625=>"000000110",
  38626=>"111111111",
  38627=>"000000110",
  38628=>"001000000",
  38629=>"010001001",
  38630=>"111000111",
  38631=>"000000000",
  38632=>"110100100",
  38633=>"000000111",
  38634=>"000100111",
  38635=>"001000010",
  38636=>"000010110",
  38637=>"111111010",
  38638=>"100111111",
  38639=>"000000000",
  38640=>"000111100",
  38641=>"111111111",
  38642=>"111111111",
  38643=>"101000100",
  38644=>"111100000",
  38645=>"111110100",
  38646=>"011000000",
  38647=>"000000000",
  38648=>"000000000",
  38649=>"000000000",
  38650=>"010110010",
  38651=>"000000000",
  38652=>"110010111",
  38653=>"001001001",
  38654=>"000001111",
  38655=>"000000000",
  38656=>"000000101",
  38657=>"001000001",
  38658=>"000000000",
  38659=>"111111000",
  38660=>"111101000",
  38661=>"101101100",
  38662=>"100111111",
  38663=>"111111011",
  38664=>"000000100",
  38665=>"101001001",
  38666=>"100101001",
  38667=>"001000000",
  38668=>"100000110",
  38669=>"100000111",
  38670=>"111111111",
  38671=>"111111000",
  38672=>"100101001",
  38673=>"100111111",
  38674=>"000000000",
  38675=>"111111111",
  38676=>"100000000",
  38677=>"100000000",
  38678=>"001001001",
  38679=>"111111100",
  38680=>"000000000",
  38681=>"111000000",
  38682=>"111001111",
  38683=>"000000000",
  38684=>"011011111",
  38685=>"000010010",
  38686=>"111000000",
  38687=>"111101111",
  38688=>"110011011",
  38689=>"101101111",
  38690=>"110111010",
  38691=>"110110011",
  38692=>"000000000",
  38693=>"000101111",
  38694=>"110111000",
  38695=>"000000000",
  38696=>"000010110",
  38697=>"000000111",
  38698=>"101100111",
  38699=>"111000011",
  38700=>"111111110",
  38701=>"001000000",
  38702=>"111111000",
  38703=>"011000000",
  38704=>"100111111",
  38705=>"000100111",
  38706=>"100100110",
  38707=>"011011110",
  38708=>"000000000",
  38709=>"111000000",
  38710=>"000111111",
  38711=>"000000000",
  38712=>"010000000",
  38713=>"000000111",
  38714=>"110110111",
  38715=>"000000110",
  38716=>"000100100",
  38717=>"000111000",
  38718=>"111101111",
  38719=>"000001111",
  38720=>"111111001",
  38721=>"111111100",
  38722=>"000001000",
  38723=>"111110000",
  38724=>"101011101",
  38725=>"000110010",
  38726=>"100000000",
  38727=>"000000001",
  38728=>"000000000",
  38729=>"111001001",
  38730=>"001000001",
  38731=>"111111000",
  38732=>"010110000",
  38733=>"011010000",
  38734=>"000000000",
  38735=>"011011011",
  38736=>"000010001",
  38737=>"111001111",
  38738=>"101111011",
  38739=>"001111111",
  38740=>"000101001",
  38741=>"000011011",
  38742=>"111001000",
  38743=>"000000000",
  38744=>"000000101",
  38745=>"000000000",
  38746=>"000000000",
  38747=>"000100111",
  38748=>"111111111",
  38749=>"000000000",
  38750=>"111101111",
  38751=>"011111000",
  38752=>"111011011",
  38753=>"000000000",
  38754=>"000111111",
  38755=>"111111111",
  38756=>"111001000",
  38757=>"001100000",
  38758=>"110110010",
  38759=>"001001111",
  38760=>"001101101",
  38761=>"011111010",
  38762=>"000001001",
  38763=>"001001000",
  38764=>"011011011",
  38765=>"000001101",
  38766=>"110000000",
  38767=>"000000111",
  38768=>"011011101",
  38769=>"111111001",
  38770=>"101111111",
  38771=>"110111111",
  38772=>"000000000",
  38773=>"100000000",
  38774=>"001011001",
  38775=>"011010000",
  38776=>"000000000",
  38777=>"111011011",
  38778=>"000000000",
  38779=>"111111111",
  38780=>"111111111",
  38781=>"001000111",
  38782=>"111100111",
  38783=>"000000110",
  38784=>"111111111",
  38785=>"100000001",
  38786=>"111001001",
  38787=>"001000000",
  38788=>"000111111",
  38789=>"000000000",
  38790=>"000000000",
  38791=>"111111111",
  38792=>"111101000",
  38793=>"001000000",
  38794=>"000000000",
  38795=>"000000111",
  38796=>"101000011",
  38797=>"001011111",
  38798=>"101000000",
  38799=>"000000000",
  38800=>"000001011",
  38801=>"111111111",
  38802=>"000000011",
  38803=>"000000000",
  38804=>"111111111",
  38805=>"010010011",
  38806=>"000000000",
  38807=>"000001101",
  38808=>"111111011",
  38809=>"111111111",
  38810=>"100111111",
  38811=>"011011111",
  38812=>"111101111",
  38813=>"101111111",
  38814=>"111111110",
  38815=>"110110111",
  38816=>"111110110",
  38817=>"100100000",
  38818=>"111101111",
  38819=>"011111111",
  38820=>"000001111",
  38821=>"110111111",
  38822=>"000000000",
  38823=>"111111100",
  38824=>"111111111",
  38825=>"000000111",
  38826=>"111000000",
  38827=>"111101100",
  38828=>"000000000",
  38829=>"111000000",
  38830=>"011111001",
  38831=>"000000100",
  38832=>"111111111",
  38833=>"000001001",
  38834=>"000000000",
  38835=>"100100111",
  38836=>"000000100",
  38837=>"101100000",
  38838=>"000110101",
  38839=>"001001001",
  38840=>"000000011",
  38841=>"111100101",
  38842=>"100000000",
  38843=>"101000000",
  38844=>"000000000",
  38845=>"101100101",
  38846=>"111111000",
  38847=>"011001001",
  38848=>"100111111",
  38849=>"000000000",
  38850=>"111011000",
  38851=>"000000000",
  38852=>"111101111",
  38853=>"111000000",
  38854=>"100000000",
  38855=>"010000000",
  38856=>"000000000",
  38857=>"000100100",
  38858=>"010000111",
  38859=>"000000111",
  38860=>"000000000",
  38861=>"000000000",
  38862=>"011101001",
  38863=>"100000010",
  38864=>"000001000",
  38865=>"111000000",
  38866=>"000000100",
  38867=>"111111111",
  38868=>"000000001",
  38869=>"000000111",
  38870=>"111000100",
  38871=>"111111000",
  38872=>"100000000",
  38873=>"100000100",
  38874=>"001000000",
  38875=>"111111111",
  38876=>"111111100",
  38877=>"110110000",
  38878=>"111111111",
  38879=>"111111111",
  38880=>"111111000",
  38881=>"111110110",
  38882=>"111011111",
  38883=>"100000000",
  38884=>"001101111",
  38885=>"011111000",
  38886=>"100000000",
  38887=>"111111111",
  38888=>"111001111",
  38889=>"111111000",
  38890=>"000000000",
  38891=>"000000001",
  38892=>"111001000",
  38893=>"100100000",
  38894=>"111001000",
  38895=>"111111111",
  38896=>"010010000",
  38897=>"111111111",
  38898=>"000000001",
  38899=>"111100000",
  38900=>"000000000",
  38901=>"000000000",
  38902=>"000111011",
  38903=>"000000000",
  38904=>"000011111",
  38905=>"000111010",
  38906=>"110100000",
  38907=>"111111111",
  38908=>"011001000",
  38909=>"000000000",
  38910=>"000000001",
  38911=>"000000000",
  38912=>"000001001",
  38913=>"000000000",
  38914=>"000000000",
  38915=>"000001000",
  38916=>"000000000",
  38917=>"011011000",
  38918=>"111111011",
  38919=>"111111111",
  38920=>"111111111",
  38921=>"000000000",
  38922=>"000111111",
  38923=>"011011001",
  38924=>"001111100",
  38925=>"111111111",
  38926=>"111001000",
  38927=>"001001000",
  38928=>"110111111",
  38929=>"000011011",
  38930=>"000000000",
  38931=>"000101111",
  38932=>"111111111",
  38933=>"000000111",
  38934=>"000000000",
  38935=>"100100100",
  38936=>"100000110",
  38937=>"111111101",
  38938=>"111101111",
  38939=>"111110000",
  38940=>"100100100",
  38941=>"011111111",
  38942=>"000111110",
  38943=>"000000111",
  38944=>"000000001",
  38945=>"010110000",
  38946=>"000000000",
  38947=>"111000111",
  38948=>"111101111",
  38949=>"111011000",
  38950=>"111111000",
  38951=>"100110000",
  38952=>"100110110",
  38953=>"111111111",
  38954=>"111111111",
  38955=>"111111111",
  38956=>"111111111",
  38957=>"001001000",
  38958=>"111111111",
  38959=>"001001001",
  38960=>"111011000",
  38961=>"111111111",
  38962=>"100100000",
  38963=>"001001000",
  38964=>"100111111",
  38965=>"010100100",
  38966=>"000000100",
  38967=>"001000100",
  38968=>"100000000",
  38969=>"111111000",
  38970=>"111111111",
  38971=>"000000001",
  38972=>"111011111",
  38973=>"000000000",
  38974=>"011111111",
  38975=>"000000111",
  38976=>"111111111",
  38977=>"111001000",
  38978=>"111111111",
  38979=>"111000100",
  38980=>"000000000",
  38981=>"011011111",
  38982=>"111000100",
  38983=>"000000000",
  38984=>"000000100",
  38985=>"000000000",
  38986=>"000000000",
  38987=>"000000111",
  38988=>"000001111",
  38989=>"000100000",
  38990=>"011000000",
  38991=>"000000000",
  38992=>"010000100",
  38993=>"010010000",
  38994=>"000000000",
  38995=>"111111111",
  38996=>"000111111",
  38997=>"110111000",
  38998=>"111110100",
  38999=>"110100111",
  39000=>"000110100",
  39001=>"111000000",
  39002=>"000000000",
  39003=>"100000100",
  39004=>"000000000",
  39005=>"000000000",
  39006=>"100111111",
  39007=>"111111000",
  39008=>"111111111",
  39009=>"000000000",
  39010=>"111011000",
  39011=>"011011010",
  39012=>"111000011",
  39013=>"110100000",
  39014=>"110111110",
  39015=>"001001001",
  39016=>"000100000",
  39017=>"010111111",
  39018=>"001001111",
  39019=>"010000000",
  39020=>"111111011",
  39021=>"001111111",
  39022=>"001111111",
  39023=>"000000000",
  39024=>"001000000",
  39025=>"000100100",
  39026=>"101100100",
  39027=>"010111111",
  39028=>"010100000",
  39029=>"101110110",
  39030=>"000000000",
  39031=>"000111111",
  39032=>"010010100",
  39033=>"100000000",
  39034=>"011011000",
  39035=>"111111111",
  39036=>"110110000",
  39037=>"111111111",
  39038=>"000000000",
  39039=>"011011001",
  39040=>"111111111",
  39041=>"000111111",
  39042=>"000000000",
  39043=>"111100110",
  39044=>"000000111",
  39045=>"000000001",
  39046=>"111000000",
  39047=>"111001000",
  39048=>"111111111",
  39049=>"111001000",
  39050=>"111111111",
  39051=>"111111111",
  39052=>"111101111",
  39053=>"111111111",
  39054=>"111110111",
  39055=>"011110000",
  39056=>"111000001",
  39057=>"000000000",
  39058=>"000100000",
  39059=>"001000000",
  39060=>"000000100",
  39061=>"110000000",
  39062=>"001001000",
  39063=>"111111000",
  39064=>"100000000",
  39065=>"111110111",
  39066=>"000000000",
  39067=>"000100000",
  39068=>"010000000",
  39069=>"001000000",
  39070=>"101101111",
  39071=>"111111110",
  39072=>"011011111",
  39073=>"111001001",
  39074=>"000000000",
  39075=>"000000000",
  39076=>"000011110",
  39077=>"000111111",
  39078=>"000000000",
  39079=>"011111111",
  39080=>"000000000",
  39081=>"011001111",
  39082=>"000000000",
  39083=>"010000000",
  39084=>"010011111",
  39085=>"100100100",
  39086=>"111111111",
  39087=>"000000000",
  39088=>"111111000",
  39089=>"110110111",
  39090=>"011111111",
  39091=>"000000000",
  39092=>"111000010",
  39093=>"111111100",
  39094=>"000001101",
  39095=>"000010000",
  39096=>"000000100",
  39097=>"111111000",
  39098=>"001111111",
  39099=>"000011000",
  39100=>"110001001",
  39101=>"100000010",
  39102=>"111110110",
  39103=>"001111111",
  39104=>"000000000",
  39105=>"001100101",
  39106=>"000000000",
  39107=>"000111110",
  39108=>"001011011",
  39109=>"001001000",
  39110=>"100000010",
  39111=>"000001111",
  39112=>"000000101",
  39113=>"111111110",
  39114=>"000000000",
  39115=>"000000000",
  39116=>"100000100",
  39117=>"000000000",
  39118=>"001000000",
  39119=>"001111100",
  39120=>"000010000",
  39121=>"110000000",
  39122=>"111111000",
  39123=>"111010000",
  39124=>"000000111",
  39125=>"111111111",
  39126=>"101000000",
  39127=>"001000000",
  39128=>"000011111",
  39129=>"111100000",
  39130=>"011001011",
  39131=>"111101000",
  39132=>"111111111",
  39133=>"000000000",
  39134=>"000000000",
  39135=>"111100000",
  39136=>"010111000",
  39137=>"000000000",
  39138=>"000000000",
  39139=>"011001001",
  39140=>"111111111",
  39141=>"011111111",
  39142=>"100111111",
  39143=>"111110111",
  39144=>"000000000",
  39145=>"111011001",
  39146=>"111111000",
  39147=>"001000000",
  39148=>"000000001",
  39149=>"000000000",
  39150=>"000010000",
  39151=>"000010000",
  39152=>"101100100",
  39153=>"111110110",
  39154=>"111101000",
  39155=>"000001001",
  39156=>"000000000",
  39157=>"110100000",
  39158=>"000110110",
  39159=>"011111000",
  39160=>"001000000",
  39161=>"000000000",
  39162=>"000100100",
  39163=>"111011011",
  39164=>"111011011",
  39165=>"001000000",
  39166=>"000000000",
  39167=>"010010010",
  39168=>"000000000",
  39169=>"110101100",
  39170=>"000000000",
  39171=>"000000000",
  39172=>"111111111",
  39173=>"000000000",
  39174=>"110110100",
  39175=>"101100100",
  39176=>"011011000",
  39177=>"000000000",
  39178=>"000000000",
  39179=>"000000100",
  39180=>"111111111",
  39181=>"000000000",
  39182=>"111111111",
  39183=>"000000101",
  39184=>"100110111",
  39185=>"000000000",
  39186=>"111101111",
  39187=>"000000000",
  39188=>"000000001",
  39189=>"000000000",
  39190=>"110101111",
  39191=>"101111100",
  39192=>"100001100",
  39193=>"111111111",
  39194=>"111111111",
  39195=>"000000000",
  39196=>"000110111",
  39197=>"000000000",
  39198=>"010010000",
  39199=>"000100111",
  39200=>"000000000",
  39201=>"011011011",
  39202=>"000000000",
  39203=>"000100110",
  39204=>"110000010",
  39205=>"011111111",
  39206=>"011011001",
  39207=>"000000000",
  39208=>"111111111",
  39209=>"000000001",
  39210=>"100100000",
  39211=>"000000000",
  39212=>"000100100",
  39213=>"000100101",
  39214=>"111000000",
  39215=>"000001000",
  39216=>"000000001",
  39217=>"000000000",
  39218=>"111111000",
  39219=>"110110111",
  39220=>"000000000",
  39221=>"000100111",
  39222=>"000110100",
  39223=>"000111111",
  39224=>"100111111",
  39225=>"100000000",
  39226=>"111111110",
  39227=>"111111111",
  39228=>"111111110",
  39229=>"000000001",
  39230=>"101000000",
  39231=>"011111111",
  39232=>"111111111",
  39233=>"000000000",
  39234=>"111110111",
  39235=>"110110111",
  39236=>"100100101",
  39237=>"000110100",
  39238=>"110111111",
  39239=>"111001000",
  39240=>"001000000",
  39241=>"000000000",
  39242=>"111001000",
  39243=>"000110110",
  39244=>"011010000",
  39245=>"000000000",
  39246=>"111000000",
  39247=>"111111111",
  39248=>"011111001",
  39249=>"100100110",
  39250=>"101001100",
  39251=>"000000000",
  39252=>"000000000",
  39253=>"011011001",
  39254=>"000000000",
  39255=>"111111100",
  39256=>"111111011",
  39257=>"000000000",
  39258=>"111111111",
  39259=>"000000000",
  39260=>"000000001",
  39261=>"001000000",
  39262=>"011011001",
  39263=>"110100101",
  39264=>"111001000",
  39265=>"111111111",
  39266=>"111111111",
  39267=>"111110000",
  39268=>"011011011",
  39269=>"000000000",
  39270=>"000000000",
  39271=>"111110000",
  39272=>"011001111",
  39273=>"000000000",
  39274=>"111111011",
  39275=>"111111000",
  39276=>"000000000",
  39277=>"000000001",
  39278=>"000011010",
  39279=>"111111100",
  39280=>"000000000",
  39281=>"011011001",
  39282=>"001111111",
  39283=>"110111001",
  39284=>"010000000",
  39285=>"010010000",
  39286=>"000000000",
  39287=>"000000100",
  39288=>"111111111",
  39289=>"000000000",
  39290=>"111111101",
  39291=>"110111011",
  39292=>"001111111",
  39293=>"111101110",
  39294=>"000000000",
  39295=>"111111111",
  39296=>"001001100",
  39297=>"000000110",
  39298=>"000000001",
  39299=>"111111111",
  39300=>"111111111",
  39301=>"000000000",
  39302=>"111111111",
  39303=>"111010000",
  39304=>"111001001",
  39305=>"000111000",
  39306=>"000000000",
  39307=>"000000000",
  39308=>"111100000",
  39309=>"111111111",
  39310=>"000100100",
  39311=>"000010011",
  39312=>"000100000",
  39313=>"010000000",
  39314=>"000000000",
  39315=>"000000001",
  39316=>"111111111",
  39317=>"000000000",
  39318=>"001000110",
  39319=>"111111110",
  39320=>"000111011",
  39321=>"010111110",
  39322=>"111101111",
  39323=>"000000000",
  39324=>"111001001",
  39325=>"011001001",
  39326=>"100000111",
  39327=>"111111111",
  39328=>"000000000",
  39329=>"001010111",
  39330=>"000100110",
  39331=>"111110111",
  39332=>"001000111",
  39333=>"000000000",
  39334=>"000000111",
  39335=>"100100100",
  39336=>"111111010",
  39337=>"110100100",
  39338=>"000000001",
  39339=>"101001000",
  39340=>"000000000",
  39341=>"000000000",
  39342=>"011001000",
  39343=>"001011111",
  39344=>"111111111",
  39345=>"001111111",
  39346=>"000100001",
  39347=>"000000000",
  39348=>"000000000",
  39349=>"111011111",
  39350=>"110000111",
  39351=>"111111111",
  39352=>"111111111",
  39353=>"000000000",
  39354=>"001000000",
  39355=>"111111111",
  39356=>"110111111",
  39357=>"000000110",
  39358=>"000111111",
  39359=>"100111110",
  39360=>"111000000",
  39361=>"111111001",
  39362=>"111111111",
  39363=>"100110000",
  39364=>"100100111",
  39365=>"001011111",
  39366=>"001011111",
  39367=>"001001111",
  39368=>"011001000",
  39369=>"111111110",
  39370=>"001001100",
  39371=>"000000000",
  39372=>"111111000",
  39373=>"000000000",
  39374=>"010100100",
  39375=>"000100000",
  39376=>"110010000",
  39377=>"000000000",
  39378=>"000000000",
  39379=>"111111111",
  39380=>"111111111",
  39381=>"011001001",
  39382=>"001000000",
  39383=>"000000000",
  39384=>"111101111",
  39385=>"100100100",
  39386=>"111111001",
  39387=>"000000000",
  39388=>"001111111",
  39389=>"001001000",
  39390=>"000000110",
  39391=>"111110100",
  39392=>"111011011",
  39393=>"111111110",
  39394=>"111111111",
  39395=>"011001111",
  39396=>"000001000",
  39397=>"000000111",
  39398=>"011111001",
  39399=>"000000000",
  39400=>"101001001",
  39401=>"000000110",
  39402=>"110000000",
  39403=>"111111111",
  39404=>"000000111",
  39405=>"111111111",
  39406=>"000000111",
  39407=>"011001101",
  39408=>"111111111",
  39409=>"000000000",
  39410=>"111111111",
  39411=>"111111111",
  39412=>"000000000",
  39413=>"100000110",
  39414=>"111111010",
  39415=>"000000010",
  39416=>"010111111",
  39417=>"001111111",
  39418=>"001000000",
  39419=>"000000111",
  39420=>"000000000",
  39421=>"111111111",
  39422=>"111111111",
  39423=>"001001001",
  39424=>"100000000",
  39425=>"011110110",
  39426=>"000000000",
  39427=>"111111111",
  39428=>"000000011",
  39429=>"111111000",
  39430=>"000000000",
  39431=>"111110111",
  39432=>"000000010",
  39433=>"111000000",
  39434=>"001001000",
  39435=>"000000111",
  39436=>"000000000",
  39437=>"100000000",
  39438=>"000000000",
  39439=>"001001001",
  39440=>"011000011",
  39441=>"111111111",
  39442=>"111110000",
  39443=>"111011011",
  39444=>"000011111",
  39445=>"000000000",
  39446=>"000000000",
  39447=>"111011000",
  39448=>"000111111",
  39449=>"000011000",
  39450=>"000000000",
  39451=>"001100100",
  39452=>"000000000",
  39453=>"000000101",
  39454=>"000000011",
  39455=>"111111111",
  39456=>"111111110",
  39457=>"101100101",
  39458=>"000000000",
  39459=>"110111111",
  39460=>"000111111",
  39461=>"111110000",
  39462=>"011111111",
  39463=>"111111111",
  39464=>"000000111",
  39465=>"000000000",
  39466=>"000000010",
  39467=>"001111111",
  39468=>"001001101",
  39469=>"000000000",
  39470=>"001111011",
  39471=>"111000000",
  39472=>"000000100",
  39473=>"001000000",
  39474=>"000000000",
  39475=>"000111111",
  39476=>"111001011",
  39477=>"111111011",
  39478=>"100000000",
  39479=>"111001000",
  39480=>"101101111",
  39481=>"000000111",
  39482=>"000000000",
  39483=>"111111111",
  39484=>"100000000",
  39485=>"111110111",
  39486=>"111111111",
  39487=>"000000000",
  39488=>"001111111",
  39489=>"110010010",
  39490=>"001011001",
  39491=>"001000100",
  39492=>"011111111",
  39493=>"000011110",
  39494=>"011000000",
  39495=>"100111111",
  39496=>"011011101",
  39497=>"111111111",
  39498=>"000110111",
  39499=>"111111101",
  39500=>"001001111",
  39501=>"111111111",
  39502=>"000100000",
  39503=>"101000000",
  39504=>"000000000",
  39505=>"011001011",
  39506=>"000000110",
  39507=>"100000000",
  39508=>"100000000",
  39509=>"000100111",
  39510=>"000000001",
  39511=>"000000000",
  39512=>"101000000",
  39513=>"111001101",
  39514=>"111111110",
  39515=>"001000011",
  39516=>"100000000",
  39517=>"100110111",
  39518=>"101100001",
  39519=>"000000000",
  39520=>"000001111",
  39521=>"000100111",
  39522=>"000010100",
  39523=>"000000111",
  39524=>"000000000",
  39525=>"000000000",
  39526=>"111111111",
  39527=>"000000100",
  39528=>"011011011",
  39529=>"000000110",
  39530=>"000000011",
  39531=>"110110000",
  39532=>"100100100",
  39533=>"111111000",
  39534=>"111111100",
  39535=>"111111111",
  39536=>"111110000",
  39537=>"000001001",
  39538=>"111011011",
  39539=>"000000001",
  39540=>"111111111",
  39541=>"000100111",
  39542=>"000000111",
  39543=>"001011011",
  39544=>"100101000",
  39545=>"001111101",
  39546=>"111110100",
  39547=>"000000000",
  39548=>"111001010",
  39549=>"111111111",
  39550=>"100100100",
  39551=>"111000000",
  39552=>"000000000",
  39553=>"011010111",
  39554=>"111111101",
  39555=>"110110001",
  39556=>"111111011",
  39557=>"000000100",
  39558=>"000000011",
  39559=>"000000100",
  39560=>"000110111",
  39561=>"011001001",
  39562=>"000000000",
  39563=>"000000000",
  39564=>"000000000",
  39565=>"001011000",
  39566=>"111111111",
  39567=>"000000000",
  39568=>"000110111",
  39569=>"101000000",
  39570=>"000100000",
  39571=>"011111011",
  39572=>"100100100",
  39573=>"111111111",
  39574=>"000000000",
  39575=>"011000000",
  39576=>"111111000",
  39577=>"111111111",
  39578=>"000000000",
  39579=>"001010000",
  39580=>"111111111",
  39581=>"111111001",
  39582=>"000000000",
  39583=>"000000000",
  39584=>"111000000",
  39585=>"000000000",
  39586=>"000110111",
  39587=>"000000000",
  39588=>"111001000",
  39589=>"000000110",
  39590=>"100100000",
  39591=>"111111000",
  39592=>"010110111",
  39593=>"100000000",
  39594=>"001000000",
  39595=>"101111111",
  39596=>"000001001",
  39597=>"111100000",
  39598=>"111110111",
  39599=>"111111000",
  39600=>"000000000",
  39601=>"000001011",
  39602=>"001001111",
  39603=>"111111000",
  39604=>"000000000",
  39605=>"111001001",
  39606=>"111111111",
  39607=>"011000000",
  39608=>"110111101",
  39609=>"000000000",
  39610=>"111000000",
  39611=>"011111011",
  39612=>"000000110",
  39613=>"111111111",
  39614=>"111111111",
  39615=>"000111111",
  39616=>"001111111",
  39617=>"111111111",
  39618=>"000000010",
  39619=>"000000000",
  39620=>"000001111",
  39621=>"111100000",
  39622=>"100000000",
  39623=>"001001000",
  39624=>"000000111",
  39625=>"000000000",
  39626=>"010000000",
  39627=>"111101100",
  39628=>"100110100",
  39629=>"000000000",
  39630=>"000000111",
  39631=>"110100100",
  39632=>"000000100",
  39633=>"000000000",
  39634=>"111111101",
  39635=>"111000000",
  39636=>"000001001",
  39637=>"001111111",
  39638=>"111111011",
  39639=>"111111111",
  39640=>"100100111",
  39641=>"000000011",
  39642=>"000001111",
  39643=>"111100100",
  39644=>"001001101",
  39645=>"000000000",
  39646=>"110100111",
  39647=>"111000000",
  39648=>"000000000",
  39649=>"000000010",
  39650=>"011110010",
  39651=>"011111111",
  39652=>"000000000",
  39653=>"000000010",
  39654=>"110000000",
  39655=>"111110000",
  39656=>"111110110",
  39657=>"111110111",
  39658=>"111110111",
  39659=>"001000000",
  39660=>"000000000",
  39661=>"010000000",
  39662=>"000011111",
  39663=>"000000000",
  39664=>"000000000",
  39665=>"111111111",
  39666=>"000000111",
  39667=>"000101111",
  39668=>"010011111",
  39669=>"000000000",
  39670=>"111111111",
  39671=>"011011111",
  39672=>"110000000",
  39673=>"111111111",
  39674=>"111111111",
  39675=>"000000111",
  39676=>"110110111",
  39677=>"001001001",
  39678=>"000000001",
  39679=>"111111111",
  39680=>"000001001",
  39681=>"001001000",
  39682=>"111111110",
  39683=>"101000000",
  39684=>"000011111",
  39685=>"101011000",
  39686=>"000000000",
  39687=>"111111111",
  39688=>"001000100",
  39689=>"011111111",
  39690=>"001111111",
  39691=>"000000000",
  39692=>"001000101",
  39693=>"010000011",
  39694=>"000000100",
  39695=>"111111111",
  39696=>"000000000",
  39697=>"000000000",
  39698=>"000001001",
  39699=>"000000000",
  39700=>"111000000",
  39701=>"000000000",
  39702=>"000100100",
  39703=>"111111000",
  39704=>"000001011",
  39705=>"111111111",
  39706=>"000000000",
  39707=>"111111111",
  39708=>"001001001",
  39709=>"000110111",
  39710=>"000000000",
  39711=>"111100000",
  39712=>"100100000",
  39713=>"111111111",
  39714=>"100111000",
  39715=>"111111111",
  39716=>"111111011",
  39717=>"000000111",
  39718=>"000000000",
  39719=>"111111111",
  39720=>"111100000",
  39721=>"110111111",
  39722=>"000000000",
  39723=>"111000000",
  39724=>"000000000",
  39725=>"100000000",
  39726=>"000000000",
  39727=>"000000000",
  39728=>"111111011",
  39729=>"000000100",
  39730=>"000000001",
  39731=>"100000000",
  39732=>"000000000",
  39733=>"111100000",
  39734=>"101111111",
  39735=>"000000000",
  39736=>"111111000",
  39737=>"111111000",
  39738=>"111100000",
  39739=>"111111111",
  39740=>"101111000",
  39741=>"111100111",
  39742=>"000001001",
  39743=>"111011000",
  39744=>"000000000",
  39745=>"011001100",
  39746=>"000000000",
  39747=>"000000000",
  39748=>"000001000",
  39749=>"001001101",
  39750=>"110000000",
  39751=>"111111111",
  39752=>"001001000",
  39753=>"111001000",
  39754=>"000110111",
  39755=>"110111010",
  39756=>"100111111",
  39757=>"000001011",
  39758=>"000000000",
  39759=>"110110110",
  39760=>"100110111",
  39761=>"011000111",
  39762=>"000000000",
  39763=>"111111000",
  39764=>"111001000",
  39765=>"111111011",
  39766=>"000100010",
  39767=>"111111111",
  39768=>"000000000",
  39769=>"111111110",
  39770=>"000000001",
  39771=>"001101000",
  39772=>"110111110",
  39773=>"111111111",
  39774=>"101111011",
  39775=>"111111111",
  39776=>"110111111",
  39777=>"000101111",
  39778=>"000011111",
  39779=>"011111111",
  39780=>"001000000",
  39781=>"000000000",
  39782=>"000000000",
  39783=>"001000111",
  39784=>"111111111",
  39785=>"110110100",
  39786=>"000000000",
  39787=>"011111111",
  39788=>"000000001",
  39789=>"000000000",
  39790=>"000000111",
  39791=>"000001000",
  39792=>"000000000",
  39793=>"000000000",
  39794=>"111010111",
  39795=>"000111110",
  39796=>"111111011",
  39797=>"000000000",
  39798=>"000000000",
  39799=>"000000011",
  39800=>"001000000",
  39801=>"011000000",
  39802=>"111000000",
  39803=>"000001010",
  39804=>"000001111",
  39805=>"000000111",
  39806=>"010010000",
  39807=>"000000000",
  39808=>"000001001",
  39809=>"000100111",
  39810=>"111111001",
  39811=>"011011110",
  39812=>"000000111",
  39813=>"000000000",
  39814=>"110000111",
  39815=>"010000111",
  39816=>"111111000",
  39817=>"000000000",
  39818=>"111111110",
  39819=>"000000011",
  39820=>"000100111",
  39821=>"111001001",
  39822=>"000100001",
  39823=>"000000100",
  39824=>"000000000",
  39825=>"011001000",
  39826=>"101100000",
  39827=>"111011001",
  39828=>"111111111",
  39829=>"000010000",
  39830=>"110100000",
  39831=>"111011011",
  39832=>"100100000",
  39833=>"000000101",
  39834=>"111111100",
  39835=>"100100000",
  39836=>"000000000",
  39837=>"111111100",
  39838=>"110000110",
  39839=>"000000000",
  39840=>"111100111",
  39841=>"111111000",
  39842=>"000000001",
  39843=>"000000111",
  39844=>"000000000",
  39845=>"000000110",
  39846=>"100100110",
  39847=>"010111001",
  39848=>"000001000",
  39849=>"000001011",
  39850=>"000010000",
  39851=>"100000000",
  39852=>"011010000",
  39853=>"111111101",
  39854=>"000000000",
  39855=>"000000000",
  39856=>"000011111",
  39857=>"111111011",
  39858=>"111000000",
  39859=>"111110100",
  39860=>"000000000",
  39861=>"000000100",
  39862=>"001000110",
  39863=>"100101111",
  39864=>"100000000",
  39865=>"001011111",
  39866=>"000000001",
  39867=>"011000111",
  39868=>"001000000",
  39869=>"000010111",
  39870=>"001000000",
  39871=>"000000000",
  39872=>"000000111",
  39873=>"000001001",
  39874=>"111111111",
  39875=>"000000000",
  39876=>"000000001",
  39877=>"100110001",
  39878=>"111100000",
  39879=>"010000000",
  39880=>"000000000",
  39881=>"100000000",
  39882=>"011011001",
  39883=>"000111000",
  39884=>"101000000",
  39885=>"000000000",
  39886=>"100100000",
  39887=>"100010010",
  39888=>"111111001",
  39889=>"000111111",
  39890=>"000000111",
  39891=>"000000110",
  39892=>"100000110",
  39893=>"010000111",
  39894=>"001000000",
  39895=>"011000000",
  39896=>"000001000",
  39897=>"110100000",
  39898=>"111111010",
  39899=>"111111011",
  39900=>"000011111",
  39901=>"100100111",
  39902=>"100100111",
  39903=>"100001001",
  39904=>"000000000",
  39905=>"111111111",
  39906=>"000000101",
  39907=>"001000000",
  39908=>"111111111",
  39909=>"111111100",
  39910=>"111111111",
  39911=>"110111111",
  39912=>"001000010",
  39913=>"100111001",
  39914=>"110000000",
  39915=>"111111000",
  39916=>"011111111",
  39917=>"111111000",
  39918=>"001101001",
  39919=>"111000010",
  39920=>"101000111",
  39921=>"000011111",
  39922=>"000000111",
  39923=>"111000000",
  39924=>"111111111",
  39925=>"100000000",
  39926=>"000111111",
  39927=>"111110000",
  39928=>"000000000",
  39929=>"000000001",
  39930=>"000000000",
  39931=>"110110111",
  39932=>"000111111",
  39933=>"000000000",
  39934=>"111111111",
  39935=>"000000001",
  39936=>"011011101",
  39937=>"111011001",
  39938=>"111111111",
  39939=>"101111111",
  39940=>"101101111",
  39941=>"100101101",
  39942=>"001001111",
  39943=>"010010010",
  39944=>"011000000",
  39945=>"110100100",
  39946=>"001100000",
  39947=>"000000011",
  39948=>"110001001",
  39949=>"101111111",
  39950=>"001000011",
  39951=>"111000100",
  39952=>"111100111",
  39953=>"001000000",
  39954=>"000000111",
  39955=>"111100000",
  39956=>"000000000",
  39957=>"100100000",
  39958=>"100111111",
  39959=>"110110111",
  39960=>"001000000",
  39961=>"011011110",
  39962=>"000101111",
  39963=>"111110110",
  39964=>"111111010",
  39965=>"100111101",
  39966=>"111111010",
  39967=>"111111000",
  39968=>"000000000",
  39969=>"110110111",
  39970=>"101000001",
  39971=>"011010010",
  39972=>"110101110",
  39973=>"000111111",
  39974=>"000000000",
  39975=>"101101111",
  39976=>"000110111",
  39977=>"100110010",
  39978=>"000000000",
  39979=>"011111111",
  39980=>"111011001",
  39981=>"101001011",
  39982=>"000100100",
  39983=>"100000000",
  39984=>"111111100",
  39985=>"000000011",
  39986=>"111111111",
  39987=>"101100100",
  39988=>"101101111",
  39989=>"111111111",
  39990=>"001011101",
  39991=>"110111111",
  39992=>"011001111",
  39993=>"111111100",
  39994=>"111100111",
  39995=>"000000001",
  39996=>"100100000",
  39997=>"100100000",
  39998=>"111011000",
  39999=>"111111110",
  40000=>"000000100",
  40001=>"100100100",
  40002=>"011111111",
  40003=>"100110111",
  40004=>"000000000",
  40005=>"010010000",
  40006=>"000000000",
  40007=>"110000000",
  40008=>"000000000",
  40009=>"000000000",
  40010=>"000101111",
  40011=>"011010110",
  40012=>"001101111",
  40013=>"111001111",
  40014=>"000100001",
  40015=>"111111111",
  40016=>"011011000",
  40017=>"100000001",
  40018=>"000000000",
  40019=>"000000011",
  40020=>"101100101",
  40021=>"111011000",
  40022=>"101101101",
  40023=>"001000111",
  40024=>"111111011",
  40025=>"000000000",
  40026=>"000110111",
  40027=>"111111111",
  40028=>"111111111",
  40029=>"000000000",
  40030=>"110111111",
  40031=>"100110100",
  40032=>"111101111",
  40033=>"100000000",
  40034=>"110110000",
  40035=>"000100110",
  40036=>"001000000",
  40037=>"111111111",
  40038=>"110110000",
  40039=>"111001001",
  40040=>"000111111",
  40041=>"110111111",
  40042=>"000000010",
  40043=>"111111111",
  40044=>"000000001",
  40045=>"000110000",
  40046=>"000000000",
  40047=>"000000000",
  40048=>"111111111",
  40049=>"111111011",
  40050=>"000000011",
  40051=>"111111011",
  40052=>"100100100",
  40053=>"111111111",
  40054=>"000000000",
  40055=>"101000000",
  40056=>"000000000",
  40057=>"000101000",
  40058=>"001000000",
  40059=>"111011111",
  40060=>"000000000",
  40061=>"110110000",
  40062=>"000000000",
  40063=>"101111111",
  40064=>"100000000",
  40065=>"000001101",
  40066=>"110010110",
  40067=>"100100110",
  40068=>"111111111",
  40069=>"000000110",
  40070=>"111111101",
  40071=>"111010000",
  40072=>"111000000",
  40073=>"000000001",
  40074=>"100100000",
  40075=>"111111111",
  40076=>"000000000",
  40077=>"111111111",
  40078=>"000000101",
  40079=>"111111111",
  40080=>"000000000",
  40081=>"100101111",
  40082=>"011111111",
  40083=>"111111111",
  40084=>"000000000",
  40085=>"100100101",
  40086=>"000000000",
  40087=>"000000000",
  40088=>"001000101",
  40089=>"000000000",
  40090=>"000000000",
  40091=>"110100000",
  40092=>"111111111",
  40093=>"111010000",
  40094=>"110100111",
  40095=>"111111111",
  40096=>"000100000",
  40097=>"100111111",
  40098=>"111101100",
  40099=>"011000101",
  40100=>"111010100",
  40101=>"111101111",
  40102=>"111111011",
  40103=>"010110110",
  40104=>"011011000",
  40105=>"100111111",
  40106=>"000001011",
  40107=>"111111111",
  40108=>"000000000",
  40109=>"101111001",
  40110=>"000100111",
  40111=>"000011111",
  40112=>"000000000",
  40113=>"100100001",
  40114=>"111001001",
  40115=>"111111111",
  40116=>"111000011",
  40117=>"111111111",
  40118=>"000000000",
  40119=>"111111111",
  40120=>"100111111",
  40121=>"111000001",
  40122=>"011011010",
  40123=>"101100001",
  40124=>"011011000",
  40125=>"111111111",
  40126=>"011000000",
  40127=>"111001101",
  40128=>"000100100",
  40129=>"001011111",
  40130=>"000101111",
  40131=>"111111111",
  40132=>"111010000",
  40133=>"111111111",
  40134=>"011111111",
  40135=>"000100101",
  40136=>"111110010",
  40137=>"000100101",
  40138=>"101111111",
  40139=>"100100000",
  40140=>"000100001",
  40141=>"000111111",
  40142=>"011110111",
  40143=>"011000000",
  40144=>"110110111",
  40145=>"000000100",
  40146=>"000111000",
  40147=>"000000000",
  40148=>"000110110",
  40149=>"000011011",
  40150=>"000000000",
  40151=>"000000100",
  40152=>"111111111",
  40153=>"000000000",
  40154=>"010000000",
  40155=>"001011111",
  40156=>"100000000",
  40157=>"001011111",
  40158=>"111111111",
  40159=>"111111111",
  40160=>"000000111",
  40161=>"101100110",
  40162=>"000111111",
  40163=>"111111111",
  40164=>"111110111",
  40165=>"111111111",
  40166=>"111111011",
  40167=>"111111111",
  40168=>"111101100",
  40169=>"000000000",
  40170=>"011001111",
  40171=>"011111111",
  40172=>"111011000",
  40173=>"000000000",
  40174=>"111111001",
  40175=>"111110000",
  40176=>"000011011",
  40177=>"000010100",
  40178=>"111111111",
  40179=>"000000000",
  40180=>"001111111",
  40181=>"001011011",
  40182=>"100100110",
  40183=>"111000000",
  40184=>"111111111",
  40185=>"101100100",
  40186=>"111111111",
  40187=>"000000110",
  40188=>"110101111",
  40189=>"111000001",
  40190=>"111000001",
  40191=>"000000000",
  40192=>"111111111",
  40193=>"001000000",
  40194=>"111111111",
  40195=>"000110111",
  40196=>"000000000",
  40197=>"100100111",
  40198=>"001010000",
  40199=>"000111111",
  40200=>"011000000",
  40201=>"111111100",
  40202=>"111111111",
  40203=>"000100111",
  40204=>"111101101",
  40205=>"000100111",
  40206=>"011111111",
  40207=>"000000000",
  40208=>"111011001",
  40209=>"001101111",
  40210=>"011001000",
  40211=>"111111111",
  40212=>"011011000",
  40213=>"000000000",
  40214=>"000000000",
  40215=>"000000000",
  40216=>"101000000",
  40217=>"111100000",
  40218=>"000001111",
  40219=>"101101101",
  40220=>"110110110",
  40221=>"100100100",
  40222=>"001111111",
  40223=>"111111111",
  40224=>"111111111",
  40225=>"011111110",
  40226=>"111111111",
  40227=>"000000111",
  40228=>"000000000",
  40229=>"011001001",
  40230=>"000000100",
  40231=>"000011100",
  40232=>"111111101",
  40233=>"010000001",
  40234=>"111011000",
  40235=>"000000000",
  40236=>"111111111",
  40237=>"100110111",
  40238=>"001011000",
  40239=>"000001101",
  40240=>"001001001",
  40241=>"111111111",
  40242=>"000000100",
  40243=>"111110100",
  40244=>"000001000",
  40245=>"000100111",
  40246=>"111111111",
  40247=>"000010111",
  40248=>"000000000",
  40249=>"000000001",
  40250=>"111111000",
  40251=>"101111001",
  40252=>"000000000",
  40253=>"100100100",
  40254=>"111111101",
  40255=>"001001001",
  40256=>"100110000",
  40257=>"000000010",
  40258=>"111101101",
  40259=>"000000000",
  40260=>"000000000",
  40261=>"111110100",
  40262=>"001000000",
  40263=>"101001001",
  40264=>"001100111",
  40265=>"110111111",
  40266=>"111111100",
  40267=>"100100100",
  40268=>"011111111",
  40269=>"000110011",
  40270=>"100100101",
  40271=>"000001000",
  40272=>"001011111",
  40273=>"000000100",
  40274=>"111000100",
  40275=>"001001000",
  40276=>"101000000",
  40277=>"000000000",
  40278=>"101111111",
  40279=>"000100000",
  40280=>"111111111",
  40281=>"000000000",
  40282=>"000101111",
  40283=>"111100111",
  40284=>"000000000",
  40285=>"100111111",
  40286=>"111101001",
  40287=>"000000011",
  40288=>"100111110",
  40289=>"000110111",
  40290=>"111111110",
  40291=>"000000001",
  40292=>"000001111",
  40293=>"000101101",
  40294=>"111111111",
  40295=>"000000011",
  40296=>"000000000",
  40297=>"000000000",
  40298=>"001011110",
  40299=>"111000000",
  40300=>"001001000",
  40301=>"110000010",
  40302=>"000000000",
  40303=>"000000000",
  40304=>"111001100",
  40305=>"000011001",
  40306=>"111000000",
  40307=>"011011001",
  40308=>"111111001",
  40309=>"111100111",
  40310=>"000010000",
  40311=>"000000000",
  40312=>"000000000",
  40313=>"100000000",
  40314=>"111111111",
  40315=>"011111111",
  40316=>"000000000",
  40317=>"001000000",
  40318=>"000000000",
  40319=>"000000000",
  40320=>"000000011",
  40321=>"001001101",
  40322=>"000010000",
  40323=>"111100100",
  40324=>"011000001",
  40325=>"000000000",
  40326=>"100000000",
  40327=>"000000000",
  40328=>"000001100",
  40329=>"111100010",
  40330=>"111101101",
  40331=>"111111111",
  40332=>"000000000",
  40333=>"111101000",
  40334=>"100111111",
  40335=>"001011000",
  40336=>"111110100",
  40337=>"111100000",
  40338=>"100111000",
  40339=>"000011000",
  40340=>"000000111",
  40341=>"001001001",
  40342=>"101111111",
  40343=>"110111111",
  40344=>"011111111",
  40345=>"111111101",
  40346=>"111111111",
  40347=>"111111111",
  40348=>"111100100",
  40349=>"111111011",
  40350=>"001001111",
  40351=>"000000000",
  40352=>"011001100",
  40353=>"000000010",
  40354=>"000000111",
  40355=>"111111111",
  40356=>"111111111",
  40357=>"101000000",
  40358=>"000001000",
  40359=>"001100100",
  40360=>"101101111",
  40361=>"000011000",
  40362=>"111111111",
  40363=>"100100110",
  40364=>"111101101",
  40365=>"100000000",
  40366=>"111010110",
  40367=>"111001000",
  40368=>"000000000",
  40369=>"111001111",
  40370=>"111111111",
  40371=>"001101100",
  40372=>"001000000",
  40373=>"100100010",
  40374=>"000110000",
  40375=>"101110000",
  40376=>"111111011",
  40377=>"111111111",
  40378=>"010011111",
  40379=>"000000000",
  40380=>"000001111",
  40381=>"000011001",
  40382=>"000000000",
  40383=>"110100011",
  40384=>"100100000",
  40385=>"100000000",
  40386=>"000000000",
  40387=>"000000000",
  40388=>"111111111",
  40389=>"000110110",
  40390=>"000110111",
  40391=>"000000000",
  40392=>"011111100",
  40393=>"111111100",
  40394=>"000101111",
  40395=>"000111111",
  40396=>"000111111",
  40397=>"111111000",
  40398=>"111111111",
  40399=>"111111111",
  40400=>"001001000",
  40401=>"111100111",
  40402=>"011011011",
  40403=>"111111111",
  40404=>"000000110",
  40405=>"000000111",
  40406=>"111111111",
  40407=>"100000110",
  40408=>"111111101",
  40409=>"101100111",
  40410=>"000111111",
  40411=>"011010011",
  40412=>"000001111",
  40413=>"001100000",
  40414=>"000000110",
  40415=>"011011111",
  40416=>"111111010",
  40417=>"010000001",
  40418=>"111111000",
  40419=>"111000000",
  40420=>"010000000",
  40421=>"010000000",
  40422=>"100001010",
  40423=>"001000000",
  40424=>"000000000",
  40425=>"111111001",
  40426=>"110000000",
  40427=>"000001000",
  40428=>"000011111",
  40429=>"000000000",
  40430=>"000000011",
  40431=>"000011001",
  40432=>"001011011",
  40433=>"001000100",
  40434=>"111000100",
  40435=>"101100101",
  40436=>"111000000",
  40437=>"001000000",
  40438=>"111111000",
  40439=>"001011011",
  40440=>"110000000",
  40441=>"000000001",
  40442=>"100000000",
  40443=>"000111111",
  40444=>"001101111",
  40445=>"001000001",
  40446=>"111111000",
  40447=>"000000111",
  40448=>"111011011",
  40449=>"000000000",
  40450=>"000000000",
  40451=>"011011001",
  40452=>"010111111",
  40453=>"000101111",
  40454=>"111111111",
  40455=>"001001000",
  40456=>"111101111",
  40457=>"110010110",
  40458=>"111111111",
  40459=>"101100000",
  40460=>"001000100",
  40461=>"001001000",
  40462=>"000000000",
  40463=>"000011000",
  40464=>"000010111",
  40465=>"000001101",
  40466=>"111111111",
  40467=>"111111111",
  40468=>"011111111",
  40469=>"011011000",
  40470=>"000000000",
  40471=>"100100101",
  40472=>"111011011",
  40473=>"000000100",
  40474=>"111011001",
  40475=>"010110100",
  40476=>"010110111",
  40477=>"111111111",
  40478=>"001001111",
  40479=>"000000100",
  40480=>"011011011",
  40481=>"111111100",
  40482=>"110110110",
  40483=>"100000000",
  40484=>"001000001",
  40485=>"111111101",
  40486=>"000000000",
  40487=>"001000000",
  40488=>"000010000",
  40489=>"000000000",
  40490=>"110100111",
  40491=>"110100110",
  40492=>"000000000",
  40493=>"101001111",
  40494=>"000000000",
  40495=>"111111111",
  40496=>"111011001",
  40497=>"000000001",
  40498=>"011111011",
  40499=>"011111100",
  40500=>"000000000",
  40501=>"000000000",
  40502=>"000000000",
  40503=>"111100111",
  40504=>"000000001",
  40505=>"011111111",
  40506=>"100111111",
  40507=>"000000000",
  40508=>"000000101",
  40509=>"001001000",
  40510=>"000000000",
  40511=>"111111111",
  40512=>"000000010",
  40513=>"111111111",
  40514=>"100001000",
  40515=>"111111100",
  40516=>"110110110",
  40517=>"101000101",
  40518=>"111000000",
  40519=>"111111001",
  40520=>"011111011",
  40521=>"000000000",
  40522=>"111001000",
  40523=>"000111111",
  40524=>"000000000",
  40525=>"111111000",
  40526=>"000001111",
  40527=>"100100000",
  40528=>"101111111",
  40529=>"111111111",
  40530=>"000000000",
  40531=>"111011000",
  40532=>"011011111",
  40533=>"000111111",
  40534=>"000000000",
  40535=>"110110111",
  40536=>"000000000",
  40537=>"000000000",
  40538=>"000000000",
  40539=>"111111111",
  40540=>"000111111",
  40541=>"000110111",
  40542=>"000010010",
  40543=>"000011000",
  40544=>"111111111",
  40545=>"111111111",
  40546=>"110111111",
  40547=>"000000000",
  40548=>"000000111",
  40549=>"000000001",
  40550=>"110110100",
  40551=>"111111000",
  40552=>"000000110",
  40553=>"111111100",
  40554=>"011001000",
  40555=>"110010011",
  40556=>"111011000",
  40557=>"000000001",
  40558=>"000000000",
  40559=>"000000000",
  40560=>"101111000",
  40561=>"000000000",
  40562=>"001011011",
  40563=>"000000000",
  40564=>"000001000",
  40565=>"111111111",
  40566=>"111111111",
  40567=>"111111110",
  40568=>"000000111",
  40569=>"111111111",
  40570=>"111101001",
  40571=>"101111111",
  40572=>"011011001",
  40573=>"111111110",
  40574=>"000000000",
  40575=>"111111111",
  40576=>"111111111",
  40577=>"011010000",
  40578=>"100000000",
  40579=>"000100000",
  40580=>"000000111",
  40581=>"000000000",
  40582=>"000000000",
  40583=>"001000000",
  40584=>"111111011",
  40585=>"001100110",
  40586=>"111110000",
  40587=>"000000000",
  40588=>"000000110",
  40589=>"111111000",
  40590=>"010010000",
  40591=>"000100100",
  40592=>"001000000",
  40593=>"001101111",
  40594=>"000000000",
  40595=>"100101100",
  40596=>"111111000",
  40597=>"001000000",
  40598=>"111111111",
  40599=>"111111010",
  40600=>"000000000",
  40601=>"000110111",
  40602=>"111111111",
  40603=>"111111111",
  40604=>"110010000",
  40605=>"111001101",
  40606=>"000000000",
  40607=>"000000000",
  40608=>"011001000",
  40609=>"000000000",
  40610=>"111111111",
  40611=>"111111111",
  40612=>"000000000",
  40613=>"011001000",
  40614=>"111111111",
  40615=>"000100111",
  40616=>"001001000",
  40617=>"000001001",
  40618=>"100000000",
  40619=>"000000000",
  40620=>"000000000",
  40621=>"111100101",
  40622=>"010111111",
  40623=>"100000000",
  40624=>"111111100",
  40625=>"000011111",
  40626=>"000001011",
  40627=>"000000101",
  40628=>"111101100",
  40629=>"101011011",
  40630=>"010111110",
  40631=>"100000100",
  40632=>"000000000",
  40633=>"000000000",
  40634=>"001000110",
  40635=>"001011000",
  40636=>"110100111",
  40637=>"111111111",
  40638=>"111000000",
  40639=>"111001011",
  40640=>"110000000",
  40641=>"100111111",
  40642=>"000111111",
  40643=>"110100100",
  40644=>"111111110",
  40645=>"000000010",
  40646=>"111101001",
  40647=>"000001111",
  40648=>"000000000",
  40649=>"000000000",
  40650=>"000000000",
  40651=>"001001000",
  40652=>"001000000",
  40653=>"111001001",
  40654=>"001001000",
  40655=>"111111111",
  40656=>"111000010",
  40657=>"111100000",
  40658=>"111100100",
  40659=>"111111000",
  40660=>"000000011",
  40661=>"001000000",
  40662=>"001000101",
  40663=>"110000110",
  40664=>"111111111",
  40665=>"000110111",
  40666=>"100000011",
  40667=>"000000000",
  40668=>"001000000",
  40669=>"100001000",
  40670=>"000000000",
  40671=>"111111111",
  40672=>"000000010",
  40673=>"000000111",
  40674=>"000000000",
  40675=>"111111000",
  40676=>"101000110",
  40677=>"000111101",
  40678=>"111111001",
  40679=>"010111111",
  40680=>"000111111",
  40681=>"000100000",
  40682=>"000000011",
  40683=>"111111001",
  40684=>"000110011",
  40685=>"000000111",
  40686=>"011010000",
  40687=>"111011000",
  40688=>"100000000",
  40689=>"111111011",
  40690=>"111111111",
  40691=>"001000100",
  40692=>"111111110",
  40693=>"000010011",
  40694=>"011111111",
  40695=>"000000111",
  40696=>"000000000",
  40697=>"000000111",
  40698=>"000111111",
  40699=>"000001101",
  40700=>"100100011",
  40701=>"000000100",
  40702=>"001111000",
  40703=>"111111110",
  40704=>"000000000",
  40705=>"000100100",
  40706=>"000000001",
  40707=>"000000000",
  40708=>"011011011",
  40709=>"110110110",
  40710=>"111111111",
  40711=>"000000000",
  40712=>"000101001",
  40713=>"100111111",
  40714=>"111111111",
  40715=>"000000000",
  40716=>"111011000",
  40717=>"000000010",
  40718=>"111111111",
  40719=>"100100111",
  40720=>"100111001",
  40721=>"000100111",
  40722=>"001001001",
  40723=>"000000100",
  40724=>"100111111",
  40725=>"000000000",
  40726=>"001100110",
  40727=>"011011000",
  40728=>"011100110",
  40729=>"111111111",
  40730=>"000000000",
  40731=>"111101111",
  40732=>"110110110",
  40733=>"000000000",
  40734=>"000000111",
  40735=>"000000111",
  40736=>"100100111",
  40737=>"000110100",
  40738=>"111111111",
  40739=>"111011000",
  40740=>"111111000",
  40741=>"110110110",
  40742=>"100000011",
  40743=>"000000011",
  40744=>"111111110",
  40745=>"111111111",
  40746=>"000000000",
  40747=>"000000000",
  40748=>"011000000",
  40749=>"011011111",
  40750=>"100111111",
  40751=>"001001001",
  40752=>"100110111",
  40753=>"000000000",
  40754=>"111111111",
  40755=>"000000000",
  40756=>"001111111",
  40757=>"011101100",
  40758=>"000001001",
  40759=>"111100000",
  40760=>"111111111",
  40761=>"111011111",
  40762=>"001001000",
  40763=>"111110100",
  40764=>"110111100",
  40765=>"000000000",
  40766=>"000000000",
  40767=>"000001000",
  40768=>"011000000",
  40769=>"000110010",
  40770=>"000111111",
  40771=>"111111111",
  40772=>"000000110",
  40773=>"000011011",
  40774=>"111111100",
  40775=>"001000000",
  40776=>"000000000",
  40777=>"111010010",
  40778=>"000000000",
  40779=>"000000100",
  40780=>"110111111",
  40781=>"000000000",
  40782=>"000000000",
  40783=>"000111001",
  40784=>"000011111",
  40785=>"001001001",
  40786=>"000110110",
  40787=>"000000000",
  40788=>"111111011",
  40789=>"011011001",
  40790=>"000011001",
  40791=>"000000000",
  40792=>"001001000",
  40793=>"000000000",
  40794=>"000000000",
  40795=>"000000000",
  40796=>"111111000",
  40797=>"110000000",
  40798=>"001111111",
  40799=>"000000000",
  40800=>"111111111",
  40801=>"111101111",
  40802=>"000000000",
  40803=>"100000000",
  40804=>"000001111",
  40805=>"000000100",
  40806=>"001000000",
  40807=>"000001011",
  40808=>"001011011",
  40809=>"111001010",
  40810=>"111000000",
  40811=>"000000101",
  40812=>"000110110",
  40813=>"000000110",
  40814=>"110010100",
  40815=>"010111011",
  40816=>"110000010",
  40817=>"001000000",
  40818=>"110111010",
  40819=>"110111011",
  40820=>"000000000",
  40821=>"000000011",
  40822=>"010000000",
  40823=>"111011000",
  40824=>"111110000",
  40825=>"000000000",
  40826=>"001001001",
  40827=>"000000000",
  40828=>"111000000",
  40829=>"000000100",
  40830=>"000111111",
  40831=>"110111111",
  40832=>"111101000",
  40833=>"111100000",
  40834=>"110110110",
  40835=>"000000000",
  40836=>"101001111",
  40837=>"000000000",
  40838=>"111111011",
  40839=>"000110100",
  40840=>"000000110",
  40841=>"110010000",
  40842=>"000000001",
  40843=>"000000000",
  40844=>"110111111",
  40845=>"111111000",
  40846=>"000010111",
  40847=>"101101111",
  40848=>"000001111",
  40849=>"001000000",
  40850=>"111111111",
  40851=>"111111111",
  40852=>"000000000",
  40853=>"011001011",
  40854=>"000000000",
  40855=>"000000111",
  40856=>"110111111",
  40857=>"111111111",
  40858=>"000000000",
  40859=>"100000000",
  40860=>"111111111",
  40861=>"110111000",
  40862=>"101111111",
  40863=>"000000100",
  40864=>"110000000",
  40865=>"110110110",
  40866=>"000110100",
  40867=>"111111010",
  40868=>"000000110",
  40869=>"110111011",
  40870=>"000000111",
  40871=>"000111111",
  40872=>"100111111",
  40873=>"010111000",
  40874=>"000000100",
  40875=>"000000000",
  40876=>"001001001",
  40877=>"011011000",
  40878=>"001000000",
  40879=>"100000000",
  40880=>"001001010",
  40881=>"110100111",
  40882=>"000011111",
  40883=>"000011111",
  40884=>"101101100",
  40885=>"000000000",
  40886=>"001011111",
  40887=>"111111111",
  40888=>"000111111",
  40889=>"000001000",
  40890=>"111111000",
  40891=>"111111101",
  40892=>"101000000",
  40893=>"111100100",
  40894=>"111101000",
  40895=>"011111000",
  40896=>"111111110",
  40897=>"001000001",
  40898=>"000000001",
  40899=>"000000000",
  40900=>"000001111",
  40901=>"110111000",
  40902=>"111111111",
  40903=>"000111111",
  40904=>"000001001",
  40905=>"011011001",
  40906=>"000000000",
  40907=>"000000000",
  40908=>"111100101",
  40909=>"001111111",
  40910=>"111110100",
  40911=>"111111000",
  40912=>"000111111",
  40913=>"000011001",
  40914=>"000001111",
  40915=>"111000000",
  40916=>"000100110",
  40917=>"011111110",
  40918=>"011001001",
  40919=>"000000011",
  40920=>"011011111",
  40921=>"001111111",
  40922=>"111000000",
  40923=>"000000000",
  40924=>"100110111",
  40925=>"000100000",
  40926=>"001000000",
  40927=>"111111111",
  40928=>"011111010",
  40929=>"000000000",
  40930=>"000000000",
  40931=>"100100101",
  40932=>"000010111",
  40933=>"101000000",
  40934=>"000000000",
  40935=>"000010010",
  40936=>"000000001",
  40937=>"111111000",
  40938=>"001001101",
  40939=>"000000001",
  40940=>"000000000",
  40941=>"000001001",
  40942=>"001001001",
  40943=>"111111111",
  40944=>"111100101",
  40945=>"011110000",
  40946=>"101000000",
  40947=>"111011001",
  40948=>"000001011",
  40949=>"111111011",
  40950=>"000000000",
  40951=>"111011011",
  40952=>"011111011",
  40953=>"010011011",
  40954=>"100000000",
  40955=>"011000000",
  40956=>"001001111",
  40957=>"011111110",
  40958=>"011011000",
  40959=>"001000000",
  40960=>"010111111",
  40961=>"000100100",
  40962=>"110000101",
  40963=>"111111000",
  40964=>"001000111",
  40965=>"111011100",
  40966=>"000000111",
  40967=>"111101111",
  40968=>"110111111",
  40969=>"111000001",
  40970=>"101001101",
  40971=>"001000001",
  40972=>"110000000",
  40973=>"000111111",
  40974=>"000000100",
  40975=>"000001000",
  40976=>"111111110",
  40977=>"111111111",
  40978=>"101111100",
  40979=>"111111111",
  40980=>"001000111",
  40981=>"001110111",
  40982=>"111110000",
  40983=>"111011000",
  40984=>"111001001",
  40985=>"001110110",
  40986=>"111111111",
  40987=>"110110111",
  40988=>"111010001",
  40989=>"100110000",
  40990=>"000000000",
  40991=>"010111010",
  40992=>"101101101",
  40993=>"000001111",
  40994=>"000000100",
  40995=>"001000011",
  40996=>"111110000",
  40997=>"000000101",
  40998=>"111111011",
  40999=>"001000001",
  41000=>"000001000",
  41001=>"000000000",
  41002=>"101100111",
  41003=>"000110110",
  41004=>"010110010",
  41005=>"100000100",
  41006=>"010000001",
  41007=>"000000000",
  41008=>"001111110",
  41009=>"000111000",
  41010=>"011011001",
  41011=>"111111111",
  41012=>"101001101",
  41013=>"100111001",
  41014=>"111111110",
  41015=>"001111100",
  41016=>"100001111",
  41017=>"111101111",
  41018=>"000000000",
  41019=>"100000111",
  41020=>"111000000",
  41021=>"000111100",
  41022=>"001111100",
  41023=>"000000000",
  41024=>"111111110",
  41025=>"001111111",
  41026=>"000000000",
  41027=>"001000000",
  41028=>"000000111",
  41029=>"000000001",
  41030=>"000011111",
  41031=>"111011111",
  41032=>"011011000",
  41033=>"000000000",
  41034=>"101000101",
  41035=>"111111111",
  41036=>"110110111",
  41037=>"101100111",
  41038=>"000000000",
  41039=>"110111110",
  41040=>"000000000",
  41041=>"111111000",
  41042=>"111001111",
  41043=>"111000010",
  41044=>"000100100",
  41045=>"100101001",
  41046=>"111111111",
  41047=>"000000000",
  41048=>"010110100",
  41049=>"111111111",
  41050=>"000000000",
  41051=>"000110000",
  41052=>"101001111",
  41053=>"111111111",
  41054=>"000110111",
  41055=>"011111100",
  41056=>"010110000",
  41057=>"000001000",
  41058=>"101000011",
  41059=>"001000000",
  41060=>"110000000",
  41061=>"101111111",
  41062=>"110111011",
  41063=>"110110110",
  41064=>"101001111",
  41065=>"111001111",
  41066=>"111000100",
  41067=>"000000000",
  41068=>"000000001",
  41069=>"000000110",
  41070=>"000110111",
  41071=>"000000111",
  41072=>"111111111",
  41073=>"001000000",
  41074=>"111100101",
  41075=>"000000000",
  41076=>"111100110",
  41077=>"110111010",
  41078=>"111000000",
  41079=>"111011000",
  41080=>"111111011",
  41081=>"111111111",
  41082=>"000001111",
  41083=>"111000000",
  41084=>"000011010",
  41085=>"111100101",
  41086=>"010111011",
  41087=>"100101100",
  41088=>"000000011",
  41089=>"111100100",
  41090=>"100110111",
  41091=>"111100100",
  41092=>"110110000",
  41093=>"111001111",
  41094=>"000111000",
  41095=>"111001000",
  41096=>"111101111",
  41097=>"111100000",
  41098=>"000001001",
  41099=>"111100101",
  41100=>"000000000",
  41101=>"111000000",
  41102=>"111011000",
  41103=>"001000000",
  41104=>"101000001",
  41105=>"100000000",
  41106=>"111000000",
  41107=>"010000000",
  41108=>"000110010",
  41109=>"111100101",
  41110=>"100000111",
  41111=>"111101111",
  41112=>"000000011",
  41113=>"111000000",
  41114=>"111111111",
  41115=>"111111011",
  41116=>"000000000",
  41117=>"111100100",
  41118=>"111101000",
  41119=>"000000111",
  41120=>"000000111",
  41121=>"101000000",
  41122=>"011010111",
  41123=>"000111010",
  41124=>"001111111",
  41125=>"111000000",
  41126=>"111111000",
  41127=>"111111000",
  41128=>"101110110",
  41129=>"010111000",
  41130=>"111111111",
  41131=>"111111100",
  41132=>"101111010",
  41133=>"110111011",
  41134=>"000000000",
  41135=>"111111111",
  41136=>"011111000",
  41137=>"000001000",
  41138=>"010111010",
  41139=>"111001000",
  41140=>"111111010",
  41141=>"111110110",
  41142=>"110010000",
  41143=>"111000000",
  41144=>"100101111",
  41145=>"001011000",
  41146=>"000000101",
  41147=>"111110000",
  41148=>"110111111",
  41149=>"000111111",
  41150=>"110000000",
  41151=>"111111111",
  41152=>"000000000",
  41153=>"001001111",
  41154=>"110110111",
  41155=>"011111000",
  41156=>"111111111",
  41157=>"111000001",
  41158=>"000101000",
  41159=>"001000100",
  41160=>"110111110",
  41161=>"111111100",
  41162=>"100000100",
  41163=>"111000111",
  41164=>"110100111",
  41165=>"000110111",
  41166=>"001111000",
  41167=>"001111111",
  41168=>"000011000",
  41169=>"111111111",
  41170=>"111111000",
  41171=>"001000000",
  41172=>"100001001",
  41173=>"111111000",
  41174=>"000000001",
  41175=>"100101100",
  41176=>"000100111",
  41177=>"000010111",
  41178=>"000000000",
  41179=>"111111010",
  41180=>"111111000",
  41181=>"111111000",
  41182=>"111111111",
  41183=>"000000101",
  41184=>"000001000",
  41185=>"111111111",
  41186=>"010000000",
  41187=>"000000000",
  41188=>"000000000",
  41189=>"010110110",
  41190=>"000000000",
  41191=>"010000011",
  41192=>"111111110",
  41193=>"001000000",
  41194=>"111010010",
  41195=>"111100100",
  41196=>"000000100",
  41197=>"111000001",
  41198=>"011000000",
  41199=>"000000101",
  41200=>"000110110",
  41201=>"111100101",
  41202=>"111100111",
  41203=>"000000101",
  41204=>"011010111",
  41205=>"000111111",
  41206=>"000000011",
  41207=>"111110000",
  41208=>"101001000",
  41209=>"000111111",
  41210=>"001011001",
  41211=>"110000000",
  41212=>"000000001",
  41213=>"110110000",
  41214=>"110110000",
  41215=>"000010000",
  41216=>"000000001",
  41217=>"111000000",
  41218=>"111111111",
  41219=>"100110110",
  41220=>"000101001",
  41221=>"111000000",
  41222=>"000000000",
  41223=>"101101111",
  41224=>"000000110",
  41225=>"001001000",
  41226=>"000100111",
  41227=>"111111011",
  41228=>"110000001",
  41229=>"111111111",
  41230=>"000101111",
  41231=>"111001111",
  41232=>"000111000",
  41233=>"111000100",
  41234=>"110000000",
  41235=>"110111001",
  41236=>"111000000",
  41237=>"000000111",
  41238=>"001011001",
  41239=>"111111111",
  41240=>"011011001",
  41241=>"001000000",
  41242=>"000000000",
  41243=>"111000111",
  41244=>"001100111",
  41245=>"001110010",
  41246=>"000000111",
  41247=>"000000101",
  41248=>"111100110",
  41249=>"001000001",
  41250=>"000001000",
  41251=>"111111111",
  41252=>"011000000",
  41253=>"000000000",
  41254=>"101100000",
  41255=>"000000100",
  41256=>"000000000",
  41257=>"010110111",
  41258=>"110000111",
  41259=>"111101000",
  41260=>"010010000",
  41261=>"111010001",
  41262=>"111011000",
  41263=>"000000000",
  41264=>"010111111",
  41265=>"111100100",
  41266=>"111111110",
  41267=>"000000110",
  41268=>"000111010",
  41269=>"000000111",
  41270=>"000000111",
  41271=>"000000110",
  41272=>"000000111",
  41273=>"000111111",
  41274=>"000000100",
  41275=>"001001000",
  41276=>"111101011",
  41277=>"110110110",
  41278=>"001111111",
  41279=>"111011111",
  41280=>"000111111",
  41281=>"111000000",
  41282=>"000000000",
  41283=>"111000000",
  41284=>"000000010",
  41285=>"000111101",
  41286=>"101001111",
  41287=>"111111001",
  41288=>"000000000",
  41289=>"111111111",
  41290=>"011000111",
  41291=>"111000000",
  41292=>"000100100",
  41293=>"110110110",
  41294=>"011000000",
  41295=>"111000101",
  41296=>"100111100",
  41297=>"111000000",
  41298=>"001000000",
  41299=>"111111101",
  41300=>"000000111",
  41301=>"011000000",
  41302=>"110110110",
  41303=>"110110000",
  41304=>"000000000",
  41305=>"011111000",
  41306=>"110111101",
  41307=>"100100111",
  41308=>"000000001",
  41309=>"111000010",
  41310=>"100000000",
  41311=>"000101001",
  41312=>"111011000",
  41313=>"101111111",
  41314=>"000000000",
  41315=>"000010000",
  41316=>"000001111",
  41317=>"111100111",
  41318=>"111101101",
  41319=>"000000100",
  41320=>"110110000",
  41321=>"000000000",
  41322=>"111111111",
  41323=>"000000110",
  41324=>"101000000",
  41325=>"100101111",
  41326=>"001011111",
  41327=>"111001111",
  41328=>"000000000",
  41329=>"000000000",
  41330=>"000110000",
  41331=>"011111001",
  41332=>"000000000",
  41333=>"000000000",
  41334=>"111101000",
  41335=>"000000000",
  41336=>"000010111",
  41337=>"011111111",
  41338=>"000000000",
  41339=>"000000010",
  41340=>"000000000",
  41341=>"111111001",
  41342=>"111111111",
  41343=>"001000011",
  41344=>"000000000",
  41345=>"110110111",
  41346=>"000000000",
  41347=>"001001111",
  41348=>"100101111",
  41349=>"000000100",
  41350=>"000000000",
  41351=>"111111111",
  41352=>"000000000",
  41353=>"111010000",
  41354=>"010111111",
  41355=>"111111110",
  41356=>"111011000",
  41357=>"111111000",
  41358=>"000000000",
  41359=>"100000001",
  41360=>"000111011",
  41361=>"011111111",
  41362=>"111000000",
  41363=>"111101100",
  41364=>"111100111",
  41365=>"000000000",
  41366=>"111001011",
  41367=>"100001011",
  41368=>"000000000",
  41369=>"110111111",
  41370=>"000111000",
  41371=>"011000000",
  41372=>"111111110",
  41373=>"111110111",
  41374=>"100000101",
  41375=>"111111111",
  41376=>"000000101",
  41377=>"111001000",
  41378=>"001001011",
  41379=>"111001000",
  41380=>"000011110",
  41381=>"010110000",
  41382=>"001111011",
  41383=>"111111110",
  41384=>"111111110",
  41385=>"111000000",
  41386=>"111000000",
  41387=>"100000101",
  41388=>"000011010",
  41389=>"110111010",
  41390=>"000000111",
  41391=>"110100111",
  41392=>"110110000",
  41393=>"111111111",
  41394=>"110001000",
  41395=>"111111111",
  41396=>"011000000",
  41397=>"001000100",
  41398=>"000111111",
  41399=>"000000000",
  41400=>"101111111",
  41401=>"111111111",
  41402=>"000000000",
  41403=>"101111111",
  41404=>"110000001",
  41405=>"111111111",
  41406=>"000000111",
  41407=>"011110000",
  41408=>"000000000",
  41409=>"111111111",
  41410=>"111111101",
  41411=>"000001111",
  41412=>"111011111",
  41413=>"000000000",
  41414=>"111111111",
  41415=>"000110111",
  41416=>"000000111",
  41417=>"000011110",
  41418=>"000000000",
  41419=>"000000000",
  41420=>"000001011",
  41421=>"001101100",
  41422=>"000010010",
  41423=>"000000111",
  41424=>"000000000",
  41425=>"011111111",
  41426=>"111111111",
  41427=>"001111111",
  41428=>"000101110",
  41429=>"100111110",
  41430=>"010010000",
  41431=>"000000000",
  41432=>"001100110",
  41433=>"100101000",
  41434=>"111111111",
  41435=>"100100111",
  41436=>"000101110",
  41437=>"001111111",
  41438=>"111110000",
  41439=>"001000111",
  41440=>"000111000",
  41441=>"001000000",
  41442=>"000000000",
  41443=>"111111111",
  41444=>"000011000",
  41445=>"100100111",
  41446=>"001000000",
  41447=>"111000000",
  41448=>"111111110",
  41449=>"000111000",
  41450=>"010011011",
  41451=>"011000000",
  41452=>"111111111",
  41453=>"011111110",
  41454=>"100111101",
  41455=>"000000000",
  41456=>"000000111",
  41457=>"111000110",
  41458=>"111111011",
  41459=>"001001000",
  41460=>"111010010",
  41461=>"000101111",
  41462=>"111001001",
  41463=>"110110010",
  41464=>"000000000",
  41465=>"000011000",
  41466=>"110010001",
  41467=>"111111111",
  41468=>"000000011",
  41469=>"111111110",
  41470=>"000100110",
  41471=>"111001011",
  41472=>"000000001",
  41473=>"000100101",
  41474=>"000111111",
  41475=>"110000000",
  41476=>"011110111",
  41477=>"111110000",
  41478=>"000000000",
  41479=>"011111111",
  41480=>"001000000",
  41481=>"111111111",
  41482=>"111111001",
  41483=>"110000000",
  41484=>"001001000",
  41485=>"010110111",
  41486=>"000000001",
  41487=>"001000000",
  41488=>"001000000",
  41489=>"111000000",
  41490=>"111111111",
  41491=>"000011111",
  41492=>"000110111",
  41493=>"000110000",
  41494=>"111111111",
  41495=>"001101000",
  41496=>"111111111",
  41497=>"000000100",
  41498=>"000000000",
  41499=>"111111111",
  41500=>"111111111",
  41501=>"111111111",
  41502=>"010111111",
  41503=>"111100000",
  41504=>"111111100",
  41505=>"000000000",
  41506=>"111111110",
  41507=>"111111110",
  41508=>"111011000",
  41509=>"000000011",
  41510=>"010000000",
  41511=>"101111111",
  41512=>"011001111",
  41513=>"000000000",
  41514=>"000111111",
  41515=>"010111110",
  41516=>"111111111",
  41517=>"111111111",
  41518=>"101000000",
  41519=>"110110111",
  41520=>"000111111",
  41521=>"100000000",
  41522=>"111110100",
  41523=>"100101110",
  41524=>"001111111",
  41525=>"000110110",
  41526=>"001001000",
  41527=>"100110111",
  41528=>"101110000",
  41529=>"000000000",
  41530=>"001001000",
  41531=>"000110110",
  41532=>"101001001",
  41533=>"011111111",
  41534=>"111111111",
  41535=>"101000000",
  41536=>"011111011",
  41537=>"000010111",
  41538=>"111111101",
  41539=>"011111000",
  41540=>"001001000",
  41541=>"000001000",
  41542=>"111111111",
  41543=>"111111111",
  41544=>"000000000",
  41545=>"111111111",
  41546=>"000000000",
  41547=>"000000000",
  41548=>"000001011",
  41549=>"111111000",
  41550=>"000101111",
  41551=>"110111111",
  41552=>"100000000",
  41553=>"010011000",
  41554=>"011111111",
  41555=>"010111111",
  41556=>"110111111",
  41557=>"000001000",
  41558=>"001000110",
  41559=>"000000000",
  41560=>"111110110",
  41561=>"000000000",
  41562=>"000000000",
  41563=>"111111111",
  41564=>"111111000",
  41565=>"110111010",
  41566=>"000000000",
  41567=>"000000000",
  41568=>"000000000",
  41569=>"000000101",
  41570=>"111110000",
  41571=>"000000000",
  41572=>"011000000",
  41573=>"000000010",
  41574=>"000000100",
  41575=>"111111111",
  41576=>"101001000",
  41577=>"111111111",
  41578=>"000000000",
  41579=>"000000000",
  41580=>"110000111",
  41581=>"000000000",
  41582=>"000000000",
  41583=>"111111111",
  41584=>"111111001",
  41585=>"110111111",
  41586=>"001111011",
  41587=>"010100100",
  41588=>"000000000",
  41589=>"001011100",
  41590=>"000000000",
  41591=>"110010000",
  41592=>"110111110",
  41593=>"111111000",
  41594=>"000000000",
  41595=>"010010111",
  41596=>"000110110",
  41597=>"000000000",
  41598=>"011110000",
  41599=>"000000000",
  41600=>"111111111",
  41601=>"111111000",
  41602=>"111111111",
  41603=>"110111110",
  41604=>"100000000",
  41605=>"000000100",
  41606=>"111110110",
  41607=>"111111100",
  41608=>"000000010",
  41609=>"111111111",
  41610=>"000000000",
  41611=>"011011011",
  41612=>"111111110",
  41613=>"000010010",
  41614=>"001011111",
  41615=>"101001011",
  41616=>"111111111",
  41617=>"111111111",
  41618=>"000000000",
  41619=>"111111111",
  41620=>"000000000",
  41621=>"110000000",
  41622=>"100111111",
  41623=>"000000100",
  41624=>"111010010",
  41625=>"010000001",
  41626=>"000110110",
  41627=>"101111111",
  41628=>"000000000",
  41629=>"101011011",
  41630=>"011111111",
  41631=>"111111011",
  41632=>"110000000",
  41633=>"010010111",
  41634=>"111111111",
  41635=>"111011000",
  41636=>"111110110",
  41637=>"111111111",
  41638=>"111111111",
  41639=>"110100110",
  41640=>"010110110",
  41641=>"111000000",
  41642=>"000000111",
  41643=>"000000000",
  41644=>"000000111",
  41645=>"000001000",
  41646=>"000000100",
  41647=>"011011000",
  41648=>"111111111",
  41649=>"100001000",
  41650=>"100111110",
  41651=>"111111000",
  41652=>"001100110",
  41653=>"110110000",
  41654=>"111110110",
  41655=>"100000000",
  41656=>"000000100",
  41657=>"111111011",
  41658=>"111111000",
  41659=>"100110000",
  41660=>"110111111",
  41661=>"000000110",
  41662=>"000000111",
  41663=>"000000000",
  41664=>"000000000",
  41665=>"001000000",
  41666=>"000000100",
  41667=>"000000000",
  41668=>"111111010",
  41669=>"101111111",
  41670=>"010011111",
  41671=>"001000111",
  41672=>"111101001",
  41673=>"101111111",
  41674=>"000000101",
  41675=>"000000000",
  41676=>"000101111",
  41677=>"101111111",
  41678=>"010111111",
  41679=>"000111111",
  41680=>"011111000",
  41681=>"000000000",
  41682=>"111000000",
  41683=>"111000000",
  41684=>"000000000",
  41685=>"110110000",
  41686=>"000000000",
  41687=>"010010000",
  41688=>"000101111",
  41689=>"111111111",
  41690=>"111101101",
  41691=>"100000000",
  41692=>"101000001",
  41693=>"111111000",
  41694=>"000000000",
  41695=>"000011111",
  41696=>"111111111",
  41697=>"000000000",
  41698=>"000000000",
  41699=>"100010110",
  41700=>"111111111",
  41701=>"111111110",
  41702=>"111111111",
  41703=>"000000000",
  41704=>"111111111",
  41705=>"111010011",
  41706=>"111010111",
  41707=>"101101111",
  41708=>"000111111",
  41709=>"000000111",
  41710=>"111111111",
  41711=>"101000000",
  41712=>"110110111",
  41713=>"000010010",
  41714=>"011011000",
  41715=>"110000000",
  41716=>"000000110",
  41717=>"000000000",
  41718=>"000000000",
  41719=>"010110010",
  41720=>"110111111",
  41721=>"000000100",
  41722=>"000000111",
  41723=>"000000000",
  41724=>"111100011",
  41725=>"111111111",
  41726=>"111111000",
  41727=>"000111000",
  41728=>"010000110",
  41729=>"011011111",
  41730=>"111111111",
  41731=>"110000000",
  41732=>"011010000",
  41733=>"101000100",
  41734=>"000000000",
  41735=>"110111111",
  41736=>"000000000",
  41737=>"010000010",
  41738=>"111111000",
  41739=>"000000000",
  41740=>"110110000",
  41741=>"101001011",
  41742=>"000000000",
  41743=>"010010000",
  41744=>"110000000",
  41745=>"001000000",
  41746=>"001101111",
  41747=>"111000000",
  41748=>"001000000",
  41749=>"000000111",
  41750=>"100110100",
  41751=>"000000000",
  41752=>"000001000",
  41753=>"101100111",
  41754=>"111111110",
  41755=>"110000000",
  41756=>"011000000",
  41757=>"000000011",
  41758=>"000000000",
  41759=>"111100111",
  41760=>"101001000",
  41761=>"111111111",
  41762=>"111111111",
  41763=>"100111111",
  41764=>"011111111",
  41765=>"011011111",
  41766=>"000010000",
  41767=>"000001100",
  41768=>"111011001",
  41769=>"111111111",
  41770=>"111111111",
  41771=>"000000000",
  41772=>"000010000",
  41773=>"010010011",
  41774=>"111111111",
  41775=>"000000000",
  41776=>"000111111",
  41777=>"000000000",
  41778=>"001111111",
  41779=>"000100111",
  41780=>"000000000",
  41781=>"111100000",
  41782=>"000010111",
  41783=>"111111110",
  41784=>"000000000",
  41785=>"000000000",
  41786=>"000000110",
  41787=>"000000000",
  41788=>"110110100",
  41789=>"000010000",
  41790=>"000000000",
  41791=>"000000000",
  41792=>"000000000",
  41793=>"000000000",
  41794=>"001000000",
  41795=>"111111111",
  41796=>"011111111",
  41797=>"110110000",
  41798=>"111101000",
  41799=>"000000000",
  41800=>"111111001",
  41801=>"000000110",
  41802=>"111010011",
  41803=>"011111111",
  41804=>"100100000",
  41805=>"010010110",
  41806=>"110110000",
  41807=>"000111111",
  41808=>"110000000",
  41809=>"110110000",
  41810=>"100110111",
  41811=>"111111111",
  41812=>"101000000",
  41813=>"001111011",
  41814=>"100111111",
  41815=>"111011100",
  41816=>"111101100",
  41817=>"100111111",
  41818=>"000000000",
  41819=>"100110100",
  41820=>"111111000",
  41821=>"001001101",
  41822=>"000001111",
  41823=>"000011111",
  41824=>"111111000",
  41825=>"000000000",
  41826=>"001011011",
  41827=>"000000000",
  41828=>"111010000",
  41829=>"000000000",
  41830=>"111111111",
  41831=>"000000010",
  41832=>"110111111",
  41833=>"000000000",
  41834=>"001111111",
  41835=>"001001000",
  41836=>"001101000",
  41837=>"010111111",
  41838=>"111011000",
  41839=>"111010111",
  41840=>"100111110",
  41841=>"111111100",
  41842=>"000000000",
  41843=>"111000000",
  41844=>"111111100",
  41845=>"000100100",
  41846=>"111111000",
  41847=>"100000100",
  41848=>"111111111",
  41849=>"100110000",
  41850=>"111111111",
  41851=>"000000000",
  41852=>"000000000",
  41853=>"111110000",
  41854=>"111111110",
  41855=>"100000100",
  41856=>"101011001",
  41857=>"111111000",
  41858=>"100000110",
  41859=>"010000000",
  41860=>"000000001",
  41861=>"100111111",
  41862=>"000000101",
  41863=>"101111111",
  41864=>"111111111",
  41865=>"000000000",
  41866=>"111111000",
  41867=>"000000000",
  41868=>"111111111",
  41869=>"000000001",
  41870=>"101111111",
  41871=>"100000000",
  41872=>"000000010",
  41873=>"010100100",
  41874=>"111010000",
  41875=>"010000000",
  41876=>"111111101",
  41877=>"011111010",
  41878=>"111110110",
  41879=>"101000100",
  41880=>"000000001",
  41881=>"001001111",
  41882=>"111111010",
  41883=>"101111111",
  41884=>"111111111",
  41885=>"001000000",
  41886=>"101001111",
  41887=>"000000000",
  41888=>"000000000",
  41889=>"001001100",
  41890=>"100110111",
  41891=>"010111111",
  41892=>"000010010",
  41893=>"110111001",
  41894=>"000000001",
  41895=>"000111100",
  41896=>"000000010",
  41897=>"110111010",
  41898=>"111111111",
  41899=>"000000110",
  41900=>"000000000",
  41901=>"100000000",
  41902=>"000111111",
  41903=>"111111111",
  41904=>"110111111",
  41905=>"000101001",
  41906=>"111000000",
  41907=>"010000000",
  41908=>"001000000",
  41909=>"000000000",
  41910=>"011111111",
  41911=>"101000001",
  41912=>"111111111",
  41913=>"000000000",
  41914=>"110110110",
  41915=>"111110110",
  41916=>"111111000",
  41917=>"100111101",
  41918=>"101111111",
  41919=>"110011001",
  41920=>"000000000",
  41921=>"111010000",
  41922=>"000000100",
  41923=>"000000000",
  41924=>"111000011",
  41925=>"100100111",
  41926=>"000000000",
  41927=>"011000000",
  41928=>"010000000",
  41929=>"100111111",
  41930=>"110111111",
  41931=>"011111111",
  41932=>"000111111",
  41933=>"010000000",
  41934=>"000000000",
  41935=>"111100000",
  41936=>"000111111",
  41937=>"111011000",
  41938=>"100111110",
  41939=>"000000000",
  41940=>"000000001",
  41941=>"110000000",
  41942=>"100000000",
  41943=>"000001001",
  41944=>"000000101",
  41945=>"100000111",
  41946=>"100001101",
  41947=>"000000000",
  41948=>"111111111",
  41949=>"111001011",
  41950=>"000000110",
  41951=>"000100001",
  41952=>"110110110",
  41953=>"001000000",
  41954=>"111111111",
  41955=>"111001010",
  41956=>"111111111",
  41957=>"000000000",
  41958=>"001110110",
  41959=>"000000111",
  41960=>"100010000",
  41961=>"000000000",
  41962=>"101000000",
  41963=>"111111000",
  41964=>"000001000",
  41965=>"011000000",
  41966=>"110000000",
  41967=>"000001001",
  41968=>"111000000",
  41969=>"000000000",
  41970=>"000000000",
  41971=>"001101111",
  41972=>"111111111",
  41973=>"000000011",
  41974=>"111111000",
  41975=>"110111110",
  41976=>"111000000",
  41977=>"000000010",
  41978=>"111000000",
  41979=>"111111111",
  41980=>"101101000",
  41981=>"111111111",
  41982=>"011000000",
  41983=>"111000000",
  41984=>"000111011",
  41985=>"000000001",
  41986=>"111111000",
  41987=>"000000111",
  41988=>"000001011",
  41989=>"000100111",
  41990=>"110000000",
  41991=>"000101101",
  41992=>"011111001",
  41993=>"000111111",
  41994=>"111000000",
  41995=>"000000000",
  41996=>"110000000",
  41997=>"100111000",
  41998=>"100001001",
  41999=>"000010010",
  42000=>"110111111",
  42001=>"010001011",
  42002=>"111111111",
  42003=>"001000000",
  42004=>"000100111",
  42005=>"111110000",
  42006=>"111110111",
  42007=>"111110110",
  42008=>"100111000",
  42009=>"100110100",
  42010=>"111111000",
  42011=>"101111111",
  42012=>"110111111",
  42013=>"000001101",
  42014=>"110000011",
  42015=>"000001000",
  42016=>"011000000",
  42017=>"111011000",
  42018=>"111111110",
  42019=>"001111110",
  42020=>"000000000",
  42021=>"000000000",
  42022=>"111111111",
  42023=>"011001000",
  42024=>"000100001",
  42025=>"111110000",
  42026=>"100000000",
  42027=>"001000001",
  42028=>"111111001",
  42029=>"000111111",
  42030=>"000010111",
  42031=>"000000000",
  42032=>"000000000",
  42033=>"110000000",
  42034=>"000000100",
  42035=>"010111110",
  42036=>"001000000",
  42037=>"111111100",
  42038=>"000000111",
  42039=>"101101101",
  42040=>"010000100",
  42041=>"100000001",
  42042=>"110000000",
  42043=>"111011011",
  42044=>"111000000",
  42045=>"110000100",
  42046=>"111111111",
  42047=>"000000000",
  42048=>"000000001",
  42049=>"000110111",
  42050=>"000110110",
  42051=>"000000000",
  42052=>"001001000",
  42053=>"111111111",
  42054=>"000000000",
  42055=>"111000001",
  42056=>"000000000",
  42057=>"111101111",
  42058=>"000111111",
  42059=>"001011011",
  42060=>"100100111",
  42061=>"011000000",
  42062=>"110100101",
  42063=>"001000000",
  42064=>"100111000",
  42065=>"001001001",
  42066=>"110111111",
  42067=>"111001101",
  42068=>"100111111",
  42069=>"000000000",
  42070=>"011111111",
  42071=>"111111110",
  42072=>"000000000",
  42073=>"111000000",
  42074=>"011011111",
  42075=>"100110111",
  42076=>"000011111",
  42077=>"111111111",
  42078=>"000001111",
  42079=>"000001011",
  42080=>"111111011",
  42081=>"100100000",
  42082=>"111001000",
  42083=>"110001011",
  42084=>"000000000",
  42085=>"001001010",
  42086=>"111111111",
  42087=>"111111111",
  42088=>"111110000",
  42089=>"000000001",
  42090=>"000010111",
  42091=>"000000000",
  42092=>"011001111",
  42093=>"000000101",
  42094=>"000000111",
  42095=>"111111001",
  42096=>"001001000",
  42097=>"111101111",
  42098=>"000101111",
  42099=>"100100111",
  42100=>"110110000",
  42101=>"111011001",
  42102=>"011010000",
  42103=>"111000000",
  42104=>"111000000",
  42105=>"111111111",
  42106=>"111000000",
  42107=>"100100100",
  42108=>"111011000",
  42109=>"110010000",
  42110=>"101100011",
  42111=>"010000000",
  42112=>"111011000",
  42113=>"110000000",
  42114=>"011001000",
  42115=>"001000000",
  42116=>"000111111",
  42117=>"111001000",
  42118=>"100111111",
  42119=>"000000000",
  42120=>"100100111",
  42121=>"000000001",
  42122=>"000000000",
  42123=>"000000000",
  42124=>"001000010",
  42125=>"000000000",
  42126=>"101100100",
  42127=>"000000000",
  42128=>"111011011",
  42129=>"000111111",
  42130=>"111101011",
  42131=>"111100000",
  42132=>"110111111",
  42133=>"100110100",
  42134=>"000111111",
  42135=>"111111111",
  42136=>"101000000",
  42137=>"111111111",
  42138=>"000101001",
  42139=>"000111010",
  42140=>"000000001",
  42141=>"000110110",
  42142=>"111000000",
  42143=>"000011111",
  42144=>"001000000",
  42145=>"111111000",
  42146=>"110010000",
  42147=>"010111111",
  42148=>"111011000",
  42149=>"000011001",
  42150=>"111100000",
  42151=>"111111111",
  42152=>"000000000",
  42153=>"000000101",
  42154=>"111111011",
  42155=>"010111111",
  42156=>"111111011",
  42157=>"000111111",
  42158=>"111101110",
  42159=>"000000010",
  42160=>"111011011",
  42161=>"110111110",
  42162=>"111010110",
  42163=>"001000111",
  42164=>"010111111",
  42165=>"001001000",
  42166=>"110000000",
  42167=>"110010001",
  42168=>"000011111",
  42169=>"111000000",
  42170=>"111001001",
  42171=>"111001000",
  42172=>"000100111",
  42173=>"000000111",
  42174=>"000000111",
  42175=>"001100100",
  42176=>"111000000",
  42177=>"110111000",
  42178=>"110100000",
  42179=>"111000000",
  42180=>"111111111",
  42181=>"001000000",
  42182=>"001101001",
  42183=>"000101000",
  42184=>"000110110",
  42185=>"000000000",
  42186=>"110000000",
  42187=>"111111111",
  42188=>"110000000",
  42189=>"000000000",
  42190=>"010000000",
  42191=>"111001001",
  42192=>"111111111",
  42193=>"010010010",
  42194=>"111111011",
  42195=>"000000000",
  42196=>"111111111",
  42197=>"110000000",
  42198=>"111010010",
  42199=>"001111111",
  42200=>"000111111",
  42201=>"000000000",
  42202=>"111111000",
  42203=>"001000111",
  42204=>"110111111",
  42205=>"111111111",
  42206=>"110100100",
  42207=>"100000111",
  42208=>"001111111",
  42209=>"001000000",
  42210=>"111111010",
  42211=>"111111001",
  42212=>"100000000",
  42213=>"010111110",
  42214=>"100111000",
  42215=>"000000000",
  42216=>"111111111",
  42217=>"101011011",
  42218=>"000000011",
  42219=>"000000110",
  42220=>"111100000",
  42221=>"011001001",
  42222=>"111001000",
  42223=>"110010000",
  42224=>"010111111",
  42225=>"111001001",
  42226=>"100000001",
  42227=>"111001000",
  42228=>"000000111",
  42229=>"001010111",
  42230=>"000111110",
  42231=>"000000000",
  42232=>"111111010",
  42233=>"111111000",
  42234=>"000000000",
  42235=>"111111111",
  42236=>"100111011",
  42237=>"100000000",
  42238=>"110000001",
  42239=>"000000011",
  42240=>"100000000",
  42241=>"110111111",
  42242=>"100000000",
  42243=>"110000000",
  42244=>"000100100",
  42245=>"001000111",
  42246=>"111111000",
  42247=>"001000000",
  42248=>"000100000",
  42249=>"010000000",
  42250=>"000110111",
  42251=>"000000000",
  42252=>"111111111",
  42253=>"000011111",
  42254=>"111111111",
  42255=>"001000000",
  42256=>"010001101",
  42257=>"110100101",
  42258=>"111100100",
  42259=>"000011111",
  42260=>"011111111",
  42261=>"001111111",
  42262=>"100100100",
  42263=>"110000010",
  42264=>"101111111",
  42265=>"111000000",
  42266=>"111111111",
  42267=>"000001111",
  42268=>"111100100",
  42269=>"001000111",
  42270=>"011011011",
  42271=>"110100000",
  42272=>"100110111",
  42273=>"000110111",
  42274=>"111111111",
  42275=>"111000100",
  42276=>"010010000",
  42277=>"110000001",
  42278=>"111000000",
  42279=>"001000111",
  42280=>"100111111",
  42281=>"110000010",
  42282=>"100000000",
  42283=>"111100100",
  42284=>"110100000",
  42285=>"001001111",
  42286=>"000111000",
  42287=>"110111010",
  42288=>"111111111",
  42289=>"000000100",
  42290=>"000000000",
  42291=>"101111100",
  42292=>"000000000",
  42293=>"100100000",
  42294=>"101111000",
  42295=>"101101010",
  42296=>"001000011",
  42297=>"001000000",
  42298=>"111110000",
  42299=>"001000111",
  42300=>"100100000",
  42301=>"110000000",
  42302=>"000000001",
  42303=>"100110111",
  42304=>"111111000",
  42305=>"110010111",
  42306=>"000000000",
  42307=>"111010000",
  42308=>"000100100",
  42309=>"000000110",
  42310=>"010000000",
  42311=>"111111110",
  42312=>"110111110",
  42313=>"000000000",
  42314=>"100100010",
  42315=>"011011011",
  42316=>"110111101",
  42317=>"111111111",
  42318=>"000000000",
  42319=>"000100100",
  42320=>"110110100",
  42321=>"111001000",
  42322=>"111111111",
  42323=>"110111111",
  42324=>"111000000",
  42325=>"001000011",
  42326=>"111111111",
  42327=>"111110000",
  42328=>"111000000",
  42329=>"010000011",
  42330=>"101100110",
  42331=>"001001111",
  42332=>"011010000",
  42333=>"000000000",
  42334=>"100100100",
  42335=>"001011001",
  42336=>"100111111",
  42337=>"111111111",
  42338=>"000001001",
  42339=>"110110110",
  42340=>"110110110",
  42341=>"100000000",
  42342=>"001101111",
  42343=>"111111111",
  42344=>"101101111",
  42345=>"001001111",
  42346=>"111001100",
  42347=>"111111110",
  42348=>"000111111",
  42349=>"111001111",
  42350=>"000000000",
  42351=>"000000010",
  42352=>"111111111",
  42353=>"000000111",
  42354=>"000000011",
  42355=>"111000000",
  42356=>"111111111",
  42357=>"100000000",
  42358=>"000111111",
  42359=>"000101100",
  42360=>"111111000",
  42361=>"000011000",
  42362=>"000000000",
  42363=>"100110000",
  42364=>"111110000",
  42365=>"000001011",
  42366=>"000000001",
  42367=>"110100111",
  42368=>"110011011",
  42369=>"001001001",
  42370=>"110111111",
  42371=>"000000000",
  42372=>"110111111",
  42373=>"011111101",
  42374=>"000110111",
  42375=>"111000001",
  42376=>"100000000",
  42377=>"000000000",
  42378=>"111111110",
  42379=>"001001001",
  42380=>"111111111",
  42381=>"111001000",
  42382=>"000000110",
  42383=>"010010000",
  42384=>"000011111",
  42385=>"111111111",
  42386=>"011110110",
  42387=>"100100110",
  42388=>"111111111",
  42389=>"000010000",
  42390=>"111000000",
  42391=>"111011011",
  42392=>"111111001",
  42393=>"111111111",
  42394=>"100000000",
  42395=>"111111111",
  42396=>"111110110",
  42397=>"000000000",
  42398=>"111111111",
  42399=>"111000000",
  42400=>"111111111",
  42401=>"100100001",
  42402=>"110000000",
  42403=>"111111010",
  42404=>"111111000",
  42405=>"000011111",
  42406=>"110110111",
  42407=>"000111111",
  42408=>"000000010",
  42409=>"111111111",
  42410=>"000001000",
  42411=>"111111000",
  42412=>"000000100",
  42413=>"111111000",
  42414=>"110000001",
  42415=>"111110110",
  42416=>"000000000",
  42417=>"000000000",
  42418=>"000010000",
  42419=>"010000000",
  42420=>"111011000",
  42421=>"111000011",
  42422=>"111000001",
  42423=>"000000000",
  42424=>"110011111",
  42425=>"000000111",
  42426=>"000000111",
  42427=>"110000000",
  42428=>"000000000",
  42429=>"110111001",
  42430=>"111100000",
  42431=>"110100000",
  42432=>"000000000",
  42433=>"110000000",
  42434=>"000000000",
  42435=>"100111000",
  42436=>"111100100",
  42437=>"000000000",
  42438=>"001000000",
  42439=>"111111111",
  42440=>"000000000",
  42441=>"101000111",
  42442=>"000000000",
  42443=>"000000111",
  42444=>"100111111",
  42445=>"010111111",
  42446=>"000111011",
  42447=>"111111111",
  42448=>"011000000",
  42449=>"010000000",
  42450=>"000111111",
  42451=>"000110100",
  42452=>"000001111",
  42453=>"100000111",
  42454=>"100100110",
  42455=>"000000000",
  42456=>"101111100",
  42457=>"100110111",
  42458=>"000110000",
  42459=>"101000000",
  42460=>"010111010",
  42461=>"000000000",
  42462=>"000000101",
  42463=>"110111011",
  42464=>"111111011",
  42465=>"000000000",
  42466=>"110000000",
  42467=>"000000000",
  42468=>"110000111",
  42469=>"000001000",
  42470=>"111111111",
  42471=>"011111111",
  42472=>"111111010",
  42473=>"010111111",
  42474=>"001111111",
  42475=>"000111111",
  42476=>"111011000",
  42477=>"011000110",
  42478=>"001000000",
  42479=>"111111100",
  42480=>"111011000",
  42481=>"111110000",
  42482=>"111110110",
  42483=>"111000000",
  42484=>"101000000",
  42485=>"000000000",
  42486=>"000000010",
  42487=>"001000110",
  42488=>"110100100",
  42489=>"100100100",
  42490=>"000000001",
  42491=>"000000000",
  42492=>"111111111",
  42493=>"111000000",
  42494=>"111111110",
  42495=>"000000000",
  42496=>"000000001",
  42497=>"000000000",
  42498=>"111111111",
  42499=>"101000000",
  42500=>"000000000",
  42501=>"011000111",
  42502=>"000000000",
  42503=>"111111111",
  42504=>"111110000",
  42505=>"111111111",
  42506=>"000000000",
  42507=>"111010000",
  42508=>"100100000",
  42509=>"111111111",
  42510=>"000100111",
  42511=>"000000000",
  42512=>"000000000",
  42513=>"011111111",
  42514=>"000100111",
  42515=>"000011111",
  42516=>"111101101",
  42517=>"000000001",
  42518=>"000000000",
  42519=>"111111111",
  42520=>"011010000",
  42521=>"001110110",
  42522=>"001000111",
  42523=>"111001111",
  42524=>"000100000",
  42525=>"000000000",
  42526=>"010011111",
  42527=>"000000000",
  42528=>"001001001",
  42529=>"111111111",
  42530=>"110001111",
  42531=>"110110010",
  42532=>"000000000",
  42533=>"001011111",
  42534=>"111111111",
  42535=>"000111111",
  42536=>"001001111",
  42537=>"000000000",
  42538=>"000000000",
  42539=>"110111111",
  42540=>"111111011",
  42541=>"111110111",
  42542=>"111000011",
  42543=>"010110111",
  42544=>"000001001",
  42545=>"001001000",
  42546=>"000111011",
  42547=>"111111111",
  42548=>"101111100",
  42549=>"110000000",
  42550=>"000000000",
  42551=>"011011111",
  42552=>"111110110",
  42553=>"111111111",
  42554=>"000000000",
  42555=>"111111000",
  42556=>"000000000",
  42557=>"101111111",
  42558=>"011101111",
  42559=>"000100000",
  42560=>"111111111",
  42561=>"000001000",
  42562=>"111111000",
  42563=>"000000110",
  42564=>"010011011",
  42565=>"011001000",
  42566=>"111001001",
  42567=>"111111111",
  42568=>"001011011",
  42569=>"000000011",
  42570=>"111111010",
  42571=>"111000000",
  42572=>"100011010",
  42573=>"111101101",
  42574=>"001000000",
  42575=>"110111100",
  42576=>"000000000",
  42577=>"001110110",
  42578=>"111100001",
  42579=>"010011111",
  42580=>"000000000",
  42581=>"011111111",
  42582=>"111000000",
  42583=>"111111111",
  42584=>"100100000",
  42585=>"001001000",
  42586=>"111111000",
  42587=>"001000001",
  42588=>"000000110",
  42589=>"111111111",
  42590=>"000000000",
  42591=>"000000000",
  42592=>"111111010",
  42593=>"111111000",
  42594=>"001101001",
  42595=>"000000111",
  42596=>"100111111",
  42597=>"011000000",
  42598=>"000001000",
  42599=>"100100101",
  42600=>"111111000",
  42601=>"111111111",
  42602=>"111111000",
  42603=>"000000000",
  42604=>"000000000",
  42605=>"101000000",
  42606=>"000101000",
  42607=>"101101001",
  42608=>"000000000",
  42609=>"111111011",
  42610=>"001001001",
  42611=>"111001001",
  42612=>"011001111",
  42613=>"000000000",
  42614=>"000000011",
  42615=>"111011001",
  42616=>"000000000",
  42617=>"000000000",
  42618=>"111111000",
  42619=>"000000000",
  42620=>"111111110",
  42621=>"111000000",
  42622=>"000000100",
  42623=>"000000000",
  42624=>"100000000",
  42625=>"000111010",
  42626=>"111111111",
  42627=>"011111100",
  42628=>"111111111",
  42629=>"000000000",
  42630=>"000000000",
  42631=>"000000000",
  42632=>"110111111",
  42633=>"001000000",
  42634=>"001110110",
  42635=>"011010000",
  42636=>"111111111",
  42637=>"000000000",
  42638=>"110111111",
  42639=>"000111000",
  42640=>"111111111",
  42641=>"000000001",
  42642=>"000000000",
  42643=>"111110000",
  42644=>"000010010",
  42645=>"000001111",
  42646=>"010111111",
  42647=>"000000000",
  42648=>"111111111",
  42649=>"000000000",
  42650=>"111001011",
  42651=>"000111111",
  42652=>"000000110",
  42653=>"000000101",
  42654=>"000010110",
  42655=>"110110111",
  42656=>"111111111",
  42657=>"111000000",
  42658=>"111101111",
  42659=>"000000011",
  42660=>"000011001",
  42661=>"000000111",
  42662=>"110010000",
  42663=>"011011011",
  42664=>"110010010",
  42665=>"010100100",
  42666=>"111111111",
  42667=>"111000100",
  42668=>"000000000",
  42669=>"000000000",
  42670=>"000000100",
  42671=>"101000000",
  42672=>"000000000",
  42673=>"001111101",
  42674=>"010000001",
  42675=>"000100110",
  42676=>"000000000",
  42677=>"111100100",
  42678=>"000000001",
  42679=>"111111000",
  42680=>"001001110",
  42681=>"000111111",
  42682=>"111111001",
  42683=>"001001001",
  42684=>"111111111",
  42685=>"000000000",
  42686=>"000000000",
  42687=>"111111111",
  42688=>"000000000",
  42689=>"100000110",
  42690=>"000000111",
  42691=>"101101111",
  42692=>"001111000",
  42693=>"111111111",
  42694=>"010010000",
  42695=>"000100000",
  42696=>"000000000",
  42697=>"011111111",
  42698=>"011011011",
  42699=>"101111111",
  42700=>"111110011",
  42701=>"000001111",
  42702=>"111100111",
  42703=>"011110000",
  42704=>"010010001",
  42705=>"000000000",
  42706=>"111111000",
  42707=>"000000000",
  42708=>"000000000",
  42709=>"111111111",
  42710=>"000000010",
  42711=>"111111011",
  42712=>"000101111",
  42713=>"111111110",
  42714=>"001001001",
  42715=>"000110111",
  42716=>"001001111",
  42717=>"111111111",
  42718=>"010110111",
  42719=>"010000000",
  42720=>"000000001",
  42721=>"000100001",
  42722=>"111001111",
  42723=>"100100001",
  42724=>"111111111",
  42725=>"111111110",
  42726=>"000000011",
  42727=>"000000100",
  42728=>"011000000",
  42729=>"101011001",
  42730=>"111110101",
  42731=>"111110111",
  42732=>"111110000",
  42733=>"000111111",
  42734=>"110110111",
  42735=>"010110111",
  42736=>"000000000",
  42737=>"111101000",
  42738=>"100101000",
  42739=>"111101001",
  42740=>"000000000",
  42741=>"000000000",
  42742=>"000000111",
  42743=>"111000000",
  42744=>"000000000",
  42745=>"000000000",
  42746=>"101001001",
  42747=>"110000000",
  42748=>"100110100",
  42749=>"110110010",
  42750=>"000000000",
  42751=>"111001100",
  42752=>"111111111",
  42753=>"011011011",
  42754=>"110000000",
  42755=>"000000000",
  42756=>"000000000",
  42757=>"000000001",
  42758=>"100100000",
  42759=>"111111000",
  42760=>"111111111",
  42761=>"111111100",
  42762=>"000000100",
  42763=>"000100111",
  42764=>"100000000",
  42765=>"111111111",
  42766=>"000000100",
  42767=>"000000000",
  42768=>"000000000",
  42769=>"111101111",
  42770=>"011000000",
  42771=>"010010000",
  42772=>"000000000",
  42773=>"111111100",
  42774=>"011111010",
  42775=>"111100111",
  42776=>"111101111",
  42777=>"000000000",
  42778=>"111111111",
  42779=>"110100000",
  42780=>"000111111",
  42781=>"101111111",
  42782=>"000000100",
  42783=>"101011111",
  42784=>"111001011",
  42785=>"111111011",
  42786=>"000000000",
  42787=>"001111111",
  42788=>"000111111",
  42789=>"111111000",
  42790=>"000000000",
  42791=>"000101101",
  42792=>"111001111",
  42793=>"001111011",
  42794=>"111111111",
  42795=>"000000000",
  42796=>"001100100",
  42797=>"110110111",
  42798=>"000111000",
  42799=>"110100110",
  42800=>"111111111",
  42801=>"111111111",
  42802=>"110111111",
  42803=>"111111111",
  42804=>"111111010",
  42805=>"110100100",
  42806=>"111010010",
  42807=>"001000000",
  42808=>"000010000",
  42809=>"111111111",
  42810=>"000000000",
  42811=>"000000000",
  42812=>"011011111",
  42813=>"001001000",
  42814=>"111100111",
  42815=>"110100000",
  42816=>"000000010",
  42817=>"111111111",
  42818=>"000011111",
  42819=>"010110000",
  42820=>"001000000",
  42821=>"111111111",
  42822=>"000011111",
  42823=>"000000000",
  42824=>"000000001",
  42825=>"111011001",
  42826=>"011000100",
  42827=>"110110000",
  42828=>"000001111",
  42829=>"111111111",
  42830=>"111111100",
  42831=>"000000110",
  42832=>"010000000",
  42833=>"100000000",
  42834=>"111111000",
  42835=>"111111111",
  42836=>"000000111",
  42837=>"111111011",
  42838=>"111111000",
  42839=>"111101111",
  42840=>"000100000",
  42841=>"111011001",
  42842=>"110111100",
  42843=>"000101011",
  42844=>"000000000",
  42845=>"000000111",
  42846=>"011111001",
  42847=>"001001111",
  42848=>"000000000",
  42849=>"111111111",
  42850=>"110110110",
  42851=>"000000001",
  42852=>"110110110",
  42853=>"000000000",
  42854=>"111110111",
  42855=>"111111111",
  42856=>"010010010",
  42857=>"111101000",
  42858=>"111111011",
  42859=>"110010111",
  42860=>"111111111",
  42861=>"111111000",
  42862=>"111011000",
  42863=>"000000001",
  42864=>"111011111",
  42865=>"111111010",
  42866=>"000000000",
  42867=>"111111111",
  42868=>"101101000",
  42869=>"100100100",
  42870=>"111111000",
  42871=>"100111110",
  42872=>"000010010",
  42873=>"000000111",
  42874=>"010000000",
  42875=>"111111111",
  42876=>"101101101",
  42877=>"001011111",
  42878=>"000000000",
  42879=>"111111111",
  42880=>"011000000",
  42881=>"000000000",
  42882=>"111110010",
  42883=>"000000000",
  42884=>"100000000",
  42885=>"000100000",
  42886=>"111111101",
  42887=>"110011001",
  42888=>"111111111",
  42889=>"111111111",
  42890=>"110111000",
  42891=>"111111111",
  42892=>"111111111",
  42893=>"000111111",
  42894=>"101111111",
  42895=>"000000000",
  42896=>"000011000",
  42897=>"101100000",
  42898=>"111111111",
  42899=>"111111011",
  42900=>"101101111",
  42901=>"000100110",
  42902=>"111111111",
  42903=>"110110110",
  42904=>"000000000",
  42905=>"000000000",
  42906=>"111111111",
  42907=>"111111111",
  42908=>"111111111",
  42909=>"000000000",
  42910=>"111111111",
  42911=>"000000000",
  42912=>"100100000",
  42913=>"111111111",
  42914=>"010001111",
  42915=>"111111001",
  42916=>"011001111",
  42917=>"100100000",
  42918=>"111111110",
  42919=>"000100111",
  42920=>"111000000",
  42921=>"110111111",
  42922=>"110000001",
  42923=>"011000000",
  42924=>"111000111",
  42925=>"000000000",
  42926=>"111111111",
  42927=>"111111111",
  42928=>"001000000",
  42929=>"000000000",
  42930=>"110111000",
  42931=>"111111111",
  42932=>"000000000",
  42933=>"111111111",
  42934=>"111111111",
  42935=>"000000100",
  42936=>"000000000",
  42937=>"000000000",
  42938=>"111101100",
  42939=>"000000000",
  42940=>"111111111",
  42941=>"111111110",
  42942=>"000000000",
  42943=>"010011011",
  42944=>"000000000",
  42945=>"000000000",
  42946=>"011010000",
  42947=>"111111000",
  42948=>"010111111",
  42949=>"110110110",
  42950=>"000000000",
  42951=>"111011010",
  42952=>"000000010",
  42953=>"000000000",
  42954=>"111111000",
  42955=>"000110111",
  42956=>"011001000",
  42957=>"111111111",
  42958=>"011111111",
  42959=>"001001111",
  42960=>"100110111",
  42961=>"111101111",
  42962=>"111111111",
  42963=>"000000100",
  42964=>"000100110",
  42965=>"111111001",
  42966=>"000000000",
  42967=>"001000001",
  42968=>"000000000",
  42969=>"000000000",
  42970=>"000001111",
  42971=>"111110000",
  42972=>"000000001",
  42973=>"111111111",
  42974=>"111111111",
  42975=>"000010000",
  42976=>"000010000",
  42977=>"111111011",
  42978=>"100100100",
  42979=>"001010111",
  42980=>"111111111",
  42981=>"111111000",
  42982=>"001001001",
  42983=>"111111111",
  42984=>"111110110",
  42985=>"000000101",
  42986=>"000000000",
  42987=>"111111011",
  42988=>"000000110",
  42989=>"001000000",
  42990=>"000100111",
  42991=>"011000110",
  42992=>"011011011",
  42993=>"111100000",
  42994=>"111100111",
  42995=>"000110100",
  42996=>"000000000",
  42997=>"000000111",
  42998=>"000001111",
  42999=>"010000000",
  43000=>"000000001",
  43001=>"100100100",
  43002=>"111011011",
  43003=>"000000000",
  43004=>"111111111",
  43005=>"000000111",
  43006=>"000000000",
  43007=>"100000000",
  43008=>"111111111",
  43009=>"111111111",
  43010=>"111000000",
  43011=>"110100111",
  43012=>"000010111",
  43013=>"000111111",
  43014=>"001111111",
  43015=>"001000000",
  43016=>"000000010",
  43017=>"111111000",
  43018=>"111011000",
  43019=>"110010010",
  43020=>"000001001",
  43021=>"111111111",
  43022=>"111111111",
  43023=>"111111111",
  43024=>"101101111",
  43025=>"010000011",
  43026=>"111111111",
  43027=>"001001001",
  43028=>"000000000",
  43029=>"000000000",
  43030=>"111000000",
  43031=>"001001011",
  43032=>"111111111",
  43033=>"000000000",
  43034=>"111000000",
  43035=>"000000110",
  43036=>"000000000",
  43037=>"111110111",
  43038=>"001101100",
  43039=>"111111111",
  43040=>"111111111",
  43041=>"111110110",
  43042=>"000000000",
  43043=>"100110110",
  43044=>"111111111",
  43045=>"000000000",
  43046=>"111111111",
  43047=>"110111111",
  43048=>"010000111",
  43049=>"000000000",
  43050=>"000000000",
  43051=>"111111110",
  43052=>"100100111",
  43053=>"100011111",
  43054=>"111111111",
  43055=>"110111111",
  43056=>"111111111",
  43057=>"000000000",
  43058=>"110111001",
  43059=>"000001011",
  43060=>"111101001",
  43061=>"011111011",
  43062=>"000000000",
  43063=>"111000000",
  43064=>"011111110",
  43065=>"000001111",
  43066=>"011010000",
  43067=>"111111111",
  43068=>"111111101",
  43069=>"111111111",
  43070=>"111111111",
  43071=>"111111111",
  43072=>"111001001",
  43073=>"000000001",
  43074=>"011011111",
  43075=>"001000000",
  43076=>"011111000",
  43077=>"111111110",
  43078=>"111110100",
  43079=>"111111111",
  43080=>"111010011",
  43081=>"111111111",
  43082=>"000000001",
  43083=>"111001000",
  43084=>"111111011",
  43085=>"000000111",
  43086=>"000111111",
  43087=>"100110111",
  43088=>"000000000",
  43089=>"000101000",
  43090=>"000000000",
  43091=>"000000001",
  43092=>"111111111",
  43093=>"000000010",
  43094=>"000000000",
  43095=>"111111111",
  43096=>"000000000",
  43097=>"111000000",
  43098=>"111111111",
  43099=>"000000001",
  43100=>"110110000",
  43101=>"000000000",
  43102=>"000101111",
  43103=>"010001000",
  43104=>"000000000",
  43105=>"000000000",
  43106=>"000000101",
  43107=>"000000001",
  43108=>"000000000",
  43109=>"111110011",
  43110=>"111111000",
  43111=>"111111111",
  43112=>"000000000",
  43113=>"000111111",
  43114=>"011000000",
  43115=>"000000000",
  43116=>"111001001",
  43117=>"111000000",
  43118=>"001111111",
  43119=>"110111000",
  43120=>"000111111",
  43121=>"011111111",
  43122=>"111111101",
  43123=>"111111111",
  43124=>"111100100",
  43125=>"010011011",
  43126=>"111100110",
  43127=>"011011111",
  43128=>"111110010",
  43129=>"000000000",
  43130=>"000000000",
  43131=>"111101000",
  43132=>"110111111",
  43133=>"000000000",
  43134=>"001001001",
  43135=>"000000000",
  43136=>"000000000",
  43137=>"111111000",
  43138=>"101001001",
  43139=>"111101001",
  43140=>"000000000",
  43141=>"111110110",
  43142=>"111110110",
  43143=>"001111111",
  43144=>"000000000",
  43145=>"111111111",
  43146=>"111111110",
  43147=>"010000000",
  43148=>"000100111",
  43149=>"000000000",
  43150=>"101000000",
  43151=>"111111101",
  43152=>"110111111",
  43153=>"111111001",
  43154=>"000000000",
  43155=>"000010000",
  43156=>"000000100",
  43157=>"000100111",
  43158=>"000000000",
  43159=>"111101000",
  43160=>"111111110",
  43161=>"110000010",
  43162=>"111011000",
  43163=>"101000101",
  43164=>"110000000",
  43165=>"000000000",
  43166=>"000000000",
  43167=>"111111111",
  43168=>"000000000",
  43169=>"000000011",
  43170=>"000000000",
  43171=>"000000100",
  43172=>"000000000",
  43173=>"000001111",
  43174=>"000000000",
  43175=>"110110110",
  43176=>"000000000",
  43177=>"000000000",
  43178=>"111111111",
  43179=>"111111111",
  43180=>"011010000",
  43181=>"111000001",
  43182=>"111111110",
  43183=>"100001001",
  43184=>"111111111",
  43185=>"000000000",
  43186=>"110111110",
  43187=>"000000010",
  43188=>"000000000",
  43189=>"001001111",
  43190=>"000000000",
  43191=>"000111111",
  43192=>"111111111",
  43193=>"111111111",
  43194=>"000000000",
  43195=>"100000111",
  43196=>"111110110",
  43197=>"111100100",
  43198=>"000000000",
  43199=>"111000101",
  43200=>"111111111",
  43201=>"001000000",
  43202=>"111111111",
  43203=>"000111110",
  43204=>"111111111",
  43205=>"111111000",
  43206=>"100100100",
  43207=>"111111110",
  43208=>"111111111",
  43209=>"000000000",
  43210=>"000000000",
  43211=>"101000000",
  43212=>"000000001",
  43213=>"100001001",
  43214=>"100001000",
  43215=>"111111111",
  43216=>"010111111",
  43217=>"000111110",
  43218=>"000111111",
  43219=>"111000111",
  43220=>"000011000",
  43221=>"001001000",
  43222=>"000000010",
  43223=>"101001000",
  43224=>"111111111",
  43225=>"011111111",
  43226=>"000000000",
  43227=>"000000000",
  43228=>"111111100",
  43229=>"000000000",
  43230=>"000011110",
  43231=>"000100000",
  43232=>"110111111",
  43233=>"000000000",
  43234=>"111111111",
  43235=>"111111111",
  43236=>"001001111",
  43237=>"000000000",
  43238=>"001111100",
  43239=>"010111111",
  43240=>"000000111",
  43241=>"000011111",
  43242=>"001000000",
  43243=>"000000100",
  43244=>"000110011",
  43245=>"000000000",
  43246=>"000000000",
  43247=>"000010111",
  43248=>"000000000",
  43249=>"111111111",
  43250=>"011111011",
  43251=>"000011000",
  43252=>"111000000",
  43253=>"000000000",
  43254=>"011000110",
  43255=>"111111111",
  43256=>"000100100",
  43257=>"110110110",
  43258=>"110000000",
  43259=>"000000000",
  43260=>"001000001",
  43261=>"100110111",
  43262=>"111111100",
  43263=>"001011111",
  43264=>"000111100",
  43265=>"000100110",
  43266=>"000000000",
  43267=>"000111111",
  43268=>"000000000",
  43269=>"000011011",
  43270=>"000000000",
  43271=>"111000000",
  43272=>"001111111",
  43273=>"111111111",
  43274=>"110100101",
  43275=>"001000001",
  43276=>"100000110",
  43277=>"111111000",
  43278=>"000000000",
  43279=>"111111100",
  43280=>"000001111",
  43281=>"000011000",
  43282=>"101111111",
  43283=>"100000010",
  43284=>"000000000",
  43285=>"001011111",
  43286=>"110111111",
  43287=>"111111100",
  43288=>"000000011",
  43289=>"111111111",
  43290=>"111111111",
  43291=>"011010000",
  43292=>"001001000",
  43293=>"000011111",
  43294=>"000000000",
  43295=>"100111001",
  43296=>"000000000",
  43297=>"111111111",
  43298=>"110110110",
  43299=>"111111110",
  43300=>"001000000",
  43301=>"100101001",
  43302=>"111100000",
  43303=>"111011011",
  43304=>"111111100",
  43305=>"111111111",
  43306=>"100000000",
  43307=>"001101011",
  43308=>"111001000",
  43309=>"000000000",
  43310=>"000000000",
  43311=>"000000000",
  43312=>"011001111",
  43313=>"111111101",
  43314=>"111111111",
  43315=>"100110000",
  43316=>"000000000",
  43317=>"000000011",
  43318=>"000000000",
  43319=>"000001001",
  43320=>"000000000",
  43321=>"000110111",
  43322=>"010110111",
  43323=>"111111111",
  43324=>"001001011",
  43325=>"110000000",
  43326=>"111111111",
  43327=>"111111000",
  43328=>"000110111",
  43329=>"110111101",
  43330=>"111111111",
  43331=>"111111111",
  43332=>"111100000",
  43333=>"110100000",
  43334=>"000000000",
  43335=>"010000000",
  43336=>"110100000",
  43337=>"111111111",
  43338=>"111111110",
  43339=>"111010001",
  43340=>"000000000",
  43341=>"111100111",
  43342=>"000000000",
  43343=>"000000000",
  43344=>"100110000",
  43345=>"001100111",
  43346=>"111000000",
  43347=>"111111111",
  43348=>"111111000",
  43349=>"001011111",
  43350=>"111000001",
  43351=>"000000000",
  43352=>"000000111",
  43353=>"111111001",
  43354=>"111011000",
  43355=>"111100100",
  43356=>"000000111",
  43357=>"111111111",
  43358=>"000001001",
  43359=>"000110100",
  43360=>"011000001",
  43361=>"000000000",
  43362=>"011000011",
  43363=>"111111111",
  43364=>"111111111",
  43365=>"000000000",
  43366=>"000100000",
  43367=>"001001101",
  43368=>"000000000",
  43369=>"110111100",
  43370=>"101110111",
  43371=>"100000000",
  43372=>"111010000",
  43373=>"000001111",
  43374=>"010111111",
  43375=>"000110000",
  43376=>"000000000",
  43377=>"000000000",
  43378=>"111111111",
  43379=>"000101111",
  43380=>"111111111",
  43381=>"011001110",
  43382=>"111111111",
  43383=>"000000000",
  43384=>"111000111",
  43385=>"000000000",
  43386=>"000000101",
  43387=>"000101111",
  43388=>"111111111",
  43389=>"111101000",
  43390=>"001001001",
  43391=>"000000000",
  43392=>"000000111",
  43393=>"011000010",
  43394=>"011011111",
  43395=>"000000000",
  43396=>"000000000",
  43397=>"111111111",
  43398=>"011000100",
  43399=>"100111111",
  43400=>"001011111",
  43401=>"111111111",
  43402=>"001000100",
  43403=>"111000000",
  43404=>"000001111",
  43405=>"111111111",
  43406=>"000111111",
  43407=>"000000000",
  43408=>"111111111",
  43409=>"110111111",
  43410=>"001011111",
  43411=>"000000000",
  43412=>"111111111",
  43413=>"000000001",
  43414=>"101001000",
  43415=>"010001011",
  43416=>"000000110",
  43417=>"111111111",
  43418=>"111111111",
  43419=>"000000001",
  43420=>"000100111",
  43421=>"010000011",
  43422=>"000000000",
  43423=>"110110111",
  43424=>"111111111",
  43425=>"001001001",
  43426=>"111100101",
  43427=>"000000110",
  43428=>"111001111",
  43429=>"001111101",
  43430=>"111111111",
  43431=>"000000110",
  43432=>"001001000",
  43433=>"000000000",
  43434=>"011000000",
  43435=>"100111011",
  43436=>"110101111",
  43437=>"111011001",
  43438=>"010111001",
  43439=>"000000111",
  43440=>"000000000",
  43441=>"111111110",
  43442=>"111111001",
  43443=>"111111111",
  43444=>"000001011",
  43445=>"001001001",
  43446=>"000011111",
  43447=>"010011111",
  43448=>"000000000",
  43449=>"000000111",
  43450=>"111111111",
  43451=>"011000000",
  43452=>"000000110",
  43453=>"000000000",
  43454=>"110101001",
  43455=>"111110111",
  43456=>"000000000",
  43457=>"111111100",
  43458=>"000010011",
  43459=>"111111111",
  43460=>"111100000",
  43461=>"010000001",
  43462=>"111000000",
  43463=>"001100101",
  43464=>"000000000",
  43465=>"000000110",
  43466=>"101000100",
  43467=>"000000000",
  43468=>"111111000",
  43469=>"100000000",
  43470=>"111111100",
  43471=>"000000111",
  43472=>"001001011",
  43473=>"000000000",
  43474=>"111111111",
  43475=>"111111110",
  43476=>"111111111",
  43477=>"111111111",
  43478=>"101101000",
  43479=>"100100110",
  43480=>"111001001",
  43481=>"101001000",
  43482=>"010000000",
  43483=>"111111000",
  43484=>"000000000",
  43485=>"110011000",
  43486=>"111111111",
  43487=>"001000000",
  43488=>"000000000",
  43489=>"111011000",
  43490=>"000000000",
  43491=>"111111111",
  43492=>"000001001",
  43493=>"000000000",
  43494=>"111111100",
  43495=>"110111111",
  43496=>"000000111",
  43497=>"111111111",
  43498=>"000011111",
  43499=>"111110100",
  43500=>"001001000",
  43501=>"100000000",
  43502=>"101111111",
  43503=>"111111110",
  43504=>"000001011",
  43505=>"001111111",
  43506=>"000000000",
  43507=>"000000000",
  43508=>"001001111",
  43509=>"111111011",
  43510=>"000000001",
  43511=>"000000000",
  43512=>"111111010",
  43513=>"100110111",
  43514=>"011011000",
  43515=>"111111010",
  43516=>"111111001",
  43517=>"111100111",
  43518=>"111111111",
  43519=>"000000000",
  43520=>"110111011",
  43521=>"110000000",
  43522=>"111111111",
  43523=>"001000100",
  43524=>"000000000",
  43525=>"111111011",
  43526=>"000100001",
  43527=>"000000111",
  43528=>"111001111",
  43529=>"000000000",
  43530=>"001000000",
  43531=>"111100100",
  43532=>"001111001",
  43533=>"111010011",
  43534=>"000110110",
  43535=>"000000111",
  43536=>"111110111",
  43537=>"000000000",
  43538=>"110111111",
  43539=>"111111111",
  43540=>"111111001",
  43541=>"111111111",
  43542=>"000111100",
  43543=>"111001001",
  43544=>"100100100",
  43545=>"001101111",
  43546=>"111111111",
  43547=>"111111000",
  43548=>"111111111",
  43549=>"110000000",
  43550=>"000111111",
  43551=>"111001000",
  43552=>"000000000",
  43553=>"111110000",
  43554=>"111011011",
  43555=>"000000000",
  43556=>"100100110",
  43557=>"111111111",
  43558=>"111110110",
  43559=>"111111111",
  43560=>"111011000",
  43561=>"111000001",
  43562=>"111000000",
  43563=>"111111111",
  43564=>"000111111",
  43565=>"000000100",
  43566=>"000100100",
  43567=>"101111101",
  43568=>"000000000",
  43569=>"100000000",
  43570=>"001001010",
  43571=>"111001000",
  43572=>"000000000",
  43573=>"000000001",
  43574=>"111101101",
  43575=>"111111111",
  43576=>"111111111",
  43577=>"000000001",
  43578=>"000000001",
  43579=>"111011011",
  43580=>"111111111",
  43581=>"100100000",
  43582=>"111111111",
  43583=>"111100000",
  43584=>"000100111",
  43585=>"100000110",
  43586=>"111111111",
  43587=>"111111111",
  43588=>"111111111",
  43589=>"000000001",
  43590=>"111111001",
  43591=>"111111111",
  43592=>"011011000",
  43593=>"000000110",
  43594=>"111000000",
  43595=>"000000110",
  43596=>"000101000",
  43597=>"010110000",
  43598=>"000010111",
  43599=>"111111111",
  43600=>"111111111",
  43601=>"000000111",
  43602=>"000000001",
  43603=>"000110000",
  43604=>"000100000",
  43605=>"111111000",
  43606=>"111000001",
  43607=>"010010110",
  43608=>"111111001",
  43609=>"000000000",
  43610=>"100100010",
  43611=>"110111111",
  43612=>"000001101",
  43613=>"011000000",
  43614=>"111001001",
  43615=>"000000000",
  43616=>"000000000",
  43617=>"000000011",
  43618=>"110111001",
  43619=>"111110000",
  43620=>"111111101",
  43621=>"000000000",
  43622=>"000010000",
  43623=>"000001111",
  43624=>"000000000",
  43625=>"000111111",
  43626=>"011000000",
  43627=>"010110000",
  43628=>"111000011",
  43629=>"111111000",
  43630=>"000111110",
  43631=>"000111010",
  43632=>"111111111",
  43633=>"110000101",
  43634=>"000000111",
  43635=>"000000000",
  43636=>"111111000",
  43637=>"000000000",
  43638=>"000000000",
  43639=>"111111001",
  43640=>"111010000",
  43641=>"000100001",
  43642=>"000100110",
  43643=>"011111011",
  43644=>"011111001",
  43645=>"000000000",
  43646=>"000000000",
  43647=>"000000000",
  43648=>"010111011",
  43649=>"000001111",
  43650=>"000000000",
  43651=>"111111111",
  43652=>"111111000",
  43653=>"111000000",
  43654=>"000000001",
  43655=>"111011000",
  43656=>"111111110",
  43657=>"000000011",
  43658=>"111111100",
  43659=>"000000111",
  43660=>"000000000",
  43661=>"010111000",
  43662=>"000110111",
  43663=>"111111111",
  43664=>"001111101",
  43665=>"110000000",
  43666=>"010111111",
  43667=>"111110111",
  43668=>"000000001",
  43669=>"000000000",
  43670=>"111111111",
  43671=>"001000000",
  43672=>"011111111",
  43673=>"101100110",
  43674=>"111111111",
  43675=>"010000001",
  43676=>"111100100",
  43677=>"110010001",
  43678=>"100100101",
  43679=>"111111111",
  43680=>"000001111",
  43681=>"110111111",
  43682=>"000000000",
  43683=>"000000000",
  43684=>"001111111",
  43685=>"001111101",
  43686=>"000111010",
  43687=>"000011011",
  43688=>"111000000",
  43689=>"100111111",
  43690=>"111111111",
  43691=>"110000001",
  43692=>"011111010",
  43693=>"111101011",
  43694=>"111111110",
  43695=>"000000111",
  43696=>"001111111",
  43697=>"100110110",
  43698=>"000000110",
  43699=>"000100000",
  43700=>"111110100",
  43701=>"111111111",
  43702=>"000110000",
  43703=>"110000011",
  43704=>"000000111",
  43705=>"111111000",
  43706=>"000000011",
  43707=>"000000001",
  43708=>"111111111",
  43709=>"000000000",
  43710=>"000000000",
  43711=>"111011011",
  43712=>"110111001",
  43713=>"111111111",
  43714=>"010000111",
  43715=>"001111111",
  43716=>"000110111",
  43717=>"011111111",
  43718=>"000000100",
  43719=>"011000000",
  43720=>"111111111",
  43721=>"111111111",
  43722=>"111111011",
  43723=>"010111111",
  43724=>"100100000",
  43725=>"111111111",
  43726=>"111001000",
  43727=>"111110000",
  43728=>"111110110",
  43729=>"010000000",
  43730=>"110000000",
  43731=>"000000001",
  43732=>"000100000",
  43733=>"001001111",
  43734=>"000011000",
  43735=>"001000000",
  43736=>"111110110",
  43737=>"111111111",
  43738=>"000000000",
  43739=>"100101111",
  43740=>"110111110",
  43741=>"000000111",
  43742=>"000000000",
  43743=>"111111111",
  43744=>"111000000",
  43745=>"111111111",
  43746=>"000000000",
  43747=>"101100000",
  43748=>"000000000",
  43749=>"000000100",
  43750=>"111100110",
  43751=>"111111000",
  43752=>"100111111",
  43753=>"111111110",
  43754=>"011000000",
  43755=>"000000000",
  43756=>"000000000",
  43757=>"111000000",
  43758=>"110110111",
  43759=>"111111111",
  43760=>"000000111",
  43761=>"000000110",
  43762=>"100110010",
  43763=>"001001111",
  43764=>"111111111",
  43765=>"110100001",
  43766=>"111111111",
  43767=>"000000110",
  43768=>"100001000",
  43769=>"010010111",
  43770=>"111111111",
  43771=>"111110110",
  43772=>"111111111",
  43773=>"100100000",
  43774=>"101101001",
  43775=>"000101111",
  43776=>"001000000",
  43777=>"110110010",
  43778=>"111010111",
  43779=>"111111111",
  43780=>"111000101",
  43781=>"100000000",
  43782=>"000110110",
  43783=>"111111101",
  43784=>"001111111",
  43785=>"000000000",
  43786=>"011100000",
  43787=>"110000000",
  43788=>"100010111",
  43789=>"000000000",
  43790=>"111111111",
  43791=>"000000111",
  43792=>"111111100",
  43793=>"100100101",
  43794=>"001001111",
  43795=>"100111110",
  43796=>"111111000",
  43797=>"000001001",
  43798=>"000000000",
  43799=>"001111111",
  43800=>"111111011",
  43801=>"100000000",
  43802=>"011111111",
  43803=>"000111111",
  43804=>"100110000",
  43805=>"110111111",
  43806=>"111111111",
  43807=>"000001111",
  43808=>"000000000",
  43809=>"000001101",
  43810=>"111100100",
  43811=>"000000111",
  43812=>"010000000",
  43813=>"011101101",
  43814=>"000000000",
  43815=>"111110100",
  43816=>"010111010",
  43817=>"101111111",
  43818=>"000000100",
  43819=>"000000000",
  43820=>"000000000",
  43821=>"000000111",
  43822=>"111111000",
  43823=>"111110010",
  43824=>"001000010",
  43825=>"000000000",
  43826=>"000000000",
  43827=>"000000001",
  43828=>"000000000",
  43829=>"111111111",
  43830=>"111000000",
  43831=>"000000000",
  43832=>"000000000",
  43833=>"111111111",
  43834=>"111111010",
  43835=>"111111000",
  43836=>"111111011",
  43837=>"001001011",
  43838=>"000000000",
  43839=>"000100000",
  43840=>"000000111",
  43841=>"101001100",
  43842=>"101100000",
  43843=>"000000000",
  43844=>"111100000",
  43845=>"100000110",
  43846=>"110111111",
  43847=>"000111111",
  43848=>"000000000",
  43849=>"000000000",
  43850=>"110111100",
  43851=>"111111110",
  43852=>"100000000",
  43853=>"100000000",
  43854=>"111111100",
  43855=>"001001000",
  43856=>"101100100",
  43857=>"111111100",
  43858=>"110010111",
  43859=>"111101111",
  43860=>"011001000",
  43861=>"111111111",
  43862=>"000000000",
  43863=>"100100100",
  43864=>"000111111",
  43865=>"001000000",
  43866=>"000000001",
  43867=>"000000100",
  43868=>"001001000",
  43869=>"110111111",
  43870=>"110100000",
  43871=>"000000000",
  43872=>"111100000",
  43873=>"110000000",
  43874=>"000001111",
  43875=>"111111110",
  43876=>"000000000",
  43877=>"111000000",
  43878=>"100000000",
  43879=>"011000000",
  43880=>"111111111",
  43881=>"000110111",
  43882=>"111000000",
  43883=>"111110000",
  43884=>"001011101",
  43885=>"000000000",
  43886=>"000000000",
  43887=>"000000000",
  43888=>"000000000",
  43889=>"001001000",
  43890=>"111111111",
  43891=>"100110110",
  43892=>"111111111",
  43893=>"000000010",
  43894=>"111111111",
  43895=>"100110111",
  43896=>"110111000",
  43897=>"111000000",
  43898=>"011000000",
  43899=>"110010111",
  43900=>"011111111",
  43901=>"111000000",
  43902=>"001000000",
  43903=>"000000111",
  43904=>"100110111",
  43905=>"011011111",
  43906=>"000000000",
  43907=>"111111111",
  43908=>"000000001",
  43909=>"000000000",
  43910=>"000000110",
  43911=>"000000000",
  43912=>"000000000",
  43913=>"111111011",
  43914=>"111111111",
  43915=>"111100100",
  43916=>"000000110",
  43917=>"011011011",
  43918=>"101100000",
  43919=>"111111111",
  43920=>"010000000",
  43921=>"111001101",
  43922=>"110110110",
  43923=>"111100000",
  43924=>"100101111",
  43925=>"111111111",
  43926=>"110111001",
  43927=>"000000001",
  43928=>"111111111",
  43929=>"010110111",
  43930=>"101101111",
  43931=>"111111111",
  43932=>"001111001",
  43933=>"101000000",
  43934=>"001000000",
  43935=>"000000000",
  43936=>"111111111",
  43937=>"110010000",
  43938=>"111000000",
  43939=>"000000000",
  43940=>"000100000",
  43941=>"110111000",
  43942=>"100110000",
  43943=>"011000000",
  43944=>"000000000",
  43945=>"111110110",
  43946=>"111000000",
  43947=>"000110000",
  43948=>"111000000",
  43949=>"111111111",
  43950=>"111111000",
  43951=>"111111000",
  43952=>"111111000",
  43953=>"110000110",
  43954=>"000000000",
  43955=>"000000000",
  43956=>"001111111",
  43957=>"000100111",
  43958=>"111100000",
  43959=>"111111001",
  43960=>"111111000",
  43961=>"000000111",
  43962=>"000001001",
  43963=>"100100110",
  43964=>"000000000",
  43965=>"101111111",
  43966=>"000000000",
  43967=>"011011011",
  43968=>"111111001",
  43969=>"111111111",
  43970=>"000010111",
  43971=>"111111011",
  43972=>"011000000",
  43973=>"001000000",
  43974=>"000000000",
  43975=>"100110110",
  43976=>"001111111",
  43977=>"000000000",
  43978=>"111111100",
  43979=>"111111000",
  43980=>"101111111",
  43981=>"111111110",
  43982=>"011000110",
  43983=>"000000111",
  43984=>"100000000",
  43985=>"000000110",
  43986=>"101000111",
  43987=>"111111111",
  43988=>"000100111",
  43989=>"000000000",
  43990=>"001011111",
  43991=>"111111110",
  43992=>"000100000",
  43993=>"111111000",
  43994=>"000011000",
  43995=>"000000000",
  43996=>"000000000",
  43997=>"000000000",
  43998=>"000000000",
  43999=>"000010000",
  44000=>"000000111",
  44001=>"000111111",
  44002=>"111111000",
  44003=>"000111111",
  44004=>"000010111",
  44005=>"101001011",
  44006=>"000000001",
  44007=>"000000000",
  44008=>"111111111",
  44009=>"111111111",
  44010=>"111111110",
  44011=>"000000000",
  44012=>"011000000",
  44013=>"111100100",
  44014=>"001111000",
  44015=>"111111100",
  44016=>"000010000",
  44017=>"000010111",
  44018=>"000001111",
  44019=>"111111100",
  44020=>"001100000",
  44021=>"111111000",
  44022=>"000000111",
  44023=>"000000011",
  44024=>"111010000",
  44025=>"100100110",
  44026=>"111111111",
  44027=>"110000000",
  44028=>"111111101",
  44029=>"000000000",
  44030=>"011000000",
  44031=>"111101000",
  44032=>"011100000",
  44033=>"000000111",
  44034=>"111111111",
  44035=>"111111011",
  44036=>"111111000",
  44037=>"001000010",
  44038=>"000000000",
  44039=>"110111111",
  44040=>"000000000",
  44041=>"110111111",
  44042=>"100000111",
  44043=>"000000000",
  44044=>"000000000",
  44045=>"011111111",
  44046=>"100000000",
  44047=>"000000111",
  44048=>"111111111",
  44049=>"000000001",
  44050=>"000000000",
  44051=>"000000010",
  44052=>"110000000",
  44053=>"000000111",
  44054=>"000001000",
  44055=>"001011011",
  44056=>"000000010",
  44057=>"111110100",
  44058=>"000000000",
  44059=>"111111011",
  44060=>"000000000",
  44061=>"000000000",
  44062=>"000000100",
  44063=>"001111000",
  44064=>"110010111",
  44065=>"110111011",
  44066=>"110111000",
  44067=>"111111011",
  44068=>"000111111",
  44069=>"100000001",
  44070=>"000001000",
  44071=>"111111111",
  44072=>"001111111",
  44073=>"000101111",
  44074=>"000000000",
  44075=>"100110111",
  44076=>"001111111",
  44077=>"000000000",
  44078=>"101100110",
  44079=>"000000000",
  44080=>"000000000",
  44081=>"000000000",
  44082=>"000011111",
  44083=>"111111111",
  44084=>"100111000",
  44085=>"010111111",
  44086=>"001000000",
  44087=>"110110111",
  44088=>"111111111",
  44089=>"000000000",
  44090=>"000001000",
  44091=>"000001000",
  44092=>"000100111",
  44093=>"111000010",
  44094=>"000000111",
  44095=>"000000000",
  44096=>"000000000",
  44097=>"100100111",
  44098=>"000000011",
  44099=>"000000111",
  44100=>"000000000",
  44101=>"000001111",
  44102=>"110101111",
  44103=>"111111110",
  44104=>"100100101",
  44105=>"000000001",
  44106=>"101000000",
  44107=>"001000110",
  44108=>"000000000",
  44109=>"000000000",
  44110=>"110110110",
  44111=>"000111111",
  44112=>"000000001",
  44113=>"000000001",
  44114=>"110010110",
  44115=>"011111100",
  44116=>"000000100",
  44117=>"111111110",
  44118=>"111000000",
  44119=>"000000011",
  44120=>"000000000",
  44121=>"111000111",
  44122=>"111011000",
  44123=>"001001001",
  44124=>"111111000",
  44125=>"000000000",
  44126=>"011000000",
  44127=>"111111011",
  44128=>"000001111",
  44129=>"011011010",
  44130=>"000000010",
  44131=>"111000100",
  44132=>"110111111",
  44133=>"111000000",
  44134=>"111000010",
  44135=>"000000001",
  44136=>"000000000",
  44137=>"111000000",
  44138=>"100100111",
  44139=>"000000000",
  44140=>"000000110",
  44141=>"010000011",
  44142=>"111111001",
  44143=>"110000000",
  44144=>"010111111",
  44145=>"000001000",
  44146=>"000000000",
  44147=>"000111111",
  44148=>"001011011",
  44149=>"000000000",
  44150=>"111111111",
  44151=>"000110000",
  44152=>"010000000",
  44153=>"000000101",
  44154=>"111001000",
  44155=>"000000000",
  44156=>"111001000",
  44157=>"010000001",
  44158=>"010010000",
  44159=>"001011111",
  44160=>"001111111",
  44161=>"000000000",
  44162=>"111101000",
  44163=>"000100000",
  44164=>"001111111",
  44165=>"001100111",
  44166=>"111110010",
  44167=>"000110110",
  44168=>"011111111",
  44169=>"111011111",
  44170=>"110000000",
  44171=>"000100111",
  44172=>"000000000",
  44173=>"111111111",
  44174=>"111111110",
  44175=>"011000000",
  44176=>"000001001",
  44177=>"100111110",
  44178=>"000111111",
  44179=>"000111110",
  44180=>"111111000",
  44181=>"000000001",
  44182=>"111100000",
  44183=>"111000000",
  44184=>"000000000",
  44185=>"000000111",
  44186=>"111111000",
  44187=>"000000000",
  44188=>"100000101",
  44189=>"111111000",
  44190=>"000000111",
  44191=>"000101101",
  44192=>"000000000",
  44193=>"110111111",
  44194=>"000111111",
  44195=>"000000000",
  44196=>"111001000",
  44197=>"111111011",
  44198=>"000101000",
  44199=>"000000000",
  44200=>"111000000",
  44201=>"010011100",
  44202=>"111111111",
  44203=>"000000000",
  44204=>"000111111",
  44205=>"110110100",
  44206=>"111110110",
  44207=>"111001111",
  44208=>"111111001",
  44209=>"111111111",
  44210=>"011111011",
  44211=>"111111000",
  44212=>"000001000",
  44213=>"010111011",
  44214=>"100111111",
  44215=>"000000110",
  44216=>"000000000",
  44217=>"110111111",
  44218=>"111111001",
  44219=>"000000000",
  44220=>"011000000",
  44221=>"000000111",
  44222=>"100100111",
  44223=>"111111111",
  44224=>"000000000",
  44225=>"000000111",
  44226=>"000010000",
  44227=>"000000000",
  44228=>"010111111",
  44229=>"111111111",
  44230=>"000000101",
  44231=>"000000100",
  44232=>"111111101",
  44233=>"011010110",
  44234=>"000000111",
  44235=>"111111001",
  44236=>"000111000",
  44237=>"110001001",
  44238=>"001011100",
  44239=>"111111111",
  44240=>"100101111",
  44241=>"000001001",
  44242=>"111001000",
  44243=>"000000000",
  44244=>"000000111",
  44245=>"110111000",
  44246=>"111011000",
  44247=>"111110111",
  44248=>"000010111",
  44249=>"110111101",
  44250=>"110010000",
  44251=>"000111111",
  44252=>"000001000",
  44253=>"000000111",
  44254=>"111111111",
  44255=>"111111110",
  44256=>"100000000",
  44257=>"110100000",
  44258=>"000100100",
  44259=>"001000000",
  44260=>"111111000",
  44261=>"100100000",
  44262=>"111011011",
  44263=>"111111111",
  44264=>"111111000",
  44265=>"001100110",
  44266=>"000111111",
  44267=>"111111100",
  44268=>"000111000",
  44269=>"110000000",
  44270=>"111111111",
  44271=>"000111111",
  44272=>"111110110",
  44273=>"000000000",
  44274=>"100111110",
  44275=>"011111001",
  44276=>"111111111",
  44277=>"011100000",
  44278=>"000000111",
  44279=>"001000001",
  44280=>"111011000",
  44281=>"000011111",
  44282=>"000000010",
  44283=>"000111111",
  44284=>"111111111",
  44285=>"000000000",
  44286=>"000010010",
  44287=>"011000000",
  44288=>"111111000",
  44289=>"001110000",
  44290=>"111111000",
  44291=>"000000000",
  44292=>"000000111",
  44293=>"000000000",
  44294=>"111111110",
  44295=>"111011000",
  44296=>"001111000",
  44297=>"111000000",
  44298=>"000001111",
  44299=>"000000000",
  44300=>"010111011",
  44301=>"100110111",
  44302=>"000000000",
  44303=>"001101111",
  44304=>"000110010",
  44305=>"111111111",
  44306=>"000000000",
  44307=>"000000100",
  44308=>"111111111",
  44309=>"000110111",
  44310=>"111111111",
  44311=>"111111111",
  44312=>"000000100",
  44313=>"111111000",
  44314=>"111111111",
  44315=>"111111111",
  44316=>"000111111",
  44317=>"111110000",
  44318=>"111111000",
  44319=>"000001000",
  44320=>"000110111",
  44321=>"111111000",
  44322=>"100000111",
  44323=>"000000100",
  44324=>"111111111",
  44325=>"111000001",
  44326=>"000111111",
  44327=>"110111111",
  44328=>"111111011",
  44329=>"110110111",
  44330=>"111111110",
  44331=>"000000000",
  44332=>"000000001",
  44333=>"000110110",
  44334=>"000000000",
  44335=>"000000110",
  44336=>"111111110",
  44337=>"000000000",
  44338=>"010111010",
  44339=>"000110111",
  44340=>"000000000",
  44341=>"100101111",
  44342=>"000000000",
  44343=>"110111111",
  44344=>"111101111",
  44345=>"000000111",
  44346=>"011000000",
  44347=>"101101101",
  44348=>"011001000",
  44349=>"000000000",
  44350=>"000111111",
  44351=>"010000111",
  44352=>"000000111",
  44353=>"110111000",
  44354=>"001001001",
  44355=>"111000010",
  44356=>"000001101",
  44357=>"000100101",
  44358=>"011011000",
  44359=>"111111000",
  44360=>"011011000",
  44361=>"000000011",
  44362=>"111111111",
  44363=>"110111111",
  44364=>"000000011",
  44365=>"000000100",
  44366=>"000111110",
  44367=>"011011001",
  44368=>"001011011",
  44369=>"111111000",
  44370=>"111111111",
  44371=>"001111111",
  44372=>"111111000",
  44373=>"001000000",
  44374=>"111111111",
  44375=>"100111001",
  44376=>"111111111",
  44377=>"001101001",
  44378=>"000011000",
  44379=>"111111111",
  44380=>"000000000",
  44381=>"000000000",
  44382=>"001001000",
  44383=>"000000000",
  44384=>"000000000",
  44385=>"000000000",
  44386=>"001011011",
  44387=>"111111111",
  44388=>"110000111",
  44389=>"111000000",
  44390=>"000000111",
  44391=>"000000000",
  44392=>"000001001",
  44393=>"111111001",
  44394=>"000110000",
  44395=>"000000001",
  44396=>"000000100",
  44397=>"111000001",
  44398=>"000000000",
  44399=>"100110110",
  44400=>"011000001",
  44401=>"001001000",
  44402=>"111111001",
  44403=>"100101111",
  44404=>"001111111",
  44405=>"010000000",
  44406=>"000000000",
  44407=>"110110000",
  44408=>"001000000",
  44409=>"000011111",
  44410=>"000000000",
  44411=>"000000000",
  44412=>"100111111",
  44413=>"111111110",
  44414=>"010011000",
  44415=>"111111111",
  44416=>"111111111",
  44417=>"111011000",
  44418=>"000011111",
  44419=>"000111000",
  44420=>"011111111",
  44421=>"111111111",
  44422=>"000100111",
  44423=>"001000000",
  44424=>"111111000",
  44425=>"011111101",
  44426=>"000000000",
  44427=>"111100111",
  44428=>"111111111",
  44429=>"000000000",
  44430=>"111111111",
  44431=>"001001001",
  44432=>"000111111",
  44433=>"000000100",
  44434=>"111110111",
  44435=>"000000000",
  44436=>"111111011",
  44437=>"111111111",
  44438=>"111001101",
  44439=>"110110100",
  44440=>"111111110",
  44441=>"111111000",
  44442=>"111111111",
  44443=>"000011111",
  44444=>"000000011",
  44445=>"000000111",
  44446=>"110111111",
  44447=>"000010000",
  44448=>"001111111",
  44449=>"111110110",
  44450=>"011001111",
  44451=>"111011000",
  44452=>"011000101",
  44453=>"000100000",
  44454=>"111001000",
  44455=>"000000000",
  44456=>"000000101",
  44457=>"111001010",
  44458=>"000000000",
  44459=>"100111111",
  44460=>"000000001",
  44461=>"011011000",
  44462=>"111111111",
  44463=>"000000000",
  44464=>"111111000",
  44465=>"111110100",
  44466=>"000100101",
  44467=>"000011111",
  44468=>"111111000",
  44469=>"111010000",
  44470=>"010000100",
  44471=>"000000110",
  44472=>"110111110",
  44473=>"111111110",
  44474=>"111111111",
  44475=>"000000001",
  44476=>"111111111",
  44477=>"111111111",
  44478=>"000100111",
  44479=>"110111110",
  44480=>"111111000",
  44481=>"000000111",
  44482=>"001001010",
  44483=>"111000101",
  44484=>"000000111",
  44485=>"011011000",
  44486=>"000000100",
  44487=>"111101111",
  44488=>"111011000",
  44489=>"111010000",
  44490=>"000000100",
  44491=>"011001000",
  44492=>"000000100",
  44493=>"000000111",
  44494=>"001100111",
  44495=>"111111111",
  44496=>"111110000",
  44497=>"000000011",
  44498=>"111110111",
  44499=>"011111111",
  44500=>"101000000",
  44501=>"000000000",
  44502=>"000000000",
  44503=>"011111101",
  44504=>"111111111",
  44505=>"111111111",
  44506=>"000000000",
  44507=>"011101001",
  44508=>"110000000",
  44509=>"111111000",
  44510=>"111111111",
  44511=>"000110111",
  44512=>"000100111",
  44513=>"100111111",
  44514=>"000000000",
  44515=>"111100000",
  44516=>"111111010",
  44517=>"100101000",
  44518=>"000000111",
  44519=>"111111000",
  44520=>"000010110",
  44521=>"001011001",
  44522=>"111111111",
  44523=>"111111010",
  44524=>"000000000",
  44525=>"101111111",
  44526=>"111111111",
  44527=>"111111000",
  44528=>"000001001",
  44529=>"000000100",
  44530=>"111111000",
  44531=>"111111000",
  44532=>"000000000",
  44533=>"000001111",
  44534=>"110110111",
  44535=>"110110111",
  44536=>"110111101",
  44537=>"000011000",
  44538=>"111111111",
  44539=>"110110111",
  44540=>"000010110",
  44541=>"000000000",
  44542=>"001111100",
  44543=>"001111111",
  44544=>"000000010",
  44545=>"100100001",
  44546=>"000000000",
  44547=>"000000000",
  44548=>"011011111",
  44549=>"001000011",
  44550=>"001000100",
  44551=>"111111111",
  44552=>"000000011",
  44553=>"000111110",
  44554=>"000000000",
  44555=>"000001111",
  44556=>"011011001",
  44557=>"000000001",
  44558=>"000000000",
  44559=>"000000000",
  44560=>"110111111",
  44561=>"000111111",
  44562=>"000000111",
  44563=>"000000000",
  44564=>"111111000",
  44565=>"001011001",
  44566=>"000000100",
  44567=>"100110000",
  44568=>"111111001",
  44569=>"111111111",
  44570=>"001000000",
  44571=>"000000000",
  44572=>"111111000",
  44573=>"110110111",
  44574=>"000000000",
  44575=>"000000001",
  44576=>"111111111",
  44577=>"000000111",
  44578=>"011111110",
  44579=>"111000000",
  44580=>"000000100",
  44581=>"111111111",
  44582=>"111111111",
  44583=>"111011011",
  44584=>"000000101",
  44585=>"100100000",
  44586=>"110110100",
  44587=>"000000011",
  44588=>"000001111",
  44589=>"100111101",
  44590=>"111111111",
  44591=>"000000000",
  44592=>"000001001",
  44593=>"111111110",
  44594=>"100110111",
  44595=>"111111111",
  44596=>"100110000",
  44597=>"000001001",
  44598=>"110110000",
  44599=>"010110010",
  44600=>"000000111",
  44601=>"000000001",
  44602=>"111111110",
  44603=>"111111111",
  44604=>"111111111",
  44605=>"111111111",
  44606=>"000110000",
  44607=>"000000111",
  44608=>"111000100",
  44609=>"101111101",
  44610=>"111000000",
  44611=>"111011000",
  44612=>"000111111",
  44613=>"000000000",
  44614=>"110110111",
  44615=>"000000111",
  44616=>"011011111",
  44617=>"011001001",
  44618=>"000000000",
  44619=>"001000110",
  44620=>"000110111",
  44621=>"111111000",
  44622=>"011000000",
  44623=>"110010000",
  44624=>"111001001",
  44625=>"011111111",
  44626=>"110110110",
  44627=>"011011111",
  44628=>"010000000",
  44629=>"000000000",
  44630=>"110000101",
  44631=>"000000011",
  44632=>"000001111",
  44633=>"111000000",
  44634=>"111111000",
  44635=>"111010010",
  44636=>"000000001",
  44637=>"101111101",
  44638=>"111111111",
  44639=>"111111110",
  44640=>"000001111",
  44641=>"011011000",
  44642=>"111111111",
  44643=>"011011111",
  44644=>"000001011",
  44645=>"000101111",
  44646=>"111111110",
  44647=>"111000000",
  44648=>"100111001",
  44649=>"001101111",
  44650=>"001011111",
  44651=>"000000100",
  44652=>"011011111",
  44653=>"111111100",
  44654=>"111001000",
  44655=>"111111110",
  44656=>"111111111",
  44657=>"000000101",
  44658=>"110111011",
  44659=>"000000111",
  44660=>"000000000",
  44661=>"000000000",
  44662=>"000000000",
  44663=>"101101111",
  44664=>"101011011",
  44665=>"000000000",
  44666=>"000001001",
  44667=>"000000000",
  44668=>"110111111",
  44669=>"111111000",
  44670=>"000000000",
  44671=>"000110001",
  44672=>"110111111",
  44673=>"010101000",
  44674=>"011111110",
  44675=>"001110110",
  44676=>"111110100",
  44677=>"000000000",
  44678=>"111110100",
  44679=>"011011011",
  44680=>"100111111",
  44681=>"000000000",
  44682=>"000000111",
  44683=>"100101111",
  44684=>"111111011",
  44685=>"111111000",
  44686=>"011001111",
  44687=>"111111000",
  44688=>"000000000",
  44689=>"001001001",
  44690=>"111100101",
  44691=>"111111111",
  44692=>"111000000",
  44693=>"111111011",
  44694=>"100111111",
  44695=>"000000100",
  44696=>"001000001",
  44697=>"000000001",
  44698=>"000000001",
  44699=>"010000110",
  44700=>"000000000",
  44701=>"100111111",
  44702=>"111111000",
  44703=>"000000110",
  44704=>"001001001",
  44705=>"100001000",
  44706=>"000000000",
  44707=>"010000100",
  44708=>"100001011",
  44709=>"001011111",
  44710=>"101111111",
  44711=>"000011011",
  44712=>"111111111",
  44713=>"000001111",
  44714=>"111111111",
  44715=>"000011011",
  44716=>"111111111",
  44717=>"001111111",
  44718=>"111001111",
  44719=>"110111111",
  44720=>"000001000",
  44721=>"110110111",
  44722=>"110111111",
  44723=>"000001111",
  44724=>"101010000",
  44725=>"011001001",
  44726=>"011000111",
  44727=>"000000100",
  44728=>"111111111",
  44729=>"000100101",
  44730=>"000000101",
  44731=>"001000000",
  44732=>"111111111",
  44733=>"001000000",
  44734=>"111011001",
  44735=>"000000111",
  44736=>"111111111",
  44737=>"011001011",
  44738=>"100101101",
  44739=>"100111111",
  44740=>"000000011",
  44741=>"000000000",
  44742=>"000111001",
  44743=>"000100111",
  44744=>"000000000",
  44745=>"111111111",
  44746=>"010110000",
  44747=>"000111111",
  44748=>"011111111",
  44749=>"010111111",
  44750=>"110110111",
  44751=>"111111000",
  44752=>"111111011",
  44753=>"010110100",
  44754=>"000111011",
  44755=>"111111111",
  44756=>"000001011",
  44757=>"001011111",
  44758=>"111100000",
  44759=>"000000000",
  44760=>"000100111",
  44761=>"011001000",
  44762=>"000000000",
  44763=>"111111100",
  44764=>"111011111",
  44765=>"000111001",
  44766=>"110111111",
  44767=>"001001001",
  44768=>"100100000",
  44769=>"100111110",
  44770=>"111111000",
  44771=>"110000000",
  44772=>"100111000",
  44773=>"111101111",
  44774=>"111111000",
  44775=>"111111111",
  44776=>"100110100",
  44777=>"000001011",
  44778=>"111011000",
  44779=>"000001001",
  44780=>"000011000",
  44781=>"000000001",
  44782=>"110000000",
  44783=>"000001111",
  44784=>"111111000",
  44785=>"000110110",
  44786=>"111111101",
  44787=>"000001111",
  44788=>"000000010",
  44789=>"110111000",
  44790=>"000000110",
  44791=>"010000000",
  44792=>"000110110",
  44793=>"000000000",
  44794=>"000001011",
  44795=>"000000000",
  44796=>"000000000",
  44797=>"000000001",
  44798=>"010111111",
  44799=>"111111100",
  44800=>"000000001",
  44801=>"001001001",
  44802=>"111111000",
  44803=>"000010000",
  44804=>"001100111",
  44805=>"000010110",
  44806=>"111111000",
  44807=>"100000000",
  44808=>"011000000",
  44809=>"000000000",
  44810=>"000000101",
  44811=>"011100101",
  44812=>"001001001",
  44813=>"001011111",
  44814=>"000010110",
  44815=>"111110000",
  44816=>"111001000",
  44817=>"000000000",
  44818=>"100100001",
  44819=>"001000100",
  44820=>"111100110",
  44821=>"011111010",
  44822=>"111111111",
  44823=>"111111111",
  44824=>"110111111",
  44825=>"000000010",
  44826=>"100000000",
  44827=>"011000001",
  44828=>"111111111",
  44829=>"011011011",
  44830=>"111110000",
  44831=>"000000001",
  44832=>"000111111",
  44833=>"000000011",
  44834=>"100100111",
  44835=>"111111111",
  44836=>"110110110",
  44837=>"111111111",
  44838=>"100111110",
  44839=>"001001000",
  44840=>"111111111",
  44841=>"000000000",
  44842=>"110111011",
  44843=>"000000000",
  44844=>"000000100",
  44845=>"000001111",
  44846=>"001000111",
  44847=>"111000111",
  44848=>"000000100",
  44849=>"111111111",
  44850=>"111111111",
  44851=>"100110010",
  44852=>"010000000",
  44853=>"010110111",
  44854=>"001001111",
  44855=>"001000000",
  44856=>"000000111",
  44857=>"000000111",
  44858=>"011000000",
  44859=>"111010010",
  44860=>"000000100",
  44861=>"111111110",
  44862=>"010000000",
  44863=>"001001111",
  44864=>"000000111",
  44865=>"111011001",
  44866=>"110100111",
  44867=>"111111111",
  44868=>"110111111",
  44869=>"000000000",
  44870=>"010011000",
  44871=>"001000111",
  44872=>"000000000",
  44873=>"000000111",
  44874=>"000000000",
  44875=>"100100101",
  44876=>"000000010",
  44877=>"000000001",
  44878=>"111111001",
  44879=>"111111111",
  44880=>"111111111",
  44881=>"011011000",
  44882=>"110010111",
  44883=>"000000000",
  44884=>"111101001",
  44885=>"000010010",
  44886=>"110111101",
  44887=>"000101001",
  44888=>"111111000",
  44889=>"111111111",
  44890=>"110000011",
  44891=>"011000000",
  44892=>"000000111",
  44893=>"000000000",
  44894=>"001001011",
  44895=>"000000000",
  44896=>"101111100",
  44897=>"000111011",
  44898=>"100100110",
  44899=>"110000000",
  44900=>"110110111",
  44901=>"000000110",
  44902=>"000000000",
  44903=>"011111111",
  44904=>"110010000",
  44905=>"111111000",
  44906=>"111111001",
  44907=>"000001111",
  44908=>"111011001",
  44909=>"000011111",
  44910=>"000000000",
  44911=>"000001100",
  44912=>"000001111",
  44913=>"111111100",
  44914=>"110110110",
  44915=>"000000110",
  44916=>"111111100",
  44917=>"111111111",
  44918=>"111000011",
  44919=>"011001111",
  44920=>"111001000",
  44921=>"111111111",
  44922=>"000001001",
  44923=>"011010111",
  44924=>"000010000",
  44925=>"000011111",
  44926=>"111101000",
  44927=>"000110111",
  44928=>"000000000",
  44929=>"011011000",
  44930=>"100000000",
  44931=>"111111000",
  44932=>"000001001",
  44933=>"000000000",
  44934=>"000001001",
  44935=>"011000000",
  44936=>"000100111",
  44937=>"000000000",
  44938=>"100000000",
  44939=>"000100110",
  44940=>"111111111",
  44941=>"011001000",
  44942=>"001111111",
  44943=>"111111001",
  44944=>"011001000",
  44945=>"000000000",
  44946=>"111110110",
  44947=>"001000000",
  44948=>"000111000",
  44949=>"000000000",
  44950=>"011111111",
  44951=>"001001011",
  44952=>"000000100",
  44953=>"000000000",
  44954=>"111000000",
  44955=>"000000000",
  44956=>"000000000",
  44957=>"000000000",
  44958=>"001000100",
  44959=>"000000000",
  44960=>"000111111",
  44961=>"010110111",
  44962=>"001000000",
  44963=>"111111111",
  44964=>"001000000",
  44965=>"000010011",
  44966=>"000000111",
  44967=>"111111111",
  44968=>"011000000",
  44969=>"111101100",
  44970=>"000000111",
  44971=>"011011000",
  44972=>"000000000",
  44973=>"001110000",
  44974=>"110111111",
  44975=>"001111111",
  44976=>"000111111",
  44977=>"000010000",
  44978=>"000011011",
  44979=>"010110110",
  44980=>"000100000",
  44981=>"111101000",
  44982=>"111101111",
  44983=>"111111111",
  44984=>"011011000",
  44985=>"111110000",
  44986=>"110010010",
  44987=>"111100100",
  44988=>"111110110",
  44989=>"110110111",
  44990=>"000001011",
  44991=>"011010010",
  44992=>"110111001",
  44993=>"111111111",
  44994=>"100101101",
  44995=>"000000001",
  44996=>"001001111",
  44997=>"000111111",
  44998=>"001001000",
  44999=>"001111111",
  45000=>"101001101",
  45001=>"011011001",
  45002=>"111111101",
  45003=>"000000000",
  45004=>"001000000",
  45005=>"111111111",
  45006=>"001000101",
  45007=>"000000000",
  45008=>"111110010",
  45009=>"011111111",
  45010=>"000000001",
  45011=>"111111100",
  45012=>"111110000",
  45013=>"000000000",
  45014=>"000001000",
  45015=>"100110100",
  45016=>"000000000",
  45017=>"111111111",
  45018=>"111111111",
  45019=>"000000101",
  45020=>"110111111",
  45021=>"000000000",
  45022=>"000000111",
  45023=>"111001001",
  45024=>"101111111",
  45025=>"000000000",
  45026=>"000111110",
  45027=>"000000001",
  45028=>"010010111",
  45029=>"100100000",
  45030=>"000110110",
  45031=>"000000000",
  45032=>"001000110",
  45033=>"000001011",
  45034=>"110010000",
  45035=>"111111111",
  45036=>"111111111",
  45037=>"000000111",
  45038=>"000000111",
  45039=>"011001111",
  45040=>"111111111",
  45041=>"010111111",
  45042=>"111111111",
  45043=>"000000000",
  45044=>"000000111",
  45045=>"001000000",
  45046=>"001111001",
  45047=>"011000000",
  45048=>"010111111",
  45049=>"001111001",
  45050=>"011011011",
  45051=>"111111000",
  45052=>"000001000",
  45053=>"000011111",
  45054=>"011100111",
  45055=>"111100111",
  45056=>"100100011",
  45057=>"100101000",
  45058=>"111111111",
  45059=>"000110111",
  45060=>"110110111",
  45061=>"101101101",
  45062=>"000000000",
  45063=>"111111111",
  45064=>"001111001",
  45065=>"111111101",
  45066=>"110010000",
  45067=>"000110110",
  45068=>"111111100",
  45069=>"110000000",
  45070=>"011011111",
  45071=>"000000000",
  45072=>"001100100",
  45073=>"110100011",
  45074=>"000101101",
  45075=>"111111111",
  45076=>"111111111",
  45077=>"010000000",
  45078=>"101001111",
  45079=>"100000000",
  45080=>"001001000",
  45081=>"011111101",
  45082=>"111101000",
  45083=>"111010111",
  45084=>"111111111",
  45085=>"000000111",
  45086=>"110000100",
  45087=>"000100000",
  45088=>"101101101",
  45089=>"100000000",
  45090=>"111001001",
  45091=>"111011011",
  45092=>"101101111",
  45093=>"111111111",
  45094=>"001111111",
  45095=>"000000001",
  45096=>"110000000",
  45097=>"100000111",
  45098=>"111111111",
  45099=>"000010100",
  45100=>"101101101",
  45101=>"000000000",
  45102=>"111100000",
  45103=>"111111111",
  45104=>"111110111",
  45105=>"000000111",
  45106=>"110111111",
  45107=>"111011111",
  45108=>"100110010",
  45109=>"101011111",
  45110=>"101001011",
  45111=>"001000100",
  45112=>"101111111",
  45113=>"010110111",
  45114=>"111111111",
  45115=>"000000000",
  45116=>"000000000",
  45117=>"111000100",
  45118=>"100000000",
  45119=>"111110110",
  45120=>"111111111",
  45121=>"001011011",
  45122=>"000100111",
  45123=>"011001000",
  45124=>"111001110",
  45125=>"000000000",
  45126=>"110110000",
  45127=>"000000000",
  45128=>"000000010",
  45129=>"000100100",
  45130=>"111111111",
  45131=>"101001000",
  45132=>"111111101",
  45133=>"100110111",
  45134=>"111110111",
  45135=>"100000110",
  45136=>"110111111",
  45137=>"000011111",
  45138=>"000000000",
  45139=>"101111011",
  45140=>"111111001",
  45141=>"000100110",
  45142=>"111111011",
  45143=>"111101111",
  45144=>"010000000",
  45145=>"111100100",
  45146=>"000000111",
  45147=>"110001001",
  45148=>"100100100",
  45149=>"000011111",
  45150=>"110110111",
  45151=>"000000000",
  45152=>"111111111",
  45153=>"101101111",
  45154=>"000000111",
  45155=>"111001000",
  45156=>"010000000",
  45157=>"100111000",
  45158=>"100000000",
  45159=>"111101101",
  45160=>"000000000",
  45161=>"000110010",
  45162=>"001111110",
  45163=>"111111111",
  45164=>"001000000",
  45165=>"001011111",
  45166=>"000000000",
  45167=>"000000000",
  45168=>"100100100",
  45169=>"001111111",
  45170=>"100100100",
  45171=>"101001001",
  45172=>"111111011",
  45173=>"100100000",
  45174=>"111111111",
  45175=>"110111111",
  45176=>"101111111",
  45177=>"101001011",
  45178=>"000111000",
  45179=>"110000000",
  45180=>"000000000",
  45181=>"000011000",
  45182=>"011111111",
  45183=>"000101101",
  45184=>"111111000",
  45185=>"001001000",
  45186=>"101000000",
  45187=>"111111111",
  45188=>"001001111",
  45189=>"101111111",
  45190=>"000110000",
  45191=>"001011000",
  45192=>"000000000",
  45193=>"000101101",
  45194=>"010000001",
  45195=>"110110111",
  45196=>"000000000",
  45197=>"001111111",
  45198=>"001000000",
  45199=>"111111111",
  45200=>"100001111",
  45201=>"111011011",
  45202=>"111111111",
  45203=>"111000000",
  45204=>"110001001",
  45205=>"000110111",
  45206=>"000000000",
  45207=>"111111000",
  45208=>"000001000",
  45209=>"111111100",
  45210=>"111111111",
  45211=>"111110111",
  45212=>"011000000",
  45213=>"101100111",
  45214=>"000000000",
  45215=>"111111111",
  45216=>"111111000",
  45217=>"000000000",
  45218=>"111110100",
  45219=>"111100111",
  45220=>"100001111",
  45221=>"000000000",
  45222=>"000000000",
  45223=>"000011111",
  45224=>"000000000",
  45225=>"111000000",
  45226=>"000000000",
  45227=>"111000101",
  45228=>"111111111",
  45229=>"000000010",
  45230=>"111111001",
  45231=>"001000000",
  45232=>"000001000",
  45233=>"001011010",
  45234=>"000000010",
  45235=>"111111111",
  45236=>"100100101",
  45237=>"001101000",
  45238=>"000111111",
  45239=>"010010110",
  45240=>"100000010",
  45241=>"111111111",
  45242=>"100000111",
  45243=>"100000111",
  45244=>"111111100",
  45245=>"000001111",
  45246=>"000110110",
  45247=>"000010111",
  45248=>"010011111",
  45249=>"110000000",
  45250=>"111001111",
  45251=>"000000000",
  45252=>"000000001",
  45253=>"000000000",
  45254=>"111001111",
  45255=>"110110110",
  45256=>"101101111",
  45257=>"100100111",
  45258=>"110110110",
  45259=>"001000000",
  45260=>"001011111",
  45261=>"110011000",
  45262=>"000000000",
  45263=>"101000111",
  45264=>"111100111",
  45265=>"111111111",
  45266=>"000000000",
  45267=>"110110111",
  45268=>"111110100",
  45269=>"000111110",
  45270=>"101101000",
  45271=>"111000000",
  45272=>"111111101",
  45273=>"111001101",
  45274=>"000000000",
  45275=>"110111000",
  45276=>"000000000",
  45277=>"000000000",
  45278=>"010000000",
  45279=>"000100111",
  45280=>"010000000",
  45281=>"001111011",
  45282=>"000111011",
  45283=>"101000000",
  45284=>"100100001",
  45285=>"001000000",
  45286=>"101111111",
  45287=>"110110000",
  45288=>"010000111",
  45289=>"000000011",
  45290=>"111111111",
  45291=>"100000000",
  45292=>"111111010",
  45293=>"000111001",
  45294=>"000001101",
  45295=>"100111111",
  45296=>"001110110",
  45297=>"001001011",
  45298=>"010000000",
  45299=>"110101111",
  45300=>"111111111",
  45301=>"000000000",
  45302=>"010000000",
  45303=>"111111001",
  45304=>"000001000",
  45305=>"001101101",
  45306=>"001000110",
  45307=>"101001101",
  45308=>"001111001",
  45309=>"100100100",
  45310=>"000000100",
  45311=>"000010000",
  45312=>"100000000",
  45313=>"100100100",
  45314=>"000000000",
  45315=>"110110000",
  45316=>"100100110",
  45317=>"111010111",
  45318=>"000010000",
  45319=>"011000100",
  45320=>"110100111",
  45321=>"000111111",
  45322=>"100100100",
  45323=>"111111000",
  45324=>"111100111",
  45325=>"101111111",
  45326=>"100101111",
  45327=>"000001110",
  45328=>"001111111",
  45329=>"001000001",
  45330=>"100000000",
  45331=>"100111011",
  45332=>"011001000",
  45333=>"000000111",
  45334=>"000110111",
  45335=>"111000001",
  45336=>"011011111",
  45337=>"111101000",
  45338=>"111001001",
  45339=>"000000000",
  45340=>"000000000",
  45341=>"000110111",
  45342=>"111000000",
  45343=>"111111111",
  45344=>"000011011",
  45345=>"101100000",
  45346=>"000000100",
  45347=>"000000000",
  45348=>"011001111",
  45349=>"111111111",
  45350=>"110111000",
  45351=>"100111110",
  45352=>"111110110",
  45353=>"001000101",
  45354=>"111001000",
  45355=>"001000101",
  45356=>"000000000",
  45357=>"111011001",
  45358=>"100111111",
  45359=>"111111111",
  45360=>"100100101",
  45361=>"111110011",
  45362=>"111111111",
  45363=>"110110111",
  45364=>"100000100",
  45365=>"000100111",
  45366=>"000111111",
  45367=>"111110010",
  45368=>"001001111",
  45369=>"111010111",
  45370=>"111010000",
  45371=>"110100000",
  45372=>"110011011",
  45373=>"110000000",
  45374=>"111111111",
  45375=>"111111001",
  45376=>"101111001",
  45377=>"111111111",
  45378=>"111110001",
  45379=>"111000000",
  45380=>"011011011",
  45381=>"011011100",
  45382=>"000111101",
  45383=>"000000001",
  45384=>"011000000",
  45385=>"111111100",
  45386=>"111011111",
  45387=>"001001001",
  45388=>"011000000",
  45389=>"000000110",
  45390=>"111111111",
  45391=>"011111011",
  45392=>"001111011",
  45393=>"000111001",
  45394=>"100000100",
  45395=>"000010111",
  45396=>"000001011",
  45397=>"011010000",
  45398=>"010111111",
  45399=>"000000100",
  45400=>"010000110",
  45401=>"011001000",
  45402=>"011000000",
  45403=>"111001001",
  45404=>"111101101",
  45405=>"000000001",
  45406=>"111100000",
  45407=>"001101001",
  45408=>"000000000",
  45409=>"000000000",
  45410=>"001111011",
  45411=>"111001111",
  45412=>"111011111",
  45413=>"110100111",
  45414=>"000111000",
  45415=>"011111001",
  45416=>"100000100",
  45417=>"111111111",
  45418=>"111011111",
  45419=>"110100100",
  45420=>"111111111",
  45421=>"110100001",
  45422=>"000010110",
  45423=>"111111111",
  45424=>"111101111",
  45425=>"111111111",
  45426=>"100101111",
  45427=>"000000101",
  45428=>"000000000",
  45429=>"000000000",
  45430=>"110100101",
  45431=>"111111000",
  45432=>"111111000",
  45433=>"110111111",
  45434=>"111111111",
  45435=>"111111111",
  45436=>"011110111",
  45437=>"111110111",
  45438=>"101111111",
  45439=>"111111111",
  45440=>"111000000",
  45441=>"110110111",
  45442=>"110000000",
  45443=>"111100111",
  45444=>"000000000",
  45445=>"000010010",
  45446=>"001000100",
  45447=>"110100111",
  45448=>"100100001",
  45449=>"111011010",
  45450=>"101101000",
  45451=>"111111110",
  45452=>"000000111",
  45453=>"011010000",
  45454=>"111111111",
  45455=>"000010000",
  45456=>"111111111",
  45457=>"001000111",
  45458=>"001011011",
  45459=>"111110100",
  45460=>"000000000",
  45461=>"010111111",
  45462=>"110100000",
  45463=>"110011011",
  45464=>"001001001",
  45465=>"111101100",
  45466=>"111111001",
  45467=>"000100011",
  45468=>"111000000",
  45469=>"101111010",
  45470=>"101111111",
  45471=>"111111011",
  45472=>"111110110",
  45473=>"100100000",
  45474=>"111101101",
  45475=>"000000001",
  45476=>"110010000",
  45477=>"000100101",
  45478=>"000000000",
  45479=>"111111001",
  45480=>"001001001",
  45481=>"100000001",
  45482=>"111110000",
  45483=>"100100111",
  45484=>"111111000",
  45485=>"000000000",
  45486=>"000010110",
  45487=>"111011111",
  45488=>"111100100",
  45489=>"000000001",
  45490=>"111111011",
  45491=>"000001111",
  45492=>"110101110",
  45493=>"111111111",
  45494=>"111111111",
  45495=>"111111111",
  45496=>"000111111",
  45497=>"111000100",
  45498=>"100111110",
  45499=>"011111010",
  45500=>"011111111",
  45501=>"000010110",
  45502=>"111001011",
  45503=>"100101100",
  45504=>"001000000",
  45505=>"000000000",
  45506=>"000000000",
  45507=>"111111111",
  45508=>"000000100",
  45509=>"011000000",
  45510=>"101000000",
  45511=>"111001001",
  45512=>"110001011",
  45513=>"100100111",
  45514=>"111110000",
  45515=>"111111111",
  45516=>"001000000",
  45517=>"111111111",
  45518=>"100000001",
  45519=>"001011100",
  45520=>"001000011",
  45521=>"011011011",
  45522=>"000000111",
  45523=>"001010000",
  45524=>"110110011",
  45525=>"000000001",
  45526=>"100110110",
  45527=>"111000000",
  45528=>"111000000",
  45529=>"111101111",
  45530=>"111111110",
  45531=>"010011111",
  45532=>"111111111",
  45533=>"110100100",
  45534=>"000101111",
  45535=>"100100100",
  45536=>"111110110",
  45537=>"000000000",
  45538=>"111111111",
  45539=>"001000010",
  45540=>"111111111",
  45541=>"001000000",
  45542=>"011001001",
  45543=>"000000111",
  45544=>"000000010",
  45545=>"001101111",
  45546=>"111100111",
  45547=>"110110110",
  45548=>"111001010",
  45549=>"001011110",
  45550=>"101001111",
  45551=>"000000000",
  45552=>"111111111",
  45553=>"011111111",
  45554=>"110000111",
  45555=>"111101111",
  45556=>"100100000",
  45557=>"000000010",
  45558=>"000000000",
  45559=>"000001000",
  45560=>"111101000",
  45561=>"111111001",
  45562=>"111001000",
  45563=>"001000000",
  45564=>"110111000",
  45565=>"111111110",
  45566=>"111111111",
  45567=>"111111000",
  45568=>"011000001",
  45569=>"101111111",
  45570=>"111101101",
  45571=>"100100000",
  45572=>"111111000",
  45573=>"111111000",
  45574=>"111111110",
  45575=>"111111111",
  45576=>"010000000",
  45577=>"000000101",
  45578=>"111111111",
  45579=>"101100101",
  45580=>"001011001",
  45581=>"000001001",
  45582=>"000000001",
  45583=>"010111000",
  45584=>"111111111",
  45585=>"000000111",
  45586=>"100001000",
  45587=>"111111111",
  45588=>"111000001",
  45589=>"001001111",
  45590=>"111011000",
  45591=>"100100110",
  45592=>"011111111",
  45593=>"110000011",
  45594=>"111111111",
  45595=>"111011011",
  45596=>"111100000",
  45597=>"000000000",
  45598=>"100000100",
  45599=>"000000000",
  45600=>"000000000",
  45601=>"000000000",
  45602=>"000000000",
  45603=>"111111111",
  45604=>"111111111",
  45605=>"111111111",
  45606=>"000000000",
  45607=>"110110111",
  45608=>"000000000",
  45609=>"000000000",
  45610=>"111111111",
  45611=>"000000000",
  45612=>"000000000",
  45613=>"000000000",
  45614=>"111111111",
  45615=>"111000100",
  45616=>"011011110",
  45617=>"000000000",
  45618=>"111111111",
  45619=>"000000000",
  45620=>"101100000",
  45621=>"110111111",
  45622=>"111100000",
  45623=>"100111001",
  45624=>"111111011",
  45625=>"000000001",
  45626=>"001111111",
  45627=>"011111111",
  45628=>"000000000",
  45629=>"001001000",
  45630=>"111111111",
  45631=>"000000111",
  45632=>"111111110",
  45633=>"111111111",
  45634=>"111111111",
  45635=>"000000000",
  45636=>"001001000",
  45637=>"111111111",
  45638=>"001111111",
  45639=>"111111111",
  45640=>"111111111",
  45641=>"111111111",
  45642=>"000000000",
  45643=>"111111111",
  45644=>"111111111",
  45645=>"000000000",
  45646=>"000000000",
  45647=>"100110111",
  45648=>"111111001",
  45649=>"110110111",
  45650=>"000000000",
  45651=>"100100000",
  45652=>"000000000",
  45653=>"111111011",
  45654=>"111001000",
  45655=>"111001000",
  45656=>"010000000",
  45657=>"000000000",
  45658=>"111111111",
  45659=>"001000000",
  45660=>"111111000",
  45661=>"000001111",
  45662=>"000000110",
  45663=>"000000000",
  45664=>"000000000",
  45665=>"110000000",
  45666=>"111100111",
  45667=>"000000000",
  45668=>"111011011",
  45669=>"000000000",
  45670=>"111111111",
  45671=>"100100111",
  45672=>"001101111",
  45673=>"000010111",
  45674=>"000000000",
  45675=>"111111111",
  45676=>"001001100",
  45677=>"100111111",
  45678=>"111111000",
  45679=>"000000000",
  45680=>"000000111",
  45681=>"000000000",
  45682=>"000000000",
  45683=>"011010011",
  45684=>"111111111",
  45685=>"000001000",
  45686=>"111111111",
  45687=>"100111111",
  45688=>"111111001",
  45689=>"001011111",
  45690=>"111111101",
  45691=>"000000000",
  45692=>"000100100",
  45693=>"111111111",
  45694=>"111111111",
  45695=>"111111111",
  45696=>"010111111",
  45697=>"000000100",
  45698=>"010000000",
  45699=>"011111111",
  45700=>"100100111",
  45701=>"111111111",
  45702=>"000000000",
  45703=>"011111111",
  45704=>"111111111",
  45705=>"111110100",
  45706=>"111111001",
  45707=>"110110111",
  45708=>"111111111",
  45709=>"000000111",
  45710=>"100101000",
  45711=>"111111111",
  45712=>"011001001",
  45713=>"000000000",
  45714=>"111111100",
  45715=>"000000000",
  45716=>"000000000",
  45717=>"000000000",
  45718=>"111111111",
  45719=>"110000011",
  45720=>"000000000",
  45721=>"111111111",
  45722=>"000000000",
  45723=>"000000111",
  45724=>"000000010",
  45725=>"111011011",
  45726=>"111111111",
  45727=>"111001101",
  45728=>"110110110",
  45729=>"101111111",
  45730=>"001001000",
  45731=>"111111010",
  45732=>"001101101",
  45733=>"010111011",
  45734=>"000000000",
  45735=>"000000000",
  45736=>"000000000",
  45737=>"000000000",
  45738=>"000000000",
  45739=>"000000000",
  45740=>"010110100",
  45741=>"111111111",
  45742=>"111111001",
  45743=>"110111111",
  45744=>"000111000",
  45745=>"000111111",
  45746=>"010000010",
  45747=>"111111000",
  45748=>"100110111",
  45749=>"111111111",
  45750=>"000111111",
  45751=>"000000000",
  45752=>"100100000",
  45753=>"001001000",
  45754=>"100110100",
  45755=>"000000000",
  45756=>"111011011",
  45757=>"010011110",
  45758=>"100111111",
  45759=>"001000000",
  45760=>"000000000",
  45761=>"110110110",
  45762=>"000000000",
  45763=>"111111100",
  45764=>"111111111",
  45765=>"111111111",
  45766=>"000000000",
  45767=>"111110111",
  45768=>"000000000",
  45769=>"000000000",
  45770=>"101111111",
  45771=>"000000000",
  45772=>"101011011",
  45773=>"000000000",
  45774=>"000010000",
  45775=>"000000111",
  45776=>"101111111",
  45777=>"001111111",
  45778=>"000010011",
  45779=>"100000000",
  45780=>"101100100",
  45781=>"110000000",
  45782=>"000000000",
  45783=>"000000000",
  45784=>"000000111",
  45785=>"100111000",
  45786=>"111111111",
  45787=>"111111110",
  45788=>"100100000",
  45789=>"000000000",
  45790=>"111111011",
  45791=>"111111111",
  45792=>"111111111",
  45793=>"010111111",
  45794=>"111111111",
  45795=>"000001000",
  45796=>"111111111",
  45797=>"011010000",
  45798=>"000100000",
  45799=>"000000000",
  45800=>"000000111",
  45801=>"000000111",
  45802=>"000000000",
  45803=>"111111111",
  45804=>"000111111",
  45805=>"000000000",
  45806=>"110110111",
  45807=>"110111111",
  45808=>"000100110",
  45809=>"100000000",
  45810=>"011011111",
  45811=>"000000000",
  45812=>"110111010",
  45813=>"101100000",
  45814=>"000000000",
  45815=>"010000000",
  45816=>"111111111",
  45817=>"110110111",
  45818=>"111111111",
  45819=>"011011000",
  45820=>"001001001",
  45821=>"111111001",
  45822=>"010100100",
  45823=>"001101001",
  45824=>"001001011",
  45825=>"001000010",
  45826=>"000100111",
  45827=>"000000001",
  45828=>"110111000",
  45829=>"111010000",
  45830=>"000000000",
  45831=>"111101001",
  45832=>"000000011",
  45833=>"000000000",
  45834=>"000100001",
  45835=>"000000010",
  45836=>"101001001",
  45837=>"000010010",
  45838=>"100000000",
  45839=>"111111111",
  45840=>"111100100",
  45841=>"000000011",
  45842=>"010110111",
  45843=>"100100000",
  45844=>"000000001",
  45845=>"000000101",
  45846=>"100111111",
  45847=>"111010110",
  45848=>"000111101",
  45849=>"000000000",
  45850=>"000000000",
  45851=>"000011111",
  45852=>"111111111",
  45853=>"000110111",
  45854=>"000000000",
  45855=>"000110110",
  45856=>"110111010",
  45857=>"000000000",
  45858=>"111000000",
  45859=>"000000000",
  45860=>"000100100",
  45861=>"000111111",
  45862=>"000111111",
  45863=>"111111001",
  45864=>"111111111",
  45865=>"110000100",
  45866=>"000100000",
  45867=>"000000000",
  45868=>"000000000",
  45869=>"111111111",
  45870=>"000000000",
  45871=>"100000000",
  45872=>"000001111",
  45873=>"000000000",
  45874=>"000110100",
  45875=>"100000001",
  45876=>"111111111",
  45877=>"110000000",
  45878=>"110110000",
  45879=>"001011001",
  45880=>"000000000",
  45881=>"000000000",
  45882=>"000000000",
  45883=>"011111111",
  45884=>"000100111",
  45885=>"000000000",
  45886=>"000000111",
  45887=>"011111001",
  45888=>"101000001",
  45889=>"111111010",
  45890=>"101001000",
  45891=>"111111101",
  45892=>"000011110",
  45893=>"000000110",
  45894=>"110110100",
  45895=>"101000000",
  45896=>"000000000",
  45897=>"000000000",
  45898=>"000000000",
  45899=>"001100100",
  45900=>"011111110",
  45901=>"011011000",
  45902=>"000000000",
  45903=>"000100100",
  45904=>"000000000",
  45905=>"111111000",
  45906=>"110110111",
  45907=>"110111000",
  45908=>"000000000",
  45909=>"011011011",
  45910=>"011000000",
  45911=>"000000000",
  45912=>"010011011",
  45913=>"111011011",
  45914=>"011011000",
  45915=>"111111111",
  45916=>"111111111",
  45917=>"001000000",
  45918=>"111111000",
  45919=>"110110110",
  45920=>"001000011",
  45921=>"000000000",
  45922=>"000011011",
  45923=>"000001010",
  45924=>"011010000",
  45925=>"000010000",
  45926=>"000000111",
  45927=>"110000000",
  45928=>"111111110",
  45929=>"000000110",
  45930=>"000000101",
  45931=>"001111111",
  45932=>"000100110",
  45933=>"100110111",
  45934=>"111110000",
  45935=>"000000000",
  45936=>"000000000",
  45937=>"110001011",
  45938=>"110110000",
  45939=>"011001001",
  45940=>"111110010",
  45941=>"000000000",
  45942=>"000000000",
  45943=>"110110110",
  45944=>"000000100",
  45945=>"000000000",
  45946=>"000010110",
  45947=>"111100000",
  45948=>"000000000",
  45949=>"111110110",
  45950=>"100100000",
  45951=>"000000001",
  45952=>"000110000",
  45953=>"111111111",
  45954=>"000111111",
  45955=>"111111011",
  45956=>"111111111",
  45957=>"000000000",
  45958=>"011001111",
  45959=>"000000000",
  45960=>"000000000",
  45961=>"010000000",
  45962=>"111000110",
  45963=>"111111000",
  45964=>"111111111",
  45965=>"101000001",
  45966=>"000000000",
  45967=>"111111111",
  45968=>"111111111",
  45969=>"110110110",
  45970=>"001111111",
  45971=>"000000111",
  45972=>"111111111",
  45973=>"000000010",
  45974=>"101101100",
  45975=>"001000000",
  45976=>"011001000",
  45977=>"000101000",
  45978=>"100000000",
  45979=>"011011000",
  45980=>"000100111",
  45981=>"000000000",
  45982=>"000000000",
  45983=>"000000100",
  45984=>"000000010",
  45985=>"110111000",
  45986=>"111111111",
  45987=>"111000000",
  45988=>"000111111",
  45989=>"000000000",
  45990=>"000000000",
  45991=>"000000000",
  45992=>"011111111",
  45993=>"111111101",
  45994=>"000000000",
  45995=>"111111111",
  45996=>"000000010",
  45997=>"100000010",
  45998=>"000000000",
  45999=>"000000101",
  46000=>"111000000",
  46001=>"111111111",
  46002=>"011011000",
  46003=>"000000000",
  46004=>"000000000",
  46005=>"000000000",
  46006=>"110111111",
  46007=>"111111111",
  46008=>"111111111",
  46009=>"111111111",
  46010=>"000100111",
  46011=>"111111111",
  46012=>"001001001",
  46013=>"111111100",
  46014=>"000000000",
  46015=>"111111101",
  46016=>"000111111",
  46017=>"000011000",
  46018=>"011001011",
  46019=>"000000000",
  46020=>"111111011",
  46021=>"110111111",
  46022=>"111111111",
  46023=>"111111001",
  46024=>"000000000",
  46025=>"111100000",
  46026=>"000000000",
  46027=>"000000000",
  46028=>"000000000",
  46029=>"000000000",
  46030=>"111111111",
  46031=>"111110110",
  46032=>"100100000",
  46033=>"111111000",
  46034=>"110111110",
  46035=>"111111111",
  46036=>"000001001",
  46037=>"000000001",
  46038=>"111111111",
  46039=>"000000000",
  46040=>"111111110",
  46041=>"011011111",
  46042=>"000000000",
  46043=>"000111000",
  46044=>"000000000",
  46045=>"111011001",
  46046=>"111111111",
  46047=>"100110110",
  46048=>"000000000",
  46049=>"000110000",
  46050=>"111111111",
  46051=>"111111111",
  46052=>"111110000",
  46053=>"010011000",
  46054=>"111000111",
  46055=>"010000000",
  46056=>"111111000",
  46057=>"110000010",
  46058=>"001000000",
  46059=>"110111100",
  46060=>"001001001",
  46061=>"111111110",
  46062=>"111011001",
  46063=>"000000000",
  46064=>"110110100",
  46065=>"000000000",
  46066=>"000000000",
  46067=>"000100100",
  46068=>"111111111",
  46069=>"111011011",
  46070=>"111111110",
  46071=>"111111111",
  46072=>"111111111",
  46073=>"111111110",
  46074=>"011111110",
  46075=>"111111111",
  46076=>"110111111",
  46077=>"111001001",
  46078=>"001010111",
  46079=>"111111000",
  46080=>"000000000",
  46081=>"000001011",
  46082=>"111111111",
  46083=>"000001111",
  46084=>"001100110",
  46085=>"010000000",
  46086=>"000000000",
  46087=>"111111111",
  46088=>"101100000",
  46089=>"000001111",
  46090=>"010000000",
  46091=>"101101100",
  46092=>"100110001",
  46093=>"000000001",
  46094=>"111110110",
  46095=>"110111110",
  46096=>"000000110",
  46097=>"000011000",
  46098=>"000000000",
  46099=>"100000000",
  46100=>"111111111",
  46101=>"100111111",
  46102=>"001111111",
  46103=>"111111111",
  46104=>"110110111",
  46105=>"010100111",
  46106=>"111111111",
  46107=>"000000111",
  46108=>"000100100",
  46109=>"000000000",
  46110=>"100101111",
  46111=>"111111011",
  46112=>"000000000",
  46113=>"111111111",
  46114=>"111100000",
  46115=>"001000000",
  46116=>"000100111",
  46117=>"111111100",
  46118=>"000000000",
  46119=>"000000101",
  46120=>"111111111",
  46121=>"000000000",
  46122=>"111111111",
  46123=>"011000000",
  46124=>"110110001",
  46125=>"111111000",
  46126=>"001000111",
  46127=>"001111001",
  46128=>"000001111",
  46129=>"110000000",
  46130=>"011011000",
  46131=>"000001000",
  46132=>"000010000",
  46133=>"000111111",
  46134=>"000110110",
  46135=>"111001011",
  46136=>"111111111",
  46137=>"011111000",
  46138=>"000000000",
  46139=>"111111111",
  46140=>"100000000",
  46141=>"101001001",
  46142=>"001001000",
  46143=>"001010000",
  46144=>"000010111",
  46145=>"000000111",
  46146=>"000000000",
  46147=>"111110000",
  46148=>"110111111",
  46149=>"001000110",
  46150=>"000000000",
  46151=>"000000000",
  46152=>"111111111",
  46153=>"111000000",
  46154=>"000000000",
  46155=>"111111111",
  46156=>"001100100",
  46157=>"000000111",
  46158=>"000000111",
  46159=>"011110110",
  46160=>"000100111",
  46161=>"000000000",
  46162=>"110000001",
  46163=>"011000001",
  46164=>"000111111",
  46165=>"000000000",
  46166=>"000000100",
  46167=>"000000000",
  46168=>"000111111",
  46169=>"100000001",
  46170=>"101111111",
  46171=>"000001001",
  46172=>"000010000",
  46173=>"010000000",
  46174=>"111001000",
  46175=>"000000100",
  46176=>"000100100",
  46177=>"111000011",
  46178=>"111111111",
  46179=>"000000111",
  46180=>"000000101",
  46181=>"000000000",
  46182=>"101000000",
  46183=>"000000000",
  46184=>"000101111",
  46185=>"110111111",
  46186=>"111111111",
  46187=>"000011000",
  46188=>"110111001",
  46189=>"011011000",
  46190=>"110100110",
  46191=>"110011011",
  46192=>"111111111",
  46193=>"000000111",
  46194=>"000000011",
  46195=>"000001001",
  46196=>"110111000",
  46197=>"111110110",
  46198=>"111000000",
  46199=>"000000000",
  46200=>"110000000",
  46201=>"111111011",
  46202=>"010010111",
  46203=>"000000000",
  46204=>"110111111",
  46205=>"000010110",
  46206=>"001000000",
  46207=>"000000000",
  46208=>"111111111",
  46209=>"111000000",
  46210=>"000100100",
  46211=>"011001011",
  46212=>"111000000",
  46213=>"000000111",
  46214=>"000000100",
  46215=>"000000001",
  46216=>"111110000",
  46217=>"010000000",
  46218=>"000011110",
  46219=>"111111111",
  46220=>"110000000",
  46221=>"111010000",
  46222=>"011001000",
  46223=>"110000000",
  46224=>"110111111",
  46225=>"001011110",
  46226=>"100010001",
  46227=>"100100111",
  46228=>"000000000",
  46229=>"000000110",
  46230=>"000100111",
  46231=>"110010000",
  46232=>"110101011",
  46233=>"110110000",
  46234=>"000000000",
  46235=>"000111111",
  46236=>"111111000",
  46237=>"000000101",
  46238=>"110110011",
  46239=>"000000000",
  46240=>"000000000",
  46241=>"000000011",
  46242=>"110100001",
  46243=>"001001000",
  46244=>"100100110",
  46245=>"111100000",
  46246=>"111111111",
  46247=>"001101111",
  46248=>"111111111",
  46249=>"000000100",
  46250=>"000000000",
  46251=>"011011000",
  46252=>"111111000",
  46253=>"100000111",
  46254=>"111100000",
  46255=>"000010111",
  46256=>"000111111",
  46257=>"100001100",
  46258=>"111111111",
  46259=>"111111100",
  46260=>"110000111",
  46261=>"111011000",
  46262=>"111111111",
  46263=>"111000000",
  46264=>"000000111",
  46265=>"001000111",
  46266=>"000111111",
  46267=>"111001001",
  46268=>"000000011",
  46269=>"011101111",
  46270=>"011000000",
  46271=>"111000000",
  46272=>"000011111",
  46273=>"111111111",
  46274=>"100111110",
  46275=>"111111111",
  46276=>"111111111",
  46277=>"001000111",
  46278=>"000100110",
  46279=>"010011000",
  46280=>"001000000",
  46281=>"111111100",
  46282=>"111001000",
  46283=>"001001001",
  46284=>"000100111",
  46285=>"000000000",
  46286=>"111011111",
  46287=>"000000000",
  46288=>"111001000",
  46289=>"000000000",
  46290=>"000000110",
  46291=>"111111010",
  46292=>"100100000",
  46293=>"111101111",
  46294=>"000000010",
  46295=>"000000000",
  46296=>"000000000",
  46297=>"111111001",
  46298=>"001000000",
  46299=>"000000000",
  46300=>"111011011",
  46301=>"000000001",
  46302=>"001011000",
  46303=>"111000000",
  46304=>"111111111",
  46305=>"100000100",
  46306=>"111111111",
  46307=>"000111111",
  46308=>"111111001",
  46309=>"000000000",
  46310=>"000000000",
  46311=>"000000000",
  46312=>"011011100",
  46313=>"111011111",
  46314=>"111000000",
  46315=>"011111001",
  46316=>"000111111",
  46317=>"000000000",
  46318=>"111111011",
  46319=>"000101111",
  46320=>"000000011",
  46321=>"111110111",
  46322=>"000000111",
  46323=>"010111110",
  46324=>"000000000",
  46325=>"100100111",
  46326=>"100000111",
  46327=>"111111000",
  46328=>"000011000",
  46329=>"011001000",
  46330=>"111111111",
  46331=>"000000000",
  46332=>"111111111",
  46333=>"111111111",
  46334=>"111111111",
  46335=>"000111110",
  46336=>"111111100",
  46337=>"000100100",
  46338=>"110111111",
  46339=>"000110101",
  46340=>"111000000",
  46341=>"111111000",
  46342=>"101100000",
  46343=>"111111111",
  46344=>"000000100",
  46345=>"000110111",
  46346=>"000001001",
  46347=>"111111111",
  46348=>"111010111",
  46349=>"011001001",
  46350=>"000000111",
  46351=>"000111111",
  46352=>"000000000",
  46353=>"111111000",
  46354=>"000000000",
  46355=>"111100000",
  46356=>"000000000",
  46357=>"000000111",
  46358=>"011000111",
  46359=>"000111111",
  46360=>"011101111",
  46361=>"100100110",
  46362=>"000000000",
  46363=>"111000000",
  46364=>"111111111",
  46365=>"111111001",
  46366=>"111000000",
  46367=>"110110111",
  46368=>"100111000",
  46369=>"000000000",
  46370=>"011011000",
  46371=>"011110011",
  46372=>"100010010",
  46373=>"000010111",
  46374=>"001111111",
  46375=>"010010111",
  46376=>"111000111",
  46377=>"000110111",
  46378=>"011000000",
  46379=>"000000000",
  46380=>"000000000",
  46381=>"001110110",
  46382=>"000111000",
  46383=>"000011111",
  46384=>"000000011",
  46385=>"000110100",
  46386=>"001111101",
  46387=>"111000000",
  46388=>"111100000",
  46389=>"000010000",
  46390=>"000000000",
  46391=>"000111011",
  46392=>"000000000",
  46393=>"000000100",
  46394=>"010110110",
  46395=>"000000100",
  46396=>"111111011",
  46397=>"100111111",
  46398=>"000111111",
  46399=>"111111111",
  46400=>"111111111",
  46401=>"111111111",
  46402=>"111111111",
  46403=>"111111111",
  46404=>"111000110",
  46405=>"000101111",
  46406=>"111111001",
  46407=>"001000000",
  46408=>"000000111",
  46409=>"111111000",
  46410=>"100001001",
  46411=>"011011011",
  46412=>"000000000",
  46413=>"111000000",
  46414=>"100111101",
  46415=>"001001011",
  46416=>"000000000",
  46417=>"000000000",
  46418=>"001000011",
  46419=>"011000001",
  46420=>"000000000",
  46421=>"011011011",
  46422=>"001011111",
  46423=>"001100000",
  46424=>"111111111",
  46425=>"000100111",
  46426=>"111000000",
  46427=>"000111000",
  46428=>"111001000",
  46429=>"110110111",
  46430=>"000000001",
  46431=>"000000101",
  46432=>"000111111",
  46433=>"001000000",
  46434=>"001100111",
  46435=>"000000001",
  46436=>"001001001",
  46437=>"000001001",
  46438=>"111010011",
  46439=>"111000001",
  46440=>"100110111",
  46441=>"100000000",
  46442=>"010110111",
  46443=>"111111111",
  46444=>"000000000",
  46445=>"000001001",
  46446=>"000000000",
  46447=>"111111111",
  46448=>"111111000",
  46449=>"111111111",
  46450=>"111011111",
  46451=>"111111100",
  46452=>"110111111",
  46453=>"111111001",
  46454=>"110000111",
  46455=>"010000001",
  46456=>"111111111",
  46457=>"111001111",
  46458=>"000001111",
  46459=>"000000000",
  46460=>"100110000",
  46461=>"111010000",
  46462=>"111011000",
  46463=>"011000110",
  46464=>"111111111",
  46465=>"001110111",
  46466=>"000100111",
  46467=>"000000000",
  46468=>"010000000",
  46469=>"000000000",
  46470=>"111111000",
  46471=>"101000000",
  46472=>"000111111",
  46473=>"111011000",
  46474=>"111111111",
  46475=>"111111011",
  46476=>"000010010",
  46477=>"001111111",
  46478=>"111111000",
  46479=>"111111111",
  46480=>"000000000",
  46481=>"000000000",
  46482=>"000000011",
  46483=>"110111100",
  46484=>"000000010",
  46485=>"000000110",
  46486=>"101000001",
  46487=>"000000001",
  46488=>"011000111",
  46489=>"000000001",
  46490=>"111100110",
  46491=>"101111111",
  46492=>"111111011",
  46493=>"111111100",
  46494=>"111011001",
  46495=>"110111111",
  46496=>"111000000",
  46497=>"110110110",
  46498=>"000001000",
  46499=>"111000000",
  46500=>"000100000",
  46501=>"111111111",
  46502=>"111111111",
  46503=>"011000000",
  46504=>"101110111",
  46505=>"111111000",
  46506=>"000000001",
  46507=>"001011001",
  46508=>"000000000",
  46509=>"001010000",
  46510=>"100110111",
  46511=>"111111111",
  46512=>"110000010",
  46513=>"000000110",
  46514=>"100000100",
  46515=>"111111000",
  46516=>"000000000",
  46517=>"000100100",
  46518=>"111000000",
  46519=>"111100111",
  46520=>"111001001",
  46521=>"111010110",
  46522=>"100100111",
  46523=>"000100111",
  46524=>"010100101",
  46525=>"111111111",
  46526=>"110100111",
  46527=>"100100111",
  46528=>"111111110",
  46529=>"111111111",
  46530=>"000000000",
  46531=>"001111111",
  46532=>"111111101",
  46533=>"000000011",
  46534=>"000000111",
  46535=>"000111000",
  46536=>"110111111",
  46537=>"000000000",
  46538=>"111111111",
  46539=>"000000000",
  46540=>"000000000",
  46541=>"110000010",
  46542=>"110010110",
  46543=>"111111111",
  46544=>"111111111",
  46545=>"100110110",
  46546=>"000000000",
  46547=>"111111110",
  46548=>"000010100",
  46549=>"000011000",
  46550=>"111110000",
  46551=>"000000000",
  46552=>"101101100",
  46553=>"111100111",
  46554=>"000000110",
  46555=>"011111111",
  46556=>"111000000",
  46557=>"000000000",
  46558=>"010000001",
  46559=>"000100000",
  46560=>"001111111",
  46561=>"001000101",
  46562=>"111111111",
  46563=>"000000000",
  46564=>"111111011",
  46565=>"000000101",
  46566=>"000000110",
  46567=>"010000000",
  46568=>"111001111",
  46569=>"010000000",
  46570=>"001001000",
  46571=>"111111111",
  46572=>"000000101",
  46573=>"001000000",
  46574=>"111000000",
  46575=>"011111100",
  46576=>"101110110",
  46577=>"000000000",
  46578=>"000000000",
  46579=>"111111101",
  46580=>"110100000",
  46581=>"000000011",
  46582=>"111110111",
  46583=>"111011001",
  46584=>"111111000",
  46585=>"001001000",
  46586=>"111111000",
  46587=>"111111000",
  46588=>"111111100",
  46589=>"000000000",
  46590=>"000000000",
  46591=>"000000001",
  46592=>"111111010",
  46593=>"000000011",
  46594=>"100000000",
  46595=>"000000001",
  46596=>"110000000",
  46597=>"000000000",
  46598=>"000101101",
  46599=>"000000000",
  46600=>"111111111",
  46601=>"010000000",
  46602=>"111011000",
  46603=>"011111111",
  46604=>"000100100",
  46605=>"000000000",
  46606=>"010010111",
  46607=>"001100100",
  46608=>"001001001",
  46609=>"111000000",
  46610=>"101000000",
  46611=>"111100000",
  46612=>"111110000",
  46613=>"111110110",
  46614=>"110100000",
  46615=>"111111111",
  46616=>"000001001",
  46617=>"111111110",
  46618=>"111000000",
  46619=>"010000000",
  46620=>"011000000",
  46621=>"000101111",
  46622=>"000000101",
  46623=>"111111111",
  46624=>"100100110",
  46625=>"011001111",
  46626=>"110111111",
  46627=>"100111111",
  46628=>"000000001",
  46629=>"000111111",
  46630=>"111111111",
  46631=>"001000100",
  46632=>"111111111",
  46633=>"000100100",
  46634=>"111111111",
  46635=>"000000000",
  46636=>"111111111",
  46637=>"111111111",
  46638=>"111111011",
  46639=>"111111111",
  46640=>"000111111",
  46641=>"111111111",
  46642=>"011011001",
  46643=>"000000000",
  46644=>"000001000",
  46645=>"011001001",
  46646=>"000001001",
  46647=>"011000000",
  46648=>"111111100",
  46649=>"000100100",
  46650=>"000000011",
  46651=>"101000000",
  46652=>"111111100",
  46653=>"011111101",
  46654=>"100000000",
  46655=>"011011000",
  46656=>"000100000",
  46657=>"001000100",
  46658=>"111011001",
  46659=>"000000000",
  46660=>"110110110",
  46661=>"000000000",
  46662=>"111111111",
  46663=>"100000100",
  46664=>"110111111",
  46665=>"000000000",
  46666=>"111111111",
  46667=>"000000000",
  46668=>"111011000",
  46669=>"111111111",
  46670=>"010000111",
  46671=>"000110100",
  46672=>"111111001",
  46673=>"110110110",
  46674=>"000100100",
  46675=>"100101100",
  46676=>"111111111",
  46677=>"000111111",
  46678=>"001111111",
  46679=>"010000000",
  46680=>"111110111",
  46681=>"111111101",
  46682=>"111111011",
  46683=>"111111001",
  46684=>"000010111",
  46685=>"110111111",
  46686=>"000110110",
  46687=>"100110110",
  46688=>"110000000",
  46689=>"110110110",
  46690=>"000010010",
  46691=>"100100110",
  46692=>"110000000",
  46693=>"000000110",
  46694=>"001011010",
  46695=>"111111111",
  46696=>"110000000",
  46697=>"001000000",
  46698=>"000000000",
  46699=>"111111111",
  46700=>"011011111",
  46701=>"111111111",
  46702=>"000000010",
  46703=>"000000000",
  46704=>"111111111",
  46705=>"000000000",
  46706=>"011001000",
  46707=>"100111000",
  46708=>"000000000",
  46709=>"001111111",
  46710=>"000001001",
  46711=>"011111111",
  46712=>"111001000",
  46713=>"111000100",
  46714=>"100100101",
  46715=>"000000000",
  46716=>"011011110",
  46717=>"011111011",
  46718=>"000000000",
  46719=>"111111111",
  46720=>"000000000",
  46721=>"000001111",
  46722=>"000000000",
  46723=>"000000000",
  46724=>"000000000",
  46725=>"000000100",
  46726=>"011111000",
  46727=>"111100110",
  46728=>"111111111",
  46729=>"000000000",
  46730=>"000000000",
  46731=>"001001000",
  46732=>"010111110",
  46733=>"110110110",
  46734=>"010000100",
  46735=>"000000000",
  46736=>"000000101",
  46737=>"111111111",
  46738=>"000000000",
  46739=>"111111011",
  46740=>"000000110",
  46741=>"000000000",
  46742=>"000100100",
  46743=>"001011011",
  46744=>"000000000",
  46745=>"000100111",
  46746=>"111110100",
  46747=>"111111111",
  46748=>"000101111",
  46749=>"011000000",
  46750=>"000000000",
  46751=>"000000100",
  46752=>"000000001",
  46753=>"011001111",
  46754=>"100100101",
  46755=>"111111000",
  46756=>"000110110",
  46757=>"000000000",
  46758=>"111111111",
  46759=>"111111111",
  46760=>"001001001",
  46761=>"001000101",
  46762=>"101101000",
  46763=>"111111111",
  46764=>"010000000",
  46765=>"001001111",
  46766=>"111111111",
  46767=>"100111111",
  46768=>"000000000",
  46769=>"111111111",
  46770=>"111111110",
  46771=>"111000111",
  46772=>"011011111",
  46773=>"111111111",
  46774=>"111111111",
  46775=>"000000000",
  46776=>"100101111",
  46777=>"111111110",
  46778=>"011100101",
  46779=>"001111111",
  46780=>"111111111",
  46781=>"000000000",
  46782=>"101001000",
  46783=>"011011011",
  46784=>"001111111",
  46785=>"011011001",
  46786=>"010111111",
  46787=>"001011011",
  46788=>"111111111",
  46789=>"000000000",
  46790=>"101111111",
  46791=>"000000000",
  46792=>"000010010",
  46793=>"000101000",
  46794=>"000000000",
  46795=>"000100111",
  46796=>"000011111",
  46797=>"111100000",
  46798=>"000000000",
  46799=>"110100000",
  46800=>"111111111",
  46801=>"011110100",
  46802=>"000000111",
  46803=>"000000000",
  46804=>"000110111",
  46805=>"000011111",
  46806=>"110010010",
  46807=>"111111001",
  46808=>"000000110",
  46809=>"111111001",
  46810=>"000000000",
  46811=>"111111111",
  46812=>"111111001",
  46813=>"111001101",
  46814=>"000000001",
  46815=>"000100110",
  46816=>"000000011",
  46817=>"110100110",
  46818=>"111111111",
  46819=>"000000000",
  46820=>"101000000",
  46821=>"111110110",
  46822=>"111111111",
  46823=>"111001101",
  46824=>"111111111",
  46825=>"110010110",
  46826=>"000011111",
  46827=>"110000111",
  46828=>"011111110",
  46829=>"001000000",
  46830=>"011000000",
  46831=>"111001111",
  46832=>"011100000",
  46833=>"111111011",
  46834=>"111111111",
  46835=>"000110111",
  46836=>"000001111",
  46837=>"011011011",
  46838=>"000000000",
  46839=>"001001101",
  46840=>"000000000",
  46841=>"111111111",
  46842=>"001111111",
  46843=>"000100111",
  46844=>"110110111",
  46845=>"110000000",
  46846=>"111111111",
  46847=>"101000000",
  46848=>"000010000",
  46849=>"111110110",
  46850=>"000000000",
  46851=>"000000000",
  46852=>"000000000",
  46853=>"011000110",
  46854=>"001001011",
  46855=>"000001101",
  46856=>"111111000",
  46857=>"100000111",
  46858=>"111111000",
  46859=>"000110111",
  46860=>"111110100",
  46861=>"111011010",
  46862=>"000000011",
  46863=>"100100110",
  46864=>"000000000",
  46865=>"000000100",
  46866=>"110000000",
  46867=>"001111111",
  46868=>"110011111",
  46869=>"111111111",
  46870=>"111101110",
  46871=>"000111111",
  46872=>"000110110",
  46873=>"111111111",
  46874=>"110111111",
  46875=>"111111111",
  46876=>"001000000",
  46877=>"000000000",
  46878=>"111011000",
  46879=>"000000000",
  46880=>"011000001",
  46881=>"000010011",
  46882=>"000110010",
  46883=>"000000000",
  46884=>"001100000",
  46885=>"000000000",
  46886=>"000000001",
  46887=>"001000000",
  46888=>"111110110",
  46889=>"111001001",
  46890=>"011111000",
  46891=>"111111010",
  46892=>"110111111",
  46893=>"111110110",
  46894=>"110000100",
  46895=>"111110110",
  46896=>"001011111",
  46897=>"001000000",
  46898=>"111110010",
  46899=>"000000000",
  46900=>"111111011",
  46901=>"000000011",
  46902=>"000000000",
  46903=>"110111111",
  46904=>"000101111",
  46905=>"000011111",
  46906=>"111111110",
  46907=>"000000111",
  46908=>"000000000",
  46909=>"011111111",
  46910=>"000010100",
  46911=>"000000111",
  46912=>"000000011",
  46913=>"111111111",
  46914=>"110010000",
  46915=>"000000000",
  46916=>"000000000",
  46917=>"000000010",
  46918=>"001001111",
  46919=>"111110111",
  46920=>"000110100",
  46921=>"111000001",
  46922=>"111111111",
  46923=>"010000000",
  46924=>"000100111",
  46925=>"000000111",
  46926=>"111111111",
  46927=>"100000000",
  46928=>"100111111",
  46929=>"111111111",
  46930=>"111111000",
  46931=>"000000000",
  46932=>"000100000",
  46933=>"000100100",
  46934=>"100000010",
  46935=>"011011111",
  46936=>"001000000",
  46937=>"000000000",
  46938=>"111111111",
  46939=>"011111110",
  46940=>"111111001",
  46941=>"100000100",
  46942=>"110110111",
  46943=>"000000001",
  46944=>"000000001",
  46945=>"111111000",
  46946=>"000000101",
  46947=>"111111011",
  46948=>"110010000",
  46949=>"000000000",
  46950=>"000000101",
  46951=>"000001000",
  46952=>"011001000",
  46953=>"001011111",
  46954=>"111110111",
  46955=>"111111110",
  46956=>"000000001",
  46957=>"000001001",
  46958=>"111000000",
  46959=>"000110110",
  46960=>"111110110",
  46961=>"111111111",
  46962=>"000000000",
  46963=>"111011011",
  46964=>"001000000",
  46965=>"110111111",
  46966=>"000000000",
  46967=>"000110111",
  46968=>"100100000",
  46969=>"000100100",
  46970=>"000100111",
  46971=>"110111110",
  46972=>"111111000",
  46973=>"000001111",
  46974=>"000000000",
  46975=>"011000000",
  46976=>"001001001",
  46977=>"000000111",
  46978=>"000000000",
  46979=>"000000000",
  46980=>"111111111",
  46981=>"011001000",
  46982=>"111111111",
  46983=>"010110111",
  46984=>"111111111",
  46985=>"111111110",
  46986=>"111111111",
  46987=>"111101000",
  46988=>"111111101",
  46989=>"000000000",
  46990=>"111111111",
  46991=>"111111111",
  46992=>"111001000",
  46993=>"111111111",
  46994=>"111111111",
  46995=>"000000000",
  46996=>"111001111",
  46997=>"010000000",
  46998=>"000000111",
  46999=>"001001001",
  47000=>"000000111",
  47001=>"111111110",
  47002=>"010000001",
  47003=>"000000000",
  47004=>"000111000",
  47005=>"000000000",
  47006=>"011111111",
  47007=>"100100000",
  47008=>"101100111",
  47009=>"011000000",
  47010=>"000100101",
  47011=>"111111000",
  47012=>"000000000",
  47013=>"111111111",
  47014=>"111100111",
  47015=>"111111111",
  47016=>"000000000",
  47017=>"000000010",
  47018=>"000000000",
  47019=>"011001001",
  47020=>"000000000",
  47021=>"001111100",
  47022=>"000000000",
  47023=>"111011000",
  47024=>"100000111",
  47025=>"000000000",
  47026=>"000000000",
  47027=>"000000101",
  47028=>"111111111",
  47029=>"000000001",
  47030=>"111100000",
  47031=>"000000010",
  47032=>"000000000",
  47033=>"000111011",
  47034=>"110110000",
  47035=>"111111111",
  47036=>"111111101",
  47037=>"111111100",
  47038=>"100111110",
  47039=>"111111011",
  47040=>"111000100",
  47041=>"000000000",
  47042=>"000000000",
  47043=>"000000000",
  47044=>"111111100",
  47045=>"110010000",
  47046=>"000000000",
  47047=>"111111111",
  47048=>"000111011",
  47049=>"100010000",
  47050=>"111000001",
  47051=>"000111111",
  47052=>"100111111",
  47053=>"001111111",
  47054=>"000101101",
  47055=>"111111111",
  47056=>"111111111",
  47057=>"000000011",
  47058=>"111111111",
  47059=>"000000000",
  47060=>"000100111",
  47061=>"111001001",
  47062=>"110110111",
  47063=>"000011001",
  47064=>"001101000",
  47065=>"111101001",
  47066=>"111111110",
  47067=>"111101100",
  47068=>"011011000",
  47069=>"001001001",
  47070=>"111111111",
  47071=>"111111011",
  47072=>"111111111",
  47073=>"111111111",
  47074=>"111000101",
  47075=>"000111111",
  47076=>"010111111",
  47077=>"001000000",
  47078=>"111111111",
  47079=>"000000000",
  47080=>"000000000",
  47081=>"001111000",
  47082=>"101110110",
  47083=>"000000000",
  47084=>"111111111",
  47085=>"100100000",
  47086=>"111111111",
  47087=>"011111111",
  47088=>"111111111",
  47089=>"111000000",
  47090=>"000000000",
  47091=>"000111101",
  47092=>"011111111",
  47093=>"101001111",
  47094=>"110000000",
  47095=>"001000000",
  47096=>"000000111",
  47097=>"100000001",
  47098=>"000000001",
  47099=>"000000000",
  47100=>"000011000",
  47101=>"001001111",
  47102=>"001001000",
  47103=>"110000111",
  47104=>"111100111",
  47105=>"001000010",
  47106=>"000000100",
  47107=>"110000000",
  47108=>"111000000",
  47109=>"111110010",
  47110=>"000010000",
  47111=>"000000000",
  47112=>"000100110",
  47113=>"001001000",
  47114=>"000001111",
  47115=>"000000111",
  47116=>"001000000",
  47117=>"111000000",
  47118=>"111110101",
  47119=>"000000000",
  47120=>"111111111",
  47121=>"000111111",
  47122=>"000000000",
  47123=>"000000000",
  47124=>"010000001",
  47125=>"000000111",
  47126=>"000000000",
  47127=>"000101111",
  47128=>"001011111",
  47129=>"110110111",
  47130=>"011011011",
  47131=>"111000000",
  47132=>"111111111",
  47133=>"000111111",
  47134=>"111111101",
  47135=>"110110111",
  47136=>"011000000",
  47137=>"000001101",
  47138=>"001001111",
  47139=>"111001111",
  47140=>"000000000",
  47141=>"000000100",
  47142=>"010111111",
  47143=>"111000000",
  47144=>"111111101",
  47145=>"000000000",
  47146=>"011011111",
  47147=>"111111111",
  47148=>"011111111",
  47149=>"111111111",
  47150=>"000000000",
  47151=>"000000110",
  47152=>"000000000",
  47153=>"000000000",
  47154=>"000000110",
  47155=>"001000000",
  47156=>"000001001",
  47157=>"111101011",
  47158=>"011111111",
  47159=>"000000000",
  47160=>"000000000",
  47161=>"111101111",
  47162=>"000000000",
  47163=>"111011111",
  47164=>"000000000",
  47165=>"001000000",
  47166=>"111111111",
  47167=>"111111111",
  47168=>"000011011",
  47169=>"000000000",
  47170=>"000110000",
  47171=>"111111011",
  47172=>"000111111",
  47173=>"111111111",
  47174=>"000000111",
  47175=>"000000101",
  47176=>"110110001",
  47177=>"000000000",
  47178=>"011011111",
  47179=>"000000001",
  47180=>"000000011",
  47181=>"000000000",
  47182=>"000010111",
  47183=>"000000000",
  47184=>"001110110",
  47185=>"000000100",
  47186=>"111111111",
  47187=>"111100111",
  47188=>"001000001",
  47189=>"000010000",
  47190=>"001001000",
  47191=>"010000000",
  47192=>"000000000",
  47193=>"000000101",
  47194=>"000110111",
  47195=>"110111001",
  47196=>"000000110",
  47197=>"000111110",
  47198=>"000000000",
  47199=>"000000000",
  47200=>"000011111",
  47201=>"000000000",
  47202=>"011111111",
  47203=>"000000000",
  47204=>"111101111",
  47205=>"000000000",
  47206=>"001011011",
  47207=>"000011111",
  47208=>"110110111",
  47209=>"111111111",
  47210=>"000110110",
  47211=>"110110111",
  47212=>"111111111",
  47213=>"000000110",
  47214=>"111111000",
  47215=>"111111111",
  47216=>"000000000",
  47217=>"000000000",
  47218=>"111111111",
  47219=>"111111111",
  47220=>"000000000",
  47221=>"101101101",
  47222=>"101101000",
  47223=>"000000111",
  47224=>"111111111",
  47225=>"110000111",
  47226=>"000111111",
  47227=>"110110110",
  47228=>"000001111",
  47229=>"110110110",
  47230=>"000000111",
  47231=>"000111001",
  47232=>"000000000",
  47233=>"000000000",
  47234=>"000100110",
  47235=>"000000000",
  47236=>"001011011",
  47237=>"000000101",
  47238=>"000000000",
  47239=>"101101000",
  47240=>"110000000",
  47241=>"000010011",
  47242=>"111111000",
  47243=>"000000000",
  47244=>"011011000",
  47245=>"000000000",
  47246=>"100100000",
  47247=>"000000000",
  47248=>"110111111",
  47249=>"111111111",
  47250=>"000000000",
  47251=>"000001001",
  47252=>"000000110",
  47253=>"011111111",
  47254=>"000000000",
  47255=>"111111110",
  47256=>"010000000",
  47257=>"111011010",
  47258=>"111111111",
  47259=>"100110111",
  47260=>"000001000",
  47261=>"011010010",
  47262=>"011111000",
  47263=>"000001001",
  47264=>"000000001",
  47265=>"011011011",
  47266=>"000000001",
  47267=>"000000111",
  47268=>"111001001",
  47269=>"000000001",
  47270=>"111111111",
  47271=>"100101110",
  47272=>"000111100",
  47273=>"001011111",
  47274=>"111111111",
  47275=>"111000000",
  47276=>"000000000",
  47277=>"001001001",
  47278=>"000000011",
  47279=>"000000001",
  47280=>"000110111",
  47281=>"000000100",
  47282=>"000111111",
  47283=>"111111111",
  47284=>"000000000",
  47285=>"111001000",
  47286=>"111111111",
  47287=>"100100000",
  47288=>"000000011",
  47289=>"111111111",
  47290=>"111111111",
  47291=>"000000000",
  47292=>"011000000",
  47293=>"111111100",
  47294=>"111111111",
  47295=>"001010111",
  47296=>"110100000",
  47297=>"001000100",
  47298=>"011111111",
  47299=>"011000000",
  47300=>"111000000",
  47301=>"001001111",
  47302=>"000100000",
  47303=>"000000000",
  47304=>"111111111",
  47305=>"001000000",
  47306=>"100100000",
  47307=>"111000000",
  47308=>"000100111",
  47309=>"000111111",
  47310=>"000100111",
  47311=>"001111000",
  47312=>"111111111",
  47313=>"000010111",
  47314=>"111000111",
  47315=>"000000000",
  47316=>"001001011",
  47317=>"000001111",
  47318=>"111111111",
  47319=>"111111000",
  47320=>"001011000",
  47321=>"111111111",
  47322=>"001111111",
  47323=>"111100001",
  47324=>"111111110",
  47325=>"000000000",
  47326=>"000000111",
  47327=>"001101111",
  47328=>"111100101",
  47329=>"000100110",
  47330=>"111111111",
  47331=>"111011000",
  47332=>"101111001",
  47333=>"000110110",
  47334=>"110111110",
  47335=>"111111111",
  47336=>"111111101",
  47337=>"001000000",
  47338=>"011000000",
  47339=>"011000000",
  47340=>"111111000",
  47341=>"111000000",
  47342=>"111111111",
  47343=>"010000000",
  47344=>"011001111",
  47345=>"000000000",
  47346=>"110111111",
  47347=>"001000001",
  47348=>"000000000",
  47349=>"001000000",
  47350=>"111111001",
  47351=>"000111111",
  47352=>"111011000",
  47353=>"011111111",
  47354=>"000000000",
  47355=>"000010111",
  47356=>"111011000",
  47357=>"111111111",
  47358=>"000000111",
  47359=>"000000000",
  47360=>"111111111",
  47361=>"010011001",
  47362=>"000000111",
  47363=>"111100011",
  47364=>"000001001",
  47365=>"000000101",
  47366=>"000111111",
  47367=>"011111100",
  47368=>"001000000",
  47369=>"111000001",
  47370=>"000000111",
  47371=>"111111100",
  47372=>"010000000",
  47373=>"000111111",
  47374=>"011111111",
  47375=>"000111111",
  47376=>"111111111",
  47377=>"011110111",
  47378=>"100101101",
  47379=>"000000010",
  47380=>"011000000",
  47381=>"000010010",
  47382=>"011011010",
  47383=>"000111111",
  47384=>"000000001",
  47385=>"110000000",
  47386=>"000000111",
  47387=>"000000100",
  47388=>"000110110",
  47389=>"000000000",
  47390=>"111111111",
  47391=>"001110111",
  47392=>"100110111",
  47393=>"000000001",
  47394=>"000000000",
  47395=>"010000000",
  47396=>"000000000",
  47397=>"000000000",
  47398=>"111111111",
  47399=>"011010110",
  47400=>"001001000",
  47401=>"000000000",
  47402=>"001000000",
  47403=>"000000000",
  47404=>"000000000",
  47405=>"011111111",
  47406=>"000111111",
  47407=>"110110000",
  47408=>"111111111",
  47409=>"011000000",
  47410=>"001001000",
  47411=>"111111111",
  47412=>"000100111",
  47413=>"101001011",
  47414=>"110111111",
  47415=>"111111001",
  47416=>"000011001",
  47417=>"001000111",
  47418=>"111111100",
  47419=>"111111111",
  47420=>"011011010",
  47421=>"000001001",
  47422=>"101111100",
  47423=>"111111111",
  47424=>"000000011",
  47425=>"000000000",
  47426=>"001000000",
  47427=>"001111111",
  47428=>"000000000",
  47429=>"111100000",
  47430=>"011001111",
  47431=>"000001001",
  47432=>"000000000",
  47433=>"011011011",
  47434=>"111010000",
  47435=>"001001111",
  47436=>"111011111",
  47437=>"010000000",
  47438=>"000000000",
  47439=>"111111100",
  47440=>"111111011",
  47441=>"000000000",
  47442=>"111111111",
  47443=>"111001000",
  47444=>"111000111",
  47445=>"000001011",
  47446=>"111010000",
  47447=>"000000000",
  47448=>"001000000",
  47449=>"011011011",
  47450=>"111100010",
  47451=>"111011011",
  47452=>"110110111",
  47453=>"111101000",
  47454=>"000000100",
  47455=>"000000000",
  47456=>"000011111",
  47457=>"000000010",
  47458=>"111111111",
  47459=>"011000000",
  47460=>"111101000",
  47461=>"000000000",
  47462=>"111111001",
  47463=>"000110010",
  47464=>"010001011",
  47465=>"000001111",
  47466=>"000011111",
  47467=>"000000111",
  47468=>"110111110",
  47469=>"110110000",
  47470=>"000000111",
  47471=>"000011001",
  47472=>"001000000",
  47473=>"000101111",
  47474=>"111000011",
  47475=>"111110100",
  47476=>"000000000",
  47477=>"001000000",
  47478=>"000110111",
  47479=>"101100111",
  47480=>"000000000",
  47481=>"110111111",
  47482=>"000000111",
  47483=>"001001000",
  47484=>"000000001",
  47485=>"011001000",
  47486=>"111011111",
  47487=>"000000000",
  47488=>"000000000",
  47489=>"001000000",
  47490=>"111111011",
  47491=>"000001000",
  47492=>"111111111",
  47493=>"000011000",
  47494=>"000000000",
  47495=>"000001011",
  47496=>"000000000",
  47497=>"000000000",
  47498=>"000000000",
  47499=>"111111111",
  47500=>"000000110",
  47501=>"101101101",
  47502=>"111111111",
  47503=>"000000000",
  47504=>"000100101",
  47505=>"000111111",
  47506=>"111111111",
  47507=>"111111111",
  47508=>"011001101",
  47509=>"111111011",
  47510=>"111111111",
  47511=>"010000001",
  47512=>"000000111",
  47513=>"001000010",
  47514=>"101111111",
  47515=>"000000000",
  47516=>"000110110",
  47517=>"001001111",
  47518=>"111111101",
  47519=>"000000000",
  47520=>"000111101",
  47521=>"111111111",
  47522=>"001110000",
  47523=>"111100000",
  47524=>"000000000",
  47525=>"111101111",
  47526=>"000100111",
  47527=>"111111111",
  47528=>"000110111",
  47529=>"010111111",
  47530=>"000000000",
  47531=>"111110111",
  47532=>"011001001",
  47533=>"000000100",
  47534=>"111000000",
  47535=>"000001111",
  47536=>"010011111",
  47537=>"000000000",
  47538=>"000110100",
  47539=>"000000001",
  47540=>"000011111",
  47541=>"111111111",
  47542=>"111110110",
  47543=>"000000000",
  47544=>"000000000",
  47545=>"000001111",
  47546=>"000001111",
  47547=>"010010000",
  47548=>"000000000",
  47549=>"000000000",
  47550=>"000010111",
  47551=>"011001001",
  47552=>"000000000",
  47553=>"111111110",
  47554=>"000000111",
  47555=>"000000011",
  47556=>"011000000",
  47557=>"001011000",
  47558=>"000100101",
  47559=>"101111111",
  47560=>"011000001",
  47561=>"111111101",
  47562=>"000000000",
  47563=>"000001000",
  47564=>"011000000",
  47565=>"001001101",
  47566=>"001001000",
  47567=>"111111111",
  47568=>"100000000",
  47569=>"000100100",
  47570=>"111111111",
  47571=>"111101111",
  47572=>"101001110",
  47573=>"000000000",
  47574=>"000111111",
  47575=>"100011011",
  47576=>"111111111",
  47577=>"011111100",
  47578=>"111011111",
  47579=>"100111001",
  47580=>"111111010",
  47581=>"000000001",
  47582=>"111111111",
  47583=>"110111100",
  47584=>"101000000",
  47585=>"100110000",
  47586=>"010011111",
  47587=>"000000111",
  47588=>"111000111",
  47589=>"001001111",
  47590=>"100111111",
  47591=>"000000000",
  47592=>"111111111",
  47593=>"000000011",
  47594=>"011011011",
  47595=>"000110111",
  47596=>"000010000",
  47597=>"100100100",
  47598=>"111111111",
  47599=>"111111111",
  47600=>"100100111",
  47601=>"000111001",
  47602=>"000000000",
  47603=>"111110110",
  47604=>"000000000",
  47605=>"000011001",
  47606=>"000000001",
  47607=>"000111111",
  47608=>"011001001",
  47609=>"011111000",
  47610=>"111111111",
  47611=>"110111111",
  47612=>"011000000",
  47613=>"111111111",
  47614=>"000011011",
  47615=>"111000000",
  47616=>"111100000",
  47617=>"111001001",
  47618=>"111111111",
  47619=>"000000100",
  47620=>"000100000",
  47621=>"111000000",
  47622=>"001000000",
  47623=>"101111111",
  47624=>"111111111",
  47625=>"110110110",
  47626=>"110111110",
  47627=>"000000011",
  47628=>"001001000",
  47629=>"000100110",
  47630=>"000011111",
  47631=>"110000000",
  47632=>"111111101",
  47633=>"001011111",
  47634=>"000010110",
  47635=>"000000001",
  47636=>"011001001",
  47637=>"001101111",
  47638=>"100000100",
  47639=>"111101001",
  47640=>"001001011",
  47641=>"111101101",
  47642=>"111000001",
  47643=>"001000000",
  47644=>"111111111",
  47645=>"000010111",
  47646=>"011011011",
  47647=>"111001001",
  47648=>"011011111",
  47649=>"111000000",
  47650=>"011001101",
  47651=>"000000000",
  47652=>"000010011",
  47653=>"010001001",
  47654=>"000000111",
  47655=>"000001100",
  47656=>"000000100",
  47657=>"001001000",
  47658=>"000000000",
  47659=>"000000100",
  47660=>"111101001",
  47661=>"110111111",
  47662=>"101001000",
  47663=>"000000001",
  47664=>"110110011",
  47665=>"110010000",
  47666=>"110100101",
  47667=>"000000000",
  47668=>"110100100",
  47669=>"110100100",
  47670=>"000011001",
  47671=>"000000100",
  47672=>"000000100",
  47673=>"001001001",
  47674=>"000000000",
  47675=>"111110110",
  47676=>"000000000",
  47677=>"100100111",
  47678=>"111111111",
  47679=>"101100100",
  47680=>"011001111",
  47681=>"001001111",
  47682=>"111111111",
  47683=>"011011111",
  47684=>"000010100",
  47685=>"000000000",
  47686=>"100000000",
  47687=>"111111110",
  47688=>"110110110",
  47689=>"010110010",
  47690=>"000001000",
  47691=>"000110011",
  47692=>"001000000",
  47693=>"001001001",
  47694=>"110110010",
  47695=>"000001001",
  47696=>"010111111",
  47697=>"110110110",
  47698=>"000010110",
  47699=>"001011011",
  47700=>"101001001",
  47701=>"001000000",
  47702=>"111111111",
  47703=>"100100100",
  47704=>"000000000",
  47705=>"001101101",
  47706=>"000000001",
  47707=>"000011000",
  47708=>"000000001",
  47709=>"111111111",
  47710=>"000101101",
  47711=>"101001011",
  47712=>"110110111",
  47713=>"100100110",
  47714=>"010000111",
  47715=>"111111111",
  47716=>"100100100",
  47717=>"000000110",
  47718=>"111110110",
  47719=>"000000001",
  47720=>"001000000",
  47721=>"001101111",
  47722=>"001001111",
  47723=>"000000000",
  47724=>"000110110",
  47725=>"100110110",
  47726=>"110110111",
  47727=>"110110110",
  47728=>"000100111",
  47729=>"011011110",
  47730=>"111111010",
  47731=>"000000000",
  47732=>"001000000",
  47733=>"000001000",
  47734=>"110000110",
  47735=>"000100110",
  47736=>"000000000",
  47737=>"111111111",
  47738=>"101000100",
  47739=>"000000000",
  47740=>"110110110",
  47741=>"000000100",
  47742=>"111001001",
  47743=>"010000000",
  47744=>"111111111",
  47745=>"010111111",
  47746=>"000001000",
  47747=>"100110110",
  47748=>"111111111",
  47749=>"111101101",
  47750=>"000111111",
  47751=>"110110000",
  47752=>"011001001",
  47753=>"111101000",
  47754=>"000000000",
  47755=>"000110100",
  47756=>"010000000",
  47757=>"000000100",
  47758=>"110110111",
  47759=>"110111010",
  47760=>"000000001",
  47761=>"001000000",
  47762=>"111111111",
  47763=>"111100100",
  47764=>"101000111",
  47765=>"111111000",
  47766=>"001101001",
  47767=>"111111111",
  47768=>"111111000",
  47769=>"000111111",
  47770=>"000000000",
  47771=>"000000001",
  47772=>"000001011",
  47773=>"000000000",
  47774=>"011111111",
  47775=>"111110111",
  47776=>"011000010",
  47777=>"111111101",
  47778=>"000001111",
  47779=>"010001000",
  47780=>"111000000",
  47781=>"000000011",
  47782=>"110110110",
  47783=>"111111111",
  47784=>"111011000",
  47785=>"011111010",
  47786=>"000000000",
  47787=>"111110000",
  47788=>"110001011",
  47789=>"000000100",
  47790=>"100111111",
  47791=>"011011001",
  47792=>"000000010",
  47793=>"111111111",
  47794=>"111111111",
  47795=>"010000111",
  47796=>"000001101",
  47797=>"000000000",
  47798=>"111000110",
  47799=>"011010111",
  47800=>"000000000",
  47801=>"111111111",
  47802=>"111001000",
  47803=>"000001101",
  47804=>"111111111",
  47805=>"110110110",
  47806=>"000010000",
  47807=>"110010010",
  47808=>"011011011",
  47809=>"101111111",
  47810=>"101101111",
  47811=>"110000000",
  47812=>"111000000",
  47813=>"100100100",
  47814=>"000000000",
  47815=>"110010111",
  47816=>"001000111",
  47817=>"001101111",
  47818=>"001011000",
  47819=>"111011011",
  47820=>"110000000",
  47821=>"000000000",
  47822=>"001001111",
  47823=>"101001000",
  47824=>"100000000",
  47825=>"110010011",
  47826=>"111110000",
  47827=>"110101111",
  47828=>"110110100",
  47829=>"001001101",
  47830=>"010110000",
  47831=>"000100111",
  47832=>"000000000",
  47833=>"001111111",
  47834=>"000010000",
  47835=>"000000100",
  47836=>"000001111",
  47837=>"011000110",
  47838=>"110000000",
  47839=>"000011111",
  47840=>"001000000",
  47841=>"111111101",
  47842=>"001101101",
  47843=>"111111111",
  47844=>"000111111",
  47845=>"011001001",
  47846=>"111111110",
  47847=>"000000000",
  47848=>"000000000",
  47849=>"001101111",
  47850=>"000000110",
  47851=>"111111111",
  47852=>"111000000",
  47853=>"111111111",
  47854=>"111011011",
  47855=>"011111111",
  47856=>"110110111",
  47857=>"111111111",
  47858=>"110000000",
  47859=>"010010011",
  47860=>"000000100",
  47861=>"100100100",
  47862=>"111111111",
  47863=>"010011111",
  47864=>"111111111",
  47865=>"110000000",
  47866=>"001101111",
  47867=>"010110110",
  47868=>"110110110",
  47869=>"001111111",
  47870=>"000100111",
  47871=>"000001111",
  47872=>"000000000",
  47873=>"011100101",
  47874=>"100111111",
  47875=>"011000100",
  47876=>"011010010",
  47877=>"000110000",
  47878=>"111011011",
  47879=>"001001001",
  47880=>"110000100",
  47881=>"001001001",
  47882=>"000001111",
  47883=>"000000111",
  47884=>"110100110",
  47885=>"111101000",
  47886=>"000000000",
  47887=>"000100111",
  47888=>"000001000",
  47889=>"100000000",
  47890=>"111100100",
  47891=>"111101111",
  47892=>"010000000",
  47893=>"001000000",
  47894=>"111001000",
  47895=>"101101111",
  47896=>"100100000",
  47897=>"111000001",
  47898=>"001001001",
  47899=>"111111010",
  47900=>"001001001",
  47901=>"111110001",
  47902=>"000001000",
  47903=>"111111100",
  47904=>"111111011",
  47905=>"000000000",
  47906=>"000010010",
  47907=>"000001111",
  47908=>"001000000",
  47909=>"000111111",
  47910=>"110110100",
  47911=>"000000000",
  47912=>"111111000",
  47913=>"010111111",
  47914=>"010100000",
  47915=>"000111111",
  47916=>"100000000",
  47917=>"111111110",
  47918=>"001011000",
  47919=>"000111111",
  47920=>"010110010",
  47921=>"010110010",
  47922=>"000000110",
  47923=>"100100000",
  47924=>"111111111",
  47925=>"100000000",
  47926=>"011000000",
  47927=>"011000000",
  47928=>"110110110",
  47929=>"101101111",
  47930=>"000000000",
  47931=>"111111011",
  47932=>"100101111",
  47933=>"001011100",
  47934=>"000000000",
  47935=>"000000000",
  47936=>"111101101",
  47937=>"011110111",
  47938=>"111001000",
  47939=>"101001001",
  47940=>"110100100",
  47941=>"011111111",
  47942=>"001000000",
  47943=>"001001001",
  47944=>"111011000",
  47945=>"001101001",
  47946=>"101111001",
  47947=>"001011011",
  47948=>"000000000",
  47949=>"010000001",
  47950=>"000000100",
  47951=>"000000110",
  47952=>"100100100",
  47953=>"001000001",
  47954=>"000111111",
  47955=>"111111111",
  47956=>"011000000",
  47957=>"011001001",
  47958=>"111001001",
  47959=>"000010010",
  47960=>"110111111",
  47961=>"110111010",
  47962=>"011111110",
  47963=>"000000100",
  47964=>"000000000",
  47965=>"111111100",
  47966=>"000001001",
  47967=>"000000100",
  47968=>"111001001",
  47969=>"110010010",
  47970=>"100000001",
  47971=>"000000000",
  47972=>"110110111",
  47973=>"000000000",
  47974=>"000110111",
  47975=>"111111111",
  47976=>"001001001",
  47977=>"000000000",
  47978=>"111101001",
  47979=>"111110111",
  47980=>"001000000",
  47981=>"001011110",
  47982=>"110111111",
  47983=>"111111101",
  47984=>"000000000",
  47985=>"010010001",
  47986=>"110010011",
  47987=>"111000000",
  47988=>"011001000",
  47989=>"000000000",
  47990=>"000010110",
  47991=>"000000001",
  47992=>"010010010",
  47993=>"011000000",
  47994=>"111000001",
  47995=>"100000000",
  47996=>"000000000",
  47997=>"111011001",
  47998=>"110110000",
  47999=>"000000000",
  48000=>"000001000",
  48001=>"111111111",
  48002=>"001100100",
  48003=>"001000000",
  48004=>"000001101",
  48005=>"001101101",
  48006=>"000000001",
  48007=>"011001001",
  48008=>"110110010",
  48009=>"000000000",
  48010=>"011001001",
  48011=>"111001011",
  48012=>"101111111",
  48013=>"111110000",
  48014=>"010000000",
  48015=>"000000000",
  48016=>"111111010",
  48017=>"011011011",
  48018=>"111101000",
  48019=>"000000100",
  48020=>"000000010",
  48021=>"000000000",
  48022=>"000000010",
  48023=>"000000000",
  48024=>"001111111",
  48025=>"000100101",
  48026=>"010000000",
  48027=>"111000000",
  48028=>"111111111",
  48029=>"000000000",
  48030=>"111111111",
  48031=>"111101000",
  48032=>"111111111",
  48033=>"111111111",
  48034=>"111111111",
  48035=>"000010010",
  48036=>"111011100",
  48037=>"000000000",
  48038=>"010010000",
  48039=>"111111110",
  48040=>"011011000",
  48041=>"111111011",
  48042=>"011011000",
  48043=>"111000000",
  48044=>"010000000",
  48045=>"000001111",
  48046=>"000111111",
  48047=>"000000001",
  48048=>"111111111",
  48049=>"101101110",
  48050=>"111111110",
  48051=>"000001111",
  48052=>"111011011",
  48053=>"000000001",
  48054=>"000001011",
  48055=>"001111001",
  48056=>"111111001",
  48057=>"111010110",
  48058=>"001000000",
  48059=>"000111100",
  48060=>"001111101",
  48061=>"000000001",
  48062=>"110110110",
  48063=>"100111100",
  48064=>"111111111",
  48065=>"110100000",
  48066=>"110110110",
  48067=>"010111111",
  48068=>"001000101",
  48069=>"110110000",
  48070=>"000000001",
  48071=>"010010000",
  48072=>"000000000",
  48073=>"000001001",
  48074=>"000000000",
  48075=>"100111111",
  48076=>"111000001",
  48077=>"000000110",
  48078=>"000000110",
  48079=>"000001001",
  48080=>"011111000",
  48081=>"011111111",
  48082=>"000000000",
  48083=>"000000001",
  48084=>"111111000",
  48085=>"111111111",
  48086=>"000000000",
  48087=>"100000100",
  48088=>"111110110",
  48089=>"111111111",
  48090=>"000000001",
  48091=>"000001000",
  48092=>"111111011",
  48093=>"000000000",
  48094=>"001000000",
  48095=>"001011111",
  48096=>"001001001",
  48097=>"000000000",
  48098=>"001001001",
  48099=>"000000111",
  48100=>"111011001",
  48101=>"000001101",
  48102=>"100000111",
  48103=>"001000000",
  48104=>"010110000",
  48105=>"011000000",
  48106=>"011011011",
  48107=>"111100111",
  48108=>"001001101",
  48109=>"111001001",
  48110=>"111000100",
  48111=>"000001000",
  48112=>"111111111",
  48113=>"110111111",
  48114=>"000010000",
  48115=>"001000110",
  48116=>"000110110",
  48117=>"011011000",
  48118=>"111001000",
  48119=>"001001001",
  48120=>"110111111",
  48121=>"110110110",
  48122=>"000000000",
  48123=>"111110110",
  48124=>"010010000",
  48125=>"111111111",
  48126=>"110000110",
  48127=>"010000110",
  48128=>"000000110",
  48129=>"111000010",
  48130=>"000000000",
  48131=>"111111111",
  48132=>"001001011",
  48133=>"000000000",
  48134=>"000000000",
  48135=>"010011111",
  48136=>"011111111",
  48137=>"111100000",
  48138=>"100000111",
  48139=>"110111111",
  48140=>"000000001",
  48141=>"011000001",
  48142=>"100110110",
  48143=>"100101111",
  48144=>"110110110",
  48145=>"000000000",
  48146=>"001001101",
  48147=>"010010000",
  48148=>"000000000",
  48149=>"111110110",
  48150=>"000000111",
  48151=>"001011011",
  48152=>"110110110",
  48153=>"100001001",
  48154=>"000000001",
  48155=>"011000000",
  48156=>"001001111",
  48157=>"000000100",
  48158=>"001001000",
  48159=>"011110110",
  48160=>"010000010",
  48161=>"110111111",
  48162=>"011110110",
  48163=>"000001001",
  48164=>"111111001",
  48165=>"001000100",
  48166=>"000000000",
  48167=>"000101111",
  48168=>"111011000",
  48169=>"101101100",
  48170=>"111111111",
  48171=>"000000000",
  48172=>"000100111",
  48173=>"011010000",
  48174=>"101101101",
  48175=>"110010000",
  48176=>"011010111",
  48177=>"001101101",
  48178=>"011000000",
  48179=>"111111000",
  48180=>"101101100",
  48181=>"000100001",
  48182=>"000001000",
  48183=>"000000000",
  48184=>"111110010",
  48185=>"010010111",
  48186=>"000000001",
  48187=>"011010010",
  48188=>"101101101",
  48189=>"111111111",
  48190=>"001010010",
  48191=>"011111111",
  48192=>"010011111",
  48193=>"111111111",
  48194=>"101111101",
  48195=>"111111010",
  48196=>"001011110",
  48197=>"000001001",
  48198=>"011010010",
  48199=>"010011111",
  48200=>"011001001",
  48201=>"110100111",
  48202=>"011111111",
  48203=>"010110010",
  48204=>"010110111",
  48205=>"111110100",
  48206=>"011010000",
  48207=>"111111111",
  48208=>"000000000",
  48209=>"111111111",
  48210=>"000001101",
  48211=>"011001000",
  48212=>"111111000",
  48213=>"010010000",
  48214=>"110100101",
  48215=>"000000101",
  48216=>"010011010",
  48217=>"000000101",
  48218=>"000001101",
  48219=>"100111100",
  48220=>"000000000",
  48221=>"111111111",
  48222=>"000001000",
  48223=>"111011011",
  48224=>"111011010",
  48225=>"111110100",
  48226=>"011010010",
  48227=>"101101101",
  48228=>"101101001",
  48229=>"110111010",
  48230=>"010011101",
  48231=>"110010010",
  48232=>"111111111",
  48233=>"000101101",
  48234=>"010011011",
  48235=>"000000000",
  48236=>"110110111",
  48237=>"101101001",
  48238=>"110111011",
  48239=>"101101101",
  48240=>"111111111",
  48241=>"001111101",
  48242=>"101001101",
  48243=>"111011010",
  48244=>"000000000",
  48245=>"010110110",
  48246=>"000000000",
  48247=>"001000000",
  48248=>"110101111",
  48249=>"111111111",
  48250=>"000000001",
  48251=>"011001011",
  48252=>"100100100",
  48253=>"000000100",
  48254=>"101101000",
  48255=>"000000101",
  48256=>"000110111",
  48257=>"000000101",
  48258=>"000000111",
  48259=>"100100100",
  48260=>"111111011",
  48261=>"011111000",
  48262=>"010000110",
  48263=>"011000000",
  48264=>"111000010",
  48265=>"000000000",
  48266=>"001001111",
  48267=>"001001001",
  48268=>"111111101",
  48269=>"001001000",
  48270=>"101101101",
  48271=>"001101000",
  48272=>"001101101",
  48273=>"111101111",
  48274=>"100100101",
  48275=>"000110101",
  48276=>"000000111",
  48277=>"101100000",
  48278=>"111111101",
  48279=>"000000000",
  48280=>"101101000",
  48281=>"101101111",
  48282=>"111101100",
  48283=>"010000000",
  48284=>"001111111",
  48285=>"110110110",
  48286=>"000001011",
  48287=>"011111111",
  48288=>"001010001",
  48289=>"001011000",
  48290=>"000000000",
  48291=>"000000110",
  48292=>"000000000",
  48293=>"000000000",
  48294=>"011111111",
  48295=>"101001100",
  48296=>"000000101",
  48297=>"001111111",
  48298=>"000000000",
  48299=>"111101111",
  48300=>"010000100",
  48301=>"000010110",
  48302=>"001001101",
  48303=>"010010010",
  48304=>"000000000",
  48305=>"101101110",
  48306=>"111111011",
  48307=>"000100100",
  48308=>"111010000",
  48309=>"110010000",
  48310=>"101000000",
  48311=>"001000001",
  48312=>"001000100",
  48313=>"000100000",
  48314=>"100101101",
  48315=>"000011010",
  48316=>"111111111",
  48317=>"000000000",
  48318=>"011011001",
  48319=>"110110110",
  48320=>"100100111",
  48321=>"010011111",
  48322=>"010111110",
  48323=>"010011111",
  48324=>"111111100",
  48325=>"010010011",
  48326=>"010010010",
  48327=>"010010000",
  48328=>"011011011",
  48329=>"010110111",
  48330=>"001001010",
  48331=>"101101101",
  48332=>"011111101",
  48333=>"101001000",
  48334=>"100111100",
  48335=>"101001001",
  48336=>"100111110",
  48337=>"111110011",
  48338=>"110000010",
  48339=>"000000000",
  48340=>"100000000",
  48341=>"000010111",
  48342=>"111000010",
  48343=>"111000000",
  48344=>"000000110",
  48345=>"001000000",
  48346=>"010000000",
  48347=>"000000001",
  48348=>"111110010",
  48349=>"000001011",
  48350=>"100001000",
  48351=>"000000001",
  48352=>"111111101",
  48353=>"111111010",
  48354=>"011011011",
  48355=>"000100111",
  48356=>"111111111",
  48357=>"101100001",
  48358=>"000100101",
  48359=>"101111101",
  48360=>"000000001",
  48361=>"010010010",
  48362=>"011111111",
  48363=>"111110100",
  48364=>"101111111",
  48365=>"000000000",
  48366=>"101111111",
  48367=>"111010010",
  48368=>"011000001",
  48369=>"000111111",
  48370=>"000111111",
  48371=>"101000111",
  48372=>"000000000",
  48373=>"111111110",
  48374=>"001001101",
  48375=>"000001101",
  48376=>"011111111",
  48377=>"000000000",
  48378=>"111111111",
  48379=>"111100100",
  48380=>"100110110",
  48381=>"110010110",
  48382=>"010110111",
  48383=>"101111101",
  48384=>"000001101",
  48385=>"100000101",
  48386=>"010010010",
  48387=>"111111111",
  48388=>"000101111",
  48389=>"101101000",
  48390=>"110110010",
  48391=>"000000010",
  48392=>"010000010",
  48393=>"101101001",
  48394=>"001101111",
  48395=>"000000000",
  48396=>"111101111",
  48397=>"101001000",
  48398=>"011011111",
  48399=>"110111111",
  48400=>"110110010",
  48401=>"001000111",
  48402=>"111001101",
  48403=>"111101100",
  48404=>"111111011",
  48405=>"101111111",
  48406=>"111111101",
  48407=>"110110110",
  48408=>"010000100",
  48409=>"000000000",
  48410=>"000111111",
  48411=>"000011011",
  48412=>"110111101",
  48413=>"110101101",
  48414=>"000001001",
  48415=>"101001010",
  48416=>"001001000",
  48417=>"100100101",
  48418=>"001010111",
  48419=>"111001100",
  48420=>"000000010",
  48421=>"010000100",
  48422=>"111100110",
  48423=>"010010010",
  48424=>"111111110",
  48425=>"001001001",
  48426=>"101101001",
  48427=>"111100000",
  48428=>"101101100",
  48429=>"000000100",
  48430=>"000000110",
  48431=>"100100101",
  48432=>"100100100",
  48433=>"010000000",
  48434=>"001111000",
  48435=>"101010000",
  48436=>"111101000",
  48437=>"000000001",
  48438=>"000000000",
  48439=>"000000000",
  48440=>"111111101",
  48441=>"101111101",
  48442=>"000101111",
  48443=>"000000001",
  48444=>"000000000",
  48445=>"001101001",
  48446=>"110010011",
  48447=>"000101111",
  48448=>"100111111",
  48449=>"111111111",
  48450=>"110000000",
  48451=>"100101101",
  48452=>"011111111",
  48453=>"000111111",
  48454=>"100101001",
  48455=>"111110111",
  48456=>"000000000",
  48457=>"010000010",
  48458=>"001000000",
  48459=>"011011011",
  48460=>"000000000",
  48461=>"000000110",
  48462=>"000000000",
  48463=>"100000100",
  48464=>"001011001",
  48465=>"011011010",
  48466=>"000100111",
  48467=>"100100111",
  48468=>"110111111",
  48469=>"001001001",
  48470=>"000000000",
  48471=>"111111111",
  48472=>"010010010",
  48473=>"111001000",
  48474=>"100110110",
  48475=>"010110010",
  48476=>"100111111",
  48477=>"101101101",
  48478=>"101000001",
  48479=>"000000000",
  48480=>"001001001",
  48481=>"111111111",
  48482=>"000110100",
  48483=>"011011010",
  48484=>"110110110",
  48485=>"000000000",
  48486=>"000000000",
  48487=>"111111111",
  48488=>"110110110",
  48489=>"110111111",
  48490=>"100000000",
  48491=>"111000101",
  48492=>"000000000",
  48493=>"000101101",
  48494=>"111001001",
  48495=>"000000111",
  48496=>"001000000",
  48497=>"000001101",
  48498=>"101101011",
  48499=>"100100100",
  48500=>"000001000",
  48501=>"001001001",
  48502=>"100000111",
  48503=>"000000010",
  48504=>"101101100",
  48505=>"111011011",
  48506=>"100101111",
  48507=>"110110000",
  48508=>"000110010",
  48509=>"010010011",
  48510=>"010010010",
  48511=>"000000001",
  48512=>"010011011",
  48513=>"010010010",
  48514=>"000100100",
  48515=>"010000000",
  48516=>"111111110",
  48517=>"010010010",
  48518=>"001101000",
  48519=>"111111011",
  48520=>"001001000",
  48521=>"000000011",
  48522=>"001000000",
  48523=>"010010000",
  48524=>"100101000",
  48525=>"101100000",
  48526=>"000000000",
  48527=>"000000001",
  48528=>"011000000",
  48529=>"100000000",
  48530=>"000001101",
  48531=>"000000100",
  48532=>"000110010",
  48533=>"000010000",
  48534=>"010000000",
  48535=>"110111110",
  48536=>"011011010",
  48537=>"010010010",
  48538=>"000000000",
  48539=>"001011111",
  48540=>"100000111",
  48541=>"110110000",
  48542=>"100100001",
  48543=>"100101000",
  48544=>"110111100",
  48545=>"001001001",
  48546=>"000011011",
  48547=>"011010111",
  48548=>"000010000",
  48549=>"111111111",
  48550=>"111111011",
  48551=>"111111000",
  48552=>"000000001",
  48553=>"001000110",
  48554=>"000000101",
  48555=>"000000101",
  48556=>"000000000",
  48557=>"101101101",
  48558=>"010110111",
  48559=>"010010011",
  48560=>"010010010",
  48561=>"111111111",
  48562=>"111111100",
  48563=>"000100100",
  48564=>"111111100",
  48565=>"111011111",
  48566=>"000000001",
  48567=>"111111101",
  48568=>"000001101",
  48569=>"010111111",
  48570=>"000000010",
  48571=>"100101101",
  48572=>"100100100",
  48573=>"101011001",
  48574=>"101101100",
  48575=>"111010000",
  48576=>"001111111",
  48577=>"100100101",
  48578=>"101011001",
  48579=>"100100100",
  48580=>"110111100",
  48581=>"100101101",
  48582=>"111110110",
  48583=>"100000101",
  48584=>"010000000",
  48585=>"011001111",
  48586=>"000000000",
  48587=>"011000000",
  48588=>"100110000",
  48589=>"010000010",
  48590=>"000000000",
  48591=>"011111111",
  48592=>"111011000",
  48593=>"100000000",
  48594=>"111110110",
  48595=>"001000111",
  48596=>"101111001",
  48597=>"111111100",
  48598=>"001001101",
  48599=>"000000100",
  48600=>"000000001",
  48601=>"111011111",
  48602=>"111010011",
  48603=>"110110110",
  48604=>"000000000",
  48605=>"000111111",
  48606=>"011011011",
  48607=>"000010110",
  48608=>"101101111",
  48609=>"010010111",
  48610=>"110110010",
  48611=>"001000100",
  48612=>"010010111",
  48613=>"111111111",
  48614=>"101000101",
  48615=>"000000000",
  48616=>"001000101",
  48617=>"110111011",
  48618=>"111111111",
  48619=>"001001001",
  48620=>"010010010",
  48621=>"000100000",
  48622=>"111000110",
  48623=>"001000001",
  48624=>"000000001",
  48625=>"011011001",
  48626=>"111000000",
  48627=>"111111101",
  48628=>"010111111",
  48629=>"000000010",
  48630=>"000011010",
  48631=>"110110010",
  48632=>"001101001",
  48633=>"101100101",
  48634=>"011111111",
  48635=>"100100100",
  48636=>"001011000",
  48637=>"010010110",
  48638=>"011001110",
  48639=>"111111101",
  48640=>"111001000",
  48641=>"111000000",
  48642=>"000001111",
  48643=>"010110010",
  48644=>"100110111",
  48645=>"111000000",
  48646=>"000000111",
  48647=>"111111111",
  48648=>"111111111",
  48649=>"000111111",
  48650=>"111111100",
  48651=>"000001001",
  48652=>"111011011",
  48653=>"100100111",
  48654=>"001111111",
  48655=>"000000000",
  48656=>"111011111",
  48657=>"000000111",
  48658=>"001011111",
  48659=>"100100111",
  48660=>"000000000",
  48661=>"111000001",
  48662=>"111111000",
  48663=>"111111111",
  48664=>"000000001",
  48665=>"101000001",
  48666=>"011000000",
  48667=>"000000000",
  48668=>"111111111",
  48669=>"111111000",
  48670=>"110111111",
  48671=>"100000111",
  48672=>"000000000",
  48673=>"111100111",
  48674=>"111111100",
  48675=>"001000000",
  48676=>"000111111",
  48677=>"111000100",
  48678=>"000000000",
  48679=>"110110000",
  48680=>"111000000",
  48681=>"000111111",
  48682=>"000010100",
  48683=>"111111111",
  48684=>"100001111",
  48685=>"000111010",
  48686=>"001111111",
  48687=>"111100111",
  48688=>"000000110",
  48689=>"100011111",
  48690=>"000100000",
  48691=>"000000001",
  48692=>"000101000",
  48693=>"111111011",
  48694=>"001001010",
  48695=>"000000111",
  48696=>"101111111",
  48697=>"101000000",
  48698=>"101100111",
  48699=>"000000000",
  48700=>"111111011",
  48701=>"000010111",
  48702=>"000000000",
  48703=>"000000111",
  48704=>"111000000",
  48705=>"000000000",
  48706=>"111111100",
  48707=>"100000000",
  48708=>"110111111",
  48709=>"111011000",
  48710=>"111001000",
  48711=>"000000000",
  48712=>"100100100",
  48713=>"000000101",
  48714=>"111111111",
  48715=>"111111000",
  48716=>"100100100",
  48717=>"111000000",
  48718=>"000000111",
  48719=>"111100000",
  48720=>"111000000",
  48721=>"111100000",
  48722=>"111001001",
  48723=>"000100100",
  48724=>"011000000",
  48725=>"000101111",
  48726=>"001000000",
  48727=>"110111000",
  48728=>"000111111",
  48729=>"101000101",
  48730=>"011111111",
  48731=>"110001000",
  48732=>"000111111",
  48733=>"000000000",
  48734=>"000111111",
  48735=>"111110000",
  48736=>"000000000",
  48737=>"101100111",
  48738=>"000100000",
  48739=>"110000111",
  48740=>"100101001",
  48741=>"111110100",
  48742=>"111110010",
  48743=>"000111100",
  48744=>"011111111",
  48745=>"111100111",
  48746=>"101000101",
  48747=>"000001111",
  48748=>"010000101",
  48749=>"000111110",
  48750=>"000111111",
  48751=>"000000011",
  48752=>"001000100",
  48753=>"100000000",
  48754=>"000101111",
  48755=>"000000001",
  48756=>"000000111",
  48757=>"000111111",
  48758=>"000000100",
  48759=>"000000000",
  48760=>"100100000",
  48761=>"101111011",
  48762=>"000111000",
  48763=>"111000000",
  48764=>"110110110",
  48765=>"000000000",
  48766=>"000111111",
  48767=>"000000000",
  48768=>"001001011",
  48769=>"001011011",
  48770=>"111000000",
  48771=>"000000100",
  48772=>"111111111",
  48773=>"000000001",
  48774=>"111111101",
  48775=>"111111111",
  48776=>"001111111",
  48777=>"000000001",
  48778=>"000000111",
  48779=>"111111111",
  48780=>"110111101",
  48781=>"000000000",
  48782=>"100000001",
  48783=>"110111110",
  48784=>"111000111",
  48785=>"000000000",
  48786=>"111000000",
  48787=>"011111111",
  48788=>"000001000",
  48789=>"110111100",
  48790=>"111000000",
  48791=>"101000000",
  48792=>"000000000",
  48793=>"111110100",
  48794=>"100111111",
  48795=>"000000001",
  48796=>"111111111",
  48797=>"111000000",
  48798=>"111111111",
  48799=>"000000000",
  48800=>"100000010",
  48801=>"000000101",
  48802=>"000000011",
  48803=>"110100100",
  48804=>"000011001",
  48805=>"111000000",
  48806=>"010110011",
  48807=>"111111011",
  48808=>"101001001",
  48809=>"000001111",
  48810=>"000000000",
  48811=>"000000111",
  48812=>"011000000",
  48813=>"100100101",
  48814=>"111111111",
  48815=>"111000000",
  48816=>"000000000",
  48817=>"000000000",
  48818=>"000110110",
  48819=>"010000111",
  48820=>"000111111",
  48821=>"111011000",
  48822=>"000000000",
  48823=>"111111111",
  48824=>"111000000",
  48825=>"000011111",
  48826=>"000000000",
  48827=>"000000000",
  48828=>"111000100",
  48829=>"111111111",
  48830=>"111111101",
  48831=>"000110110",
  48832=>"111111000",
  48833=>"100000000",
  48834=>"011000000",
  48835=>"000110110",
  48836=>"110111111",
  48837=>"111000000",
  48838=>"000000001",
  48839=>"101000000",
  48840=>"000111111",
  48841=>"111000000",
  48842=>"111100100",
  48843=>"000010011",
  48844=>"111000000",
  48845=>"110110000",
  48846=>"111000000",
  48847=>"111011000",
  48848=>"000000000",
  48849=>"110110111",
  48850=>"000000100",
  48851=>"110000000",
  48852=>"111111001",
  48853=>"001000111",
  48854=>"000011000",
  48855=>"010000100",
  48856=>"000111111",
  48857=>"000000011",
  48858=>"111111100",
  48859=>"111111111",
  48860=>"000000111",
  48861=>"001111000",
  48862=>"000111111",
  48863=>"111111100",
  48864=>"000000000",
  48865=>"000000000",
  48866=>"111111000",
  48867=>"101001000",
  48868=>"111111101",
  48869=>"110111111",
  48870=>"111110001",
  48871=>"100111111",
  48872=>"001000101",
  48873=>"111000000",
  48874=>"001111100",
  48875=>"100000111",
  48876=>"111000000",
  48877=>"111000000",
  48878=>"000000111",
  48879=>"110000010",
  48880=>"110110110",
  48881=>"001000111",
  48882=>"000001111",
  48883=>"001000000",
  48884=>"111111111",
  48885=>"001111000",
  48886=>"010111000",
  48887=>"111000000",
  48888=>"000000000",
  48889=>"000000000",
  48890=>"000000000",
  48891=>"000101001",
  48892=>"000111011",
  48893=>"100100001",
  48894=>"111000000",
  48895=>"010000000",
  48896=>"111000000",
  48897=>"111000000",
  48898=>"000000000",
  48899=>"000000000",
  48900=>"100000000",
  48901=>"000000111",
  48902=>"000111110",
  48903=>"000010111",
  48904=>"111111111",
  48905=>"000101111",
  48906=>"111100100",
  48907=>"111111110",
  48908=>"110000110",
  48909=>"000000000",
  48910=>"111111111",
  48911=>"111011000",
  48912=>"111101000",
  48913=>"100000000",
  48914=>"111111000",
  48915=>"111000000",
  48916=>"000000111",
  48917=>"111010000",
  48918=>"111111111",
  48919=>"100000111",
  48920=>"000000111",
  48921=>"111111000",
  48922=>"001111110",
  48923=>"000000000",
  48924=>"100100001",
  48925=>"010000111",
  48926=>"111000000",
  48927=>"111111110",
  48928=>"111000000",
  48929=>"111000000",
  48930=>"001000011",
  48931=>"000111111",
  48932=>"010000100",
  48933=>"111010111",
  48934=>"110111000",
  48935=>"111011100",
  48936=>"100100111",
  48937=>"000000110",
  48938=>"111111100",
  48939=>"111111100",
  48940=>"111100101",
  48941=>"110111111",
  48942=>"000000111",
  48943=>"000101000",
  48944=>"000000000",
  48945=>"111111011",
  48946=>"111101111",
  48947=>"100000101",
  48948=>"111100000",
  48949=>"111011011",
  48950=>"000000110",
  48951=>"111011001",
  48952=>"000001000",
  48953=>"111001111",
  48954=>"110100000",
  48955=>"111000000",
  48956=>"111011111",
  48957=>"001100100",
  48958=>"000000111",
  48959=>"100000000",
  48960=>"000111111",
  48961=>"000000001",
  48962=>"001011111",
  48963=>"000100000",
  48964=>"100000000",
  48965=>"000000111",
  48966=>"000011001",
  48967=>"000000111",
  48968=>"110110000",
  48969=>"000111111",
  48970=>"111000000",
  48971=>"000000111",
  48972=>"111111111",
  48973=>"111111011",
  48974=>"111111111",
  48975=>"111001000",
  48976=>"111111000",
  48977=>"111011000",
  48978=>"111010010",
  48979=>"100100000",
  48980=>"111110000",
  48981=>"001011011",
  48982=>"111111000",
  48983=>"000000001",
  48984=>"111111111",
  48985=>"111011010",
  48986=>"000111111",
  48987=>"000000101",
  48988=>"111111111",
  48989=>"111000100",
  48990=>"111110010",
  48991=>"100111001",
  48992=>"111000000",
  48993=>"001000001",
  48994=>"000111111",
  48995=>"111111111",
  48996=>"000101111",
  48997=>"111000101",
  48998=>"111111000",
  48999=>"100111110",
  49000=>"100111111",
  49001=>"111111001",
  49002=>"010000100",
  49003=>"100111101",
  49004=>"100111110",
  49005=>"111001111",
  49006=>"111111011",
  49007=>"000000000",
  49008=>"111011111",
  49009=>"011000000",
  49010=>"101100111",
  49011=>"000111111",
  49012=>"111111111",
  49013=>"000000110",
  49014=>"111111111",
  49015=>"111010000",
  49016=>"111000000",
  49017=>"000000111",
  49018=>"110111111",
  49019=>"111000111",
  49020=>"011011111",
  49021=>"000100001",
  49022=>"111011000",
  49023=>"110000111",
  49024=>"000001011",
  49025=>"000111111",
  49026=>"111111001",
  49027=>"000000000",
  49028=>"011000000",
  49029=>"000000000",
  49030=>"010011111",
  49031=>"000000111",
  49032=>"000000001",
  49033=>"111111000",
  49034=>"111111000",
  49035=>"111111001",
  49036=>"101000100",
  49037=>"011011111",
  49038=>"111111111",
  49039=>"001111111",
  49040=>"000000000",
  49041=>"111101111",
  49042=>"111111000",
  49043=>"111111111",
  49044=>"111111111",
  49045=>"000000000",
  49046=>"000000100",
  49047=>"000000111",
  49048=>"000010111",
  49049=>"000001000",
  49050=>"000000001",
  49051=>"111001000",
  49052=>"000000111",
  49053=>"010100111",
  49054=>"000000100",
  49055=>"000000001",
  49056=>"000001111",
  49057=>"100110010",
  49058=>"100110001",
  49059=>"111111111",
  49060=>"111111000",
  49061=>"000111110",
  49062=>"000000000",
  49063=>"111000000",
  49064=>"000000000",
  49065=>"111000000",
  49066=>"111000000",
  49067=>"000000000",
  49068=>"111110000",
  49069=>"000100011",
  49070=>"111100000",
  49071=>"000000011",
  49072=>"111011100",
  49073=>"000000111",
  49074=>"111111000",
  49075=>"000111000",
  49076=>"000100111",
  49077=>"100110000",
  49078=>"100100111",
  49079=>"111000111",
  49080=>"111000000",
  49081=>"111000000",
  49082=>"000000001",
  49083=>"101111111",
  49084=>"111101001",
  49085=>"000001111",
  49086=>"000000100",
  49087=>"111100000",
  49088=>"000000100",
  49089=>"111111000",
  49090=>"110000111",
  49091=>"000000111",
  49092=>"000000000",
  49093=>"111111111",
  49094=>"000110100",
  49095=>"111111110",
  49096=>"001000111",
  49097=>"111111111",
  49098=>"000000000",
  49099=>"111111111",
  49100=>"111000000",
  49101=>"001000000",
  49102=>"111111111",
  49103=>"111111111",
  49104=>"000000111",
  49105=>"000111111",
  49106=>"110110111",
  49107=>"111111010",
  49108=>"111011000",
  49109=>"000000001",
  49110=>"100000000",
  49111=>"000000100",
  49112=>"101000101",
  49113=>"111111100",
  49114=>"111000000",
  49115=>"001000001",
  49116=>"010010000",
  49117=>"111010000",
  49118=>"011001000",
  49119=>"111100000",
  49120=>"110100111",
  49121=>"111111110",
  49122=>"111100111",
  49123=>"001110111",
  49124=>"111111111",
  49125=>"111111000",
  49126=>"100110111",
  49127=>"001000111",
  49128=>"111111101",
  49129=>"111000000",
  49130=>"001000000",
  49131=>"100101000",
  49132=>"111111111",
  49133=>"000000000",
  49134=>"000111111",
  49135=>"000111111",
  49136=>"000000001",
  49137=>"110111111",
  49138=>"100100100",
  49139=>"000000000",
  49140=>"111111100",
  49141=>"111011111",
  49142=>"111111000",
  49143=>"100100001",
  49144=>"010111111",
  49145=>"100111100",
  49146=>"000000000",
  49147=>"111000000",
  49148=>"100100111",
  49149=>"101111111",
  49150=>"000000000",
  49151=>"000000111",
  49152=>"100000010",
  49153=>"101000000",
  49154=>"001000111",
  49155=>"000001001",
  49156=>"110110110",
  49157=>"001000000",
  49158=>"110110111",
  49159=>"111111111",
  49160=>"111100100",
  49161=>"000000111",
  49162=>"111101100",
  49163=>"100111101",
  49164=>"100110110",
  49165=>"000000000",
  49166=>"011001011",
  49167=>"110111111",
  49168=>"110110000",
  49169=>"011010101",
  49170=>"010000000",
  49171=>"010000000",
  49172=>"000000000",
  49173=>"100101111",
  49174=>"000101111",
  49175=>"111111100",
  49176=>"100000000",
  49177=>"110110110",
  49178=>"111111111",
  49179=>"110111111",
  49180=>"001001001",
  49181=>"001101000",
  49182=>"101101101",
  49183=>"101000000",
  49184=>"111110111",
  49185=>"111111011",
  49186=>"110110110",
  49187=>"000000000",
  49188=>"111111000",
  49189=>"000001001",
  49190=>"000000000",
  49191=>"100111111",
  49192=>"000000111",
  49193=>"100100000",
  49194=>"000100111",
  49195=>"000000000",
  49196=>"000000000",
  49197=>"000100111",
  49198=>"111001000",
  49199=>"000000000",
  49200=>"000001001",
  49201=>"100100100",
  49202=>"011011001",
  49203=>"000010001",
  49204=>"101101101",
  49205=>"110010100",
  49206=>"011001000",
  49207=>"000111010",
  49208=>"111111000",
  49209=>"000000000",
  49210=>"010011111",
  49211=>"101000000",
  49212=>"000000000",
  49213=>"010111011",
  49214=>"100000000",
  49215=>"000000000",
  49216=>"000000000",
  49217=>"100101101",
  49218=>"111010010",
  49219=>"111111111",
  49220=>"110110110",
  49221=>"111111110",
  49222=>"111000111",
  49223=>"111111101",
  49224=>"011011011",
  49225=>"000000000",
  49226=>"110100100",
  49227=>"111110000",
  49228=>"111100100",
  49229=>"000000000",
  49230=>"000000111",
  49231=>"000100100",
  49232=>"000010111",
  49233=>"000000000",
  49234=>"111111001",
  49235=>"010000001",
  49236=>"000001001",
  49237=>"100100100",
  49238=>"011000110",
  49239=>"111111000",
  49240=>"000000000",
  49241=>"101101111",
  49242=>"000001111",
  49243=>"110100000",
  49244=>"110000000",
  49245=>"001000000",
  49246=>"000000110",
  49247=>"000000000",
  49248=>"000000000",
  49249=>"001111111",
  49250=>"110111111",
  49251=>"111101101",
  49252=>"111110010",
  49253=>"111001001",
  49254=>"000001111",
  49255=>"111101000",
  49256=>"001001000",
  49257=>"000000101",
  49258=>"000000000",
  49259=>"000000111",
  49260=>"110110000",
  49261=>"111111110",
  49262=>"000000101",
  49263=>"011010011",
  49264=>"111111111",
  49265=>"011000001",
  49266=>"001001001",
  49267=>"001001110",
  49268=>"100100000",
  49269=>"110110110",
  49270=>"000000101",
  49271=>"111011000",
  49272=>"110000000",
  49273=>"110110111",
  49274=>"111000000",
  49275=>"011011000",
  49276=>"001000101",
  49277=>"000111111",
  49278=>"001110000",
  49279=>"011111111",
  49280=>"100000000",
  49281=>"001001000",
  49282=>"111101101",
  49283=>"010010011",
  49284=>"001001001",
  49285=>"000000000",
  49286=>"111100000",
  49287=>"101000000",
  49288=>"000000001",
  49289=>"011111111",
  49290=>"000000101",
  49291=>"011111100",
  49292=>"111111111",
  49293=>"111111100",
  49294=>"001100000",
  49295=>"110111110",
  49296=>"111101101",
  49297=>"101001001",
  49298=>"100111101",
  49299=>"101100100",
  49300=>"000000100",
  49301=>"111110000",
  49302=>"000000000",
  49303=>"000000001",
  49304=>"000000000",
  49305=>"010111111",
  49306=>"110110110",
  49307=>"101100101",
  49308=>"111111111",
  49309=>"111111111",
  49310=>"001000000",
  49311=>"010111010",
  49312=>"000100000",
  49313=>"001111111",
  49314=>"111111111",
  49315=>"111111110",
  49316=>"110010011",
  49317=>"111111111",
  49318=>"100101111",
  49319=>"100100111",
  49320=>"000010010",
  49321=>"111101101",
  49322=>"111001001",
  49323=>"100101101",
  49324=>"000111111",
  49325=>"000000111",
  49326=>"111111110",
  49327=>"001000000",
  49328=>"010000010",
  49329=>"111110001",
  49330=>"101111111",
  49331=>"001001111",
  49332=>"110100111",
  49333=>"000001100",
  49334=>"111011000",
  49335=>"111111111",
  49336=>"111111111",
  49337=>"111111110",
  49338=>"111111110",
  49339=>"110110110",
  49340=>"111111111",
  49341=>"000000100",
  49342=>"000000000",
  49343=>"110111110",
  49344=>"100000000",
  49345=>"110110110",
  49346=>"110110110",
  49347=>"101011000",
  49348=>"111000000",
  49349=>"000000001",
  49350=>"000000100",
  49351=>"111111001",
  49352=>"011111110",
  49353=>"110100111",
  49354=>"010111001",
  49355=>"000000000",
  49356=>"101111111",
  49357=>"100001000",
  49358=>"010001001",
  49359=>"111010110",
  49360=>"111111111",
  49361=>"111101111",
  49362=>"111000001",
  49363=>"110110110",
  49364=>"000000000",
  49365=>"111111000",
  49366=>"001000000",
  49367=>"110110100",
  49368=>"000000000",
  49369=>"111111110",
  49370=>"111111101",
  49371=>"100111011",
  49372=>"000000000",
  49373=>"011001000",
  49374=>"001000000",
  49375=>"000000110",
  49376=>"000000111",
  49377=>"001000100",
  49378=>"000000000",
  49379=>"010111010",
  49380=>"000000111",
  49381=>"000001001",
  49382=>"111111000",
  49383=>"111111111",
  49384=>"100111110",
  49385=>"110000001",
  49386=>"110110110",
  49387=>"111111111",
  49388=>"000000001",
  49389=>"000000000",
  49390=>"111101101",
  49391=>"111000011",
  49392=>"000010000",
  49393=>"110110110",
  49394=>"000000000",
  49395=>"111111101",
  49396=>"111111100",
  49397=>"000000000",
  49398=>"100100101",
  49399=>"111011011",
  49400=>"111011101",
  49401=>"101000000",
  49402=>"110110110",
  49403=>"111000000",
  49404=>"001000000",
  49405=>"110110100",
  49406=>"000101000",
  49407=>"110000000",
  49408=>"000000000",
  49409=>"000000100",
  49410=>"010111111",
  49411=>"101101100",
  49412=>"000000000",
  49413=>"000000111",
  49414=>"111111111",
  49415=>"110110111",
  49416=>"001000000",
  49417=>"000111111",
  49418=>"000000000",
  49419=>"111111011",
  49420=>"100000000",
  49421=>"000001000",
  49422=>"000000101",
  49423=>"010000000",
  49424=>"000100111",
  49425=>"011111111",
  49426=>"011011011",
  49427=>"001111111",
  49428=>"110110111",
  49429=>"111101001",
  49430=>"111110110",
  49431=>"100000000",
  49432=>"000100110",
  49433=>"111110000",
  49434=>"000000000",
  49435=>"000110010",
  49436=>"100110111",
  49437=>"100111111",
  49438=>"000000000",
  49439=>"111001000",
  49440=>"111111000",
  49441=>"000111010",
  49442=>"000111101",
  49443=>"000000111",
  49444=>"110001101",
  49445=>"000000101",
  49446=>"010011011",
  49447=>"111000000",
  49448=>"111100000",
  49449=>"111111010",
  49450=>"010111111",
  49451=>"000000111",
  49452=>"111010100",
  49453=>"111110110",
  49454=>"101000111",
  49455=>"000000100",
  49456=>"110110110",
  49457=>"000010010",
  49458=>"101111111",
  49459=>"000100000",
  49460=>"111111111",
  49461=>"111100111",
  49462=>"111110101",
  49463=>"000000000",
  49464=>"011000000",
  49465=>"000000111",
  49466=>"000000000",
  49467=>"000001100",
  49468=>"100000000",
  49469=>"011111111",
  49470=>"100000100",
  49471=>"000000000",
  49472=>"111111111",
  49473=>"000001001",
  49474=>"110111110",
  49475=>"000000001",
  49476=>"001001001",
  49477=>"000000100",
  49478=>"111111110",
  49479=>"000000000",
  49480=>"101001000",
  49481=>"100000001",
  49482=>"000100110",
  49483=>"110010000",
  49484=>"000000111",
  49485=>"000011111",
  49486=>"111000000",
  49487=>"000011111",
  49488=>"010010011",
  49489=>"000000100",
  49490=>"111111110",
  49491=>"110100000",
  49492=>"001011011",
  49493=>"111011001",
  49494=>"110111111",
  49495=>"101101101",
  49496=>"000000000",
  49497=>"001000001",
  49498=>"011111111",
  49499=>"000000000",
  49500=>"010100000",
  49501=>"001001110",
  49502=>"000000111",
  49503=>"011000000",
  49504=>"101111111",
  49505=>"111001001",
  49506=>"111111101",
  49507=>"101101001",
  49508=>"111111001",
  49509=>"111100000",
  49510=>"111111111",
  49511=>"110010000",
  49512=>"001001001",
  49513=>"111100000",
  49514=>"100000000",
  49515=>"110100111",
  49516=>"110110110",
  49517=>"000011111",
  49518=>"110111111",
  49519=>"111100101",
  49520=>"000000111",
  49521=>"101101101",
  49522=>"101000000",
  49523=>"111111000",
  49524=>"100100000",
  49525=>"110110000",
  49526=>"111100001",
  49527=>"111111001",
  49528=>"101000000",
  49529=>"111101101",
  49530=>"001001111",
  49531=>"000000000",
  49532=>"111100000",
  49533=>"000000111",
  49534=>"010111011",
  49535=>"111101111",
  49536=>"000000001",
  49537=>"111111100",
  49538=>"110111111",
  49539=>"100000000",
  49540=>"001001111",
  49541=>"000000101",
  49542=>"100100111",
  49543=>"111101101",
  49544=>"001000111",
  49545=>"100110000",
  49546=>"101000000",
  49547=>"000000000",
  49548=>"000011111",
  49549=>"010010010",
  49550=>"011001000",
  49551=>"000000000",
  49552=>"101000000",
  49553=>"010000000",
  49554=>"011111000",
  49555=>"001000111",
  49556=>"111111111",
  49557=>"110110010",
  49558=>"100010000",
  49559=>"010011111",
  49560=>"000000011",
  49561=>"110110111",
  49562=>"101101101",
  49563=>"000000000",
  49564=>"000000000",
  49565=>"011010011",
  49566=>"100111111",
  49567=>"110110000",
  49568=>"111111110",
  49569=>"011001001",
  49570=>"011000000",
  49571=>"111111111",
  49572=>"000000000",
  49573=>"110100111",
  49574=>"101000101",
  49575=>"001000000",
  49576=>"111101001",
  49577=>"110000000",
  49578=>"000001001",
  49579=>"000000111",
  49580=>"111100000",
  49581=>"101101000",
  49582=>"000000000",
  49583=>"111101100",
  49584=>"111111111",
  49585=>"100000000",
  49586=>"000000000",
  49587=>"000000000",
  49588=>"111111111",
  49589=>"001011001",
  49590=>"010010000",
  49591=>"111110010",
  49592=>"000101101",
  49593=>"110111111",
  49594=>"011101100",
  49595=>"000001000",
  49596=>"111001000",
  49597=>"111111110",
  49598=>"111111010",
  49599=>"001010010",
  49600=>"000010111",
  49601=>"001001111",
  49602=>"000000001",
  49603=>"001000111",
  49604=>"111110110",
  49605=>"000001100",
  49606=>"001100100",
  49607=>"000000000",
  49608=>"001000000",
  49609=>"001000001",
  49610=>"011110110",
  49611=>"000111111",
  49612=>"011000001",
  49613=>"111111011",
  49614=>"101101001",
  49615=>"100100000",
  49616=>"111111111",
  49617=>"000000011",
  49618=>"000000100",
  49619=>"111001001",
  49620=>"000000000",
  49621=>"011111000",
  49622=>"011010000",
  49623=>"011011011",
  49624=>"000000000",
  49625=>"110000000",
  49626=>"111001111",
  49627=>"111111111",
  49628=>"100001111",
  49629=>"111110111",
  49630=>"111001111",
  49631=>"001101100",
  49632=>"101001001",
  49633=>"001000000",
  49634=>"111111111",
  49635=>"000000000",
  49636=>"101001010",
  49637=>"100110000",
  49638=>"000000111",
  49639=>"000000000",
  49640=>"010000000",
  49641=>"000010010",
  49642=>"100100000",
  49643=>"111011011",
  49644=>"100000010",
  49645=>"110110110",
  49646=>"111111111",
  49647=>"000000100",
  49648=>"001001111",
  49649=>"000010010",
  49650=>"111111110",
  49651=>"111111111",
  49652=>"000000100",
  49653=>"000000000",
  49654=>"110110000",
  49655=>"000000100",
  49656=>"011000000",
  49657=>"100010000",
  49658=>"110000000",
  49659=>"110101101",
  49660=>"001000100",
  49661=>"000000111",
  49662=>"001000000",
  49663=>"111111111",
  49664=>"001111110",
  49665=>"110000000",
  49666=>"000011010",
  49667=>"100000000",
  49668=>"000000100",
  49669=>"100110011",
  49670=>"111111000",
  49671=>"000111111",
  49672=>"100111100",
  49673=>"101100000",
  49674=>"111000000",
  49675=>"111111000",
  49676=>"111011011",
  49677=>"111000000",
  49678=>"000000000",
  49679=>"000111111",
  49680=>"001001001",
  49681=>"111111111",
  49682=>"111111100",
  49683=>"000111111",
  49684=>"000000110",
  49685=>"011110111",
  49686=>"000000111",
  49687=>"000000001",
  49688=>"000000000",
  49689=>"011011011",
  49690=>"000000000",
  49691=>"010000001",
  49692=>"000000000",
  49693=>"000001011",
  49694=>"000011011",
  49695=>"001000000",
  49696=>"000111111",
  49697=>"010000001",
  49698=>"111111011",
  49699=>"000101111",
  49700=>"000000011",
  49701=>"001001000",
  49702=>"000110111",
  49703=>"100111101",
  49704=>"000101111",
  49705=>"000000111",
  49706=>"000000000",
  49707=>"000000111",
  49708=>"100001011",
  49709=>"000111111",
  49710=>"110100110",
  49711=>"111101110",
  49712=>"110000011",
  49713=>"111000000",
  49714=>"000000011",
  49715=>"000010000",
  49716=>"000001011",
  49717=>"100000011",
  49718=>"011001001",
  49719=>"000100000",
  49720=>"011111000",
  49721=>"000000000",
  49722=>"111000000",
  49723=>"000000010",
  49724=>"111000111",
  49725=>"000111111",
  49726=>"011101111",
  49727=>"111111000",
  49728=>"111111011",
  49729=>"000000000",
  49730=>"000111000",
  49731=>"111111111",
  49732=>"111001011",
  49733=>"000000100",
  49734=>"111000000",
  49735=>"111111111",
  49736=>"111010110",
  49737=>"000000000",
  49738=>"111111000",
  49739=>"111011111",
  49740=>"110100000",
  49741=>"111000000",
  49742=>"111000000",
  49743=>"101000000",
  49744=>"111111111",
  49745=>"000000111",
  49746=>"000000000",
  49747=>"000110000",
  49748=>"111111111",
  49749=>"000000000",
  49750=>"111000000",
  49751=>"111111110",
  49752=>"011011000",
  49753=>"111001000",
  49754=>"101111111",
  49755=>"110110110",
  49756=>"111111001",
  49757=>"000100111",
  49758=>"001100111",
  49759=>"000010011",
  49760=>"000000000",
  49761=>"000111111",
  49762=>"000000110",
  49763=>"010000100",
  49764=>"000000000",
  49765=>"110010000",
  49766=>"111111111",
  49767=>"111111100",
  49768=>"000000000",
  49769=>"111000000",
  49770=>"100100111",
  49771=>"111111000",
  49772=>"000111111",
  49773=>"111111111",
  49774=>"000000000",
  49775=>"000111111",
  49776=>"111001000",
  49777=>"010110100",
  49778=>"001000000",
  49779=>"000111111",
  49780=>"111111111",
  49781=>"000001111",
  49782=>"000000000",
  49783=>"000000111",
  49784=>"110000010",
  49785=>"111111000",
  49786=>"011001011",
  49787=>"000000000",
  49788=>"011011111",
  49789=>"000011000",
  49790=>"001000000",
  49791=>"011001000",
  49792=>"000000110",
  49793=>"111110110",
  49794=>"111111111",
  49795=>"010010000",
  49796=>"111100110",
  49797=>"000000000",
  49798=>"110100000",
  49799=>"111111010",
  49800=>"101000011",
  49801=>"111000000",
  49802=>"000000000",
  49803=>"111100000",
  49804=>"000011011",
  49805=>"100000111",
  49806=>"000000000",
  49807=>"111100111",
  49808=>"000111111",
  49809=>"111011111",
  49810=>"101111111",
  49811=>"111111000",
  49812=>"000000000",
  49813=>"111111110",
  49814=>"111111000",
  49815=>"111111000",
  49816=>"000000000",
  49817=>"111101111",
  49818=>"000000000",
  49819=>"000010011",
  49820=>"100111111",
  49821=>"000111111",
  49822=>"000000000",
  49823=>"000100000",
  49824=>"111000000",
  49825=>"111111110",
  49826=>"001000000",
  49827=>"111100000",
  49828=>"110100100",
  49829=>"111111000",
  49830=>"000000011",
  49831=>"011011111",
  49832=>"011111000",
  49833=>"111110110",
  49834=>"111111111",
  49835=>"111111111",
  49836=>"000000011",
  49837=>"101101110",
  49838=>"111111011",
  49839=>"100000111",
  49840=>"000000001",
  49841=>"100111111",
  49842=>"000010111",
  49843=>"011111000",
  49844=>"110111100",
  49845=>"111111011",
  49846=>"000000111",
  49847=>"011111111",
  49848=>"000000001",
  49849=>"000110111",
  49850=>"111000101",
  49851=>"000111011",
  49852=>"000000111",
  49853=>"100111111",
  49854=>"000101011",
  49855=>"001001001",
  49856=>"000001111",
  49857=>"000000000",
  49858=>"000000000",
  49859=>"000000001",
  49860=>"000000011",
  49861=>"000111011",
  49862=>"000000000",
  49863=>"111111010",
  49864=>"000000100",
  49865=>"000000000",
  49866=>"000010111",
  49867=>"111111101",
  49868=>"101000000",
  49869=>"000000000",
  49870=>"001001000",
  49871=>"100000000",
  49872=>"000000100",
  49873=>"010000000",
  49874=>"000001001",
  49875=>"000000000",
  49876=>"110000000",
  49877=>"110111001",
  49878=>"000111111",
  49879=>"110110111",
  49880=>"000010111",
  49881=>"000111111",
  49882=>"000000111",
  49883=>"001001000",
  49884=>"111000111",
  49885=>"111000000",
  49886=>"010111111",
  49887=>"100000001",
  49888=>"111000000",
  49889=>"000000110",
  49890=>"000101110",
  49891=>"111101000",
  49892=>"010011000",
  49893=>"011011011",
  49894=>"001001111",
  49895=>"111000000",
  49896=>"000001001",
  49897=>"000111111",
  49898=>"111111011",
  49899=>"011000000",
  49900=>"000111111",
  49901=>"010111111",
  49902=>"000110111",
  49903=>"111111111",
  49904=>"100010000",
  49905=>"111111111",
  49906=>"000111111",
  49907=>"111000100",
  49908=>"000101100",
  49909=>"000000111",
  49910=>"000000110",
  49911=>"000111111",
  49912=>"000011111",
  49913=>"000100110",
  49914=>"000000100",
  49915=>"000000000",
  49916=>"000001001",
  49917=>"000110111",
  49918=>"111111111",
  49919=>"111111101",
  49920=>"000111000",
  49921=>"000000010",
  49922=>"110000000",
  49923=>"100111111",
  49924=>"001011111",
  49925=>"110010000",
  49926=>"101001111",
  49927=>"001111110",
  49928=>"111100000",
  49929=>"010110100",
  49930=>"111111001",
  49931=>"000000000",
  49932=>"000000000",
  49933=>"001001101",
  49934=>"100001111",
  49935=>"000000011",
  49936=>"000111111",
  49937=>"111000000",
  49938=>"100000000",
  49939=>"000000111",
  49940=>"000000000",
  49941=>"111111111",
  49942=>"000000001",
  49943=>"111111000",
  49944=>"000100111",
  49945=>"111011101",
  49946=>"100100110",
  49947=>"001111111",
  49948=>"011100011",
  49949=>"110000110",
  49950=>"111100000",
  49951=>"111111011",
  49952=>"101110111",
  49953=>"000000010",
  49954=>"111000001",
  49955=>"111111000",
  49956=>"110111011",
  49957=>"000011001",
  49958=>"110100110",
  49959=>"000010111",
  49960=>"011011000",
  49961=>"100101111",
  49962=>"110111111",
  49963=>"111111000",
  49964=>"111000101",
  49965=>"000111111",
  49966=>"111011000",
  49967=>"000000110",
  49968=>"100110111",
  49969=>"100111011",
  49970=>"110000000",
  49971=>"000001111",
  49972=>"010100111",
  49973=>"000100111",
  49974=>"110000000",
  49975=>"111111010",
  49976=>"011111000",
  49977=>"111111000",
  49978=>"000010000",
  49979=>"000110000",
  49980=>"100100100",
  49981=>"001001001",
  49982=>"110110110",
  49983=>"000000010",
  49984=>"000000011",
  49985=>"100110111",
  49986=>"000000000",
  49987=>"000010111",
  49988=>"000111000",
  49989=>"000110100",
  49990=>"111111111",
  49991=>"111000000",
  49992=>"000001111",
  49993=>"110000011",
  49994=>"100110000",
  49995=>"110110010",
  49996=>"001101111",
  49997=>"000111000",
  49998=>"000000111",
  49999=>"000110111",
  50000=>"000110110",
  50001=>"100111111",
  50002=>"000000111",
  50003=>"101000000",
  50004=>"000000000",
  50005=>"111100100",
  50006=>"100001111",
  50007=>"000000111",
  50008=>"111010101",
  50009=>"111001111",
  50010=>"111111111",
  50011=>"111111000",
  50012=>"000000110",
  50013=>"111111111",
  50014=>"110010010",
  50015=>"111111011",
  50016=>"100111111",
  50017=>"001111111",
  50018=>"000100110",
  50019=>"000000011",
  50020=>"111011001",
  50021=>"001111111",
  50022=>"100111111",
  50023=>"000000000",
  50024=>"011110000",
  50025=>"000000111",
  50026=>"100000110",
  50027=>"010011010",
  50028=>"111110100",
  50029=>"000000111",
  50030=>"001001111",
  50031=>"000110000",
  50032=>"111111010",
  50033=>"111101111",
  50034=>"000000001",
  50035=>"000001101",
  50036=>"000000000",
  50037=>"000000000",
  50038=>"101111000",
  50039=>"010000111",
  50040=>"111111111",
  50041=>"000000000",
  50042=>"110010001",
  50043=>"000000000",
  50044=>"111000000",
  50045=>"000000111",
  50046=>"100110100",
  50047=>"111110100",
  50048=>"100001111",
  50049=>"111111111",
  50050=>"100001111",
  50051=>"000110110",
  50052=>"111000000",
  50053=>"000000111",
  50054=>"000111111",
  50055=>"000011000",
  50056=>"000010110",
  50057=>"111010110",
  50058=>"111011000",
  50059=>"111010000",
  50060=>"111111111",
  50061=>"000000000",
  50062=>"111111111",
  50063=>"011010010",
  50064=>"000000101",
  50065=>"101001000",
  50066=>"100100111",
  50067=>"100000111",
  50068=>"111111000",
  50069=>"000000000",
  50070=>"000000111",
  50071=>"100000111",
  50072=>"111000000",
  50073=>"111011011",
  50074=>"111100111",
  50075=>"111110110",
  50076=>"100000000",
  50077=>"000000011",
  50078=>"000000001",
  50079=>"000000000",
  50080=>"100101000",
  50081=>"001111111",
  50082=>"000000111",
  50083=>"110111101",
  50084=>"011110110",
  50085=>"000000111",
  50086=>"111100111",
  50087=>"110111111",
  50088=>"010100000",
  50089=>"010010011",
  50090=>"110011000",
  50091=>"110000000",
  50092=>"000111000",
  50093=>"111110111",
  50094=>"110000011",
  50095=>"111111000",
  50096=>"111000011",
  50097=>"000000000",
  50098=>"000000000",
  50099=>"111111000",
  50100=>"111111111",
  50101=>"000000010",
  50102=>"000000000",
  50103=>"000000000",
  50104=>"000000011",
  50105=>"001111111",
  50106=>"111101100",
  50107=>"110000000",
  50108=>"111000000",
  50109=>"111111110",
  50110=>"100100000",
  50111=>"011001011",
  50112=>"001111110",
  50113=>"000000111",
  50114=>"010111111",
  50115=>"000000000",
  50116=>"111100000",
  50117=>"000000000",
  50118=>"101111011",
  50119=>"000000000",
  50120=>"011000000",
  50121=>"111111110",
  50122=>"100000000",
  50123=>"111111000",
  50124=>"000000111",
  50125=>"001000111",
  50126=>"100100000",
  50127=>"011111001",
  50128=>"100000000",
  50129=>"000001111",
  50130=>"000111001",
  50131=>"000000100",
  50132=>"111011010",
  50133=>"111111111",
  50134=>"000000000",
  50135=>"100111110",
  50136=>"000000111",
  50137=>"111111111",
  50138=>"111110111",
  50139=>"101000000",
  50140=>"111011111",
  50141=>"111111111",
  50142=>"000000101",
  50143=>"001011100",
  50144=>"010110011",
  50145=>"111100000",
  50146=>"000100111",
  50147=>"011111111",
  50148=>"111100000",
  50149=>"000000000",
  50150=>"010000000",
  50151=>"101100111",
  50152=>"100100010",
  50153=>"000000111",
  50154=>"111011111",
  50155=>"000000011",
  50156=>"100000011",
  50157=>"111011001",
  50158=>"011000000",
  50159=>"000000111",
  50160=>"100111111",
  50161=>"100000000",
  50162=>"111111011",
  50163=>"000000000",
  50164=>"111111000",
  50165=>"100100110",
  50166=>"000010110",
  50167=>"000000111",
  50168=>"000000111",
  50169=>"100110011",
  50170=>"011110000",
  50171=>"111111111",
  50172=>"100000000",
  50173=>"111111111",
  50174=>"111111000",
  50175=>"000000000",
  50176=>"000000000",
  50177=>"000010011",
  50178=>"111111111",
  50179=>"000000111",
  50180=>"000000001",
  50181=>"111000000",
  50182=>"000000000",
  50183=>"101111111",
  50184=>"000010011",
  50185=>"011111000",
  50186=>"111111111",
  50187=>"111001001",
  50188=>"010100000",
  50189=>"000000000",
  50190=>"011111011",
  50191=>"111111111",
  50192=>"111111111",
  50193=>"000000011",
  50194=>"000000111",
  50195=>"111111111",
  50196=>"011111111",
  50197=>"101111111",
  50198=>"000000011",
  50199=>"000100000",
  50200=>"001001111",
  50201=>"001000010",
  50202=>"000000111",
  50203=>"011100111",
  50204=>"111111111",
  50205=>"111111111",
  50206=>"110111111",
  50207=>"111111111",
  50208=>"000000111",
  50209=>"011000001",
  50210=>"001000010",
  50211=>"111111000",
  50212=>"110111111",
  50213=>"111111111",
  50214=>"100100000",
  50215=>"100000001",
  50216=>"000000100",
  50217=>"011010011",
  50218=>"111111111",
  50219=>"111111111",
  50220=>"000000000",
  50221=>"000000000",
  50222=>"100001001",
  50223=>"000000000",
  50224=>"000000000",
  50225=>"110111111",
  50226=>"001001011",
  50227=>"000000000",
  50228=>"111100000",
  50229=>"110110000",
  50230=>"000000000",
  50231=>"000000110",
  50232=>"001111111",
  50233=>"111000000",
  50234=>"000000000",
  50235=>"111111111",
  50236=>"000000000",
  50237=>"010010111",
  50238=>"000000000",
  50239=>"111011111",
  50240=>"000000001",
  50241=>"111010010",
  50242=>"000111011",
  50243=>"111000000",
  50244=>"111100101",
  50245=>"110110010",
  50246=>"000000101",
  50247=>"000011111",
  50248=>"110100000",
  50249=>"111111111",
  50250=>"000100110",
  50251=>"001001001",
  50252=>"011011111",
  50253=>"100100011",
  50254=>"111110000",
  50255=>"000001111",
  50256=>"000000010",
  50257=>"110000000",
  50258=>"010000000",
  50259=>"011111111",
  50260=>"101000000",
  50261=>"000000000",
  50262=>"111000111",
  50263=>"000000000",
  50264=>"100000000",
  50265=>"000000000",
  50266=>"111111111",
  50267=>"010010011",
  50268=>"000000000",
  50269=>"111111111",
  50270=>"000100110",
  50271=>"110000000",
  50272=>"000000000",
  50273=>"110000000",
  50274=>"000000111",
  50275=>"000000001",
  50276=>"000000000",
  50277=>"001001111",
  50278=>"111000001",
  50279=>"001000000",
  50280=>"000000000",
  50281=>"111111000",
  50282=>"111011000",
  50283=>"111111110",
  50284=>"111011000",
  50285=>"000000000",
  50286=>"111111111",
  50287=>"000000000",
  50288=>"000001000",
  50289=>"111111111",
  50290=>"000110000",
  50291=>"110111110",
  50292=>"111100100",
  50293=>"111111000",
  50294=>"000111000",
  50295=>"111111101",
  50296=>"111111111",
  50297=>"000100111",
  50298=>"000001111",
  50299=>"111111111",
  50300=>"000000000",
  50301=>"111111111",
  50302=>"000000000",
  50303=>"000000000",
  50304=>"010110110",
  50305=>"001111000",
  50306=>"000000000",
  50307=>"010000100",
  50308=>"001001001",
  50309=>"000000100",
  50310=>"111110110",
  50311=>"000111111",
  50312=>"000001111",
  50313=>"000000000",
  50314=>"111111110",
  50315=>"000000000",
  50316=>"110110111",
  50317=>"111111000",
  50318=>"000011011",
  50319=>"010000000",
  50320=>"000000111",
  50321=>"111111111",
  50322=>"000000000",
  50323=>"000000000",
  50324=>"000000111",
  50325=>"000011011",
  50326=>"001111111",
  50327=>"110000000",
  50328=>"000000000",
  50329=>"110110000",
  50330=>"100100000",
  50331=>"111111111",
  50332=>"100000000",
  50333=>"011111111",
  50334=>"111111000",
  50335=>"000111111",
  50336=>"000000000",
  50337=>"000000000",
  50338=>"111111111",
  50339=>"111011000",
  50340=>"000110111",
  50341=>"011011111",
  50342=>"111111111",
  50343=>"111011000",
  50344=>"111111000",
  50345=>"010000000",
  50346=>"000000000",
  50347=>"111111000",
  50348=>"111011000",
  50349=>"000000110",
  50350=>"100000111",
  50351=>"000000000",
  50352=>"111111110",
  50353=>"111111011",
  50354=>"111111111",
  50355=>"111111000",
  50356=>"000100000",
  50357=>"000000100",
  50358=>"111010011",
  50359=>"000000000",
  50360=>"111111101",
  50361=>"000000111",
  50362=>"000000000",
  50363=>"000000000",
  50364=>"101111100",
  50365=>"000000000",
  50366=>"000000100",
  50367=>"000000000",
  50368=>"000000000",
  50369=>"100000000",
  50370=>"000000001",
  50371=>"111111111",
  50372=>"000000001",
  50373=>"011111001",
  50374=>"000000000",
  50375=>"111111111",
  50376=>"111000000",
  50377=>"011000001",
  50378=>"000000000",
  50379=>"111111111",
  50380=>"000000000",
  50381=>"000100001",
  50382=>"111111111",
  50383=>"000000000",
  50384=>"000000000",
  50385=>"100000000",
  50386=>"000000000",
  50387=>"000000000",
  50388=>"000000111",
  50389=>"111111000",
  50390=>"000000111",
  50391=>"001111111",
  50392=>"001000111",
  50393=>"000010111",
  50394=>"000000110",
  50395=>"111000000",
  50396=>"000000000",
  50397=>"111111111",
  50398=>"111000000",
  50399=>"010001000",
  50400=>"110111101",
  50401=>"000000000",
  50402=>"111000000",
  50403=>"000010000",
  50404=>"000000000",
  50405=>"000011111",
  50406=>"001011111",
  50407=>"111111111",
  50408=>"110111111",
  50409=>"111111111",
  50410=>"111001111",
  50411=>"000000000",
  50412=>"000000000",
  50413=>"000000000",
  50414=>"000000000",
  50415=>"000000000",
  50416=>"111110000",
  50417=>"111011011",
  50418=>"000000000",
  50419=>"000000001",
  50420=>"111111111",
  50421=>"000000001",
  50422=>"110010111",
  50423=>"111111111",
  50424=>"111001000",
  50425=>"000000000",
  50426=>"111000000",
  50427=>"000100100",
  50428=>"011111111",
  50429=>"100000000",
  50430=>"000011011",
  50431=>"111111111",
  50432=>"111111111",
  50433=>"000110000",
  50434=>"010110100",
  50435=>"111111110",
  50436=>"111010111",
  50437=>"111111100",
  50438=>"110100110",
  50439=>"000000011",
  50440=>"000000000",
  50441=>"000000000",
  50442=>"001011111",
  50443=>"111111111",
  50444=>"000000111",
  50445=>"100000000",
  50446=>"111010001",
  50447=>"111111110",
  50448=>"010000000",
  50449=>"000000000",
  50450=>"000000000",
  50451=>"111011111",
  50452=>"000000000",
  50453=>"000000000",
  50454=>"000000000",
  50455=>"111111000",
  50456=>"111111111",
  50457=>"000000110",
  50458=>"101100000",
  50459=>"111111111",
  50460=>"111011001",
  50461=>"000000000",
  50462=>"111111111",
  50463=>"011010110",
  50464=>"000000111",
  50465=>"000001111",
  50466=>"000000000",
  50467=>"011111111",
  50468=>"000000111",
  50469=>"111111111",
  50470=>"000001011",
  50471=>"000011010",
  50472=>"000000000",
  50473=>"110000000",
  50474=>"111111101",
  50475=>"000100100",
  50476=>"111111111",
  50477=>"001011000",
  50478=>"111111111",
  50479=>"111111111",
  50480=>"000000001",
  50481=>"111011001",
  50482=>"101000000",
  50483=>"111010010",
  50484=>"000011000",
  50485=>"110000000",
  50486=>"001000100",
  50487=>"000000000",
  50488=>"110110010",
  50489=>"111111111",
  50490=>"001111111",
  50491=>"001111111",
  50492=>"111111111",
  50493=>"111111111",
  50494=>"011001000",
  50495=>"000000110",
  50496=>"000000000",
  50497=>"111111111",
  50498=>"111111011",
  50499=>"000001111",
  50500=>"111111111",
  50501=>"001000000",
  50502=>"000000000",
  50503=>"001000000",
  50504=>"111111111",
  50505=>"111111111",
  50506=>"000000111",
  50507=>"000000101",
  50508=>"111111111",
  50509=>"000000000",
  50510=>"000010011",
  50511=>"001011000",
  50512=>"111000000",
  50513=>"011000100",
  50514=>"100000000",
  50515=>"000000010",
  50516=>"001111011",
  50517=>"011000001",
  50518=>"000000000",
  50519=>"000000000",
  50520=>"000111111",
  50521=>"000100100",
  50522=>"000001000",
  50523=>"000000000",
  50524=>"111111111",
  50525=>"110110010",
  50526=>"000000000",
  50527=>"111100110",
  50528=>"001001001",
  50529=>"111001001",
  50530=>"110111110",
  50531=>"111111111",
  50532=>"111111111",
  50533=>"000000000",
  50534=>"000000000",
  50535=>"011011111",
  50536=>"000000000",
  50537=>"010000000",
  50538=>"000000000",
  50539=>"111111111",
  50540=>"001001011",
  50541=>"010110111",
  50542=>"111111100",
  50543=>"000111011",
  50544=>"111111111",
  50545=>"000010001",
  50546=>"000000000",
  50547=>"011001111",
  50548=>"000111111",
  50549=>"111110100",
  50550=>"111111011",
  50551=>"000000000",
  50552=>"110001011",
  50553=>"000000000",
  50554=>"000000000",
  50555=>"000111111",
  50556=>"000000000",
  50557=>"100000011",
  50558=>"000010000",
  50559=>"111101000",
  50560=>"110010111",
  50561=>"110111111",
  50562=>"000001001",
  50563=>"000000000",
  50564=>"000000000",
  50565=>"000000000",
  50566=>"110001101",
  50567=>"000000011",
  50568=>"111111111",
  50569=>"000000000",
  50570=>"111111111",
  50571=>"111111111",
  50572=>"101000001",
  50573=>"001001000",
  50574=>"000000001",
  50575=>"001001000",
  50576=>"000000000",
  50577=>"000000110",
  50578=>"000011111",
  50579=>"111111110",
  50580=>"000000000",
  50581=>"000000000",
  50582=>"110100101",
  50583=>"000000000",
  50584=>"000011011",
  50585=>"111111011",
  50586=>"111111100",
  50587=>"111111111",
  50588=>"001000000",
  50589=>"010000000",
  50590=>"000000000",
  50591=>"000010111",
  50592=>"001000000",
  50593=>"010010000",
  50594=>"111001011",
  50595=>"111000000",
  50596=>"111000000",
  50597=>"001111110",
  50598=>"101101101",
  50599=>"110011000",
  50600=>"100100100",
  50601=>"111111111",
  50602=>"011000000",
  50603=>"000000001",
  50604=>"110010000",
  50605=>"000000000",
  50606=>"000001111",
  50607=>"001100000",
  50608=>"111111111",
  50609=>"111001000",
  50610=>"000000000",
  50611=>"111111111",
  50612=>"111111111",
  50613=>"111111111",
  50614=>"000111111",
  50615=>"000011111",
  50616=>"111111001",
  50617=>"011000111",
  50618=>"010000010",
  50619=>"111000000",
  50620=>"000110111",
  50621=>"110110000",
  50622=>"000000000",
  50623=>"110100110",
  50624=>"111111111",
  50625=>"111111111",
  50626=>"000001000",
  50627=>"000000000",
  50628=>"110000000",
  50629=>"101110110",
  50630=>"000000000",
  50631=>"110111111",
  50632=>"011000100",
  50633=>"000000010",
  50634=>"001000000",
  50635=>"111111111",
  50636=>"100100000",
  50637=>"000000000",
  50638=>"000000000",
  50639=>"010111111",
  50640=>"000000111",
  50641=>"111111111",
  50642=>"000001001",
  50643=>"000000000",
  50644=>"111100000",
  50645=>"000110111",
  50646=>"000000001",
  50647=>"100000000",
  50648=>"111100111",
  50649=>"000000000",
  50650=>"111110000",
  50651=>"000000000",
  50652=>"000000000",
  50653=>"111111111",
  50654=>"111111111",
  50655=>"110111000",
  50656=>"000001001",
  50657=>"000000000",
  50658=>"111111111",
  50659=>"010010000",
  50660=>"000000001",
  50661=>"001000111",
  50662=>"111111111",
  50663=>"000000111",
  50664=>"000000000",
  50665=>"001000000",
  50666=>"010010110",
  50667=>"010111010",
  50668=>"111111111",
  50669=>"011001000",
  50670=>"111111111",
  50671=>"111111111",
  50672=>"110111111",
  50673=>"000000000",
  50674=>"001001000",
  50675=>"000000000",
  50676=>"000000111",
  50677=>"111110111",
  50678=>"010010010",
  50679=>"100100000",
  50680=>"000000000",
  50681=>"011001011",
  50682=>"000000010",
  50683=>"111111101",
  50684=>"011000100",
  50685=>"110110111",
  50686=>"000000000",
  50687=>"000000000",
  50688=>"011011111",
  50689=>"100110010",
  50690=>"111000000",
  50691=>"111111100",
  50692=>"010000000",
  50693=>"001000000",
  50694=>"101111111",
  50695=>"110000100",
  50696=>"011111011",
  50697=>"001111111",
  50698=>"111111100",
  50699=>"110111000",
  50700=>"001011011",
  50701=>"110000000",
  50702=>"110000000",
  50703=>"001000101",
  50704=>"010000000",
  50705=>"000111111",
  50706=>"000111111",
  50707=>"100100110",
  50708=>"111000000",
  50709=>"111111000",
  50710=>"000000001",
  50711=>"100000000",
  50712=>"011011000",
  50713=>"001001100",
  50714=>"111111000",
  50715=>"111000000",
  50716=>"000000000",
  50717=>"000000110",
  50718=>"001001111",
  50719=>"101000000",
  50720=>"000000000",
  50721=>"011001000",
  50722=>"000111110",
  50723=>"110000000",
  50724=>"111111111",
  50725=>"111111111",
  50726=>"000000011",
  50727=>"101100101",
  50728=>"000000000",
  50729=>"111111111",
  50730=>"000000000",
  50731=>"011000001",
  50732=>"110111111",
  50733=>"000111111",
  50734=>"000000000",
  50735=>"000000111",
  50736=>"110100100",
  50737=>"001001001",
  50738=>"100100100",
  50739=>"000000110",
  50740=>"000000000",
  50741=>"110100001",
  50742=>"100000100",
  50743=>"000010000",
  50744=>"101111011",
  50745=>"100000111",
  50746=>"111111111",
  50747=>"000000111",
  50748=>"100100100",
  50749=>"000000000",
  50750=>"011111111",
  50751=>"100000111",
  50752=>"000000100",
  50753=>"000000110",
  50754=>"111001000",
  50755=>"111001011",
  50756=>"011011011",
  50757=>"001011111",
  50758=>"111000000",
  50759=>"011111111",
  50760=>"000100010",
  50761=>"000000000",
  50762=>"111100000",
  50763=>"000000011",
  50764=>"101111001",
  50765=>"101001111",
  50766=>"000000000",
  50767=>"000000001",
  50768=>"000111111",
  50769=>"111110110",
  50770=>"111000000",
  50771=>"100000000",
  50772=>"101111111",
  50773=>"111111110",
  50774=>"111011111",
  50775=>"000000000",
  50776=>"001001000",
  50777=>"111000100",
  50778=>"111100000",
  50779=>"001111111",
  50780=>"111111101",
  50781=>"000000000",
  50782=>"011001000",
  50783=>"011011011",
  50784=>"010001010",
  50785=>"000000000",
  50786=>"000000000",
  50787=>"010011111",
  50788=>"011110110",
  50789=>"000010011",
  50790=>"111111110",
  50791=>"100111100",
  50792=>"011111111",
  50793=>"000000100",
  50794=>"111111111",
  50795=>"000000001",
  50796=>"111011000",
  50797=>"000000101",
  50798=>"000000100",
  50799=>"000111111",
  50800=>"111111111",
  50801=>"111001001",
  50802=>"000100111",
  50803=>"100000000",
  50804=>"000110100",
  50805=>"111101111",
  50806=>"001111111",
  50807=>"111111111",
  50808=>"010000001",
  50809=>"011000000",
  50810=>"100100100",
  50811=>"000000000",
  50812=>"111111101",
  50813=>"000000000",
  50814=>"100000000",
  50815=>"000001111",
  50816=>"000000001",
  50817=>"111010110",
  50818=>"111000001",
  50819=>"100100110",
  50820=>"000111111",
  50821=>"111001111",
  50822=>"000000000",
  50823=>"111111111",
  50824=>"001000111",
  50825=>"110000001",
  50826=>"111111000",
  50827=>"111111010",
  50828=>"010111111",
  50829=>"100000000",
  50830=>"011011111",
  50831=>"000111011",
  50832=>"111101001",
  50833=>"111111101",
  50834=>"111101101",
  50835=>"000000000",
  50836=>"000000011",
  50837=>"000000000",
  50838=>"000110111",
  50839=>"111111000",
  50840=>"000000101",
  50841=>"111111010",
  50842=>"000000001",
  50843=>"000000000",
  50844=>"100111011",
  50845=>"000000001",
  50846=>"111000000",
  50847=>"000100100",
  50848=>"111111111",
  50849=>"111111000",
  50850=>"111101101",
  50851=>"111111111",
  50852=>"111001111",
  50853=>"111000101",
  50854=>"111111000",
  50855=>"001010010",
  50856=>"000000000",
  50857=>"000000001",
  50858=>"001001000",
  50859=>"000000000",
  50860=>"000011111",
  50861=>"111111000",
  50862=>"110110110",
  50863=>"000000000",
  50864=>"000111111",
  50865=>"100111011",
  50866=>"001101001",
  50867=>"111101101",
  50868=>"011100101",
  50869=>"111011001",
  50870=>"111111111",
  50871=>"100100010",
  50872=>"000011010",
  50873=>"000111010",
  50874=>"110100111",
  50875=>"100001111",
  50876=>"011011000",
  50877=>"000000000",
  50878=>"111111101",
  50879=>"000110100",
  50880=>"000000111",
  50881=>"011011000",
  50882=>"000000000",
  50883=>"000000000",
  50884=>"010111111",
  50885=>"000000010",
  50886=>"000000000",
  50887=>"111011101",
  50888=>"101111111",
  50889=>"000001111",
  50890=>"000000000",
  50891=>"000000111",
  50892=>"011000000",
  50893=>"000111111",
  50894=>"000000100",
  50895=>"110110111",
  50896=>"111111101",
  50897=>"000001111",
  50898=>"101101101",
  50899=>"000000110",
  50900=>"111111111",
  50901=>"100000000",
  50902=>"001001001",
  50903=>"000000000",
  50904=>"000001000",
  50905=>"000111111",
  50906=>"000000111",
  50907=>"111111011",
  50908=>"111100000",
  50909=>"110000000",
  50910=>"001000000",
  50911=>"001000000",
  50912=>"001000010",
  50913=>"000111111",
  50914=>"110111110",
  50915=>"111111111",
  50916=>"110010000",
  50917=>"100110111",
  50918=>"000100111",
  50919=>"111111111",
  50920=>"111111100",
  50921=>"011111111",
  50922=>"111111111",
  50923=>"000000001",
  50924=>"100100111",
  50925=>"000000000",
  50926=>"110000010",
  50927=>"101101100",
  50928=>"110011011",
  50929=>"111101111",
  50930=>"100101111",
  50931=>"111101101",
  50932=>"000000111",
  50933=>"101100100",
  50934=>"100100101",
  50935=>"000011000",
  50936=>"111110010",
  50937=>"000100000",
  50938=>"100000001",
  50939=>"011011011",
  50940=>"100111000",
  50941=>"000000000",
  50942=>"100000111",
  50943=>"000111111",
  50944=>"101111111",
  50945=>"011010110",
  50946=>"111011000",
  50947=>"111111000",
  50948=>"111111111",
  50949=>"001001101",
  50950=>"000000000",
  50951=>"101100001",
  50952=>"110100100",
  50953=>"000000000",
  50954=>"111100100",
  50955=>"010101111",
  50956=>"000000000",
  50957=>"100001101",
  50958=>"000000000",
  50959=>"111000000",
  50960=>"101001000",
  50961=>"111100101",
  50962=>"000000000",
  50963=>"000000000",
  50964=>"001001000",
  50965=>"110111111",
  50966=>"000111111",
  50967=>"000000000",
  50968=>"000000111",
  50969=>"111101011",
  50970=>"000000010",
  50971=>"101111111",
  50972=>"001001000",
  50973=>"111111111",
  50974=>"001111111",
  50975=>"111111100",
  50976=>"100100110",
  50977=>"100000000",
  50978=>"100111111",
  50979=>"111110000",
  50980=>"000010111",
  50981=>"000000000",
  50982=>"000110010",
  50983=>"011001010",
  50984=>"010000101",
  50985=>"100100101",
  50986=>"000101000",
  50987=>"100000000",
  50988=>"000000000",
  50989=>"011010110",
  50990=>"111111111",
  50991=>"000000111",
  50992=>"111111111",
  50993=>"000000100",
  50994=>"111000000",
  50995=>"111111000",
  50996=>"000000000",
  50997=>"011111100",
  50998=>"110011011",
  50999=>"000111001",
  51000=>"011110000",
  51001=>"111000000",
  51002=>"000000000",
  51003=>"100000111",
  51004=>"101100100",
  51005=>"111111110",
  51006=>"000111001",
  51007=>"111100000",
  51008=>"111111000",
  51009=>"100100100",
  51010=>"000000000",
  51011=>"010010010",
  51012=>"000000001",
  51013=>"110011111",
  51014=>"010010000",
  51015=>"111100000",
  51016=>"001000000",
  51017=>"001000000",
  51018=>"111110000",
  51019=>"000000000",
  51020=>"001111111",
  51021=>"000000111",
  51022=>"101000000",
  51023=>"000000101",
  51024=>"000000001",
  51025=>"111110111",
  51026=>"111111000",
  51027=>"000001011",
  51028=>"000110000",
  51029=>"111110111",
  51030=>"111000000",
  51031=>"100110111",
  51032=>"000000000",
  51033=>"001001001",
  51034=>"111001000",
  51035=>"110000111",
  51036=>"111111110",
  51037=>"101100101",
  51038=>"010000001",
  51039=>"111111110",
  51040=>"000000111",
  51041=>"000111111",
  51042=>"000110111",
  51043=>"111111000",
  51044=>"000001111",
  51045=>"111000000",
  51046=>"000100100",
  51047=>"000111110",
  51048=>"011010010",
  51049=>"000011011",
  51050=>"001111111",
  51051=>"101100000",
  51052=>"011011011",
  51053=>"111100100",
  51054=>"000011011",
  51055=>"111101111",
  51056=>"111111000",
  51057=>"111111000",
  51058=>"100111111",
  51059=>"001100100",
  51060=>"000000000",
  51061=>"000000000",
  51062=>"000000000",
  51063=>"111111110",
  51064=>"000000000",
  51065=>"000111001",
  51066=>"111011000",
  51067=>"101001001",
  51068=>"000000111",
  51069=>"000100110",
  51070=>"000000000",
  51071=>"001010010",
  51072=>"001001101",
  51073=>"000001000",
  51074=>"100100011",
  51075=>"000111000",
  51076=>"000010111",
  51077=>"000000000",
  51078=>"000000000",
  51079=>"010010111",
  51080=>"111111011",
  51081=>"000000000",
  51082=>"011011011",
  51083=>"000010000",
  51084=>"000000001",
  51085=>"110000000",
  51086=>"000000111",
  51087=>"000000111",
  51088=>"111111111",
  51089=>"111100101",
  51090=>"000111111",
  51091=>"000101111",
  51092=>"111111000",
  51093=>"000110110",
  51094=>"000000000",
  51095=>"111100000",
  51096=>"000001001",
  51097=>"111001001",
  51098=>"110100000",
  51099=>"111111111",
  51100=>"101001100",
  51101=>"000010100",
  51102=>"111000100",
  51103=>"011111111",
  51104=>"000100000",
  51105=>"101100100",
  51106=>"000000000",
  51107=>"111011000",
  51108=>"000000000",
  51109=>"001111110",
  51110=>"111000000",
  51111=>"111011000",
  51112=>"110110000",
  51113=>"100110111",
  51114=>"000000000",
  51115=>"111000000",
  51116=>"011111111",
  51117=>"111111011",
  51118=>"111111111",
  51119=>"111000000",
  51120=>"111100000",
  51121=>"101101000",
  51122=>"000111111",
  51123=>"111101111",
  51124=>"111100100",
  51125=>"000000000",
  51126=>"000000000",
  51127=>"000000000",
  51128=>"101111111",
  51129=>"111000101",
  51130=>"000000101",
  51131=>"000100110",
  51132=>"111101100",
  51133=>"000000000",
  51134=>"000001000",
  51135=>"000000011",
  51136=>"111111111",
  51137=>"000000110",
  51138=>"111000000",
  51139=>"000111000",
  51140=>"100000000",
  51141=>"011001000",
  51142=>"001000000",
  51143=>"000000000",
  51144=>"110110100",
  51145=>"100000000",
  51146=>"100000010",
  51147=>"000000110",
  51148=>"100111000",
  51149=>"111000111",
  51150=>"100000001",
  51151=>"111011111",
  51152=>"111000001",
  51153=>"111100000",
  51154=>"000011011",
  51155=>"000001001",
  51156=>"111100100",
  51157=>"111110111",
  51158=>"000000000",
  51159=>"100110110",
  51160=>"111101101",
  51161=>"111111111",
  51162=>"000001111",
  51163=>"111001000",
  51164=>"000111000",
  51165=>"110111101",
  51166=>"000011111",
  51167=>"000000010",
  51168=>"011001011",
  51169=>"000000111",
  51170=>"110111111",
  51171=>"111111000",
  51172=>"111111000",
  51173=>"000000001",
  51174=>"000100111",
  51175=>"111111111",
  51176=>"000111111",
  51177=>"111111011",
  51178=>"000111110",
  51179=>"000000100",
  51180=>"101000001",
  51181=>"111110100",
  51182=>"111111000",
  51183=>"100000000",
  51184=>"111101101",
  51185=>"000000000",
  51186=>"000100100",
  51187=>"001000000",
  51188=>"110111000",
  51189=>"000000001",
  51190=>"110001001",
  51191=>"001001001",
  51192=>"000000000",
  51193=>"000000000",
  51194=>"000000001",
  51195=>"111111101",
  51196=>"101111111",
  51197=>"100000000",
  51198=>"101000111",
  51199=>"000010111",
  51200=>"000000000",
  51201=>"110100110",
  51202=>"111001111",
  51203=>"111111111",
  51204=>"111000100",
  51205=>"000100000",
  51206=>"011111111",
  51207=>"000000000",
  51208=>"111111000",
  51209=>"001001111",
  51210=>"011000001",
  51211=>"000000000",
  51212=>"100100100",
  51213=>"111111101",
  51214=>"111110100",
  51215=>"000110110",
  51216=>"000000111",
  51217=>"000000000",
  51218=>"001001000",
  51219=>"000001001",
  51220=>"000000000",
  51221=>"111001111",
  51222=>"101111111",
  51223=>"000000000",
  51224=>"011001000",
  51225=>"111111100",
  51226=>"000000000",
  51227=>"000000101",
  51228=>"100000000",
  51229=>"000000000",
  51230=>"100000000",
  51231=>"111111000",
  51232=>"000000100",
  51233=>"111111111",
  51234=>"101101001",
  51235=>"111111111",
  51236=>"000000110",
  51237=>"111000000",
  51238=>"000000000",
  51239=>"000000000",
  51240=>"000000100",
  51241=>"101111111",
  51242=>"000000000",
  51243=>"111111111",
  51244=>"000000111",
  51245=>"000000000",
  51246=>"111100001",
  51247=>"111111111",
  51248=>"111110110",
  51249=>"000001001",
  51250=>"111111111",
  51251=>"000000100",
  51252=>"000000000",
  51253=>"111111111",
  51254=>"001100100",
  51255=>"101000000",
  51256=>"111111111",
  51257=>"000000000",
  51258=>"111111011",
  51259=>"111111110",
  51260=>"100000000",
  51261=>"001001000",
  51262=>"111111111",
  51263=>"111100111",
  51264=>"011111111",
  51265=>"100111111",
  51266=>"000111111",
  51267=>"000000000",
  51268=>"111111111",
  51269=>"111111111",
  51270=>"000000000",
  51271=>"111111111",
  51272=>"000000000",
  51273=>"111111111",
  51274=>"111111111",
  51275=>"000000000",
  51276=>"000000111",
  51277=>"000000011",
  51278=>"000100000",
  51279=>"111111111",
  51280=>"111111110",
  51281=>"000000000",
  51282=>"000000100",
  51283=>"000000000",
  51284=>"111111111",
  51285=>"001001111",
  51286=>"100110111",
  51287=>"111111111",
  51288=>"001000001",
  51289=>"100000101",
  51290=>"111111111",
  51291=>"101000000",
  51292=>"011111111",
  51293=>"111111110",
  51294=>"110111110",
  51295=>"111100000",
  51296=>"110111111",
  51297=>"001101111",
  51298=>"011001111",
  51299=>"000110111",
  51300=>"000000000",
  51301=>"000000000",
  51302=>"001000000",
  51303=>"111110011",
  51304=>"000001101",
  51305=>"110111111",
  51306=>"000000000",
  51307=>"111011111",
  51308=>"111111111",
  51309=>"001000000",
  51310=>"000101111",
  51311=>"011011011",
  51312=>"111000000",
  51313=>"011001101",
  51314=>"000000001",
  51315=>"000010011",
  51316=>"000000000",
  51317=>"000000000",
  51318=>"000000001",
  51319=>"001001011",
  51320=>"010111110",
  51321=>"000000001",
  51322=>"000000000",
  51323=>"111111111",
  51324=>"110000010",
  51325=>"000010010",
  51326=>"000000000",
  51327=>"000000000",
  51328=>"000000000",
  51329=>"000000000",
  51330=>"000011001",
  51331=>"100000000",
  51332=>"000000000",
  51333=>"101101111",
  51334=>"001111111",
  51335=>"011111000",
  51336=>"111111111",
  51337=>"111010111",
  51338=>"111111111",
  51339=>"111001001",
  51340=>"111111111",
  51341=>"000000001",
  51342=>"101101100",
  51343=>"001000000",
  51344=>"000110110",
  51345=>"000000000",
  51346=>"000000001",
  51347=>"000000000",
  51348=>"000000000",
  51349=>"000100000",
  51350=>"011001000",
  51351=>"000000000",
  51352=>"111110110",
  51353=>"111111111",
  51354=>"000111111",
  51355=>"000000000",
  51356=>"001000000",
  51357=>"010010001",
  51358=>"100000100",
  51359=>"000000000",
  51360=>"001000000",
  51361=>"011111111",
  51362=>"000000000",
  51363=>"000000000",
  51364=>"000100000",
  51365=>"000000111",
  51366=>"100100100",
  51367=>"110000000",
  51368=>"111111111",
  51369=>"000100110",
  51370=>"000111100",
  51371=>"111011000",
  51372=>"000000000",
  51373=>"101100110",
  51374=>"111100100",
  51375=>"000000000",
  51376=>"111111111",
  51377=>"111111011",
  51378=>"110100000",
  51379=>"000000101",
  51380=>"111010110",
  51381=>"111111100",
  51382=>"100110110",
  51383=>"111111111",
  51384=>"011011001",
  51385=>"111111111",
  51386=>"000000000",
  51387=>"100101001",
  51388=>"000010011",
  51389=>"001000000",
  51390=>"111111111",
  51391=>"111000000",
  51392=>"111111111",
  51393=>"000100100",
  51394=>"000000000",
  51395=>"111111110",
  51396=>"000010111",
  51397=>"000000000",
  51398=>"000001001",
  51399=>"111000110",
  51400=>"011010000",
  51401=>"111101101",
  51402=>"000000000",
  51403=>"000001001",
  51404=>"100110011",
  51405=>"000100100",
  51406=>"000000000",
  51407=>"000000000",
  51408=>"100100000",
  51409=>"001000000",
  51410=>"000000000",
  51411=>"000000100",
  51412=>"111111111",
  51413=>"000000110",
  51414=>"000100111",
  51415=>"001101111",
  51416=>"111000000",
  51417=>"111110000",
  51418=>"000000000",
  51419=>"111111111",
  51420=>"001000000",
  51421=>"110110111",
  51422=>"000001111",
  51423=>"000000000",
  51424=>"111001011",
  51425=>"000000000",
  51426=>"110111110",
  51427=>"011001000",
  51428=>"000000000",
  51429=>"111110100",
  51430=>"000001011",
  51431=>"111111111",
  51432=>"111011001",
  51433=>"000000000",
  51434=>"000000000",
  51435=>"001001000",
  51436=>"011111111",
  51437=>"000000000",
  51438=>"000111111",
  51439=>"000000001",
  51440=>"100000000",
  51441=>"000000000",
  51442=>"001001111",
  51443=>"100000000",
  51444=>"011010000",
  51445=>"001111111",
  51446=>"000000001",
  51447=>"000000000",
  51448=>"111111000",
  51449=>"111111100",
  51450=>"000000000",
  51451=>"100000000",
  51452=>"011110111",
  51453=>"000000000",
  51454=>"000000111",
  51455=>"111111111",
  51456=>"000000000",
  51457=>"100100111",
  51458=>"000000000",
  51459=>"000001001",
  51460=>"111111111",
  51461=>"111111111",
  51462=>"100000000",
  51463=>"101000000",
  51464=>"011000000",
  51465=>"000000000",
  51466=>"111111111",
  51467=>"111111111",
  51468=>"110100000",
  51469=>"111101111",
  51470=>"000000000",
  51471=>"110000100",
  51472=>"000000000",
  51473=>"001001000",
  51474=>"000000000",
  51475=>"110111111",
  51476=>"000000000",
  51477=>"011000010",
  51478=>"000100111",
  51479=>"100100111",
  51480=>"000101000",
  51481=>"111110000",
  51482=>"000000000",
  51483=>"111011000",
  51484=>"110111111",
  51485=>"111111001",
  51486=>"000000000",
  51487=>"011111001",
  51488=>"011111001",
  51489=>"011111111",
  51490=>"000000000",
  51491=>"000000000",
  51492=>"111011011",
  51493=>"001111111",
  51494=>"111111111",
  51495=>"001001001",
  51496=>"010000011",
  51497=>"111111111",
  51498=>"011101101",
  51499=>"111111111",
  51500=>"101111000",
  51501=>"011011000",
  51502=>"111111000",
  51503=>"110110100",
  51504=>"000000000",
  51505=>"110100000",
  51506=>"000000000",
  51507=>"111111111",
  51508=>"000000000",
  51509=>"001101001",
  51510=>"100110011",
  51511=>"011000000",
  51512=>"101000000",
  51513=>"000000000",
  51514=>"000000000",
  51515=>"111111001",
  51516=>"001111110",
  51517=>"000000000",
  51518=>"000000000",
  51519=>"111111000",
  51520=>"000000000",
  51521=>"111011000",
  51522=>"000000000",
  51523=>"111111111",
  51524=>"111110110",
  51525=>"100100000",
  51526=>"000000000",
  51527=>"111011000",
  51528=>"100000000",
  51529=>"110000100",
  51530=>"111111000",
  51531=>"110110100",
  51532=>"000000000",
  51533=>"111111010",
  51534=>"111111111",
  51535=>"110110110",
  51536=>"000001000",
  51537=>"011000000",
  51538=>"000000011",
  51539=>"000000000",
  51540=>"000000000",
  51541=>"001001011",
  51542=>"111111111",
  51543=>"000000000",
  51544=>"111000000",
  51545=>"111111111",
  51546=>"000000000",
  51547=>"000000000",
  51548=>"000000110",
  51549=>"000011001",
  51550=>"110101101",
  51551=>"000000000",
  51552=>"110111111",
  51553=>"111111011",
  51554=>"000000000",
  51555=>"111000000",
  51556=>"000000010",
  51557=>"001001000",
  51558=>"000000000",
  51559=>"000000000",
  51560=>"111111111",
  51561=>"001111111",
  51562=>"000000000",
  51563=>"011000000",
  51564=>"000000111",
  51565=>"010000000",
  51566=>"111000000",
  51567=>"110110111",
  51568=>"111111010",
  51569=>"111111111",
  51570=>"000000000",
  51571=>"111111111",
  51572=>"000000000",
  51573=>"000000000",
  51574=>"000000000",
  51575=>"111111000",
  51576=>"111000000",
  51577=>"111001000",
  51578=>"000000000",
  51579=>"000111111",
  51580=>"000000000",
  51581=>"111110111",
  51582=>"011011011",
  51583=>"000000000",
  51584=>"111111111",
  51585=>"000000000",
  51586=>"111111111",
  51587=>"111111111",
  51588=>"111111111",
  51589=>"000110110",
  51590=>"000001011",
  51591=>"111111101",
  51592=>"000000000",
  51593=>"011011111",
  51594=>"111110111",
  51595=>"000110110",
  51596=>"100111111",
  51597=>"000110110",
  51598=>"000000110",
  51599=>"111111111",
  51600=>"000000001",
  51601=>"101000000",
  51602=>"000110000",
  51603=>"110001011",
  51604=>"111111010",
  51605=>"000000000",
  51606=>"000100111",
  51607=>"110110110",
  51608=>"001101111",
  51609=>"111111110",
  51610=>"111000000",
  51611=>"111111110",
  51612=>"000000000",
  51613=>"000000000",
  51614=>"111100000",
  51615=>"000000011",
  51616=>"011100111",
  51617=>"111100110",
  51618=>"111101111",
  51619=>"000000001",
  51620=>"111000000",
  51621=>"111011011",
  51622=>"111111111",
  51623=>"000000010",
  51624=>"001000000",
  51625=>"111111111",
  51626=>"000000000",
  51627=>"111011000",
  51628=>"110110100",
  51629=>"101100110",
  51630=>"000010111",
  51631=>"000000000",
  51632=>"011011111",
  51633=>"000111001",
  51634=>"111111000",
  51635=>"000110000",
  51636=>"000000000",
  51637=>"100000000",
  51638=>"000000000",
  51639=>"111111001",
  51640=>"100000111",
  51641=>"010111111",
  51642=>"111111011",
  51643=>"111000000",
  51644=>"111011011",
  51645=>"000100111",
  51646=>"000000101",
  51647=>"000000100",
  51648=>"111111111",
  51649=>"111001000",
  51650=>"000000111",
  51651=>"111100100",
  51652=>"111111111",
  51653=>"000000100",
  51654=>"111111111",
  51655=>"111101101",
  51656=>"111101100",
  51657=>"000000000",
  51658=>"100100100",
  51659=>"000100100",
  51660=>"000000000",
  51661=>"001000000",
  51662=>"111111110",
  51663=>"000000111",
  51664=>"000000000",
  51665=>"111111111",
  51666=>"000000000",
  51667=>"101000000",
  51668=>"110110100",
  51669=>"011000001",
  51670=>"100000000",
  51671=>"000000100",
  51672=>"100110111",
  51673=>"111111111",
  51674=>"100000001",
  51675=>"000000101",
  51676=>"100111111",
  51677=>"111111111",
  51678=>"000000000",
  51679=>"001101111",
  51680=>"000100111",
  51681=>"011011011",
  51682=>"010000000",
  51683=>"111001001",
  51684=>"011000000",
  51685=>"000011111",
  51686=>"000000000",
  51687=>"111111000",
  51688=>"000001111",
  51689=>"010111100",
  51690=>"111111111",
  51691=>"111111111",
  51692=>"000000000",
  51693=>"111111111",
  51694=>"000001001",
  51695=>"111111001",
  51696=>"000000000",
  51697=>"010111111",
  51698=>"001011001",
  51699=>"000000000",
  51700=>"001000000",
  51701=>"111111111",
  51702=>"111111111",
  51703=>"000000110",
  51704=>"000000000",
  51705=>"000000000",
  51706=>"011011001",
  51707=>"111111111",
  51708=>"000000000",
  51709=>"111111111",
  51710=>"001001111",
  51711=>"111111111",
  51712=>"010110110",
  51713=>"000000000",
  51714=>"111111111",
  51715=>"011000000",
  51716=>"100000000",
  51717=>"000001001",
  51718=>"011001001",
  51719=>"111100111",
  51720=>"000100000",
  51721=>"000000000",
  51722=>"000000001",
  51723=>"111100111",
  51724=>"111101101",
  51725=>"111110100",
  51726=>"010111011",
  51727=>"000000000",
  51728=>"010000001",
  51729=>"011111000",
  51730=>"011111110",
  51731=>"111001000",
  51732=>"000000000",
  51733=>"001000100",
  51734=>"000110110",
  51735=>"001011111",
  51736=>"110000000",
  51737=>"001001001",
  51738=>"000000000",
  51739=>"011001001",
  51740=>"100100100",
  51741=>"011000010",
  51742=>"000001011",
  51743=>"000000111",
  51744=>"101100000",
  51745=>"110111111",
  51746=>"000000111",
  51747=>"000000011",
  51748=>"000000110",
  51749=>"000111111",
  51750=>"111111110",
  51751=>"111000000",
  51752=>"100101111",
  51753=>"111111111",
  51754=>"001001000",
  51755=>"111110100",
  51756=>"011111000",
  51757=>"000001000",
  51758=>"000000001",
  51759=>"000100111",
  51760=>"101111011",
  51761=>"111111101",
  51762=>"001001001",
  51763=>"000000110",
  51764=>"010011100",
  51765=>"111100000",
  51766=>"111111110",
  51767=>"000000100",
  51768=>"111001000",
  51769=>"101000000",
  51770=>"111111111",
  51771=>"000000000",
  51772=>"110111100",
  51773=>"011011100",
  51774=>"110111111",
  51775=>"111000000",
  51776=>"111000001",
  51777=>"110110110",
  51778=>"000111111",
  51779=>"101000000",
  51780=>"100111001",
  51781=>"001001001",
  51782=>"000000000",
  51783=>"111101111",
  51784=>"011111110",
  51785=>"111111110",
  51786=>"111111111",
  51787=>"111111010",
  51788=>"000000000",
  51789=>"000100100",
  51790=>"000000000",
  51791=>"011111111",
  51792=>"000011110",
  51793=>"110111011",
  51794=>"100000100",
  51795=>"001111111",
  51796=>"001000000",
  51797=>"111111111",
  51798=>"101001111",
  51799=>"000110110",
  51800=>"001000001",
  51801=>"000000100",
  51802=>"000000011",
  51803=>"100100000",
  51804=>"111111111",
  51805=>"000000000",
  51806=>"111111101",
  51807=>"110111000",
  51808=>"000000000",
  51809=>"010111000",
  51810=>"001101111",
  51811=>"000000000",
  51812=>"110111111",
  51813=>"111111010",
  51814=>"000000111",
  51815=>"000001111",
  51816=>"000001011",
  51817=>"100000000",
  51818=>"111111100",
  51819=>"111111111",
  51820=>"111100100",
  51821=>"001101111",
  51822=>"111111111",
  51823=>"110111101",
  51824=>"000000001",
  51825=>"000000000",
  51826=>"000000100",
  51827=>"111111111",
  51828=>"011000111",
  51829=>"111111000",
  51830=>"000000000",
  51831=>"111111111",
  51832=>"000000000",
  51833=>"000000111",
  51834=>"111111011",
  51835=>"111101000",
  51836=>"110110001",
  51837=>"110000110",
  51838=>"111001000",
  51839=>"111111111",
  51840=>"000111100",
  51841=>"111111111",
  51842=>"111111110",
  51843=>"000000000",
  51844=>"101111111",
  51845=>"111101111",
  51846=>"100000000",
  51847=>"000000000",
  51848=>"101111111",
  51849=>"100000111",
  51850=>"111111111",
  51851=>"001000000",
  51852=>"011001001",
  51853=>"001000111",
  51854=>"111100000",
  51855=>"000111111",
  51856=>"011001000",
  51857=>"111111100",
  51858=>"000000011",
  51859=>"100110111",
  51860=>"111111111",
  51861=>"110111011",
  51862=>"000111111",
  51863=>"111000000",
  51864=>"011000000",
  51865=>"001011110",
  51866=>"111101111",
  51867=>"000111000",
  51868=>"111100100",
  51869=>"100111000",
  51870=>"111011011",
  51871=>"000000000",
  51872=>"011000110",
  51873=>"000101111",
  51874=>"111111011",
  51875=>"011111111",
  51876=>"111111010",
  51877=>"111111100",
  51878=>"111111111",
  51879=>"110110110",
  51880=>"111000100",
  51881=>"000011000",
  51882=>"111101001",
  51883=>"011011010",
  51884=>"101100100",
  51885=>"111111111",
  51886=>"000011110",
  51887=>"011000000",
  51888=>"111000001",
  51889=>"100100110",
  51890=>"111111000",
  51891=>"000000000",
  51892=>"100111111",
  51893=>"011000000",
  51894=>"111111111",
  51895=>"111111011",
  51896=>"110111111",
  51897=>"110000000",
  51898=>"100111110",
  51899=>"010010110",
  51900=>"000000000",
  51901=>"110100000",
  51902=>"000111111",
  51903=>"111111111",
  51904=>"111111111",
  51905=>"110000000",
  51906=>"100100101",
  51907=>"111111111",
  51908=>"111111110",
  51909=>"100000000",
  51910=>"010111010",
  51911=>"011000000",
  51912=>"111111100",
  51913=>"111111001",
  51914=>"101100101",
  51915=>"111111111",
  51916=>"100100100",
  51917=>"111111000",
  51918=>"111111111",
  51919=>"111111111",
  51920=>"000001001",
  51921=>"000111000",
  51922=>"000011000",
  51923=>"011111111",
  51924=>"100111111",
  51925=>"111111111",
  51926=>"000001000",
  51927=>"111110111",
  51928=>"111111000",
  51929=>"110110110",
  51930=>"000000000",
  51931=>"000100110",
  51932=>"111000111",
  51933=>"000000011",
  51934=>"100000011",
  51935=>"000000000",
  51936=>"111011000",
  51937=>"011111000",
  51938=>"000000000",
  51939=>"111100100",
  51940=>"101111111",
  51941=>"011000000",
  51942=>"111000111",
  51943=>"001101111",
  51944=>"110111000",
  51945=>"111111111",
  51946=>"111111100",
  51947=>"001101011",
  51948=>"100100000",
  51949=>"000000000",
  51950=>"101100000",
  51951=>"000000000",
  51952=>"111110110",
  51953=>"111010000",
  51954=>"011011111",
  51955=>"111000000",
  51956=>"111111100",
  51957=>"000000000",
  51958=>"011011011",
  51959=>"000000000",
  51960=>"011111111",
  51961=>"000000000",
  51962=>"111000000",
  51963=>"000000011",
  51964=>"000000111",
  51965=>"111110000",
  51966=>"111111111",
  51967=>"000111100",
  51968=>"010000011",
  51969=>"000000110",
  51970=>"101000001",
  51971=>"111111111",
  51972=>"111011001",
  51973=>"010110000",
  51974=>"001011111",
  51975=>"000000000",
  51976=>"101000000",
  51977=>"110110100",
  51978=>"000000001",
  51979=>"100100111",
  51980=>"000000000",
  51981=>"111011111",
  51982=>"000000000",
  51983=>"000000000",
  51984=>"001000000",
  51985=>"001000000",
  51986=>"111111001",
  51987=>"000100111",
  51988=>"000110000",
  51989=>"011000000",
  51990=>"001000101",
  51991=>"110000111",
  51992=>"111011001",
  51993=>"111111111",
  51994=>"000010111",
  51995=>"000000000",
  51996=>"100100100",
  51997=>"111000000",
  51998=>"000001001",
  51999=>"000000000",
  52000=>"000001101",
  52001=>"111000001",
  52002=>"111111111",
  52003=>"111111111",
  52004=>"111001000",
  52005=>"000011111",
  52006=>"000000110",
  52007=>"001001011",
  52008=>"000000011",
  52009=>"001111111",
  52010=>"111111111",
  52011=>"000000000",
  52012=>"111101100",
  52013=>"110111111",
  52014=>"000000000",
  52015=>"111111110",
  52016=>"011111001",
  52017=>"111000000",
  52018=>"000000011",
  52019=>"111111011",
  52020=>"000000000",
  52021=>"000000001",
  52022=>"111111111",
  52023=>"100000000",
  52024=>"011111111",
  52025=>"111111111",
  52026=>"000011111",
  52027=>"011111011",
  52028=>"000000111",
  52029=>"001011111",
  52030=>"100111111",
  52031=>"000010010",
  52032=>"111111101",
  52033=>"111111111",
  52034=>"000010110",
  52035=>"000000111",
  52036=>"000000000",
  52037=>"000000000",
  52038=>"000000101",
  52039=>"000000000",
  52040=>"111010000",
  52041=>"000000000",
  52042=>"000010011",
  52043=>"100100110",
  52044=>"000001000",
  52045=>"000110111",
  52046=>"111101111",
  52047=>"100010011",
  52048=>"111000000",
  52049=>"001101111",
  52050=>"000000100",
  52051=>"001000110",
  52052=>"000111111",
  52053=>"111001111",
  52054=>"111110101",
  52055=>"000000101",
  52056=>"111111101",
  52057=>"000000000",
  52058=>"110111010",
  52059=>"111001011",
  52060=>"000000000",
  52061=>"111011000",
  52062=>"000111000",
  52063=>"011111111",
  52064=>"001011011",
  52065=>"111101111",
  52066=>"000000101",
  52067=>"000000000",
  52068=>"000010100",
  52069=>"000000000",
  52070=>"000000000",
  52071=>"111000110",
  52072=>"000000110",
  52073=>"111001000",
  52074=>"000001011",
  52075=>"110110111",
  52076=>"111111111",
  52077=>"111011001",
  52078=>"000000101",
  52079=>"111100000",
  52080=>"111110000",
  52081=>"110100111",
  52082=>"010110011",
  52083=>"011011000",
  52084=>"001000000",
  52085=>"100100100",
  52086=>"110000000",
  52087=>"000000000",
  52088=>"000011001",
  52089=>"000000000",
  52090=>"000000000",
  52091=>"011111111",
  52092=>"111111011",
  52093=>"000101110",
  52094=>"000000000",
  52095=>"000000000",
  52096=>"100100100",
  52097=>"111110111",
  52098=>"111111011",
  52099=>"000000000",
  52100=>"111001000",
  52101=>"111111010",
  52102=>"110110000",
  52103=>"000000011",
  52104=>"000111000",
  52105=>"000000011",
  52106=>"111001001",
  52107=>"110011000",
  52108=>"111000001",
  52109=>"110110110",
  52110=>"000000111",
  52111=>"100101000",
  52112=>"100100100",
  52113=>"000000000",
  52114=>"000110111",
  52115=>"000000111",
  52116=>"011111111",
  52117=>"000011111",
  52118=>"111101011",
  52119=>"011000000",
  52120=>"001001001",
  52121=>"100111111",
  52122=>"000000000",
  52123=>"111111111",
  52124=>"001000000",
  52125=>"000000000",
  52126=>"100000000",
  52127=>"010000000",
  52128=>"000110111",
  52129=>"001001111",
  52130=>"111100100",
  52131=>"111101101",
  52132=>"111111110",
  52133=>"111111111",
  52134=>"000000000",
  52135=>"110100001",
  52136=>"000100111",
  52137=>"000000110",
  52138=>"111111111",
  52139=>"000000000",
  52140=>"000110110",
  52141=>"111111111",
  52142=>"110110111",
  52143=>"111111100",
  52144=>"111100000",
  52145=>"000001001",
  52146=>"000010000",
  52147=>"000000000",
  52148=>"010011000",
  52149=>"011000000",
  52150=>"100100110",
  52151=>"000000111",
  52152=>"110000000",
  52153=>"101001011",
  52154=>"100000001",
  52155=>"000000000",
  52156=>"000000000",
  52157=>"101001101",
  52158=>"000000000",
  52159=>"100000110",
  52160=>"001101111",
  52161=>"110011111",
  52162=>"111111110",
  52163=>"110100111",
  52164=>"001000111",
  52165=>"000000100",
  52166=>"011110111",
  52167=>"000000000",
  52168=>"011000000",
  52169=>"000000000",
  52170=>"000000100",
  52171=>"000000000",
  52172=>"000000000",
  52173=>"000111111",
  52174=>"000111110",
  52175=>"000000001",
  52176=>"000000110",
  52177=>"100111111",
  52178=>"111111111",
  52179=>"010000000",
  52180=>"000000000",
  52181=>"111111111",
  52182=>"111111111",
  52183=>"001011011",
  52184=>"111001001",
  52185=>"111001000",
  52186=>"000000000",
  52187=>"111000100",
  52188=>"111110000",
  52189=>"111111111",
  52190=>"111010000",
  52191=>"010110110",
  52192=>"000000000",
  52193=>"111001000",
  52194=>"000000001",
  52195=>"100000111",
  52196=>"111111111",
  52197=>"000000000",
  52198=>"010111011",
  52199=>"111111000",
  52200=>"000000000",
  52201=>"111111111",
  52202=>"101101111",
  52203=>"011111000",
  52204=>"000110000",
  52205=>"111111000",
  52206=>"110111110",
  52207=>"111111000",
  52208=>"100100100",
  52209=>"001001000",
  52210=>"000000111",
  52211=>"110111111",
  52212=>"111111110",
  52213=>"000100100",
  52214=>"000000000",
  52215=>"011000100",
  52216=>"111111100",
  52217=>"111111110",
  52218=>"111110111",
  52219=>"000001101",
  52220=>"111111111",
  52221=>"101110111",
  52222=>"101001111",
  52223=>"000000000",
  52224=>"000000000",
  52225=>"000111111",
  52226=>"000000000",
  52227=>"000111000",
  52228=>"000000101",
  52229=>"111111011",
  52230=>"100100000",
  52231=>"000000000",
  52232=>"111010111",
  52233=>"111001000",
  52234=>"001001000",
  52235=>"111111010",
  52236=>"000000011",
  52237=>"000100000",
  52238=>"000000000",
  52239=>"111001111",
  52240=>"000111111",
  52241=>"001111111",
  52242=>"111111100",
  52243=>"000000001",
  52244=>"110000000",
  52245=>"110110111",
  52246=>"000110110",
  52247=>"011001001",
  52248=>"000100000",
  52249=>"011111111",
  52250=>"000000000",
  52251=>"111111001",
  52252=>"111111111",
  52253=>"000000010",
  52254=>"111111110",
  52255=>"111111111",
  52256=>"001000000",
  52257=>"010000000",
  52258=>"111111111",
  52259=>"111111010",
  52260=>"001001000",
  52261=>"110111111",
  52262=>"111111111",
  52263=>"110111111",
  52264=>"000000001",
  52265=>"000000000",
  52266=>"111111111",
  52267=>"000111111",
  52268=>"110111101",
  52269=>"011001000",
  52270=>"111111111",
  52271=>"001001001",
  52272=>"010110011",
  52273=>"111111101",
  52274=>"011011011",
  52275=>"110000000",
  52276=>"010110000",
  52277=>"000000000",
  52278=>"000000000",
  52279=>"000111011",
  52280=>"111111000",
  52281=>"000111110",
  52282=>"111000101",
  52283=>"011000000",
  52284=>"111111111",
  52285=>"000000000",
  52286=>"000000011",
  52287=>"111011000",
  52288=>"111111010",
  52289=>"000110000",
  52290=>"100100111",
  52291=>"110111111",
  52292=>"000000000",
  52293=>"101000101",
  52294=>"000111110",
  52295=>"011000000",
  52296=>"011001011",
  52297=>"100110110",
  52298=>"000010111",
  52299=>"010110010",
  52300=>"000111111",
  52301=>"001011001",
  52302=>"011000000",
  52303=>"000100000",
  52304=>"110000000",
  52305=>"000000000",
  52306=>"000000010",
  52307=>"111101111",
  52308=>"111111111",
  52309=>"000000000",
  52310=>"111111110",
  52311=>"001100000",
  52312=>"111111111",
  52313=>"000000000",
  52314=>"111010000",
  52315=>"000010000",
  52316=>"000000000",
  52317=>"100000000",
  52318=>"110111111",
  52319=>"100110100",
  52320=>"000000110",
  52321=>"000000000",
  52322=>"111111001",
  52323=>"110111111",
  52324=>"110010100",
  52325=>"011111000",
  52326=>"011111111",
  52327=>"111111101",
  52328=>"000000110",
  52329=>"000000000",
  52330=>"110110000",
  52331=>"010111111",
  52332=>"010000000",
  52333=>"000000000",
  52334=>"000000001",
  52335=>"011111111",
  52336=>"110100111",
  52337=>"110111110",
  52338=>"011110110",
  52339=>"111100111",
  52340=>"111111111",
  52341=>"001001001",
  52342=>"111111111",
  52343=>"000001000",
  52344=>"000000000",
  52345=>"000000000",
  52346=>"000101111",
  52347=>"111110000",
  52348=>"011011011",
  52349=>"000010011",
  52350=>"000000000",
  52351=>"000111000",
  52352=>"111000111",
  52353=>"111111111",
  52354=>"111111111",
  52355=>"000000000",
  52356=>"111111111",
  52357=>"001001011",
  52358=>"000000000",
  52359=>"000000000",
  52360=>"111101000",
  52361=>"111011011",
  52362=>"111111111",
  52363=>"000011111",
  52364=>"010010000",
  52365=>"011001011",
  52366=>"000000000",
  52367=>"011000000",
  52368=>"000000000",
  52369=>"110110111",
  52370=>"111111011",
  52371=>"100100000",
  52372=>"000111000",
  52373=>"011011111",
  52374=>"110000010",
  52375=>"000000000",
  52376=>"100110111",
  52377=>"111111111",
  52378=>"000000011",
  52379=>"000011000",
  52380=>"111111111",
  52381=>"011111111",
  52382=>"110010000",
  52383=>"000000010",
  52384=>"000110110",
  52385=>"111110000",
  52386=>"011111110",
  52387=>"111011011",
  52388=>"000110111",
  52389=>"101000001",
  52390=>"000000000",
  52391=>"111110110",
  52392=>"000010111",
  52393=>"111111111",
  52394=>"111111111",
  52395=>"111110110",
  52396=>"111101111",
  52397=>"010010000",
  52398=>"110111111",
  52399=>"000100000",
  52400=>"000000001",
  52401=>"111111110",
  52402=>"000000000",
  52403=>"000000000",
  52404=>"000000011",
  52405=>"101011001",
  52406=>"111101111",
  52407=>"000000100",
  52408=>"000000000",
  52409=>"000000000",
  52410=>"000000100",
  52411=>"001000000",
  52412=>"000000000",
  52413=>"100000000",
  52414=>"111111111",
  52415=>"000000000",
  52416=>"000000000",
  52417=>"101111011",
  52418=>"110111110",
  52419=>"111111110",
  52420=>"011100000",
  52421=>"001000000",
  52422=>"001111111",
  52423=>"111011000",
  52424=>"000000000",
  52425=>"000000010",
  52426=>"000000011",
  52427=>"011011111",
  52428=>"000000000",
  52429=>"011111111",
  52430=>"011101001",
  52431=>"111111000",
  52432=>"010010111",
  52433=>"000001011",
  52434=>"001000000",
  52435=>"000000001",
  52436=>"001000000",
  52437=>"010110110",
  52438=>"000000000",
  52439=>"000000000",
  52440=>"000000000",
  52441=>"000000000",
  52442=>"110110111",
  52443=>"000000000",
  52444=>"010110111",
  52445=>"000000110",
  52446=>"011111111",
  52447=>"000000000",
  52448=>"000000001",
  52449=>"000001111",
  52450=>"000000111",
  52451=>"111000111",
  52452=>"111111111",
  52453=>"100000000",
  52454=>"000000000",
  52455=>"101000000",
  52456=>"111111111",
  52457=>"001001001",
  52458=>"111011000",
  52459=>"000000000",
  52460=>"000000000",
  52461=>"111111111",
  52462=>"111101101",
  52463=>"000000000",
  52464=>"101000011",
  52465=>"000000110",
  52466=>"000000000",
  52467=>"111100000",
  52468=>"010011111",
  52469=>"010000010",
  52470=>"100100111",
  52471=>"000000000",
  52472=>"110000100",
  52473=>"000000000",
  52474=>"010000111",
  52475=>"011011001",
  52476=>"111111100",
  52477=>"100000100",
  52478=>"111111111",
  52479=>"001001000",
  52480=>"000001001",
  52481=>"001010000",
  52482=>"000001111",
  52483=>"000000111",
  52484=>"111111111",
  52485=>"000110111",
  52486=>"100110000",
  52487=>"000000100",
  52488=>"111110111",
  52489=>"100110111",
  52490=>"110111011",
  52491=>"100000000",
  52492=>"000000000",
  52493=>"111101101",
  52494=>"000000000",
  52495=>"000001001",
  52496=>"111110010",
  52497=>"101101001",
  52498=>"100000111",
  52499=>"011111101",
  52500=>"000011000",
  52501=>"011111101",
  52502=>"000000000",
  52503=>"110100101",
  52504=>"101101101",
  52505=>"000000000",
  52506=>"000000000",
  52507=>"111111011",
  52508=>"110110010",
  52509=>"111110111",
  52510=>"111111111",
  52511=>"000110100",
  52512=>"110110101",
  52513=>"000111111",
  52514=>"110110110",
  52515=>"110010001",
  52516=>"101101100",
  52517=>"000111111",
  52518=>"000000100",
  52519=>"111111101",
  52520=>"000010000",
  52521=>"111111111",
  52522=>"011111011",
  52523=>"111111011",
  52524=>"110110111",
  52525=>"111111011",
  52526=>"000000000",
  52527=>"110110000",
  52528=>"111111011",
  52529=>"001111111",
  52530=>"000000000",
  52531=>"000001111",
  52532=>"000010000",
  52533=>"001011011",
  52534=>"011010010",
  52535=>"000111011",
  52536=>"000010000",
  52537=>"010010010",
  52538=>"000111111",
  52539=>"101111111",
  52540=>"111110011",
  52541=>"000000000",
  52542=>"100000000",
  52543=>"000000000",
  52544=>"000000000",
  52545=>"011110000",
  52546=>"011010000",
  52547=>"101111101",
  52548=>"000000000",
  52549=>"000000010",
  52550=>"111111111",
  52551=>"001011011",
  52552=>"111110111",
  52553=>"000100000",
  52554=>"011000010",
  52555=>"000010000",
  52556=>"111011011",
  52557=>"111111111",
  52558=>"110110010",
  52559=>"101101111",
  52560=>"111000100",
  52561=>"111111111",
  52562=>"000000010",
  52563=>"010000000",
  52564=>"010010000",
  52565=>"111111111",
  52566=>"111111111",
  52567=>"111100111",
  52568=>"000000000",
  52569=>"000000000",
  52570=>"000001000",
  52571=>"100000011",
  52572=>"111111110",
  52573=>"100101111",
  52574=>"000000000",
  52575=>"111111111",
  52576=>"111111110",
  52577=>"111101101",
  52578=>"101111011",
  52579=>"000011011",
  52580=>"011111111",
  52581=>"001001111",
  52582=>"111111111",
  52583=>"000000000",
  52584=>"011000000",
  52585=>"010000011",
  52586=>"111111011",
  52587=>"000000000",
  52588=>"111111111",
  52589=>"001111111",
  52590=>"100000000",
  52591=>"000000000",
  52592=>"001000000",
  52593=>"000000111",
  52594=>"000100000",
  52595=>"011010010",
  52596=>"100000111",
  52597=>"111111111",
  52598=>"111111111",
  52599=>"100001001",
  52600=>"111111111",
  52601=>"111111110",
  52602=>"001000000",
  52603=>"011011000",
  52604=>"100100101",
  52605=>"111111011",
  52606=>"111100000",
  52607=>"000010010",
  52608=>"011011001",
  52609=>"111111110",
  52610=>"000000000",
  52611=>"000000000",
  52612=>"111111111",
  52613=>"000000000",
  52614=>"001111111",
  52615=>"001001111",
  52616=>"000000100",
  52617=>"100010100",
  52618=>"111111011",
  52619=>"000101001",
  52620=>"110000111",
  52621=>"010010110",
  52622=>"100100110",
  52623=>"110111111",
  52624=>"000000000",
  52625=>"000000100",
  52626=>"111111111",
  52627=>"111111100",
  52628=>"000000111",
  52629=>"101101101",
  52630=>"001001001",
  52631=>"010001000",
  52632=>"111111111",
  52633=>"110111111",
  52634=>"000000000",
  52635=>"100111000",
  52636=>"000000000",
  52637=>"000000000",
  52638=>"000000000",
  52639=>"110111111",
  52640=>"101000000",
  52641=>"001011011",
  52642=>"010010000",
  52643=>"000000011",
  52644=>"010110110",
  52645=>"111111001",
  52646=>"000000000",
  52647=>"000000111",
  52648=>"100000000",
  52649=>"110110100",
  52650=>"000000111",
  52651=>"011010010",
  52652=>"100000100",
  52653=>"111111111",
  52654=>"100000011",
  52655=>"000110110",
  52656=>"000000110",
  52657=>"111111011",
  52658=>"000000001",
  52659=>"000000000",
  52660=>"000111111",
  52661=>"111110100",
  52662=>"111111111",
  52663=>"110111111",
  52664=>"000000000",
  52665=>"000000010",
  52666=>"111101111",
  52667=>"111110000",
  52668=>"010000000",
  52669=>"100111111",
  52670=>"111100000",
  52671=>"000010000",
  52672=>"000000000",
  52673=>"000000000",
  52674=>"000000000",
  52675=>"000000111",
  52676=>"000000110",
  52677=>"000110110",
  52678=>"011111000",
  52679=>"010000000",
  52680=>"000101001",
  52681=>"110110111",
  52682=>"110110010",
  52683=>"000000111",
  52684=>"000000000",
  52685=>"000001111",
  52686=>"000111010",
  52687=>"111111111",
  52688=>"111111111",
  52689=>"110110110",
  52690=>"000000000",
  52691=>"111111111",
  52692=>"000000001",
  52693=>"111001100",
  52694=>"000000000",
  52695=>"011000111",
  52696=>"000000000",
  52697=>"111111111",
  52698=>"110111111",
  52699=>"111100000",
  52700=>"111111111",
  52701=>"111111000",
  52702=>"110110110",
  52703=>"001011011",
  52704=>"000110110",
  52705=>"000000000",
  52706=>"100110010",
  52707=>"001000010",
  52708=>"111110111",
  52709=>"011000000",
  52710=>"000000111",
  52711=>"111100111",
  52712=>"110100100",
  52713=>"111111111",
  52714=>"000000000",
  52715=>"000111111",
  52716=>"000010000",
  52717=>"001000000",
  52718=>"111111111",
  52719=>"000000000",
  52720=>"000100100",
  52721=>"110110111",
  52722=>"111111010",
  52723=>"000010000",
  52724=>"110110000",
  52725=>"101101101",
  52726=>"000000000",
  52727=>"010111001",
  52728=>"000000000",
  52729=>"100100110",
  52730=>"111111111",
  52731=>"000000000",
  52732=>"110010000",
  52733=>"111111111",
  52734=>"111111111",
  52735=>"000000001",
  52736=>"001100111",
  52737=>"000000000",
  52738=>"000000101",
  52739=>"000111111",
  52740=>"111000101",
  52741=>"000000011",
  52742=>"100100100",
  52743=>"111000000",
  52744=>"000000000",
  52745=>"001001001",
  52746=>"000000000",
  52747=>"111111110",
  52748=>"111111111",
  52749=>"111000011",
  52750=>"111010011",
  52751=>"001000100",
  52752=>"100110100",
  52753=>"111111101",
  52754=>"000111111",
  52755=>"000000000",
  52756=>"111111001",
  52757=>"111000000",
  52758=>"000111111",
  52759=>"111000100",
  52760=>"000011111",
  52761=>"111111110",
  52762=>"000000000",
  52763=>"000000111",
  52764=>"000111111",
  52765=>"100101100",
  52766=>"111111000",
  52767=>"111010000",
  52768=>"000111111",
  52769=>"111111111",
  52770=>"111111111",
  52771=>"111001001",
  52772=>"111111111",
  52773=>"110000011",
  52774=>"000000000",
  52775=>"000000100",
  52776=>"000000001",
  52777=>"001001101",
  52778=>"110000000",
  52779=>"111111000",
  52780=>"111110100",
  52781=>"110000010",
  52782=>"000000000",
  52783=>"111110111",
  52784=>"000001001",
  52785=>"000111111",
  52786=>"110000000",
  52787=>"111111000",
  52788=>"000000001",
  52789=>"000111111",
  52790=>"111111100",
  52791=>"001111000",
  52792=>"001000111",
  52793=>"000000001",
  52794=>"111011000",
  52795=>"111100000",
  52796=>"000000000",
  52797=>"101111111",
  52798=>"111111001",
  52799=>"000010010",
  52800=>"111001100",
  52801=>"000000101",
  52802=>"011110110",
  52803=>"101000111",
  52804=>"111000001",
  52805=>"011111110",
  52806=>"000000111",
  52807=>"000000111",
  52808=>"000001011",
  52809=>"111111111",
  52810=>"111111001",
  52811=>"111111111",
  52812=>"000000110",
  52813=>"000000001",
  52814=>"111111000",
  52815=>"111011111",
  52816=>"000000000",
  52817=>"001100101",
  52818=>"100000000",
  52819=>"111111001",
  52820=>"111111011",
  52821=>"000000000",
  52822=>"111001111",
  52823=>"111111111",
  52824=>"001000000",
  52825=>"101111111",
  52826=>"010000101",
  52827=>"100100000",
  52828=>"000000001",
  52829=>"000000000",
  52830=>"000000000",
  52831=>"111111000",
  52832=>"010000000",
  52833=>"000101111",
  52834=>"111111111",
  52835=>"100100111",
  52836=>"011000000",
  52837=>"111111111",
  52838=>"000000000",
  52839=>"000001001",
  52840=>"000000101",
  52841=>"110111111",
  52842=>"000000000",
  52843=>"111111000",
  52844=>"000000000",
  52845=>"111111000",
  52846=>"111000111",
  52847=>"100111111",
  52848=>"111000000",
  52849=>"000000000",
  52850=>"000010111",
  52851=>"011001111",
  52852=>"110000000",
  52853=>"111111000",
  52854=>"000000000",
  52855=>"111111011",
  52856=>"000000000",
  52857=>"111110110",
  52858=>"111111000",
  52859=>"000000001",
  52860=>"000000000",
  52861=>"000000111",
  52862=>"111001000",
  52863=>"111111111",
  52864=>"000000011",
  52865=>"100000111",
  52866=>"100000000",
  52867=>"111101000",
  52868=>"000000001",
  52869=>"000001111",
  52870=>"000111111",
  52871=>"110000000",
  52872=>"100000000",
  52873=>"111111111",
  52874=>"011111011",
  52875=>"000111111",
  52876=>"111111000",
  52877=>"111011000",
  52878=>"100100101",
  52879=>"111111111",
  52880=>"000111111",
  52881=>"000000000",
  52882=>"000001111",
  52883=>"111111001",
  52884=>"001111111",
  52885=>"111111000",
  52886=>"111000100",
  52887=>"111000111",
  52888=>"000000000",
  52889=>"111111111",
  52890=>"000000111",
  52891=>"000000000",
  52892=>"001110000",
  52893=>"001000000",
  52894=>"110100111",
  52895=>"000000000",
  52896=>"111101100",
  52897=>"111111111",
  52898=>"111000000",
  52899=>"000000000",
  52900=>"000010000",
  52901=>"000000100",
  52902=>"111111110",
  52903=>"100000001",
  52904=>"000000000",
  52905=>"000000000",
  52906=>"111000000",
  52907=>"000000000",
  52908=>"100000110",
  52909=>"111110000",
  52910=>"011000000",
  52911=>"111000001",
  52912=>"010111010",
  52913=>"000010111",
  52914=>"011101000",
  52915=>"111101000",
  52916=>"000000111",
  52917=>"000001111",
  52918=>"000000011",
  52919=>"111000000",
  52920=>"000000100",
  52921=>"111000010",
  52922=>"000000000",
  52923=>"100111111",
  52924=>"000000100",
  52925=>"111111111",
  52926=>"000000111",
  52927=>"111001001",
  52928=>"101000000",
  52929=>"000000000",
  52930=>"000000001",
  52931=>"000001111",
  52932=>"001111111",
  52933=>"000000000",
  52934=>"000000000",
  52935=>"011001000",
  52936=>"000100110",
  52937=>"100000000",
  52938=>"111011001",
  52939=>"000000111",
  52940=>"100100100",
  52941=>"111111101",
  52942=>"001101111",
  52943=>"000110111",
  52944=>"001000000",
  52945=>"000000000",
  52946=>"100101001",
  52947=>"000000000",
  52948=>"000000000",
  52949=>"111000000",
  52950=>"000000000",
  52951=>"000000000",
  52952=>"111111001",
  52953=>"111110111",
  52954=>"101000111",
  52955=>"111101000",
  52956=>"000000000",
  52957=>"111100000",
  52958=>"010111011",
  52959=>"001000111",
  52960=>"111000000",
  52961=>"001001111",
  52962=>"000001000",
  52963=>"111001000",
  52964=>"101111111",
  52965=>"011001000",
  52966=>"110110111",
  52967=>"100000111",
  52968=>"110111000",
  52969=>"000111111",
  52970=>"001000000",
  52971=>"111000101",
  52972=>"111000000",
  52973=>"000110000",
  52974=>"000101111",
  52975=>"111000000",
  52976=>"111111011",
  52977=>"111010000",
  52978=>"111001101",
  52979=>"011100000",
  52980=>"000010011",
  52981=>"111111000",
  52982=>"110000000",
  52983=>"111111111",
  52984=>"111111111",
  52985=>"100110110",
  52986=>"111010000",
  52987=>"111111111",
  52988=>"100000001",
  52989=>"111111110",
  52990=>"000100111",
  52991=>"001001111",
  52992=>"100111010",
  52993=>"001000011",
  52994=>"111111111",
  52995=>"111111111",
  52996=>"111111000",
  52997=>"111010000",
  52998=>"111010000",
  52999=>"111111111",
  53000=>"111111110",
  53001=>"000111111",
  53002=>"000000000",
  53003=>"000001111",
  53004=>"100100110",
  53005=>"000111010",
  53006=>"000000000",
  53007=>"110111111",
  53008=>"000000000",
  53009=>"001000011",
  53010=>"000000000",
  53011=>"000000001",
  53012=>"100111111",
  53013=>"111100001",
  53014=>"001000000",
  53015=>"000111111",
  53016=>"111000100",
  53017=>"111000010",
  53018=>"000000110",
  53019=>"000000000",
  53020=>"111111111",
  53021=>"001000001",
  53022=>"101111111",
  53023=>"000000000",
  53024=>"111111001",
  53025=>"000000111",
  53026=>"111111000",
  53027=>"000000111",
  53028=>"000000101",
  53029=>"000000001",
  53030=>"000110000",
  53031=>"111111111",
  53032=>"000000000",
  53033=>"111111101",
  53034=>"000000001",
  53035=>"000101001",
  53036=>"111111000",
  53037=>"000000111",
  53038=>"000010000",
  53039=>"111010000",
  53040=>"011000001",
  53041=>"111111111",
  53042=>"111110010",
  53043=>"111111000",
  53044=>"111001001",
  53045=>"111100000",
  53046=>"111000000",
  53047=>"001001000",
  53048=>"000000001",
  53049=>"111011111",
  53050=>"000000111",
  53051=>"111111111",
  53052=>"000000110",
  53053=>"000000000",
  53054=>"110010000",
  53055=>"000000111",
  53056=>"001001111",
  53057=>"000001101",
  53058=>"111111000",
  53059=>"000000111",
  53060=>"000000000",
  53061=>"000000111",
  53062=>"000000000",
  53063=>"111111111",
  53064=>"000000000",
  53065=>"000000000",
  53066=>"111111111",
  53067=>"110000000",
  53068=>"110111000",
  53069=>"111111110",
  53070=>"000000000",
  53071=>"000000000",
  53072=>"110110100",
  53073=>"000100111",
  53074=>"101110111",
  53075=>"101001111",
  53076=>"000011111",
  53077=>"001011001",
  53078=>"111111111",
  53079=>"111101111",
  53080=>"100000000",
  53081=>"000000001",
  53082=>"100100000",
  53083=>"111001000",
  53084=>"101000001",
  53085=>"000001111",
  53086=>"000001000",
  53087=>"010010000",
  53088=>"000000000",
  53089=>"000001111",
  53090=>"111111100",
  53091=>"000000011",
  53092=>"010011111",
  53093=>"000000001",
  53094=>"000000000",
  53095=>"000000000",
  53096=>"111000000",
  53097=>"111111111",
  53098=>"111000100",
  53099=>"111111111",
  53100=>"111111111",
  53101=>"111111111",
  53102=>"000101000",
  53103=>"000000111",
  53104=>"000111111",
  53105=>"000000111",
  53106=>"000000000",
  53107=>"100000010",
  53108=>"111111001",
  53109=>"000000000",
  53110=>"000011000",
  53111=>"110000000",
  53112=>"111000000",
  53113=>"100000001",
  53114=>"000000000",
  53115=>"111010000",
  53116=>"011010010",
  53117=>"111000101",
  53118=>"000111111",
  53119=>"010111111",
  53120=>"010000000",
  53121=>"111111110",
  53122=>"110111111",
  53123=>"111111111",
  53124=>"111100111",
  53125=>"110111111",
  53126=>"111100111",
  53127=>"000100101",
  53128=>"111000000",
  53129=>"111000011",
  53130=>"111111001",
  53131=>"000010111",
  53132=>"111111111",
  53133=>"111111110",
  53134=>"111010000",
  53135=>"000000000",
  53136=>"000000000",
  53137=>"111000000",
  53138=>"001000101",
  53139=>"000000000",
  53140=>"111111101",
  53141=>"000000000",
  53142=>"000001111",
  53143=>"110111101",
  53144=>"111111011",
  53145=>"000000000",
  53146=>"111111000",
  53147=>"111111111",
  53148=>"111000111",
  53149=>"111111000",
  53150=>"110100000",
  53151=>"000000100",
  53152=>"101001000",
  53153=>"000000011",
  53154=>"001111111",
  53155=>"000111110",
  53156=>"000101111",
  53157=>"111001011",
  53158=>"000010000",
  53159=>"000000001",
  53160=>"000001001",
  53161=>"111111101",
  53162=>"001111111",
  53163=>"000011010",
  53164=>"000000000",
  53165=>"000000101",
  53166=>"000000110",
  53167=>"010110110",
  53168=>"111000000",
  53169=>"000000000",
  53170=>"111000000",
  53171=>"000000001",
  53172=>"000000100",
  53173=>"111011111",
  53174=>"111111111",
  53175=>"000100111",
  53176=>"000000111",
  53177=>"110111100",
  53178=>"001000001",
  53179=>"000000000",
  53180=>"111111110",
  53181=>"111111111",
  53182=>"000000001",
  53183=>"001000000",
  53184=>"000000000",
  53185=>"100000000",
  53186=>"111100000",
  53187=>"000000000",
  53188=>"000000000",
  53189=>"000000111",
  53190=>"000000001",
  53191=>"000000000",
  53192=>"000000000",
  53193=>"111000000",
  53194=>"111111011",
  53195=>"111000000",
  53196=>"011000000",
  53197=>"100000110",
  53198=>"111111000",
  53199=>"111111111",
  53200=>"000000000",
  53201=>"110011000",
  53202=>"001111100",
  53203=>"001000111",
  53204=>"111111110",
  53205=>"000000001",
  53206=>"000001001",
  53207=>"110111011",
  53208=>"000000000",
  53209=>"000001001",
  53210=>"000110000",
  53211=>"111100000",
  53212=>"111111111",
  53213=>"111111111",
  53214=>"000000000",
  53215=>"100000101",
  53216=>"111101100",
  53217=>"001001001",
  53218=>"101111111",
  53219=>"001101111",
  53220=>"000011111",
  53221=>"011011011",
  53222=>"000111000",
  53223=>"111000000",
  53224=>"111000000",
  53225=>"100000101",
  53226=>"100000010",
  53227=>"000000001",
  53228=>"100000000",
  53229=>"111111111",
  53230=>"000001111",
  53231=>"000010011",
  53232=>"110000110",
  53233=>"001001111",
  53234=>"111011011",
  53235=>"000001101",
  53236=>"111111000",
  53237=>"111010000",
  53238=>"000001111",
  53239=>"000000001",
  53240=>"000011111",
  53241=>"110000000",
  53242=>"001001011",
  53243=>"000000110",
  53244=>"111001111",
  53245=>"000000100",
  53246=>"000000000",
  53247=>"111111110",
  53248=>"111111000",
  53249=>"111111111",
  53250=>"000111111",
  53251=>"000110110",
  53252=>"110110000",
  53253=>"101001001",
  53254=>"110111011",
  53255=>"000000111",
  53256=>"111111000",
  53257=>"111000000",
  53258=>"000000100",
  53259=>"000000000",
  53260=>"000110000",
  53261=>"000000000",
  53262=>"001111000",
  53263=>"000000000",
  53264=>"001001001",
  53265=>"110110000",
  53266=>"000111100",
  53267=>"110111111",
  53268=>"110100111",
  53269=>"000111111",
  53270=>"000000001",
  53271=>"111100000",
  53272=>"000110000",
  53273=>"000000111",
  53274=>"101101111",
  53275=>"110000000",
  53276=>"111111100",
  53277=>"000000111",
  53278=>"111000010",
  53279=>"001001111",
  53280=>"101011000",
  53281=>"101000100",
  53282=>"100000000",
  53283=>"000000111",
  53284=>"010111111",
  53285=>"101000101",
  53286=>"000000000",
  53287=>"000000000",
  53288=>"111111000",
  53289=>"100111111",
  53290=>"001000111",
  53291=>"111111101",
  53292=>"000000000",
  53293=>"111111000",
  53294=>"011011111",
  53295=>"110111111",
  53296=>"001001000",
  53297=>"000000000",
  53298=>"111111111",
  53299=>"000000000",
  53300=>"011111010",
  53301=>"001000011",
  53302=>"111111111",
  53303=>"111000001",
  53304=>"101110000",
  53305=>"111010110",
  53306=>"011000111",
  53307=>"001011000",
  53308=>"101111101",
  53309=>"111110000",
  53310=>"000000110",
  53311=>"100100111",
  53312=>"011011111",
  53313=>"010010000",
  53314=>"000010110",
  53315=>"000011111",
  53316=>"001101101",
  53317=>"000000101",
  53318=>"111111001",
  53319=>"111110111",
  53320=>"101101011",
  53321=>"110111111",
  53322=>"111111001",
  53323=>"000000000",
  53324=>"001001111",
  53325=>"000000110",
  53326=>"111110010",
  53327=>"000001001",
  53328=>"000000010",
  53329=>"111000000",
  53330=>"001000111",
  53331=>"000100000",
  53332=>"000000000",
  53333=>"000000111",
  53334=>"101000101",
  53335=>"101001000",
  53336=>"000100111",
  53337=>"000000111",
  53338=>"110110000",
  53339=>"111011010",
  53340=>"000000100",
  53341=>"111010000",
  53342=>"000000001",
  53343=>"011000000",
  53344=>"111110111",
  53345=>"000000111",
  53346=>"101000001",
  53347=>"001000000",
  53348=>"110111000",
  53349=>"101111111",
  53350=>"111111000",
  53351=>"111111111",
  53352=>"000100001",
  53353=>"111111111",
  53354=>"111000000",
  53355=>"000000010",
  53356=>"110000000",
  53357=>"111111000",
  53358=>"111111111",
  53359=>"000111000",
  53360=>"111111111",
  53361=>"000000000",
  53362=>"000000000",
  53363=>"111111100",
  53364=>"000001111",
  53365=>"000111111",
  53366=>"000101111",
  53367=>"000110000",
  53368=>"111000000",
  53369=>"000000111",
  53370=>"111000000",
  53371=>"010111111",
  53372=>"100000000",
  53373=>"100110110",
  53374=>"011000101",
  53375=>"000100111",
  53376=>"101001000",
  53377=>"001111111",
  53378=>"111111001",
  53379=>"110111110",
  53380=>"111111111",
  53381=>"111000000",
  53382=>"001000000",
  53383=>"111101000",
  53384=>"000111111",
  53385=>"100000000",
  53386=>"000000000",
  53387=>"000000111",
  53388=>"001000111",
  53389=>"000000111",
  53390=>"011111011",
  53391=>"111111010",
  53392=>"001000100",
  53393=>"111111000",
  53394=>"010000011",
  53395=>"110110111",
  53396=>"111111001",
  53397=>"001011000",
  53398=>"111010000",
  53399=>"001011111",
  53400=>"101101111",
  53401=>"111111001",
  53402=>"100100000",
  53403=>"000011111",
  53404=>"111111111",
  53405=>"000000011",
  53406=>"111010000",
  53407=>"110100010",
  53408=>"111111000",
  53409=>"111100111",
  53410=>"000000101",
  53411=>"111111010",
  53412=>"000110100",
  53413=>"001000001",
  53414=>"111111111",
  53415=>"000001011",
  53416=>"000000000",
  53417=>"000000111",
  53418=>"001000101",
  53419=>"000000000",
  53420=>"101000000",
  53421=>"011111100",
  53422=>"000111111",
  53423=>"000111111",
  53424=>"111000111",
  53425=>"000100110",
  53426=>"110111010",
  53427=>"111001000",
  53428=>"000000110",
  53429=>"001111100",
  53430=>"100111100",
  53431=>"000000000",
  53432=>"001000101",
  53433=>"110111111",
  53434=>"111000000",
  53435=>"001001111",
  53436=>"111111110",
  53437=>"111000000",
  53438=>"000010101",
  53439=>"000000011",
  53440=>"111111111",
  53441=>"001011111",
  53442=>"111001111",
  53443=>"111001101",
  53444=>"000000000",
  53445=>"001001001",
  53446=>"111111110",
  53447=>"001101000",
  53448=>"111110000",
  53449=>"000001000",
  53450=>"000000000",
  53451=>"101100111",
  53452=>"000000001",
  53453=>"110110000",
  53454=>"000000000",
  53455=>"000000000",
  53456=>"000110110",
  53457=>"001000000",
  53458=>"110000000",
  53459=>"001000111",
  53460=>"100000000",
  53461=>"000000000",
  53462=>"110111000",
  53463=>"000001111",
  53464=>"001000101",
  53465=>"111111111",
  53466=>"111000000",
  53467=>"111000000",
  53468=>"110000000",
  53469=>"000000111",
  53470=>"000111011",
  53471=>"101101101",
  53472=>"000000000",
  53473=>"000110111",
  53474=>"111111111",
  53475=>"000100111",
  53476=>"011111111",
  53477=>"110111000",
  53478=>"111111111",
  53479=>"000000000",
  53480=>"000101001",
  53481=>"111111000",
  53482=>"111111111",
  53483=>"111111101",
  53484=>"111111011",
  53485=>"000010000",
  53486=>"111010001",
  53487=>"111111111",
  53488=>"000000111",
  53489=>"000000111",
  53490=>"000000000",
  53491=>"000000101",
  53492=>"001000101",
  53493=>"110101101",
  53494=>"011111000",
  53495=>"111011000",
  53496=>"111111111",
  53497=>"111111111",
  53498=>"001000111",
  53499=>"110000000",
  53500=>"000010000",
  53501=>"111111110",
  53502=>"111111000",
  53503=>"000000000",
  53504=>"110000000",
  53505=>"111111110",
  53506=>"111111111",
  53507=>"000100000",
  53508=>"111100100",
  53509=>"100100000",
  53510=>"111111111",
  53511=>"100110111",
  53512=>"111111000",
  53513=>"111010000",
  53514=>"000100000",
  53515=>"111111000",
  53516=>"111000111",
  53517=>"001000001",
  53518=>"001000000",
  53519=>"110000000",
  53520=>"100110000",
  53521=>"000100111",
  53522=>"000000111",
  53523=>"000000000",
  53524=>"000111111",
  53525=>"010111000",
  53526=>"111111111",
  53527=>"111111000",
  53528=>"000000110",
  53529=>"000000000",
  53530=>"111010000",
  53531=>"000001111",
  53532=>"110111110",
  53533=>"000010011",
  53534=>"000000111",
  53535=>"000111111",
  53536=>"000011000",
  53537=>"110111011",
  53538=>"000111010",
  53539=>"110000110",
  53540=>"111110100",
  53541=>"110100000",
  53542=>"000000100",
  53543=>"111111000",
  53544=>"110111111",
  53545=>"101111111",
  53546=>"000000000",
  53547=>"000000111",
  53548=>"111100000",
  53549=>"000101111",
  53550=>"011000000",
  53551=>"000000000",
  53552=>"111011111",
  53553=>"000000000",
  53554=>"111111010",
  53555=>"111111010",
  53556=>"000000000",
  53557=>"001010010",
  53558=>"000111111",
  53559=>"001111111",
  53560=>"010010000",
  53561=>"000000111",
  53562=>"000000111",
  53563=>"111011111",
  53564=>"101011001",
  53565=>"000001111",
  53566=>"000001111",
  53567=>"111001000",
  53568=>"001111111",
  53569=>"000100110",
  53570=>"000000111",
  53571=>"000111111",
  53572=>"000001000",
  53573=>"001000100",
  53574=>"000111111",
  53575=>"100001000",
  53576=>"110110000",
  53577=>"100000000",
  53578=>"011001111",
  53579=>"010110111",
  53580=>"000000000",
  53581=>"000000110",
  53582=>"000000111",
  53583=>"111000111",
  53584=>"110010000",
  53585=>"001111011",
  53586=>"111000111",
  53587=>"100000000",
  53588=>"001001000",
  53589=>"011011011",
  53590=>"111011001",
  53591=>"111000000",
  53592=>"111011011",
  53593=>"001111110",
  53594=>"001000000",
  53595=>"000111001",
  53596=>"000000110",
  53597=>"000100110",
  53598=>"110111111",
  53599=>"001001010",
  53600=>"101000101",
  53601=>"001000000",
  53602=>"111001111",
  53603=>"111000000",
  53604=>"111111110",
  53605=>"111111010",
  53606=>"111111000",
  53607=>"110111111",
  53608=>"000000111",
  53609=>"000000011",
  53610=>"000000000",
  53611=>"001011101",
  53612=>"110010000",
  53613=>"101001000",
  53614=>"111000010",
  53615=>"000000000",
  53616=>"111100000",
  53617=>"000000000",
  53618=>"111111111",
  53619=>"111000000",
  53620=>"111001000",
  53621=>"000000000",
  53622=>"000000111",
  53623=>"011000001",
  53624=>"111101000",
  53625=>"111100111",
  53626=>"000000000",
  53627=>"100100011",
  53628=>"000100110",
  53629=>"111000111",
  53630=>"111111110",
  53631=>"000000111",
  53632=>"001110111",
  53633=>"001101001",
  53634=>"001001101",
  53635=>"100110111",
  53636=>"000000000",
  53637=>"011111111",
  53638=>"011011010",
  53639=>"001000000",
  53640=>"110000000",
  53641=>"000000011",
  53642=>"000000001",
  53643=>"111111011",
  53644=>"101101111",
  53645=>"000001111",
  53646=>"111111000",
  53647=>"110111010",
  53648=>"110111110",
  53649=>"000001111",
  53650=>"001000000",
  53651=>"000100000",
  53652=>"111000010",
  53653=>"010010000",
  53654=>"011001100",
  53655=>"110111111",
  53656=>"111111001",
  53657=>"110000000",
  53658=>"111111111",
  53659=>"011000000",
  53660=>"000000000",
  53661=>"000011010",
  53662=>"000000000",
  53663=>"110111111",
  53664=>"000000000",
  53665=>"101110111",
  53666=>"111111000",
  53667=>"000000000",
  53668=>"111111111",
  53669=>"001001111",
  53670=>"111111000",
  53671=>"000000011",
  53672=>"111111100",
  53673=>"000111111",
  53674=>"000000000",
  53675=>"100110111",
  53676=>"001111111",
  53677=>"110100001",
  53678=>"111000000",
  53679=>"111101000",
  53680=>"111010101",
  53681=>"000000001",
  53682=>"000000111",
  53683=>"000000111",
  53684=>"001001001",
  53685=>"001111101",
  53686=>"111111010",
  53687=>"110111000",
  53688=>"000000111",
  53689=>"111101110",
  53690=>"101101101",
  53691=>"110111111",
  53692=>"001111111",
  53693=>"111111010",
  53694=>"111111111",
  53695=>"111111001",
  53696=>"000000000",
  53697=>"111111000",
  53698=>"111001010",
  53699=>"111110111",
  53700=>"111000111",
  53701=>"101111111",
  53702=>"000111111",
  53703=>"111101101",
  53704=>"111101111",
  53705=>"100111111",
  53706=>"000000101",
  53707=>"000001111",
  53708=>"001001000",
  53709=>"000011111",
  53710=>"001000100",
  53711=>"111000100",
  53712=>"000110111",
  53713=>"101000111",
  53714=>"111111111",
  53715=>"111111000",
  53716=>"111101111",
  53717=>"110100100",
  53718=>"000011011",
  53719=>"010010000",
  53720=>"100110110",
  53721=>"001001111",
  53722=>"111111111",
  53723=>"111111010",
  53724=>"000000000",
  53725=>"100000000",
  53726=>"001000000",
  53727=>"111111111",
  53728=>"000001000",
  53729=>"110111111",
  53730=>"110110000",
  53731=>"000010100",
  53732=>"100000001",
  53733=>"111111100",
  53734=>"110111011",
  53735=>"000000011",
  53736=>"110101000",
  53737=>"111001000",
  53738=>"000110010",
  53739=>"111111011",
  53740=>"101111111",
  53741=>"110111000",
  53742=>"100000001",
  53743=>"111110000",
  53744=>"111110000",
  53745=>"111010000",
  53746=>"001000111",
  53747=>"111110000",
  53748=>"011111011",
  53749=>"000000000",
  53750=>"111111111",
  53751=>"111111111",
  53752=>"011111111",
  53753=>"111111001",
  53754=>"110111000",
  53755=>"101111100",
  53756=>"000101001",
  53757=>"111111111",
  53758=>"000000000",
  53759=>"101001000",
  53760=>"111111111",
  53761=>"011000000",
  53762=>"111000000",
  53763=>"111111111",
  53764=>"000000000",
  53765=>"001000000",
  53766=>"111101111",
  53767=>"001000101",
  53768=>"111111000",
  53769=>"111000000",
  53770=>"000000110",
  53771=>"000000000",
  53772=>"111110110",
  53773=>"010000000",
  53774=>"011111000",
  53775=>"000100000",
  53776=>"010111111",
  53777=>"000000011",
  53778=>"011001001",
  53779=>"000010010",
  53780=>"000000000",
  53781=>"111111011",
  53782=>"111111111",
  53783=>"001011011",
  53784=>"111111111",
  53785=>"001001111",
  53786=>"110111111",
  53787=>"000100000",
  53788=>"100100110",
  53789=>"111101110",
  53790=>"000000000",
  53791=>"110000000",
  53792=>"000000001",
  53793=>"001001000",
  53794=>"111111111",
  53795=>"111111111",
  53796=>"011011001",
  53797=>"011110000",
  53798=>"000000000",
  53799=>"110000000",
  53800=>"011011000",
  53801=>"000000100",
  53802=>"000111111",
  53803=>"000000000",
  53804=>"000100111",
  53805=>"000000000",
  53806=>"000011111",
  53807=>"010000000",
  53808=>"111000000",
  53809=>"000000000",
  53810=>"111111011",
  53811=>"000000000",
  53812=>"011011001",
  53813=>"001001001",
  53814=>"000111111",
  53815=>"100101000",
  53816=>"110111000",
  53817=>"000000110",
  53818=>"111111000",
  53819=>"111111111",
  53820=>"000000111",
  53821=>"000110000",
  53822=>"101101111",
  53823=>"111111111",
  53824=>"000010000",
  53825=>"000000000",
  53826=>"110000111",
  53827=>"000110111",
  53828=>"110111011",
  53829=>"011011110",
  53830=>"110000110",
  53831=>"000000000",
  53832=>"100101000",
  53833=>"111100110",
  53834=>"001000000",
  53835=>"000000001",
  53836=>"000110110",
  53837=>"000000011",
  53838=>"111110110",
  53839=>"000000011",
  53840=>"011111111",
  53841=>"111111111",
  53842=>"000000000",
  53843=>"100110011",
  53844=>"111101001",
  53845=>"111001100",
  53846=>"100100000",
  53847=>"111111111",
  53848=>"000000000",
  53849=>"101101100",
  53850=>"111111100",
  53851=>"100110110",
  53852=>"100000000",
  53853=>"111111000",
  53854=>"000000000",
  53855=>"000011101",
  53856=>"000000000",
  53857=>"111000100",
  53858=>"000000000",
  53859=>"000000001",
  53860=>"001101011",
  53861=>"110000011",
  53862=>"000000110",
  53863=>"111111111",
  53864=>"000000100",
  53865=>"000000010",
  53866=>"000000110",
  53867=>"111111010",
  53868=>"110110111",
  53869=>"111101111",
  53870=>"000000000",
  53871=>"000000000",
  53872=>"001000000",
  53873=>"000101000",
  53874=>"000000000",
  53875=>"000000000",
  53876=>"111111111",
  53877=>"001000000",
  53878=>"111111111",
  53879=>"111111111",
  53880=>"111111111",
  53881=>"011001110",
  53882=>"001000000",
  53883=>"000111101",
  53884=>"110000000",
  53885=>"000000000",
  53886=>"000000000",
  53887=>"000111111",
  53888=>"111111110",
  53889=>"000000000",
  53890=>"111111111",
  53891=>"000000101",
  53892=>"000100000",
  53893=>"100101011",
  53894=>"001101111",
  53895=>"101000000",
  53896=>"000000000",
  53897=>"111111111",
  53898=>"110000111",
  53899=>"111001000",
  53900=>"111001111",
  53901=>"101111111",
  53902=>"000100000",
  53903=>"111111111",
  53904=>"111000000",
  53905=>"000000000",
  53906=>"000000000",
  53907=>"111111110",
  53908=>"000000100",
  53909=>"000000000",
  53910=>"000000000",
  53911=>"111111000",
  53912=>"111111111",
  53913=>"001111000",
  53914=>"000100101",
  53915=>"111000000",
  53916=>"000111111",
  53917=>"001001001",
  53918=>"101101000",
  53919=>"111100100",
  53920=>"011111111",
  53921=>"111110111",
  53922=>"000000000",
  53923=>"000000000",
  53924=>"010000000",
  53925=>"000000000",
  53926=>"110110110",
  53927=>"000000000",
  53928=>"000000000",
  53929=>"111110110",
  53930=>"001001101",
  53931=>"000001111",
  53932=>"111111111",
  53933=>"000000000",
  53934=>"001100110",
  53935=>"000110000",
  53936=>"111111111",
  53937=>"111001011",
  53938=>"000011000",
  53939=>"110111111",
  53940=>"111110111",
  53941=>"111111111",
  53942=>"111111010",
  53943=>"110100000",
  53944=>"000000101",
  53945=>"111111111",
  53946=>"000010110",
  53947=>"000000100",
  53948=>"100100110",
  53949=>"000000100",
  53950=>"011011011",
  53951=>"111000000",
  53952=>"111000110",
  53953=>"111111111",
  53954=>"011001000",
  53955=>"111110000",
  53956=>"111111111",
  53957=>"000000100",
  53958=>"111111111",
  53959=>"111111111",
  53960=>"011001001",
  53961=>"111111111",
  53962=>"111110000",
  53963=>"000000100",
  53964=>"111110000",
  53965=>"000000000",
  53966=>"000000001",
  53967=>"001001111",
  53968=>"011000000",
  53969=>"110000000",
  53970=>"000000000",
  53971=>"000000000",
  53972=>"001000000",
  53973=>"000000000",
  53974=>"000000011",
  53975=>"100000101",
  53976=>"111111111",
  53977=>"010011000",
  53978=>"101111110",
  53979=>"110111111",
  53980=>"110110000",
  53981=>"111110111",
  53982=>"000000000",
  53983=>"000110110",
  53984=>"100100100",
  53985=>"000000000",
  53986=>"111111111",
  53987=>"100000101",
  53988=>"111101101",
  53989=>"011011011",
  53990=>"000100111",
  53991=>"111000000",
  53992=>"111111111",
  53993=>"111111011",
  53994=>"111111111",
  53995=>"000100111",
  53996=>"111111000",
  53997=>"000000010",
  53998=>"000000100",
  53999=>"111000000",
  54000=>"111110100",
  54001=>"000000000",
  54002=>"111110110",
  54003=>"110111101",
  54004=>"111101111",
  54005=>"000110110",
  54006=>"111111111",
  54007=>"111111000",
  54008=>"110000000",
  54009=>"111111001",
  54010=>"000010000",
  54011=>"110111111",
  54012=>"111001000",
  54013=>"111000101",
  54014=>"000000000",
  54015=>"001111001",
  54016=>"111111111",
  54017=>"111111111",
  54018=>"011001000",
  54019=>"111111110",
  54020=>"111111111",
  54021=>"111111100",
  54022=>"000001001",
  54023=>"110111111",
  54024=>"111101111",
  54025=>"000000000",
  54026=>"111011111",
  54027=>"000001001",
  54028=>"011011000",
  54029=>"000000000",
  54030=>"011011000",
  54031=>"000000000",
  54032=>"000000000",
  54033=>"000000100",
  54034=>"000000000",
  54035=>"111111111",
  54036=>"011111100",
  54037=>"111111000",
  54038=>"000010011",
  54039=>"000000000",
  54040=>"011011111",
  54041=>"111011000",
  54042=>"000000000",
  54043=>"011111110",
  54044=>"000011011",
  54045=>"010111111",
  54046=>"111111111",
  54047=>"101011111",
  54048=>"111111111",
  54049=>"000010000",
  54050=>"111111111",
  54051=>"000000000",
  54052=>"000000100",
  54053=>"111110100",
  54054=>"111111111",
  54055=>"000000011",
  54056=>"111001101",
  54057=>"111111101",
  54058=>"011100000",
  54059=>"000000000",
  54060=>"111111000",
  54061=>"111111111",
  54062=>"000000000",
  54063=>"000000011",
  54064=>"111111001",
  54065=>"000000000",
  54066=>"111111111",
  54067=>"000000000",
  54068=>"000000000",
  54069=>"000100100",
  54070=>"111111111",
  54071=>"111111111",
  54072=>"000000000",
  54073=>"000000000",
  54074=>"000000111",
  54075=>"000000000",
  54076=>"100111101",
  54077=>"000010100",
  54078=>"111000100",
  54079=>"000000000",
  54080=>"100000000",
  54081=>"000000000",
  54082=>"000000000",
  54083=>"001000000",
  54084=>"001001000",
  54085=>"000000001",
  54086=>"011000000",
  54087=>"110110111",
  54088=>"100100000",
  54089=>"000110010",
  54090=>"000000000",
  54091=>"011010001",
  54092=>"000011011",
  54093=>"111011111",
  54094=>"000100110",
  54095=>"111111011",
  54096=>"000000000",
  54097=>"111111100",
  54098=>"000001001",
  54099=>"000010111",
  54100=>"001000000",
  54101=>"001011011",
  54102=>"111111100",
  54103=>"100000000",
  54104=>"111000000",
  54105=>"000111111",
  54106=>"100100000",
  54107=>"111101110",
  54108=>"000000100",
  54109=>"110110010",
  54110=>"110111000",
  54111=>"000011000",
  54112=>"000000100",
  54113=>"000000011",
  54114=>"100110100",
  54115=>"111111111",
  54116=>"001001001",
  54117=>"110111111",
  54118=>"111000000",
  54119=>"001111110",
  54120=>"001011000",
  54121=>"111101000",
  54122=>"000000111",
  54123=>"100111111",
  54124=>"000000001",
  54125=>"000000100",
  54126=>"001000000",
  54127=>"000000000",
  54128=>"110111100",
  54129=>"000000000",
  54130=>"001001101",
  54131=>"100100001",
  54132=>"110111111",
  54133=>"000000000",
  54134=>"000000000",
  54135=>"000000000",
  54136=>"000000000",
  54137=>"000000111",
  54138=>"111000000",
  54139=>"000000000",
  54140=>"011000000",
  54141=>"001001001",
  54142=>"111111000",
  54143=>"000000000",
  54144=>"111111111",
  54145=>"000000000",
  54146=>"110111001",
  54147=>"111111111",
  54148=>"111111111",
  54149=>"001001001",
  54150=>"000000011",
  54151=>"000100100",
  54152=>"000000000",
  54153=>"001111111",
  54154=>"000100000",
  54155=>"000011010",
  54156=>"111111111",
  54157=>"000000000",
  54158=>"110110000",
  54159=>"011111111",
  54160=>"000100000",
  54161=>"000001001",
  54162=>"000010000",
  54163=>"111001000",
  54164=>"010111000",
  54165=>"001000001",
  54166=>"100100000",
  54167=>"000000000",
  54168=>"110010000",
  54169=>"000000000",
  54170=>"000111000",
  54171=>"000100111",
  54172=>"010001101",
  54173=>"010011010",
  54174=>"011011011",
  54175=>"111111111",
  54176=>"000000000",
  54177=>"000000000",
  54178=>"110000000",
  54179=>"110111111",
  54180=>"111111111",
  54181=>"010111010",
  54182=>"000000000",
  54183=>"011110111",
  54184=>"111110111",
  54185=>"000000000",
  54186=>"110000000",
  54187=>"011010011",
  54188=>"111111111",
  54189=>"000000000",
  54190=>"000010010",
  54191=>"000100100",
  54192=>"011111011",
  54193=>"001101111",
  54194=>"000111111",
  54195=>"000010000",
  54196=>"111111111",
  54197=>"000000000",
  54198=>"001000011",
  54199=>"011011000",
  54200=>"000000111",
  54201=>"111111111",
  54202=>"000000000",
  54203=>"000100111",
  54204=>"111111111",
  54205=>"111111111",
  54206=>"111111111",
  54207=>"000000000",
  54208=>"000000000",
  54209=>"100110110",
  54210=>"000000000",
  54211=>"000101000",
  54212=>"000110011",
  54213=>"011000000",
  54214=>"100111000",
  54215=>"110111110",
  54216=>"000000000",
  54217=>"111111100",
  54218=>"000000000",
  54219=>"000110011",
  54220=>"100000000",
  54221=>"111000000",
  54222=>"001111111",
  54223=>"100100001",
  54224=>"110111111",
  54225=>"100100000",
  54226=>"000000000",
  54227=>"111101101",
  54228=>"111111011",
  54229=>"010111011",
  54230=>"010110110",
  54231=>"100100000",
  54232=>"111111111",
  54233=>"011011000",
  54234=>"110111111",
  54235=>"111111110",
  54236=>"101001110",
  54237=>"100111111",
  54238=>"111000000",
  54239=>"111111111",
  54240=>"000000010",
  54241=>"111000100",
  54242=>"111111111",
  54243=>"111001000",
  54244=>"000000000",
  54245=>"111111001",
  54246=>"010000000",
  54247=>"000000000",
  54248=>"111111111",
  54249=>"111001001",
  54250=>"000000111",
  54251=>"000000000",
  54252=>"000000011",
  54253=>"000000010",
  54254=>"111111111",
  54255=>"111111111",
  54256=>"000000000",
  54257=>"001000100",
  54258=>"111111111",
  54259=>"000000000",
  54260=>"110111111",
  54261=>"011011000",
  54262=>"111111000",
  54263=>"000000110",
  54264=>"111111011",
  54265=>"000000000",
  54266=>"000100111",
  54267=>"000000000",
  54268=>"111111111",
  54269=>"000000000",
  54270=>"000000001",
  54271=>"101000000",
  54272=>"111001000",
  54273=>"001000000",
  54274=>"000000000",
  54275=>"000000000",
  54276=>"001111111",
  54277=>"111011111",
  54278=>"101000000",
  54279=>"111111111",
  54280=>"111111111",
  54281=>"101000000",
  54282=>"110011110",
  54283=>"001001001",
  54284=>"000100101",
  54285=>"001000100",
  54286=>"111111111",
  54287=>"111111111",
  54288=>"111111111",
  54289=>"111111010",
  54290=>"111111000",
  54291=>"111111111",
  54292=>"111111111",
  54293=>"000001010",
  54294=>"000000010",
  54295=>"111111000",
  54296=>"000001111",
  54297=>"011111100",
  54298=>"000000000",
  54299=>"100000011",
  54300=>"101101101",
  54301=>"111111000",
  54302=>"000000000",
  54303=>"000000001",
  54304=>"111111111",
  54305=>"001001001",
  54306=>"000000000",
  54307=>"000000010",
  54308=>"000000000",
  54309=>"000000111",
  54310=>"101000111",
  54311=>"001111111",
  54312=>"000000000",
  54313=>"000000000",
  54314=>"000000111",
  54315=>"111111011",
  54316=>"111111100",
  54317=>"111111111",
  54318=>"100000011",
  54319=>"111111111",
  54320=>"011110110",
  54321=>"000000000",
  54322=>"001001001",
  54323=>"001111111",
  54324=>"000000000",
  54325=>"001001000",
  54326=>"000000000",
  54327=>"001000000",
  54328=>"011111111",
  54329=>"000010010",
  54330=>"000000000",
  54331=>"000000000",
  54332=>"111101000",
  54333=>"000011111",
  54334=>"011011011",
  54335=>"111001001",
  54336=>"000001000",
  54337=>"100100100",
  54338=>"001000000",
  54339=>"000111000",
  54340=>"000000000",
  54341=>"110111111",
  54342=>"000000111",
  54343=>"111111000",
  54344=>"000000000",
  54345=>"000000011",
  54346=>"000000000",
  54347=>"111111000",
  54348=>"111111100",
  54349=>"011000000",
  54350=>"111110111",
  54351=>"111101000",
  54352=>"000011010",
  54353=>"000000000",
  54354=>"000000111",
  54355=>"111100000",
  54356=>"000001111",
  54357=>"000111111",
  54358=>"000000000",
  54359=>"000000000",
  54360=>"000000000",
  54361=>"111000111",
  54362=>"111111111",
  54363=>"110110111",
  54364=>"001001111",
  54365=>"100100000",
  54366=>"101101101",
  54367=>"000000000",
  54368=>"000000111",
  54369=>"111111110",
  54370=>"000011001",
  54371=>"100000111",
  54372=>"000100111",
  54373=>"111111111",
  54374=>"111111111",
  54375=>"111111100",
  54376=>"000101001",
  54377=>"000000111",
  54378=>"111010110",
  54379=>"000000001",
  54380=>"111100100",
  54381=>"001001000",
  54382=>"000110110",
  54383=>"000000000",
  54384=>"111001000",
  54385=>"000010000",
  54386=>"011111111",
  54387=>"001001001",
  54388=>"001000000",
  54389=>"111111111",
  54390=>"111000000",
  54391=>"000111111",
  54392=>"111111000",
  54393=>"111111111",
  54394=>"100000010",
  54395=>"010000000",
  54396=>"111111000",
  54397=>"011111111",
  54398=>"111111111",
  54399=>"000000000",
  54400=>"000000000",
  54401=>"101111100",
  54402=>"000000111",
  54403=>"011011001",
  54404=>"000000111",
  54405=>"000001111",
  54406=>"100110010",
  54407=>"111111000",
  54408=>"000111000",
  54409=>"000000011",
  54410=>"000000110",
  54411=>"110000000",
  54412=>"001011011",
  54413=>"000000000",
  54414=>"101100100",
  54415=>"000100110",
  54416=>"000000000",
  54417=>"000000100",
  54418=>"111110000",
  54419=>"000000000",
  54420=>"111111110",
  54421=>"001000110",
  54422=>"000000000",
  54423=>"111101101",
  54424=>"001101110",
  54425=>"000110100",
  54426=>"001111110",
  54427=>"110100000",
  54428=>"100100000",
  54429=>"110000111",
  54430=>"000100111",
  54431=>"000000001",
  54432=>"110110000",
  54433=>"000000000",
  54434=>"000000111",
  54435=>"111111111",
  54436=>"001111100",
  54437=>"001001000",
  54438=>"001000000",
  54439=>"000000000",
  54440=>"111111111",
  54441=>"000000000",
  54442=>"111111110",
  54443=>"101101101",
  54444=>"000000110",
  54445=>"000100110",
  54446=>"101110111",
  54447=>"000001111",
  54448=>"111111110",
  54449=>"110100100",
  54450=>"010001000",
  54451=>"110100000",
  54452=>"110010000",
  54453=>"000000001",
  54454=>"000000111",
  54455=>"111111111",
  54456=>"110110111",
  54457=>"111111111",
  54458=>"000000001",
  54459=>"101111000",
  54460=>"011111011",
  54461=>"111101000",
  54462=>"111001011",
  54463=>"111111111",
  54464=>"111001000",
  54465=>"011111111",
  54466=>"111111111",
  54467=>"011111000",
  54468=>"000000000",
  54469=>"011111011",
  54470=>"111111111",
  54471=>"000000111",
  54472=>"000000000",
  54473=>"101001001",
  54474=>"001001001",
  54475=>"111111111",
  54476=>"000000100",
  54477=>"000001111",
  54478=>"000000000",
  54479=>"001000000",
  54480=>"000000001",
  54481=>"100000111",
  54482=>"001000000",
  54483=>"000000011",
  54484=>"111111011",
  54485=>"111111011",
  54486=>"000011011",
  54487=>"010000000",
  54488=>"000000111",
  54489=>"110110101",
  54490=>"000010000",
  54491=>"000000000",
  54492=>"001000110",
  54493=>"111111111",
  54494=>"001101000",
  54495=>"000110111",
  54496=>"001001111",
  54497=>"110110111",
  54498=>"000111111",
  54499=>"011011000",
  54500=>"001000000",
  54501=>"001011100",
  54502=>"111111111",
  54503=>"111111100",
  54504=>"001111111",
  54505=>"010000110",
  54506=>"111111111",
  54507=>"001111010",
  54508=>"000001111",
  54509=>"111111111",
  54510=>"111111111",
  54511=>"000111111",
  54512=>"000111111",
  54513=>"000000000",
  54514=>"000010000",
  54515=>"101101110",
  54516=>"000111111",
  54517=>"000000000",
  54518=>"000010011",
  54519=>"111100000",
  54520=>"000111000",
  54521=>"001011010",
  54522=>"111111110",
  54523=>"101100111",
  54524=>"000001000",
  54525=>"001001001",
  54526=>"111111111",
  54527=>"000000010",
  54528=>"001000110",
  54529=>"011011000",
  54530=>"000000111",
  54531=>"001001111",
  54532=>"011001000",
  54533=>"111111111",
  54534=>"011010000",
  54535=>"001011111",
  54536=>"000110010",
  54537=>"110111010",
  54538=>"111101111",
  54539=>"111110100",
  54540=>"001001001",
  54541=>"001101110",
  54542=>"111111111",
  54543=>"110111000",
  54544=>"000000001",
  54545=>"000001111",
  54546=>"111001111",
  54547=>"100000111",
  54548=>"111111010",
  54549=>"111111111",
  54550=>"001000000",
  54551=>"111111111",
  54552=>"101111111",
  54553=>"011100100",
  54554=>"000011000",
  54555=>"011111111",
  54556=>"100110110",
  54557=>"000000001",
  54558=>"010111111",
  54559=>"000000000",
  54560=>"001000000",
  54561=>"111110100",
  54562=>"111001011",
  54563=>"000000000",
  54564=>"000111110",
  54565=>"111111111",
  54566=>"100000000",
  54567=>"111011001",
  54568=>"111000000",
  54569=>"000000000",
  54570=>"110000000",
  54571=>"010000000",
  54572=>"110110010",
  54573=>"000000001",
  54574=>"000000111",
  54575=>"011111111",
  54576=>"110000100",
  54577=>"000011111",
  54578=>"000001110",
  54579=>"010011111",
  54580=>"111100111",
  54581=>"000000001",
  54582=>"000010000",
  54583=>"000000010",
  54584=>"000100000",
  54585=>"011000101",
  54586=>"000010000",
  54587=>"000000000",
  54588=>"001011000",
  54589=>"111111111",
  54590=>"111100100",
  54591=>"010011000",
  54592=>"001001101",
  54593=>"111111111",
  54594=>"011010000",
  54595=>"000000111",
  54596=>"010110110",
  54597=>"000000000",
  54598=>"000011111",
  54599=>"101111111",
  54600=>"000111000",
  54601=>"011000001",
  54602=>"111001011",
  54603=>"011001001",
  54604=>"001011111",
  54605=>"111111111",
  54606=>"101000001",
  54607=>"110110110",
  54608=>"001111011",
  54609=>"101000001",
  54610=>"000111111",
  54611=>"000000000",
  54612=>"111000000",
  54613=>"011011000",
  54614=>"111111111",
  54615=>"000000111",
  54616=>"111001001",
  54617=>"111011111",
  54618=>"011011000",
  54619=>"110111111",
  54620=>"111111111",
  54621=>"110000000",
  54622=>"000111111",
  54623=>"111111110",
  54624=>"000011111",
  54625=>"000100111",
  54626=>"000000000",
  54627=>"000011111",
  54628=>"000000000",
  54629=>"001011000",
  54630=>"000000001",
  54631=>"000111111",
  54632=>"111110100",
  54633=>"000000000",
  54634=>"000000000",
  54635=>"111111111",
  54636=>"000100100",
  54637=>"101000000",
  54638=>"001000000",
  54639=>"001011000",
  54640=>"000000101",
  54641=>"100000000",
  54642=>"111111110",
  54643=>"110111111",
  54644=>"001000000",
  54645=>"100101111",
  54646=>"000100100",
  54647=>"000000000",
  54648=>"000000110",
  54649=>"000000000",
  54650=>"001000001",
  54651=>"001011111",
  54652=>"111001000",
  54653=>"111111111",
  54654=>"000000000",
  54655=>"001000000",
  54656=>"000000100",
  54657=>"001011001",
  54658=>"111111111",
  54659=>"000000000",
  54660=>"000000111",
  54661=>"100100111",
  54662=>"111111111",
  54663=>"111001000",
  54664=>"111111111",
  54665=>"100000000",
  54666=>"111111111",
  54667=>"001000111",
  54668=>"111111111",
  54669=>"100111111",
  54670=>"000111111",
  54671=>"000000010",
  54672=>"000000111",
  54673=>"011111100",
  54674=>"000011011",
  54675=>"000110110",
  54676=>"000100111",
  54677=>"000000000",
  54678=>"001000010",
  54679=>"111111100",
  54680=>"111111000",
  54681=>"000011111",
  54682=>"001010110",
  54683=>"000000000",
  54684=>"011000100",
  54685=>"110100000",
  54686=>"101111111",
  54687=>"000011001",
  54688=>"000001000",
  54689=>"101110111",
  54690=>"111111100",
  54691=>"000000000",
  54692=>"000000000",
  54693=>"000000000",
  54694=>"000000000",
  54695=>"111110111",
  54696=>"110111110",
  54697=>"000000000",
  54698=>"111111111",
  54699=>"001001111",
  54700=>"000000000",
  54701=>"000000000",
  54702=>"011011111",
  54703=>"110111011",
  54704=>"000010111",
  54705=>"000000000",
  54706=>"110110000",
  54707=>"111011000",
  54708=>"111011010",
  54709=>"000000110",
  54710=>"000100100",
  54711=>"000000100",
  54712=>"001001110",
  54713=>"111011000",
  54714=>"111001000",
  54715=>"111111111",
  54716=>"111000000",
  54717=>"111100100",
  54718=>"000000001",
  54719=>"011001001",
  54720=>"011011110",
  54721=>"111111000",
  54722=>"011011011",
  54723=>"110111111",
  54724=>"000110111",
  54725=>"001011000",
  54726=>"100000001",
  54727=>"010000011",
  54728=>"000110111",
  54729=>"000011011",
  54730=>"001111111",
  54731=>"001111111",
  54732=>"111111111",
  54733=>"000001011",
  54734=>"101011111",
  54735=>"111111111",
  54736=>"000101111",
  54737=>"111111011",
  54738=>"111111110",
  54739=>"000000011",
  54740=>"000000000",
  54741=>"111111011",
  54742=>"111111111",
  54743=>"100100000",
  54744=>"111010000",
  54745=>"101000000",
  54746=>"111111111",
  54747=>"111000000",
  54748=>"000000111",
  54749=>"111011011",
  54750=>"000000101",
  54751=>"000011111",
  54752=>"111111100",
  54753=>"101101111",
  54754=>"111111110",
  54755=>"000000000",
  54756=>"100000000",
  54757=>"100111011",
  54758=>"000101111",
  54759=>"000000000",
  54760=>"111111111",
  54761=>"001001000",
  54762=>"000000000",
  54763=>"100000000",
  54764=>"000001111",
  54765=>"000011011",
  54766=>"111111110",
  54767=>"110000011",
  54768=>"000100101",
  54769=>"111111000",
  54770=>"100111111",
  54771=>"000001111",
  54772=>"100111111",
  54773=>"111111111",
  54774=>"111111111",
  54775=>"100000000",
  54776=>"110111101",
  54777=>"000001001",
  54778=>"000000110",
  54779=>"111111011",
  54780=>"111001111",
  54781=>"001000100",
  54782=>"000000110",
  54783=>"000000011",
  54784=>"110110110",
  54785=>"000110111",
  54786=>"101001001",
  54787=>"010001111",
  54788=>"000111111",
  54789=>"001001001",
  54790=>"111000000",
  54791=>"111001001",
  54792=>"011011111",
  54793=>"000101000",
  54794=>"110110101",
  54795=>"111110000",
  54796=>"111101001",
  54797=>"110111111",
  54798=>"011111111",
  54799=>"111111111",
  54800=>"100110111",
  54801=>"111000001",
  54802=>"110111000",
  54803=>"000001111",
  54804=>"000000111",
  54805=>"101001001",
  54806=>"111000001",
  54807=>"110110110",
  54808=>"111011111",
  54809=>"011111111",
  54810=>"101111111",
  54811=>"000001001",
  54812=>"010010010",
  54813=>"000000111",
  54814=>"010110111",
  54815=>"000011111",
  54816=>"011001000",
  54817=>"010010010",
  54818=>"000000000",
  54819=>"101101001",
  54820=>"000000000",
  54821=>"000110110",
  54822=>"011000000",
  54823=>"001001111",
  54824=>"110110111",
  54825=>"101101101",
  54826=>"001001000",
  54827=>"110111011",
  54828=>"111000000",
  54829=>"111111101",
  54830=>"011001000",
  54831=>"100111111",
  54832=>"111111111",
  54833=>"000111111",
  54834=>"000010111",
  54835=>"110011010",
  54836=>"100000110",
  54837=>"110110110",
  54838=>"010010001",
  54839=>"001000001",
  54840=>"110111111",
  54841=>"000001001",
  54842=>"001001001",
  54843=>"001000111",
  54844=>"001111010",
  54845=>"010000000",
  54846=>"011110100",
  54847=>"001111011",
  54848=>"000000111",
  54849=>"101110000",
  54850=>"110111011",
  54851=>"111101111",
  54852=>"000000001",
  54853=>"001000000",
  54854=>"111000000",
  54855=>"111111111",
  54856=>"110111111",
  54857=>"111001001",
  54858=>"111000000",
  54859=>"111000001",
  54860=>"111001011",
  54861=>"111000111",
  54862=>"000111111",
  54863=>"011111111",
  54864=>"000000111",
  54865=>"001001001",
  54866=>"000000111",
  54867=>"111111110",
  54868=>"110111111",
  54869=>"000010010",
  54870=>"000001000",
  54871=>"010000000",
  54872=>"000000000",
  54873=>"111101111",
  54874=>"111111111",
  54875=>"001001001",
  54876=>"000000000",
  54877=>"111111100",
  54878=>"000000000",
  54879=>"011001000",
  54880=>"000010010",
  54881=>"110101101",
  54882=>"111000000",
  54883=>"000000000",
  54884=>"000111110",
  54885=>"111101001",
  54886=>"000000000",
  54887=>"111111000",
  54888=>"000000010",
  54889=>"000000001",
  54890=>"000000000",
  54891=>"110110000",
  54892=>"010000000",
  54893=>"000110010",
  54894=>"000000110",
  54895=>"101000000",
  54896=>"000001001",
  54897=>"111110100",
  54898=>"001111111",
  54899=>"000001111",
  54900=>"000000000",
  54901=>"000000111",
  54902=>"111111000",
  54903=>"010011000",
  54904=>"001001000",
  54905=>"000001000",
  54906=>"100000000",
  54907=>"100101111",
  54908=>"100111110",
  54909=>"110000000",
  54910=>"000000000",
  54911=>"111000000",
  54912=>"000000000",
  54913=>"111110110",
  54914=>"111111111",
  54915=>"101001000",
  54916=>"001001101",
  54917=>"110100000",
  54918=>"101101011",
  54919=>"000111111",
  54920=>"110111111",
  54921=>"000000000",
  54922=>"000111000",
  54923=>"111111111",
  54924=>"111110111",
  54925=>"111000001",
  54926=>"001001111",
  54927=>"100110111",
  54928=>"001001001",
  54929=>"000100111",
  54930=>"111001001",
  54931=>"000000010",
  54932=>"001111110",
  54933=>"110110000",
  54934=>"000001001",
  54935=>"001000101",
  54936=>"001000000",
  54937=>"000001111",
  54938=>"110111000",
  54939=>"000101111",
  54940=>"000000001",
  54941=>"001001000",
  54942=>"001001100",
  54943=>"000000000",
  54944=>"000000001",
  54945=>"000010111",
  54946=>"000111110",
  54947=>"000110011",
  54948=>"111011000",
  54949=>"010111011",
  54950=>"111111010",
  54951=>"011111111",
  54952=>"111111111",
  54953=>"010111111",
  54954=>"000000000",
  54955=>"111111111",
  54956=>"100101111",
  54957=>"000000000",
  54958=>"111111000",
  54959=>"000010101",
  54960=>"000000000",
  54961=>"110111111",
  54962=>"111111110",
  54963=>"000100111",
  54964=>"111111000",
  54965=>"110111111",
  54966=>"110100000",
  54967=>"010111010",
  54968=>"000101111",
  54969=>"000000000",
  54970=>"010000001",
  54971=>"010000011",
  54972=>"000000111",
  54973=>"001000000",
  54974=>"000111111",
  54975=>"000110111",
  54976=>"000000000",
  54977=>"010111110",
  54978=>"110010110",
  54979=>"111101000",
  54980=>"000001001",
  54981=>"111111101",
  54982=>"111111111",
  54983=>"000000000",
  54984=>"001001001",
  54985=>"111011001",
  54986=>"010111000",
  54987=>"111110111",
  54988=>"000000101",
  54989=>"111010111",
  54990=>"000001010",
  54991=>"010010110",
  54992=>"111101001",
  54993=>"000000000",
  54994=>"010111101",
  54995=>"111010000",
  54996=>"111111111",
  54997=>"001001001",
  54998=>"100000100",
  54999=>"001111111",
  55000=>"000001000",
  55001=>"000110011",
  55002=>"000000000",
  55003=>"110100000",
  55004=>"100000000",
  55005=>"111111111",
  55006=>"100111011",
  55007=>"010001011",
  55008=>"001001011",
  55009=>"101111111",
  55010=>"111110100",
  55011=>"000000000",
  55012=>"010000000",
  55013=>"000000100",
  55014=>"010000001",
  55015=>"110111111",
  55016=>"100110110",
  55017=>"000001111",
  55018=>"000110111",
  55019=>"101101101",
  55020=>"110111110",
  55021=>"111111111",
  55022=>"110110000",
  55023=>"001000000",
  55024=>"010110000",
  55025=>"000000000",
  55026=>"000100111",
  55027=>"110110000",
  55028=>"001000011",
  55029=>"111110000",
  55030=>"110100100",
  55031=>"001000101",
  55032=>"101101100",
  55033=>"111000000",
  55034=>"100000110",
  55035=>"110000000",
  55036=>"000000000",
  55037=>"011111111",
  55038=>"110111111",
  55039=>"000000011",
  55040=>"001001001",
  55041=>"000111111",
  55042=>"111111111",
  55043=>"000001111",
  55044=>"000100101",
  55045=>"001111110",
  55046=>"110111110",
  55047=>"110001111",
  55048=>"000011011",
  55049=>"001000000",
  55050=>"000000101",
  55051=>"010111111",
  55052=>"011111111",
  55053=>"110011001",
  55054=>"111111000",
  55055=>"111111100",
  55056=>"001000001",
  55057=>"001001110",
  55058=>"100001111",
  55059=>"010010001",
  55060=>"000101000",
  55061=>"000000111",
  55062=>"001001011",
  55063=>"000001000",
  55064=>"011110110",
  55065=>"111000111",
  55066=>"100000000",
  55067=>"000000111",
  55068=>"111111111",
  55069=>"000000000",
  55070=>"000000111",
  55071=>"000000000",
  55072=>"010111111",
  55073=>"111111000",
  55074=>"110000000",
  55075=>"000101000",
  55076=>"100110110",
  55077=>"100000000",
  55078=>"110010110",
  55079=>"111111001",
  55080=>"000000000",
  55081=>"111010010",
  55082=>"111100100",
  55083=>"001001111",
  55084=>"100111100",
  55085=>"000000001",
  55086=>"000000000",
  55087=>"110111111",
  55088=>"011001011",
  55089=>"111101101",
  55090=>"000000001",
  55091=>"111111000",
  55092=>"110110000",
  55093=>"000111111",
  55094=>"101101101",
  55095=>"111000000",
  55096=>"000000000",
  55097=>"101111011",
  55098=>"010000000",
  55099=>"000000100",
  55100=>"111100000",
  55101=>"110010111",
  55102=>"110111111",
  55103=>"000100111",
  55104=>"001001111",
  55105=>"111111111",
  55106=>"000000001",
  55107=>"101000000",
  55108=>"111101001",
  55109=>"111101001",
  55110=>"001001000",
  55111=>"111111000",
  55112=>"010111111",
  55113=>"100000100",
  55114=>"101001010",
  55115=>"111111011",
  55116=>"001000000",
  55117=>"000101011",
  55118=>"000000000",
  55119=>"000000100",
  55120=>"000000001",
  55121=>"010000110",
  55122=>"110111110",
  55123=>"000000000",
  55124=>"110001011",
  55125=>"011111010",
  55126=>"000110110",
  55127=>"111000000",
  55128=>"110111000",
  55129=>"111111111",
  55130=>"000000111",
  55131=>"000000011",
  55132=>"111001000",
  55133=>"001000001",
  55134=>"001000100",
  55135=>"000001111",
  55136=>"000000000",
  55137=>"111011011",
  55138=>"010011110",
  55139=>"100000000",
  55140=>"010010000",
  55141=>"000000000",
  55142=>"111101111",
  55143=>"011111111",
  55144=>"111111101",
  55145=>"101001100",
  55146=>"110110101",
  55147=>"010010100",
  55148=>"001011001",
  55149=>"011000001",
  55150=>"000001101",
  55151=>"111111111",
  55152=>"000000000",
  55153=>"000000000",
  55154=>"111001001",
  55155=>"111011011",
  55156=>"000001000",
  55157=>"000111101",
  55158=>"000011011",
  55159=>"000000001",
  55160=>"000000000",
  55161=>"000000000",
  55162=>"111111101",
  55163=>"000000001",
  55164=>"101111001",
  55165=>"110000001",
  55166=>"011000110",
  55167=>"000000000",
  55168=>"011011011",
  55169=>"100001011",
  55170=>"100000001",
  55171=>"001111111",
  55172=>"000001111",
  55173=>"111111000",
  55174=>"101101111",
  55175=>"000000100",
  55176=>"001101101",
  55177=>"000110000",
  55178=>"101000001",
  55179=>"000000101",
  55180=>"001001000",
  55181=>"011111011",
  55182=>"000100101",
  55183=>"101101111",
  55184=>"100111110",
  55185=>"110000000",
  55186=>"101111111",
  55187=>"000001001",
  55188=>"110111111",
  55189=>"000000000",
  55190=>"111011111",
  55191=>"110000000",
  55192=>"000000101",
  55193=>"001010110",
  55194=>"110010000",
  55195=>"001001000",
  55196=>"111111111",
  55197=>"000000101",
  55198=>"110110110",
  55199=>"111011111",
  55200=>"000000000",
  55201=>"000000000",
  55202=>"000000001",
  55203=>"111100100",
  55204=>"110110110",
  55205=>"111110000",
  55206=>"111111111",
  55207=>"000000000",
  55208=>"000000000",
  55209=>"111101001",
  55210=>"000100100",
  55211=>"110111110",
  55212=>"000000000",
  55213=>"011000101",
  55214=>"000000101",
  55215=>"011110110",
  55216=>"111111111",
  55217=>"000000000",
  55218=>"000000110",
  55219=>"000000101",
  55220=>"101000110",
  55221=>"111111000",
  55222=>"001011001",
  55223=>"111111111",
  55224=>"111000000",
  55225=>"111111111",
  55226=>"111000000",
  55227=>"111000000",
  55228=>"010110101",
  55229=>"000000000",
  55230=>"111001111",
  55231=>"010010001",
  55232=>"111111110",
  55233=>"110110110",
  55234=>"001001001",
  55235=>"000000000",
  55236=>"011111000",
  55237=>"001001101",
  55238=>"001001101",
  55239=>"001001111",
  55240=>"111110001",
  55241=>"000001011",
  55242=>"111001000",
  55243=>"111001001",
  55244=>"000101111",
  55245=>"111111111",
  55246=>"111001101",
  55247=>"010000000",
  55248=>"000001001",
  55249=>"000110111",
  55250=>"000000000",
  55251=>"101111111",
  55252=>"100100100",
  55253=>"110111101",
  55254=>"001111111",
  55255=>"111110100",
  55256=>"111001100",
  55257=>"000000000",
  55258=>"000000000",
  55259=>"000000000",
  55260=>"111111111",
  55261=>"110100110",
  55262=>"000000000",
  55263=>"110110011",
  55264=>"111101101",
  55265=>"000000111",
  55266=>"000000000",
  55267=>"111100000",
  55268=>"000010111",
  55269=>"101101111",
  55270=>"000111111",
  55271=>"000000100",
  55272=>"110110000",
  55273=>"100000111",
  55274=>"001000000",
  55275=>"111110000",
  55276=>"000011011",
  55277=>"011000011",
  55278=>"101111111",
  55279=>"000000000",
  55280=>"000000000",
  55281=>"111111111",
  55282=>"000111000",
  55283=>"000011001",
  55284=>"110110000",
  55285=>"010000010",
  55286=>"111011011",
  55287=>"110011011",
  55288=>"000110111",
  55289=>"000000000",
  55290=>"000000000",
  55291=>"101001101",
  55292=>"111111111",
  55293=>"000000111",
  55294=>"001000000",
  55295=>"000011000",
  55296=>"000000000",
  55297=>"111000101",
  55298=>"111111111",
  55299=>"110000000",
  55300=>"100000111",
  55301=>"111000011",
  55302=>"000000000",
  55303=>"111111111",
  55304=>"111111010",
  55305=>"001011111",
  55306=>"000000111",
  55307=>"111110111",
  55308=>"001011000",
  55309=>"000000110",
  55310=>"000011011",
  55311=>"111111000",
  55312=>"101000000",
  55313=>"101100111",
  55314=>"111101000",
  55315=>"111111111",
  55316=>"000100011",
  55317=>"000001000",
  55318=>"111001000",
  55319=>"100111111",
  55320=>"000110110",
  55321=>"000000000",
  55322=>"000000111",
  55323=>"110000101",
  55324=>"000001000",
  55325=>"000101111",
  55326=>"001001011",
  55327=>"111111000",
  55328=>"100000000",
  55329=>"111001001",
  55330=>"111100100",
  55331=>"000111111",
  55332=>"001100000",
  55333=>"010011111",
  55334=>"000000001",
  55335=>"100111111",
  55336=>"001101001",
  55337=>"011111111",
  55338=>"000000000",
  55339=>"111110111",
  55340=>"000000000",
  55341=>"111111111",
  55342=>"011011111",
  55343=>"100110110",
  55344=>"100110111",
  55345=>"000001000",
  55346=>"001111100",
  55347=>"000000000",
  55348=>"001011000",
  55349=>"101001000",
  55350=>"111111111",
  55351=>"110000111",
  55352=>"100000000",
  55353=>"111001111",
  55354=>"000011011",
  55355=>"110110000",
  55356=>"101000000",
  55357=>"100000000",
  55358=>"111111111",
  55359=>"010000000",
  55360=>"001001111",
  55361=>"000000110",
  55362=>"111111111",
  55363=>"111111111",
  55364=>"111000100",
  55365=>"001001001",
  55366=>"111010000",
  55367=>"000000000",
  55368=>"000000000",
  55369=>"011111111",
  55370=>"111111110",
  55371=>"000000111",
  55372=>"000110111",
  55373=>"100100001",
  55374=>"111011111",
  55375=>"000000000",
  55376=>"111110111",
  55377=>"010000100",
  55378=>"001011000",
  55379=>"100000000",
  55380=>"000000000",
  55381=>"111111111",
  55382=>"100111111",
  55383=>"110110110",
  55384=>"010111111",
  55385=>"111111111",
  55386=>"111111110",
  55387=>"110111111",
  55388=>"000000000",
  55389=>"000000000",
  55390=>"110111011",
  55391=>"111111111",
  55392=>"010000000",
  55393=>"000000000",
  55394=>"111110111",
  55395=>"100000000",
  55396=>"001111101",
  55397=>"100000000",
  55398=>"100100111",
  55399=>"111111111",
  55400=>"010010000",
  55401=>"000000000",
  55402=>"101101000",
  55403=>"000000000",
  55404=>"011111111",
  55405=>"000000100",
  55406=>"110111111",
  55407=>"000000000",
  55408=>"000000000",
  55409=>"111111111",
  55410=>"011001000",
  55411=>"111111111",
  55412=>"111111111",
  55413=>"111001000",
  55414=>"000110111",
  55415=>"000000000",
  55416=>"000000000",
  55417=>"001001001",
  55418=>"111000000",
  55419=>"000000000",
  55420=>"111100100",
  55421=>"110100110",
  55422=>"111111000",
  55423=>"000000000",
  55424=>"000111111",
  55425=>"101000000",
  55426=>"000000111",
  55427=>"111011011",
  55428=>"111111111",
  55429=>"000010000",
  55430=>"111110110",
  55431=>"111111111",
  55432=>"111111111",
  55433=>"111010000",
  55434=>"000000001",
  55435=>"000111011",
  55436=>"000000000",
  55437=>"001000000",
  55438=>"000000011",
  55439=>"000111111",
  55440=>"101111111",
  55441=>"111111000",
  55442=>"001111110",
  55443=>"001111111",
  55444=>"110111111",
  55445=>"100100100",
  55446=>"000000000",
  55447=>"100111011",
  55448=>"000000110",
  55449=>"111111111",
  55450=>"101100000",
  55451=>"000000000",
  55452=>"111000000",
  55453=>"110110111",
  55454=>"000000011",
  55455=>"011111000",
  55456=>"000000100",
  55457=>"010111111",
  55458=>"000000100",
  55459=>"000000000",
  55460=>"111111100",
  55461=>"111110100",
  55462=>"110100000",
  55463=>"001001001",
  55464=>"111111111",
  55465=>"110110100",
  55466=>"000000000",
  55467=>"111011111",
  55468=>"111111000",
  55469=>"001000000",
  55470=>"011000000",
  55471=>"000000000",
  55472=>"111011011",
  55473=>"011000000",
  55474=>"001001000",
  55475=>"011000000",
  55476=>"000000110",
  55477=>"111000000",
  55478=>"110000000",
  55479=>"000000000",
  55480=>"001000001",
  55481=>"000000000",
  55482=>"111101100",
  55483=>"110100110",
  55484=>"111100110",
  55485=>"001000000",
  55486=>"111111111",
  55487=>"000000010",
  55488=>"001000001",
  55489=>"010000000",
  55490=>"011111111",
  55491=>"111100111",
  55492=>"111001111",
  55493=>"111111111",
  55494=>"111111111",
  55495=>"000000001",
  55496=>"110000000",
  55497=>"111000000",
  55498=>"111111101",
  55499=>"100000000",
  55500=>"111111111",
  55501=>"000111111",
  55502=>"110000100",
  55503=>"111100000",
  55504=>"000100111",
  55505=>"110111111",
  55506=>"100100110",
  55507=>"111101000",
  55508=>"000000000",
  55509=>"011001000",
  55510=>"001111111",
  55511=>"111001111",
  55512=>"111111001",
  55513=>"000010011",
  55514=>"001001111",
  55515=>"000000000",
  55516=>"100000110",
  55517=>"111111111",
  55518=>"001111011",
  55519=>"110100010",
  55520=>"010010100",
  55521=>"000010010",
  55522=>"111111111",
  55523=>"100000000",
  55524=>"101111111",
  55525=>"011110110",
  55526=>"111111111",
  55527=>"111111111",
  55528=>"100100000",
  55529=>"111111101",
  55530=>"111111111",
  55531=>"110111011",
  55532=>"000110000",
  55533=>"000000100",
  55534=>"001011111",
  55535=>"000001111",
  55536=>"011000000",
  55537=>"000000111",
  55538=>"100101101",
  55539=>"000000000",
  55540=>"000000000",
  55541=>"111111111",
  55542=>"001011011",
  55543=>"110111110",
  55544=>"000101100",
  55545=>"111000000",
  55546=>"000000111",
  55547=>"000000111",
  55548=>"110110100",
  55549=>"001011000",
  55550=>"111111111",
  55551=>"000000100",
  55552=>"000000001",
  55553=>"001001001",
  55554=>"100111000",
  55555=>"111100111",
  55556=>"000000000",
  55557=>"011011011",
  55558=>"001111111",
  55559=>"111101111",
  55560=>"000011011",
  55561=>"000000000",
  55562=>"010100100",
  55563=>"100000000",
  55564=>"111100000",
  55565=>"000000000",
  55566=>"100101001",
  55567=>"010000000",
  55568=>"111111001",
  55569=>"000000011",
  55570=>"111111111",
  55571=>"111001000",
  55572=>"011000000",
  55573=>"110100111",
  55574=>"101001000",
  55575=>"001000000",
  55576=>"010000000",
  55577=>"110000110",
  55578=>"100000000",
  55579=>"111111111",
  55580=>"000010110",
  55581=>"100000011",
  55582=>"111111111",
  55583=>"000000111",
  55584=>"011111110",
  55585=>"100000010",
  55586=>"100100100",
  55587=>"110111111",
  55588=>"000000000",
  55589=>"111111111",
  55590=>"111111111",
  55591=>"011111000",
  55592=>"000000111",
  55593=>"000000000",
  55594=>"111100000",
  55595=>"000000000",
  55596=>"111111100",
  55597=>"000010000",
  55598=>"110010000",
  55599=>"100001001",
  55600=>"011000111",
  55601=>"000111111",
  55602=>"010000000",
  55603=>"000000111",
  55604=>"110000000",
  55605=>"000000000",
  55606=>"111111001",
  55607=>"100100110",
  55608=>"000000000",
  55609=>"111000000",
  55610=>"000101000",
  55611=>"000001000",
  55612=>"001111111",
  55613=>"111110100",
  55614=>"000101111",
  55615=>"011000000",
  55616=>"000000000",
  55617=>"111100000",
  55618=>"111111111",
  55619=>"000000000",
  55620=>"010000010",
  55621=>"001000000",
  55622=>"111111000",
  55623=>"000000000",
  55624=>"111001101",
  55625=>"011000111",
  55626=>"111100100",
  55627=>"111111111",
  55628=>"110000110",
  55629=>"111111111",
  55630=>"110111111",
  55631=>"111111111",
  55632=>"011111111",
  55633=>"111100111",
  55634=>"000110101",
  55635=>"000000000",
  55636=>"111111000",
  55637=>"000001001",
  55638=>"110111111",
  55639=>"000000000",
  55640=>"000000000",
  55641=>"111010010",
  55642=>"011000000",
  55643=>"111111011",
  55644=>"111110000",
  55645=>"100000000",
  55646=>"110110100",
  55647=>"101001001",
  55648=>"100000111",
  55649=>"000000000",
  55650=>"111110001",
  55651=>"001111111",
  55652=>"000000000",
  55653=>"111101000",
  55654=>"011111111",
  55655=>"111111111",
  55656=>"000000011",
  55657=>"111111111",
  55658=>"111111100",
  55659=>"001011011",
  55660=>"011101100",
  55661=>"111111000",
  55662=>"111000000",
  55663=>"000000000",
  55664=>"110010000",
  55665=>"100000000",
  55666=>"100000000",
  55667=>"111111111",
  55668=>"000100000",
  55669=>"000010001",
  55670=>"000011011",
  55671=>"110110000",
  55672=>"111000000",
  55673=>"111100000",
  55674=>"001001011",
  55675=>"000111111",
  55676=>"101000000",
  55677=>"000000000",
  55678=>"110000000",
  55679=>"111101111",
  55680=>"111100100",
  55681=>"111101101",
  55682=>"100111110",
  55683=>"111000000",
  55684=>"111111111",
  55685=>"010110010",
  55686=>"110110110",
  55687=>"000010000",
  55688=>"000000001",
  55689=>"000000111",
  55690=>"111111111",
  55691=>"111010110",
  55692=>"000110111",
  55693=>"000000000",
  55694=>"110100111",
  55695=>"000000000",
  55696=>"111111011",
  55697=>"111000000",
  55698=>"111110111",
  55699=>"110111111",
  55700=>"100100100",
  55701=>"000000000",
  55702=>"111100001",
  55703=>"101111110",
  55704=>"100101111",
  55705=>"111101101",
  55706=>"010111111",
  55707=>"110111111",
  55708=>"100100111",
  55709=>"111111111",
  55710=>"110100000",
  55711=>"000000000",
  55712=>"000001000",
  55713=>"000000000",
  55714=>"111111111",
  55715=>"111000000",
  55716=>"110111111",
  55717=>"111111111",
  55718=>"000000000",
  55719=>"000000101",
  55720=>"000111000",
  55721=>"111111111",
  55722=>"000000000",
  55723=>"100000000",
  55724=>"110111111",
  55725=>"000110000",
  55726=>"001001001",
  55727=>"111111111",
  55728=>"000000000",
  55729=>"000000110",
  55730=>"000011111",
  55731=>"000000000",
  55732=>"000000000",
  55733=>"110100111",
  55734=>"011001001",
  55735=>"110000000",
  55736=>"110000101",
  55737=>"111111111",
  55738=>"111000111",
  55739=>"011111110",
  55740=>"101000000",
  55741=>"000000000",
  55742=>"011011011",
  55743=>"100001000",
  55744=>"000000000",
  55745=>"010111111",
  55746=>"000001000",
  55747=>"111111111",
  55748=>"110111111",
  55749=>"111111001",
  55750=>"111101000",
  55751=>"111100100",
  55752=>"100100111",
  55753=>"111111101",
  55754=>"111110110",
  55755=>"000111111",
  55756=>"100000000",
  55757=>"011111111",
  55758=>"100100100",
  55759=>"111101000",
  55760=>"010000011",
  55761=>"000100000",
  55762=>"000000000",
  55763=>"000110111",
  55764=>"000000111",
  55765=>"101111111",
  55766=>"000000011",
  55767=>"000000000",
  55768=>"110000000",
  55769=>"000000000",
  55770=>"000000100",
  55771=>"100101111",
  55772=>"001001011",
  55773=>"100100111",
  55774=>"111111111",
  55775=>"110111111",
  55776=>"011000000",
  55777=>"111110111",
  55778=>"010111110",
  55779=>"011111000",
  55780=>"000000001",
  55781=>"101111110",
  55782=>"010111110",
  55783=>"100110110",
  55784=>"110000100",
  55785=>"000001111",
  55786=>"000000000",
  55787=>"000001000",
  55788=>"100111111",
  55789=>"111111011",
  55790=>"000000000",
  55791=>"111111111",
  55792=>"000000000",
  55793=>"010000110",
  55794=>"111100000",
  55795=>"100011111",
  55796=>"111111100",
  55797=>"100100111",
  55798=>"001111111",
  55799=>"000000001",
  55800=>"111111111",
  55801=>"111000000",
  55802=>"110000000",
  55803=>"000000000",
  55804=>"111111111",
  55805=>"000000000",
  55806=>"000000000",
  55807=>"111111111",
  55808=>"000000011",
  55809=>"111110000",
  55810=>"111111111",
  55811=>"111110000",
  55812=>"000000000",
  55813=>"101100100",
  55814=>"111111111",
  55815=>"111111111",
  55816=>"001000000",
  55817=>"011110111",
  55818=>"100111111",
  55819=>"111111110",
  55820=>"111111111",
  55821=>"001100100",
  55822=>"000000000",
  55823=>"000000111",
  55824=>"001111111",
  55825=>"011000111",
  55826=>"001000101",
  55827=>"000000000",
  55828=>"000100000",
  55829=>"000001100",
  55830=>"001000111",
  55831=>"000000001",
  55832=>"100110100",
  55833=>"100000000",
  55834=>"000000000",
  55835=>"100010000",
  55836=>"000000000",
  55837=>"000000111",
  55838=>"110000000",
  55839=>"101111001",
  55840=>"000000000",
  55841=>"110000000",
  55842=>"000001111",
  55843=>"100000011",
  55844=>"110100100",
  55845=>"001001001",
  55846=>"100111101",
  55847=>"101000111",
  55848=>"001100100",
  55849=>"000000000",
  55850=>"000000000",
  55851=>"000000001",
  55852=>"000100111",
  55853=>"000000000",
  55854=>"000010000",
  55855=>"110000101",
  55856=>"000000000",
  55857=>"111000000",
  55858=>"010011001",
  55859=>"000000011",
  55860=>"000110110",
  55861=>"111111001",
  55862=>"111111101",
  55863=>"111111101",
  55864=>"000000000",
  55865=>"011010111",
  55866=>"000000101",
  55867=>"111111111",
  55868=>"111111110",
  55869=>"000100100",
  55870=>"110110100",
  55871=>"111000110",
  55872=>"000000000",
  55873=>"000000000",
  55874=>"110001000",
  55875=>"000000110",
  55876=>"100101101",
  55877=>"000000111",
  55878=>"111111110",
  55879=>"111111111",
  55880=>"111111001",
  55881=>"000000000",
  55882=>"000000000",
  55883=>"111111111",
  55884=>"110110100",
  55885=>"000000000",
  55886=>"000111111",
  55887=>"111111010",
  55888=>"000000000",
  55889=>"110110000",
  55890=>"111111111",
  55891=>"001001000",
  55892=>"001000000",
  55893=>"011110110",
  55894=>"111111000",
  55895=>"111111000",
  55896=>"111111111",
  55897=>"000000111",
  55898=>"000000111",
  55899=>"000000000",
  55900=>"000000001",
  55901=>"100100111",
  55902=>"111100100",
  55903=>"000001000",
  55904=>"111000111",
  55905=>"000000100",
  55906=>"111111001",
  55907=>"111111111",
  55908=>"111111011",
  55909=>"000111111",
  55910=>"010000111",
  55911=>"111111001",
  55912=>"000000000",
  55913=>"111111111",
  55914=>"111111111",
  55915=>"000000000",
  55916=>"001001011",
  55917=>"000000000",
  55918=>"001000000",
  55919=>"000000000",
  55920=>"100111111",
  55921=>"110010011",
  55922=>"000000111",
  55923=>"100100000",
  55924=>"111111111",
  55925=>"011101111",
  55926=>"000000000",
  55927=>"011101100",
  55928=>"000000000",
  55929=>"101111111",
  55930=>"001000000",
  55931=>"000000011",
  55932=>"111111111",
  55933=>"000100110",
  55934=>"111000010",
  55935=>"000100000",
  55936=>"000000000",
  55937=>"011000111",
  55938=>"000000000",
  55939=>"111100000",
  55940=>"000000000",
  55941=>"111111010",
  55942=>"000100100",
  55943=>"111100100",
  55944=>"011011001",
  55945=>"111111111",
  55946=>"101000000",
  55947=>"000000000",
  55948=>"000011000",
  55949=>"111111111",
  55950=>"111110111",
  55951=>"001000000",
  55952=>"000000111",
  55953=>"100100100",
  55954=>"000101111",
  55955=>"111111111",
  55956=>"111110111",
  55957=>"111111111",
  55958=>"000000000",
  55959=>"111111111",
  55960=>"110111111",
  55961=>"000000000",
  55962=>"000000000",
  55963=>"111111011",
  55964=>"111001111",
  55965=>"000010000",
  55966=>"111101111",
  55967=>"111111111",
  55968=>"111100011",
  55969=>"111111001",
  55970=>"011000000",
  55971=>"101101011",
  55972=>"011011111",
  55973=>"011111111",
  55974=>"111111111",
  55975=>"111111111",
  55976=>"101111111",
  55977=>"000011111",
  55978=>"000000000",
  55979=>"000110110",
  55980=>"001000000",
  55981=>"111101000",
  55982=>"101111111",
  55983=>"110111111",
  55984=>"000010111",
  55985=>"111000000",
  55986=>"110000010",
  55987=>"000000000",
  55988=>"111100100",
  55989=>"111111111",
  55990=>"111111111",
  55991=>"111111111",
  55992=>"000000000",
  55993=>"000000000",
  55994=>"101001000",
  55995=>"001011111",
  55996=>"001001111",
  55997=>"010011010",
  55998=>"101111101",
  55999=>"000000001",
  56000=>"000000000",
  56001=>"111111111",
  56002=>"111111111",
  56003=>"100111111",
  56004=>"111110111",
  56005=>"111111100",
  56006=>"111111100",
  56007=>"111110100",
  56008=>"010111110",
  56009=>"111010000",
  56010=>"000000000",
  56011=>"111111111",
  56012=>"000100101",
  56013=>"111111101",
  56014=>"100100101",
  56015=>"101000000",
  56016=>"000000000",
  56017=>"000000000",
  56018=>"001011011",
  56019=>"111111011",
  56020=>"111001111",
  56021=>"011000101",
  56022=>"111111111",
  56023=>"111111111",
  56024=>"110110100",
  56025=>"000000100",
  56026=>"111111111",
  56027=>"000011111",
  56028=>"111111111",
  56029=>"000000011",
  56030=>"001001001",
  56031=>"111000000",
  56032=>"000000000",
  56033=>"011001000",
  56034=>"111111111",
  56035=>"111111111",
  56036=>"001000000",
  56037=>"000000000",
  56038=>"111100000",
  56039=>"111110010",
  56040=>"001000000",
  56041=>"110111111",
  56042=>"110000100",
  56043=>"000000000",
  56044=>"000110010",
  56045=>"111111111",
  56046=>"111111111",
  56047=>"010011011",
  56048=>"000000000",
  56049=>"111000000",
  56050=>"000011011",
  56051=>"111111111",
  56052=>"110100101",
  56053=>"110010010",
  56054=>"001011001",
  56055=>"000000000",
  56056=>"111111111",
  56057=>"000000110",
  56058=>"110110111",
  56059=>"000111001",
  56060=>"011011011",
  56061=>"001000000",
  56062=>"000000000",
  56063=>"000000000",
  56064=>"111000000",
  56065=>"000001000",
  56066=>"101100110",
  56067=>"011011000",
  56068=>"100100100",
  56069=>"110111111",
  56070=>"111111111",
  56071=>"111110111",
  56072=>"000000000",
  56073=>"000000000",
  56074=>"000000000",
  56075=>"000000110",
  56076=>"110100000",
  56077=>"111001000",
  56078=>"111110000",
  56079=>"000000011",
  56080=>"000111101",
  56081=>"111111111",
  56082=>"000000011",
  56083=>"000001001",
  56084=>"111111111",
  56085=>"001000001",
  56086=>"001001001",
  56087=>"111111011",
  56088=>"111001001",
  56089=>"000000000",
  56090=>"110111111",
  56091=>"110000000",
  56092=>"100110100",
  56093=>"100000000",
  56094=>"100000000",
  56095=>"000111011",
  56096=>"001001001",
  56097=>"001111110",
  56098=>"111111110",
  56099=>"111111110",
  56100=>"100100101",
  56101=>"000000101",
  56102=>"100100100",
  56103=>"111110000",
  56104=>"111001001",
  56105=>"111111111",
  56106=>"101111101",
  56107=>"111111111",
  56108=>"111011110",
  56109=>"011011001",
  56110=>"011001000",
  56111=>"000000000",
  56112=>"001000100",
  56113=>"111111110",
  56114=>"000100101",
  56115=>"111111111",
  56116=>"000011000",
  56117=>"000100111",
  56118=>"001101111",
  56119=>"011111111",
  56120=>"000000000",
  56121=>"100000000",
  56122=>"000000111",
  56123=>"010111111",
  56124=>"111001011",
  56125=>"100100000",
  56126=>"111111111",
  56127=>"000000100",
  56128=>"111000011",
  56129=>"100000001",
  56130=>"100000000",
  56131=>"001111111",
  56132=>"000000000",
  56133=>"000000000",
  56134=>"111000000",
  56135=>"000001000",
  56136=>"000010011",
  56137=>"000110111",
  56138=>"100000000",
  56139=>"100111100",
  56140=>"001001001",
  56141=>"110000000",
  56142=>"000000000",
  56143=>"111111111",
  56144=>"101100100",
  56145=>"001011011",
  56146=>"000000011",
  56147=>"000001011",
  56148=>"100000000",
  56149=>"011001011",
  56150=>"000100111",
  56151=>"100111111",
  56152=>"000000000",
  56153=>"000000000",
  56154=>"111001001",
  56155=>"111100100",
  56156=>"010111111",
  56157=>"111111111",
  56158=>"000000111",
  56159=>"100101000",
  56160=>"111111111",
  56161=>"000111111",
  56162=>"010010010",
  56163=>"000000000",
  56164=>"111111111",
  56165=>"001000000",
  56166=>"011111111",
  56167=>"001011111",
  56168=>"001001000",
  56169=>"110000011",
  56170=>"000000000",
  56171=>"000000000",
  56172=>"111111001",
  56173=>"101001101",
  56174=>"100100000",
  56175=>"111111111",
  56176=>"000000000",
  56177=>"000000111",
  56178=>"000111111",
  56179=>"000100111",
  56180=>"111111000",
  56181=>"011110000",
  56182=>"110110110",
  56183=>"100110000",
  56184=>"111111111",
  56185=>"000000000",
  56186=>"000101100",
  56187=>"101110111",
  56188=>"111001000",
  56189=>"000000000",
  56190=>"000000110",
  56191=>"000000000",
  56192=>"010000100",
  56193=>"111111100",
  56194=>"011010110",
  56195=>"111111111",
  56196=>"111111111",
  56197=>"000000000",
  56198=>"000001111",
  56199=>"101111111",
  56200=>"000000111",
  56201=>"010111111",
  56202=>"011010011",
  56203=>"111111110",
  56204=>"111111111",
  56205=>"000000000",
  56206=>"000010110",
  56207=>"010000000",
  56208=>"000000010",
  56209=>"000000001",
  56210=>"000010111",
  56211=>"000000000",
  56212=>"000000000",
  56213=>"110110111",
  56214=>"001000000",
  56215=>"011000000",
  56216=>"000111111",
  56217=>"111101000",
  56218=>"000000000",
  56219=>"001000101",
  56220=>"111000000",
  56221=>"111101111",
  56222=>"111100101",
  56223=>"110011001",
  56224=>"111110111",
  56225=>"111111111",
  56226=>"000000000",
  56227=>"111111110",
  56228=>"111100100",
  56229=>"100000000",
  56230=>"000000000",
  56231=>"000000000",
  56232=>"111111111",
  56233=>"000001001",
  56234=>"000011111",
  56235=>"110000000",
  56236=>"000000000",
  56237=>"111111111",
  56238=>"111111011",
  56239=>"100000100",
  56240=>"111111100",
  56241=>"100010000",
  56242=>"000000101",
  56243=>"000001000",
  56244=>"101111111",
  56245=>"111101101",
  56246=>"000011011",
  56247=>"100110110",
  56248=>"111111011",
  56249=>"000001101",
  56250=>"100111111",
  56251=>"001101111",
  56252=>"000000000",
  56253=>"111111110",
  56254=>"111111011",
  56255=>"011001000",
  56256=>"110000000",
  56257=>"000000000",
  56258=>"000000010",
  56259=>"111111111",
  56260=>"011011001",
  56261=>"100100111",
  56262=>"100110111",
  56263=>"000111011",
  56264=>"000110000",
  56265=>"111110000",
  56266=>"000100111",
  56267=>"000000000",
  56268=>"100000000",
  56269=>"111111111",
  56270=>"000110110",
  56271=>"111010000",
  56272=>"111011111",
  56273=>"111101001",
  56274=>"000000000",
  56275=>"000000000",
  56276=>"111010010",
  56277=>"000110111",
  56278=>"000000000",
  56279=>"111000101",
  56280=>"100101111",
  56281=>"111111111",
  56282=>"111111111",
  56283=>"111111111",
  56284=>"100101001",
  56285=>"000000110",
  56286=>"100111011",
  56287=>"111011111",
  56288=>"000000000",
  56289=>"000000100",
  56290=>"100100111",
  56291=>"000000100",
  56292=>"111111111",
  56293=>"000000000",
  56294=>"001111100",
  56295=>"011000001",
  56296=>"001000110",
  56297=>"000111110",
  56298=>"111000000",
  56299=>"111110000",
  56300=>"000011001",
  56301=>"100100110",
  56302=>"001000000",
  56303=>"111000000",
  56304=>"000000000",
  56305=>"111111101",
  56306=>"111100000",
  56307=>"000111011",
  56308=>"100000000",
  56309=>"111111101",
  56310=>"111111111",
  56311=>"011000000",
  56312=>"000000000",
  56313=>"101100110",
  56314=>"111111011",
  56315=>"000000000",
  56316=>"001100000",
  56317=>"000000011",
  56318=>"000000000",
  56319=>"001000000",
  56320=>"011011011",
  56321=>"111000000",
  56322=>"111111010",
  56323=>"111000011",
  56324=>"010000110",
  56325=>"100010010",
  56326=>"001000000",
  56327=>"111111111",
  56328=>"000000000",
  56329=>"011100000",
  56330=>"000000110",
  56331=>"111000010",
  56332=>"000000000",
  56333=>"111000100",
  56334=>"000000111",
  56335=>"000000000",
  56336=>"111010000",
  56337=>"011111000",
  56338=>"010000000",
  56339=>"111111111",
  56340=>"000111111",
  56341=>"000111000",
  56342=>"000100111",
  56343=>"000010100",
  56344=>"111111111",
  56345=>"111111110",
  56346=>"111111001",
  56347=>"011010011",
  56348=>"000000111",
  56349=>"000110111",
  56350=>"110111111",
  56351=>"111110000",
  56352=>"000000000",
  56353=>"000000111",
  56354=>"110100000",
  56355=>"000000110",
  56356=>"111011000",
  56357=>"111111000",
  56358=>"000000000",
  56359=>"000000101",
  56360=>"111111111",
  56361=>"000000000",
  56362=>"111111111",
  56363=>"000111111",
  56364=>"110110110",
  56365=>"010000111",
  56366=>"101001100",
  56367=>"001100111",
  56368=>"000010000",
  56369=>"111110100",
  56370=>"010010011",
  56371=>"000000011",
  56372=>"000000111",
  56373=>"000011011",
  56374=>"111111000",
  56375=>"000000000",
  56376=>"000000000",
  56377=>"000000001",
  56378=>"000000000",
  56379=>"111111111",
  56380=>"000000000",
  56381=>"000010111",
  56382=>"000001100",
  56383=>"111001011",
  56384=>"001000100",
  56385=>"101111110",
  56386=>"111111111",
  56387=>"111111111",
  56388=>"011000000",
  56389=>"001111111",
  56390=>"111110011",
  56391=>"000000000",
  56392=>"000000111",
  56393=>"000010011",
  56394=>"001101000",
  56395=>"011000101",
  56396=>"000000110",
  56397=>"110111111",
  56398=>"000100111",
  56399=>"000001011",
  56400=>"000000001",
  56401=>"000011110",
  56402=>"111111011",
  56403=>"010001110",
  56404=>"000000000",
  56405=>"111111000",
  56406=>"000000100",
  56407=>"000111111",
  56408=>"111111000",
  56409=>"000000101",
  56410=>"111101111",
  56411=>"111001001",
  56412=>"111111000",
  56413=>"111111011",
  56414=>"000000100",
  56415=>"110010110",
  56416=>"000000111",
  56417=>"111000100",
  56418=>"000000011",
  56419=>"011001111",
  56420=>"000000100",
  56421=>"111000000",
  56422=>"111000000",
  56423=>"000000000",
  56424=>"000000101",
  56425=>"010110111",
  56426=>"000000111",
  56427=>"011111000",
  56428=>"000011111",
  56429=>"000000000",
  56430=>"111011001",
  56431=>"010110110",
  56432=>"000000111",
  56433=>"000000000",
  56434=>"101101111",
  56435=>"110000000",
  56436=>"000010000",
  56437=>"011111111",
  56438=>"010000000",
  56439=>"000000000",
  56440=>"010000000",
  56441=>"000111001",
  56442=>"111000000",
  56443=>"111000000",
  56444=>"000001011",
  56445=>"000000000",
  56446=>"111000000",
  56447=>"000101101",
  56448=>"110000000",
  56449=>"000000110",
  56450=>"110110111",
  56451=>"000000000",
  56452=>"000000000",
  56453=>"111001100",
  56454=>"111111111",
  56455=>"010011011",
  56456=>"011001000",
  56457=>"011011001",
  56458=>"111000000",
  56459=>"000000010",
  56460=>"111110010",
  56461=>"111000000",
  56462=>"111111111",
  56463=>"111111100",
  56464=>"111111111",
  56465=>"000000111",
  56466=>"111111000",
  56467=>"100110000",
  56468=>"000000000",
  56469=>"100010110",
  56470=>"111111001",
  56471=>"111001111",
  56472=>"000000110",
  56473=>"111000000",
  56474=>"000000000",
  56475=>"000000001",
  56476=>"111111000",
  56477=>"111000000",
  56478=>"100000111",
  56479=>"111110000",
  56480=>"000111111",
  56481=>"111111111",
  56482=>"000011000",
  56483=>"001000000",
  56484=>"000000000",
  56485=>"111111110",
  56486=>"000111111",
  56487=>"100100111",
  56488=>"000000111",
  56489=>"010111111",
  56490=>"111100000",
  56491=>"111010011",
  56492=>"111111101",
  56493=>"110111100",
  56494=>"011000001",
  56495=>"111111000",
  56496=>"000111000",
  56497=>"111111011",
  56498=>"111111111",
  56499=>"111111111",
  56500=>"111111011",
  56501=>"000000000",
  56502=>"111111000",
  56503=>"000000101",
  56504=>"000111111",
  56505=>"000111111",
  56506=>"000001001",
  56507=>"000000111",
  56508=>"000000001",
  56509=>"111111001",
  56510=>"000000110",
  56511=>"111110000",
  56512=>"000000000",
  56513=>"000001111",
  56514=>"011001001",
  56515=>"000111111",
  56516=>"010111111",
  56517=>"101101111",
  56518=>"000000001",
  56519=>"010110010",
  56520=>"111111000",
  56521=>"000000000",
  56522=>"111000001",
  56523=>"000000111",
  56524=>"000000001",
  56525=>"100111111",
  56526=>"000000000",
  56527=>"000000000",
  56528=>"111000001",
  56529=>"110111111",
  56530=>"000010001",
  56531=>"000000000",
  56532=>"000000000",
  56533=>"111111111",
  56534=>"000000111",
  56535=>"000000011",
  56536=>"000111000",
  56537=>"000000100",
  56538=>"000000111",
  56539=>"011111000",
  56540=>"111111111",
  56541=>"001001111",
  56542=>"000010000",
  56543=>"010000100",
  56544=>"000000000",
  56545=>"000011000",
  56546=>"100000000",
  56547=>"101100000",
  56548=>"111111101",
  56549=>"000000100",
  56550=>"111011011",
  56551=>"100110111",
  56552=>"111111111",
  56553=>"000101111",
  56554=>"000100111",
  56555=>"010010011",
  56556=>"111010000",
  56557=>"000000000",
  56558=>"111111111",
  56559=>"111111100",
  56560=>"100000010",
  56561=>"101111001",
  56562=>"000111111",
  56563=>"000000010",
  56564=>"111111000",
  56565=>"001000111",
  56566=>"111111000",
  56567=>"010011001",
  56568=>"000110111",
  56569=>"111111001",
  56570=>"000000000",
  56571=>"000000000",
  56572=>"001001011",
  56573=>"111011111",
  56574=>"000000001",
  56575=>"111111111",
  56576=>"000000111",
  56577=>"000000111",
  56578=>"110111011",
  56579=>"000001001",
  56580=>"111111000",
  56581=>"000111000",
  56582=>"000111111",
  56583=>"110110111",
  56584=>"000000000",
  56585=>"000000111",
  56586=>"111111011",
  56587=>"000000010",
  56588=>"011001001",
  56589=>"000000111",
  56590=>"111111010",
  56591=>"111001000",
  56592=>"110110100",
  56593=>"000000000",
  56594=>"111111001",
  56595=>"001000000",
  56596=>"000000000",
  56597=>"011001000",
  56598=>"000000001",
  56599=>"111000000",
  56600=>"001001000",
  56601=>"000000000",
  56602=>"111000000",
  56603=>"100000000",
  56604=>"000000111",
  56605=>"111110000",
  56606=>"111111111",
  56607=>"000000000",
  56608=>"100100001",
  56609=>"111011010",
  56610=>"000000001",
  56611=>"111111111",
  56612=>"000010110",
  56613=>"000000001",
  56614=>"000000100",
  56615=>"101101101",
  56616=>"111111110",
  56617=>"000000000",
  56618=>"000000111",
  56619=>"000000111",
  56620=>"000000111",
  56621=>"000001001",
  56622=>"000000111",
  56623=>"000000111",
  56624=>"110111010",
  56625=>"000000010",
  56626=>"000111111",
  56627=>"101111011",
  56628=>"000011000",
  56629=>"000001001",
  56630=>"111111010",
  56631=>"000000001",
  56632=>"110111000",
  56633=>"000001000",
  56634=>"011011000",
  56635=>"001000000",
  56636=>"111111000",
  56637=>"111111001",
  56638=>"110110101",
  56639=>"111110101",
  56640=>"111000000",
  56641=>"111110111",
  56642=>"011111111",
  56643=>"111000101",
  56644=>"111111111",
  56645=>"111110111",
  56646=>"000011111",
  56647=>"001101110",
  56648=>"000111111",
  56649=>"000110111",
  56650=>"000000001",
  56651=>"000011111",
  56652=>"111110000",
  56653=>"111010011",
  56654=>"000110111",
  56655=>"111001100",
  56656=>"011011011",
  56657=>"111000100",
  56658=>"000110111",
  56659=>"111101101",
  56660=>"000000111",
  56661=>"001100010",
  56662=>"000000001",
  56663=>"111111001",
  56664=>"000000111",
  56665=>"000000111",
  56666=>"111111111",
  56667=>"000000110",
  56668=>"011011001",
  56669=>"110111000",
  56670=>"111000000",
  56671=>"000000000",
  56672=>"100000000",
  56673=>"111111000",
  56674=>"101011011",
  56675=>"111000000",
  56676=>"000011111",
  56677=>"000000000",
  56678=>"011010000",
  56679=>"110111110",
  56680=>"100100111",
  56681=>"000100000",
  56682=>"000000000",
  56683=>"110001101",
  56684=>"000011000",
  56685=>"000011001",
  56686=>"000000000",
  56687=>"111111111",
  56688=>"111010000",
  56689=>"111101000",
  56690=>"000000111",
  56691=>"001111111",
  56692=>"011011000",
  56693=>"100000010",
  56694=>"111111100",
  56695=>"111111000",
  56696=>"000000111",
  56697=>"000110111",
  56698=>"111011000",
  56699=>"111000111",
  56700=>"011000111",
  56701=>"111111111",
  56702=>"001010111",
  56703=>"000011001",
  56704=>"110111011",
  56705=>"111111111",
  56706=>"100111111",
  56707=>"000111111",
  56708=>"010010000",
  56709=>"000100000",
  56710=>"000111111",
  56711=>"000001110",
  56712=>"111111111",
  56713=>"110100000",
  56714=>"111000000",
  56715=>"000111111",
  56716=>"111111110",
  56717=>"001011001",
  56718=>"000000000",
  56719=>"111001000",
  56720=>"010111111",
  56721=>"011001000",
  56722=>"011011000",
  56723=>"111111111",
  56724=>"000000000",
  56725=>"000000000",
  56726=>"000000111",
  56727=>"000000000",
  56728=>"111111000",
  56729=>"111101000",
  56730=>"111111000",
  56731=>"100111111",
  56732=>"000010110",
  56733=>"011011111",
  56734=>"011000001",
  56735=>"110110111",
  56736=>"011111110",
  56737=>"110100010",
  56738=>"001000101",
  56739=>"011111111",
  56740=>"000100111",
  56741=>"110100000",
  56742=>"011111001",
  56743=>"111111000",
  56744=>"000100000",
  56745=>"110111010",
  56746=>"000000000",
  56747=>"000000001",
  56748=>"000111110",
  56749=>"000000000",
  56750=>"111111110",
  56751=>"000000000",
  56752=>"111000000",
  56753=>"111111011",
  56754=>"111000000",
  56755=>"000111110",
  56756=>"000111011",
  56757=>"000000011",
  56758=>"111111111",
  56759=>"000000011",
  56760=>"111111111",
  56761=>"111111111",
  56762=>"000110110",
  56763=>"000000000",
  56764=>"000111111",
  56765=>"111111111",
  56766=>"100101111",
  56767=>"110100001",
  56768=>"100100111",
  56769=>"000000011",
  56770=>"111111111",
  56771=>"111111111",
  56772=>"101100110",
  56773=>"010000101",
  56774=>"111111111",
  56775=>"000000000",
  56776=>"111111011",
  56777=>"101100000",
  56778=>"000000111",
  56779=>"111111111",
  56780=>"111111001",
  56781=>"111000000",
  56782=>"000000110",
  56783=>"111111111",
  56784=>"111111000",
  56785=>"111111100",
  56786=>"111001011",
  56787=>"000110111",
  56788=>"011100110",
  56789=>"111111111",
  56790=>"000000111",
  56791=>"000000010",
  56792=>"100000011",
  56793=>"000000110",
  56794=>"000000000",
  56795=>"111111111",
  56796=>"000000000",
  56797=>"100100100",
  56798=>"011011111",
  56799=>"111110100",
  56800=>"000000111",
  56801=>"000000000",
  56802=>"110111000",
  56803=>"111111110",
  56804=>"110110111",
  56805=>"111000111",
  56806=>"111001000",
  56807=>"000000000",
  56808=>"000111111",
  56809=>"011111111",
  56810=>"000010000",
  56811=>"110101000",
  56812=>"111101111",
  56813=>"001011000",
  56814=>"111111111",
  56815=>"000000010",
  56816=>"011000000",
  56817=>"000111111",
  56818=>"111000101",
  56819=>"000000111",
  56820=>"111110000",
  56821=>"000000110",
  56822=>"000011011",
  56823=>"000001000",
  56824=>"110000000",
  56825=>"001001000",
  56826=>"111111000",
  56827=>"111111000",
  56828=>"000001111",
  56829=>"011001001",
  56830=>"000000000",
  56831=>"000111111",
  56832=>"100000000",
  56833=>"100000000",
  56834=>"110010000",
  56835=>"111000000",
  56836=>"000000000",
  56837=>"000000000",
  56838=>"110111111",
  56839=>"111110111",
  56840=>"111111000",
  56841=>"111111000",
  56842=>"001111110",
  56843=>"111111111",
  56844=>"111111111",
  56845=>"000011000",
  56846=>"001101111",
  56847=>"011000000",
  56848=>"100100000",
  56849=>"000001011",
  56850=>"000000000",
  56851=>"000000010",
  56852=>"111111111",
  56853=>"011111000",
  56854=>"111111000",
  56855=>"110110100",
  56856=>"111000000",
  56857=>"000000010",
  56858=>"000111111",
  56859=>"111011001",
  56860=>"100111111",
  56861=>"001000100",
  56862=>"000001001",
  56863=>"111111111",
  56864=>"010000000",
  56865=>"000000000",
  56866=>"011111111",
  56867=>"111111100",
  56868=>"000111111",
  56869=>"111111000",
  56870=>"111110110",
  56871=>"111000000",
  56872=>"000000000",
  56873=>"111000110",
  56874=>"111000101",
  56875=>"111111111",
  56876=>"000000101",
  56877=>"111000000",
  56878=>"000000000",
  56879=>"101011001",
  56880=>"000000000",
  56881=>"100000000",
  56882=>"000000100",
  56883=>"111011001",
  56884=>"000000111",
  56885=>"100111111",
  56886=>"111111000",
  56887=>"011001001",
  56888=>"001000000",
  56889=>"001000000",
  56890=>"011000000",
  56891=>"000111111",
  56892=>"111111111",
  56893=>"001001111",
  56894=>"111100111",
  56895=>"111111111",
  56896=>"111010110",
  56897=>"000110100",
  56898=>"100000000",
  56899=>"110000000",
  56900=>"000000000",
  56901=>"000000110",
  56902=>"101101010",
  56903=>"011000000",
  56904=>"111111110",
  56905=>"111111100",
  56906=>"000000000",
  56907=>"001011111",
  56908=>"001001111",
  56909=>"001111010",
  56910=>"000000011",
  56911=>"111111111",
  56912=>"000000111",
  56913=>"001000000",
  56914=>"000000111",
  56915=>"110110000",
  56916=>"111110101",
  56917=>"000000000",
  56918=>"111111100",
  56919=>"110000000",
  56920=>"111000000",
  56921=>"111001111",
  56922=>"000000000",
  56923=>"000001011",
  56924=>"110100111",
  56925=>"000000100",
  56926=>"111111110",
  56927=>"111100100",
  56928=>"111111101",
  56929=>"000000111",
  56930=>"000000111",
  56931=>"000000000",
  56932=>"010110110",
  56933=>"000101000",
  56934=>"001001111",
  56935=>"000111111",
  56936=>"000110010",
  56937=>"111111111",
  56938=>"000000000",
  56939=>"111000000",
  56940=>"111111111",
  56941=>"111111111",
  56942=>"111111100",
  56943=>"111111111",
  56944=>"000000000",
  56945=>"001011000",
  56946=>"000111111",
  56947=>"110111111",
  56948=>"000000000",
  56949=>"000000110",
  56950=>"111111111",
  56951=>"000000011",
  56952=>"110110110",
  56953=>"111111110",
  56954=>"000111111",
  56955=>"000000110",
  56956=>"100100111",
  56957=>"111111111",
  56958=>"110000000",
  56959=>"111111101",
  56960=>"111111000",
  56961=>"111000100",
  56962=>"111000000",
  56963=>"110110000",
  56964=>"001001111",
  56965=>"000000000",
  56966=>"001111111",
  56967=>"011111110",
  56968=>"001000000",
  56969=>"111000000",
  56970=>"101111111",
  56971=>"111111000",
  56972=>"000000000",
  56973=>"000000000",
  56974=>"001111001",
  56975=>"000000111",
  56976=>"000000000",
  56977=>"000000000",
  56978=>"111111111",
  56979=>"000000111",
  56980=>"100000000",
  56981=>"000000101",
  56982=>"111111111",
  56983=>"111111000",
  56984=>"110000110",
  56985=>"000100100",
  56986=>"100000000",
  56987=>"000111110",
  56988=>"111111111",
  56989=>"110000110",
  56990=>"000111100",
  56991=>"111000000",
  56992=>"100111111",
  56993=>"101100000",
  56994=>"000000000",
  56995=>"000111000",
  56996=>"101101100",
  56997=>"001001001",
  56998=>"000000000",
  56999=>"000001111",
  57000=>"100000111",
  57001=>"100000000",
  57002=>"111111000",
  57003=>"111111111",
  57004=>"111011111",
  57005=>"100001011",
  57006=>"111000010",
  57007=>"111111111",
  57008=>"111111111",
  57009=>"001001001",
  57010=>"000110111",
  57011=>"111101000",
  57012=>"100111100",
  57013=>"000000111",
  57014=>"000000011",
  57015=>"000101001",
  57016=>"101001100",
  57017=>"000000111",
  57018=>"000100111",
  57019=>"110110111",
  57020=>"001101111",
  57021=>"111000000",
  57022=>"110111111",
  57023=>"111111000",
  57024=>"111110100",
  57025=>"111111110",
  57026=>"001000110",
  57027=>"111111111",
  57028=>"111111110",
  57029=>"000001001",
  57030=>"000000000",
  57031=>"010000111",
  57032=>"110111111",
  57033=>"111111111",
  57034=>"110100000",
  57035=>"111111111",
  57036=>"000111111",
  57037=>"000000111",
  57038=>"111111111",
  57039=>"101000111",
  57040=>"111111000",
  57041=>"110111111",
  57042=>"111110111",
  57043=>"000110111",
  57044=>"111000000",
  57045=>"000011111",
  57046=>"111111111",
  57047=>"000000110",
  57048=>"000000110",
  57049=>"000000110",
  57050=>"111011010",
  57051=>"000010110",
  57052=>"111111101",
  57053=>"111000000",
  57054=>"000000011",
  57055=>"111011000",
  57056=>"000000001",
  57057=>"000011001",
  57058=>"000111111",
  57059=>"111000010",
  57060=>"100111111",
  57061=>"001010100",
  57062=>"000000111",
  57063=>"000000001",
  57064=>"000000100",
  57065=>"000000000",
  57066=>"111000111",
  57067=>"100000000",
  57068=>"111001000",
  57069=>"111001111",
  57070=>"000110111",
  57071=>"010000000",
  57072=>"111110000",
  57073=>"111111010",
  57074=>"000000001",
  57075=>"110111111",
  57076=>"110110010",
  57077=>"111001101",
  57078=>"001001001",
  57079=>"000111111",
  57080=>"000111111",
  57081=>"001000111",
  57082=>"000000000",
  57083=>"000000000",
  57084=>"000111000",
  57085=>"111111111",
  57086=>"000000000",
  57087=>"111111111",
  57088=>"000111110",
  57089=>"011011011",
  57090=>"110000000",
  57091=>"000000000",
  57092=>"001011100",
  57093=>"000110110",
  57094=>"101011011",
  57095=>"111111100",
  57096=>"111111101",
  57097=>"111000000",
  57098=>"000000000",
  57099=>"111011000",
  57100=>"110000111",
  57101=>"000000110",
  57102=>"111111111",
  57103=>"000111111",
  57104=>"001000000",
  57105=>"001001111",
  57106=>"111111000",
  57107=>"000000000",
  57108=>"111000000",
  57109=>"001001011",
  57110=>"000110111",
  57111=>"111111000",
  57112=>"000000000",
  57113=>"111110000",
  57114=>"111011000",
  57115=>"111111010",
  57116=>"000000000",
  57117=>"000000000",
  57118=>"011000000",
  57119=>"100000110",
  57120=>"000000111",
  57121=>"100000111",
  57122=>"111111111",
  57123=>"101111110",
  57124=>"000110110",
  57125=>"000001111",
  57126=>"001001111",
  57127=>"000000000",
  57128=>"001011011",
  57129=>"101001001",
  57130=>"100000111",
  57131=>"111101111",
  57132=>"100100100",
  57133=>"000001000",
  57134=>"000000000",
  57135=>"111000011",
  57136=>"010110110",
  57137=>"001000000",
  57138=>"111111111",
  57139=>"111100000",
  57140=>"111111110",
  57141=>"111111111",
  57142=>"011000100",
  57143=>"010000000",
  57144=>"111111000",
  57145=>"000000101",
  57146=>"000000000",
  57147=>"010111111",
  57148=>"000001100",
  57149=>"000000111",
  57150=>"000000000",
  57151=>"000111111",
  57152=>"111101000",
  57153=>"010110000",
  57154=>"000000000",
  57155=>"101000000",
  57156=>"001001000",
  57157=>"000000000",
  57158=>"111110111",
  57159=>"111000000",
  57160=>"010000000",
  57161=>"111000000",
  57162=>"111111011",
  57163=>"001001111",
  57164=>"000111110",
  57165=>"000111111",
  57166=>"111000000",
  57167=>"100111111",
  57168=>"001000000",
  57169=>"101100000",
  57170=>"101000111",
  57171=>"000000111",
  57172=>"011111010",
  57173=>"001101111",
  57174=>"111001001",
  57175=>"111011111",
  57176=>"111000001",
  57177=>"111000000",
  57178=>"110010111",
  57179=>"000000100",
  57180=>"000000111",
  57181=>"111111111",
  57182=>"100011011",
  57183=>"000101111",
  57184=>"011000101",
  57185=>"000011010",
  57186=>"000000111",
  57187=>"000000010",
  57188=>"000000001",
  57189=>"100000010",
  57190=>"001111100",
  57191=>"011111100",
  57192=>"111110100",
  57193=>"000000110",
  57194=>"000000000",
  57195=>"111111011",
  57196=>"100110100",
  57197=>"001001001",
  57198=>"111111110",
  57199=>"110110000",
  57200=>"000000000",
  57201=>"000000000",
  57202=>"111111111",
  57203=>"001011001",
  57204=>"010110000",
  57205=>"111011111",
  57206=>"010000000",
  57207=>"111001001",
  57208=>"000000000",
  57209=>"000110111",
  57210=>"110101111",
  57211=>"111111111",
  57212=>"011000000",
  57213=>"000000000",
  57214=>"111111100",
  57215=>"010111111",
  57216=>"000100000",
  57217=>"000000010",
  57218=>"000000111",
  57219=>"000001100",
  57220=>"000111111",
  57221=>"011010000",
  57222=>"000011000",
  57223=>"111110000",
  57224=>"111111111",
  57225=>"000000000",
  57226=>"000000100",
  57227=>"111111111",
  57228=>"111111101",
  57229=>"000001001",
  57230=>"000000000",
  57231=>"111111110",
  57232=>"000000110",
  57233=>"000000000",
  57234=>"111110111",
  57235=>"000000000",
  57236=>"000111111",
  57237=>"010000000",
  57238=>"110001000",
  57239=>"110100000",
  57240=>"110111111",
  57241=>"111101000",
  57242=>"110100111",
  57243=>"111111111",
  57244=>"000000000",
  57245=>"000000000",
  57246=>"000100100",
  57247=>"000000000",
  57248=>"001001000",
  57249=>"011010000",
  57250=>"111111100",
  57251=>"111000000",
  57252=>"101101000",
  57253=>"000000000",
  57254=>"111001000",
  57255=>"111100111",
  57256=>"100000000",
  57257=>"000000000",
  57258=>"111101000",
  57259=>"111111111",
  57260=>"110000000",
  57261=>"000000001",
  57262=>"001111100",
  57263=>"000000000",
  57264=>"101000100",
  57265=>"110100000",
  57266=>"110101000",
  57267=>"111000101",
  57268=>"000000111",
  57269=>"100000110",
  57270=>"000111111",
  57271=>"000111111",
  57272=>"000110111",
  57273=>"111111111",
  57274=>"000000000",
  57275=>"111111000",
  57276=>"111001000",
  57277=>"001000000",
  57278=>"000000000",
  57279=>"111111111",
  57280=>"111111000",
  57281=>"111111000",
  57282=>"000000000",
  57283=>"111111111",
  57284=>"111000000",
  57285=>"000000100",
  57286=>"011001011",
  57287=>"110000000",
  57288=>"111000100",
  57289=>"110111010",
  57290=>"111110110",
  57291=>"001000000",
  57292=>"000000111",
  57293=>"111111111",
  57294=>"010111111",
  57295=>"111111000",
  57296=>"000000000",
  57297=>"000111111",
  57298=>"110111111",
  57299=>"001000111",
  57300=>"000000001",
  57301=>"001000000",
  57302=>"000110111",
  57303=>"101111110",
  57304=>"001111110",
  57305=>"000000111",
  57306=>"001000000",
  57307=>"011000000",
  57308=>"000000000",
  57309=>"111111111",
  57310=>"111000110",
  57311=>"011011011",
  57312=>"000000111",
  57313=>"000000000",
  57314=>"111111111",
  57315=>"000000000",
  57316=>"110111011",
  57317=>"001111110",
  57318=>"111111111",
  57319=>"111000000",
  57320=>"000000000",
  57321=>"000000000",
  57322=>"000100000",
  57323=>"111111000",
  57324=>"110110111",
  57325=>"001011110",
  57326=>"110000000",
  57327=>"100111111",
  57328=>"110000111",
  57329=>"000100111",
  57330=>"100111000",
  57331=>"110111111",
  57332=>"000000000",
  57333=>"011011000",
  57334=>"101001000",
  57335=>"110100001",
  57336=>"000000111",
  57337=>"101111001",
  57338=>"000000000",
  57339=>"111111110",
  57340=>"000000111",
  57341=>"110100000",
  57342=>"111111111",
  57343=>"100111111",
  57344=>"000111111",
  57345=>"110000000",
  57346=>"111111111",
  57347=>"111111000",
  57348=>"000111111",
  57349=>"100101111",
  57350=>"000010000",
  57351=>"000000000",
  57352=>"100100111",
  57353=>"000001000",
  57354=>"111110100",
  57355=>"111111011",
  57356=>"000000000",
  57357=>"111110100",
  57358=>"111111011",
  57359=>"011011000",
  57360=>"000000111",
  57361=>"111111011",
  57362=>"000000111",
  57363=>"000000111",
  57364=>"111000111",
  57365=>"111111100",
  57366=>"111111100",
  57367=>"111111111",
  57368=>"111111111",
  57369=>"011011000",
  57370=>"101000000",
  57371=>"001001011",
  57372=>"000110100",
  57373=>"111110000",
  57374=>"111110100",
  57375=>"000100110",
  57376=>"111111001",
  57377=>"010110100",
  57378=>"000000100",
  57379=>"000000100",
  57380=>"000000000",
  57381=>"000000110",
  57382=>"101111100",
  57383=>"011111111",
  57384=>"000001101",
  57385=>"000001000",
  57386=>"111111111",
  57387=>"001000000",
  57388=>"001001000",
  57389=>"111111111",
  57390=>"001001001",
  57391=>"110010111",
  57392=>"000000111",
  57393=>"000000000",
  57394=>"111011000",
  57395=>"000000000",
  57396=>"001000000",
  57397=>"010010000",
  57398=>"000000011",
  57399=>"000001111",
  57400=>"111111011",
  57401=>"111000000",
  57402=>"000000000",
  57403=>"100000000",
  57404=>"000000000",
  57405=>"111100111",
  57406=>"111110100",
  57407=>"111111111",
  57408=>"000111111",
  57409=>"100100000",
  57410=>"111100000",
  57411=>"011110111",
  57412=>"110110110",
  57413=>"000000110",
  57414=>"010000010",
  57415=>"111111111",
  57416=>"110110110",
  57417=>"111111111",
  57418=>"001000000",
  57419=>"001000000",
  57420=>"100000011",
  57421=>"000000000",
  57422=>"110110111",
  57423=>"101000000",
  57424=>"110001000",
  57425=>"101111111",
  57426=>"000000000",
  57427=>"111000000",
  57428=>"001000000",
  57429=>"000010000",
  57430=>"001001000",
  57431=>"000001111",
  57432=>"011111111",
  57433=>"000100110",
  57434=>"100000000",
  57435=>"001001001",
  57436=>"000000000",
  57437=>"000000000",
  57438=>"011010100",
  57439=>"100000000",
  57440=>"110111010",
  57441=>"000000000",
  57442=>"110111100",
  57443=>"111101111",
  57444=>"011111111",
  57445=>"001001000",
  57446=>"000000000",
  57447=>"110110111",
  57448=>"000000000",
  57449=>"000000000",
  57450=>"000000000",
  57451=>"111111111",
  57452=>"011011011",
  57453=>"000000000",
  57454=>"111111111",
  57455=>"011011000",
  57456=>"010111000",
  57457=>"011111111",
  57458=>"111111100",
  57459=>"111110111",
  57460=>"111011011",
  57461=>"000001001",
  57462=>"000000000",
  57463=>"011011011",
  57464=>"011111111",
  57465=>"000110010",
  57466=>"111111111",
  57467=>"111111111",
  57468=>"111110110",
  57469=>"100000000",
  57470=>"111111111",
  57471=>"011000000",
  57472=>"000011011",
  57473=>"000000000",
  57474=>"111111000",
  57475=>"000000101",
  57476=>"111111111",
  57477=>"000000000",
  57478=>"000000000",
  57479=>"011011110",
  57480=>"000110101",
  57481=>"011011011",
  57482=>"001000100",
  57483=>"000000000",
  57484=>"001011111",
  57485=>"000100110",
  57486=>"111111111",
  57487=>"110110000",
  57488=>"111100111",
  57489=>"111111111",
  57490=>"000000000",
  57491=>"111111111",
  57492=>"000000001",
  57493=>"000000000",
  57494=>"111111111",
  57495=>"111000000",
  57496=>"110000000",
  57497=>"011010100",
  57498=>"000000111",
  57499=>"111111110",
  57500=>"011001110",
  57501=>"010000000",
  57502=>"111111111",
  57503=>"100111111",
  57504=>"110000011",
  57505=>"111000000",
  57506=>"111111111",
  57507=>"010000000",
  57508=>"111011011",
  57509=>"000000011",
  57510=>"101000000",
  57511=>"100100100",
  57512=>"000000000",
  57513=>"000000000",
  57514=>"110000000",
  57515=>"110111111",
  57516=>"111011111",
  57517=>"111111111",
  57518=>"000010000",
  57519=>"000000000",
  57520=>"000000000",
  57521=>"000000010",
  57522=>"111111111",
  57523=>"111101101",
  57524=>"110111110",
  57525=>"111000111",
  57526=>"000000000",
  57527=>"111111100",
  57528=>"111010000",
  57529=>"000000111",
  57530=>"001000000",
  57531=>"000000111",
  57532=>"000000000",
  57533=>"011111111",
  57534=>"000000000",
  57535=>"111101101",
  57536=>"000000100",
  57537=>"000000000",
  57538=>"001111111",
  57539=>"110111010",
  57540=>"100111111",
  57541=>"000000001",
  57542=>"000011001",
  57543=>"111111111",
  57544=>"010000000",
  57545=>"111111111",
  57546=>"000000000",
  57547=>"000000100",
  57548=>"111111001",
  57549=>"000000000",
  57550=>"000000000",
  57551=>"111110000",
  57552=>"000000001",
  57553=>"000100111",
  57554=>"010000000",
  57555=>"000000111",
  57556=>"011011111",
  57557=>"110110111",
  57558=>"000000111",
  57559=>"110000000",
  57560=>"111111011",
  57561=>"001000100",
  57562=>"111111010",
  57563=>"000000000",
  57564=>"111000111",
  57565=>"110110000",
  57566=>"100111111",
  57567=>"111011000",
  57568=>"100100000",
  57569=>"000000000",
  57570=>"000000000",
  57571=>"000000000",
  57572=>"010011011",
  57573=>"100000000",
  57574=>"111111101",
  57575=>"000000000",
  57576=>"111111111",
  57577=>"111111100",
  57578=>"111101101",
  57579=>"111011011",
  57580=>"000000000",
  57581=>"000000111",
  57582=>"110110111",
  57583=>"110010101",
  57584=>"111111011",
  57585=>"111111011",
  57586=>"001001011",
  57587=>"011111100",
  57588=>"111000000",
  57589=>"000000000",
  57590=>"001111101",
  57591=>"000011010",
  57592=>"100110111",
  57593=>"000000000",
  57594=>"001111111",
  57595=>"101111111",
  57596=>"001001000",
  57597=>"001000000",
  57598=>"000000000",
  57599=>"010111111",
  57600=>"011001110",
  57601=>"111111011",
  57602=>"110000000",
  57603=>"110000011",
  57604=>"000011111",
  57605=>"000000000",
  57606=>"000000101",
  57607=>"001111111",
  57608=>"000000000",
  57609=>"000000000",
  57610=>"110010111",
  57611=>"111111110",
  57612=>"111111111",
  57613=>"000000000",
  57614=>"011111000",
  57615=>"000000000",
  57616=>"000000110",
  57617=>"000000001",
  57618=>"000000111",
  57619=>"000000000",
  57620=>"111111110",
  57621=>"000110100",
  57622=>"000000000",
  57623=>"110110000",
  57624=>"111111111",
  57625=>"111111001",
  57626=>"110000000",
  57627=>"110100001",
  57628=>"011001111",
  57629=>"000000101",
  57630=>"000000000",
  57631=>"111111100",
  57632=>"111111001",
  57633=>"111111101",
  57634=>"000000000",
  57635=>"000000000",
  57636=>"111011011",
  57637=>"010000000",
  57638=>"010000000",
  57639=>"011011000",
  57640=>"111111111",
  57641=>"111111111",
  57642=>"111111111",
  57643=>"100100100",
  57644=>"101000000",
  57645=>"011111011",
  57646=>"000000000",
  57647=>"000000000",
  57648=>"111011111",
  57649=>"111111000",
  57650=>"000000000",
  57651=>"000000011",
  57652=>"110111110",
  57653=>"111111111",
  57654=>"000000000",
  57655=>"111000000",
  57656=>"111111000",
  57657=>"111111000",
  57658=>"101101110",
  57659=>"000000111",
  57660=>"111100110",
  57661=>"000000110",
  57662=>"000000000",
  57663=>"001001001",
  57664=>"000000000",
  57665=>"111111011",
  57666=>"000000000",
  57667=>"010000011",
  57668=>"000000000",
  57669=>"110000000",
  57670=>"000000000",
  57671=>"110000000",
  57672=>"100100111",
  57673=>"000000000",
  57674=>"111100000",
  57675=>"100110110",
  57676=>"000000000",
  57677=>"011001000",
  57678=>"011000100",
  57679=>"001101010",
  57680=>"000000100",
  57681=>"000110000",
  57682=>"111110000",
  57683=>"111111111",
  57684=>"000100111",
  57685=>"011011011",
  57686=>"101111111",
  57687=>"000001000",
  57688=>"011111111",
  57689=>"111101101",
  57690=>"000001111",
  57691=>"000000000",
  57692=>"000000110",
  57693=>"111111111",
  57694=>"101001000",
  57695=>"000000000",
  57696=>"001111000",
  57697=>"000000011",
  57698=>"011101000",
  57699=>"111111111",
  57700=>"000111111",
  57701=>"000000000",
  57702=>"000000000",
  57703=>"000001001",
  57704=>"011111111",
  57705=>"000010000",
  57706=>"011000000",
  57707=>"000010010",
  57708=>"011011011",
  57709=>"000000000",
  57710=>"000010010",
  57711=>"000000100",
  57712=>"000000100",
  57713=>"000000000",
  57714=>"001001000",
  57715=>"000000000",
  57716=>"111111111",
  57717=>"000000000",
  57718=>"000000000",
  57719=>"000000000",
  57720=>"000000011",
  57721=>"111111000",
  57722=>"000000000",
  57723=>"011000000",
  57724=>"111111001",
  57725=>"000000000",
  57726=>"011111010",
  57727=>"000000000",
  57728=>"111011001",
  57729=>"000000100",
  57730=>"111111111",
  57731=>"000000110",
  57732=>"000011111",
  57733=>"000000000",
  57734=>"010000000",
  57735=>"111111111",
  57736=>"111111111",
  57737=>"010000110",
  57738=>"110110111",
  57739=>"111111011",
  57740=>"111111111",
  57741=>"001001001",
  57742=>"000000110",
  57743=>"000000000",
  57744=>"000000000",
  57745=>"111011111",
  57746=>"111111110",
  57747=>"111111011",
  57748=>"111111000",
  57749=>"000010000",
  57750=>"110110000",
  57751=>"011000000",
  57752=>"111111111",
  57753=>"111000000",
  57754=>"111111111",
  57755=>"111111111",
  57756=>"111110110",
  57757=>"000001001",
  57758=>"111000000",
  57759=>"010111010",
  57760=>"111011011",
  57761=>"111111000",
  57762=>"001011111",
  57763=>"000000000",
  57764=>"000111000",
  57765=>"101110110",
  57766=>"000000111",
  57767=>"111010011",
  57768=>"000100111",
  57769=>"000100100",
  57770=>"001000100",
  57771=>"111111011",
  57772=>"000000110",
  57773=>"000111111",
  57774=>"000000000",
  57775=>"111111000",
  57776=>"111111111",
  57777=>"000111111",
  57778=>"111100101",
  57779=>"000010000",
  57780=>"111111111",
  57781=>"110110110",
  57782=>"100111111",
  57783=>"000000000",
  57784=>"111011000",
  57785=>"000111111",
  57786=>"000000000",
  57787=>"010000111",
  57788=>"111111110",
  57789=>"111111111",
  57790=>"111111100",
  57791=>"001111111",
  57792=>"000000000",
  57793=>"000000000",
  57794=>"001001001",
  57795=>"111111111",
  57796=>"000000000",
  57797=>"100110000",
  57798=>"000000000",
  57799=>"000000000",
  57800=>"111101100",
  57801=>"000000000",
  57802=>"011011000",
  57803=>"000000111",
  57804=>"111000000",
  57805=>"111111111",
  57806=>"111011011",
  57807=>"111111111",
  57808=>"010000110",
  57809=>"000000011",
  57810=>"000000000",
  57811=>"000000000",
  57812=>"001001001",
  57813=>"100000110",
  57814=>"000000000",
  57815=>"000000001",
  57816=>"011111111",
  57817=>"000000000",
  57818=>"001000000",
  57819=>"010110000",
  57820=>"110111111",
  57821=>"111111111",
  57822=>"100100111",
  57823=>"001011010",
  57824=>"001000000",
  57825=>"100001000",
  57826=>"000001001",
  57827=>"000111111",
  57828=>"000000011",
  57829=>"100000000",
  57830=>"111000000",
  57831=>"111111111",
  57832=>"000011011",
  57833=>"001011011",
  57834=>"100111111",
  57835=>"111111010",
  57836=>"100000000",
  57837=>"101100100",
  57838=>"110100000",
  57839=>"001000000",
  57840=>"001000001",
  57841=>"000011011",
  57842=>"000000000",
  57843=>"010010000",
  57844=>"111111111",
  57845=>"000000000",
  57846=>"010011011",
  57847=>"100110000",
  57848=>"000000100",
  57849=>"010000110",
  57850=>"111101000",
  57851=>"111111101",
  57852=>"000000010",
  57853=>"000000000",
  57854=>"000000000",
  57855=>"000000010",
  57856=>"001111111",
  57857=>"111010000",
  57858=>"111000000",
  57859=>"000100110",
  57860=>"111110100",
  57861=>"101111000",
  57862=>"000000000",
  57863=>"000000000",
  57864=>"111111111",
  57865=>"011110101",
  57866=>"000000000",
  57867=>"111111111",
  57868=>"001011111",
  57869=>"001000000",
  57870=>"001000000",
  57871=>"111111111",
  57872=>"111111111",
  57873=>"000000010",
  57874=>"001001000",
  57875=>"000000101",
  57876=>"111111111",
  57877=>"111111011",
  57878=>"101000000",
  57879=>"110110110",
  57880=>"011101101",
  57881=>"111101001",
  57882=>"011000000",
  57883=>"111001000",
  57884=>"000000000",
  57885=>"111111111",
  57886=>"000000011",
  57887=>"000000000",
  57888=>"111111011",
  57889=>"111111110",
  57890=>"011011011",
  57891=>"010110010",
  57892=>"111010000",
  57893=>"111110111",
  57894=>"001111111",
  57895=>"100100000",
  57896=>"000000000",
  57897=>"000000000",
  57898=>"000000000",
  57899=>"010010011",
  57900=>"111100000",
  57901=>"111111111",
  57902=>"111010010",
  57903=>"111111111",
  57904=>"111111111",
  57905=>"000000000",
  57906=>"110110111",
  57907=>"111111111",
  57908=>"000010011",
  57909=>"000000001",
  57910=>"000000001",
  57911=>"110011001",
  57912=>"011011001",
  57913=>"001100110",
  57914=>"000000000",
  57915=>"000000000",
  57916=>"111101101",
  57917=>"000001110",
  57918=>"110100001",
  57919=>"111001001",
  57920=>"000000101",
  57921=>"110100101",
  57922=>"000000000",
  57923=>"111111111",
  57924=>"111110111",
  57925=>"111111111",
  57926=>"111111010",
  57927=>"111111111",
  57928=>"111110110",
  57929=>"111000101",
  57930=>"111111010",
  57931=>"001011110",
  57932=>"000000000",
  57933=>"100100000",
  57934=>"000111111",
  57935=>"111011001",
  57936=>"001001111",
  57937=>"000000110",
  57938=>"000000000",
  57939=>"000100000",
  57940=>"000000110",
  57941=>"111110100",
  57942=>"000001111",
  57943=>"111111111",
  57944=>"000000000",
  57945=>"000000000",
  57946=>"101111111",
  57947=>"110100100",
  57948=>"000000000",
  57949=>"000000000",
  57950=>"110000100",
  57951=>"000000000",
  57952=>"000000000",
  57953=>"011000000",
  57954=>"111111111",
  57955=>"000000111",
  57956=>"001011000",
  57957=>"010010011",
  57958=>"000001111",
  57959=>"101000000",
  57960=>"110111010",
  57961=>"000000000",
  57962=>"001000000",
  57963=>"000001101",
  57964=>"111111110",
  57965=>"111100100",
  57966=>"111111111",
  57967=>"111000000",
  57968=>"111010000",
  57969=>"001000000",
  57970=>"110100000",
  57971=>"011110110",
  57972=>"111111000",
  57973=>"111011000",
  57974=>"011000000",
  57975=>"110100110",
  57976=>"111101101",
  57977=>"011000000",
  57978=>"000001111",
  57979=>"111110000",
  57980=>"110100100",
  57981=>"000000000",
  57982=>"001000101",
  57983=>"000000010",
  57984=>"000111111",
  57985=>"000110111",
  57986=>"000000000",
  57987=>"111111100",
  57988=>"111101111",
  57989=>"000000101",
  57990=>"000100000",
  57991=>"011111000",
  57992=>"111111111",
  57993=>"000000000",
  57994=>"000000000",
  57995=>"111100100",
  57996=>"110000111",
  57997=>"000000000",
  57998=>"111111111",
  57999=>"001001111",
  58000=>"000101000",
  58001=>"110010010",
  58002=>"010000000",
  58003=>"111000000",
  58004=>"111111111",
  58005=>"111000000",
  58006=>"111111000",
  58007=>"111000000",
  58008=>"111110111",
  58009=>"111011000",
  58010=>"111001000",
  58011=>"110110011",
  58012=>"111111111",
  58013=>"011111111",
  58014=>"101101111",
  58015=>"111111111",
  58016=>"111000000",
  58017=>"100000000",
  58018=>"011011001",
  58019=>"111111111",
  58020=>"000110111",
  58021=>"011000000",
  58022=>"111111110",
  58023=>"000000000",
  58024=>"011111111",
  58025=>"000000001",
  58026=>"111000000",
  58027=>"111111111",
  58028=>"111111111",
  58029=>"000000000",
  58030=>"111001000",
  58031=>"000110111",
  58032=>"000111111",
  58033=>"110010110",
  58034=>"111111111",
  58035=>"111101001",
  58036=>"000000001",
  58037=>"111100001",
  58038=>"000011001",
  58039=>"111111111",
  58040=>"111110000",
  58041=>"000111111",
  58042=>"000011111",
  58043=>"000000000",
  58044=>"000000000",
  58045=>"111111111",
  58046=>"111111011",
  58047=>"001001111",
  58048=>"000000000",
  58049=>"111111000",
  58050=>"000100001",
  58051=>"000111111",
  58052=>"000000111",
  58053=>"000000000",
  58054=>"000000000",
  58055=>"110100100",
  58056=>"100101001",
  58057=>"111111001",
  58058=>"100001000",
  58059=>"111101111",
  58060=>"111000000",
  58061=>"000000000",
  58062=>"000000000",
  58063=>"000000000",
  58064=>"000111111",
  58065=>"000100000",
  58066=>"001000000",
  58067=>"000000000",
  58068=>"111001000",
  58069=>"001101111",
  58070=>"000111111",
  58071=>"010010000",
  58072=>"011110010",
  58073=>"000000000",
  58074=>"000001000",
  58075=>"011010000",
  58076=>"111000000",
  58077=>"111000000",
  58078=>"101111111",
  58079=>"000000100",
  58080=>"000000000",
  58081=>"000010010",
  58082=>"000000000",
  58083=>"101000000",
  58084=>"101101101",
  58085=>"111101101",
  58086=>"000000011",
  58087=>"001001000",
  58088=>"000011111",
  58089=>"111110100",
  58090=>"001000000",
  58091=>"111101101",
  58092=>"000000110",
  58093=>"111111111",
  58094=>"010101100",
  58095=>"111111111",
  58096=>"011110101",
  58097=>"111111111",
  58098=>"111111111",
  58099=>"101111111",
  58100=>"000000000",
  58101=>"011001011",
  58102=>"000010000",
  58103=>"010000000",
  58104=>"111111000",
  58105=>"111111111",
  58106=>"001000010",
  58107=>"000111111",
  58108=>"011011011",
  58109=>"101111111",
  58110=>"001001111",
  58111=>"000010111",
  58112=>"010111111",
  58113=>"000001111",
  58114=>"111010110",
  58115=>"000000111",
  58116=>"111111000",
  58117=>"101000000",
  58118=>"011001000",
  58119=>"000111111",
  58120=>"111000000",
  58121=>"111010111",
  58122=>"111111000",
  58123=>"110111111",
  58124=>"111000000",
  58125=>"111111100",
  58126=>"111111000",
  58127=>"000000000",
  58128=>"000001111",
  58129=>"000000000",
  58130=>"111001000",
  58131=>"000001011",
  58132=>"000000000",
  58133=>"100111000",
  58134=>"001001011",
  58135=>"111111111",
  58136=>"111001111",
  58137=>"110110110",
  58138=>"010110110",
  58139=>"111111110",
  58140=>"001011111",
  58141=>"110110010",
  58142=>"000000000",
  58143=>"011001000",
  58144=>"110111000",
  58145=>"111110110",
  58146=>"111000000",
  58147=>"111000000",
  58148=>"111010010",
  58149=>"100000111",
  58150=>"100000000",
  58151=>"111111000",
  58152=>"000000000",
  58153=>"111111011",
  58154=>"000000000",
  58155=>"000000000",
  58156=>"101000000",
  58157=>"011011111",
  58158=>"111111111",
  58159=>"000000000",
  58160=>"000100111",
  58161=>"000000010",
  58162=>"111111000",
  58163=>"111111111",
  58164=>"110000010",
  58165=>"000010100",
  58166=>"000000000",
  58167=>"111111111",
  58168=>"111111111",
  58169=>"111111000",
  58170=>"101000000",
  58171=>"000000000",
  58172=>"010110110",
  58173=>"000000000",
  58174=>"000000000",
  58175=>"111111111",
  58176=>"000000000",
  58177=>"110100110",
  58178=>"001011011",
  58179=>"000000000",
  58180=>"111111111",
  58181=>"111000000",
  58182=>"111000000",
  58183=>"111111011",
  58184=>"000111111",
  58185=>"111000000",
  58186=>"000000000",
  58187=>"000001001",
  58188=>"100100001",
  58189=>"000000000",
  58190=>"111101101",
  58191=>"111100000",
  58192=>"000100100",
  58193=>"000000000",
  58194=>"000000000",
  58195=>"000000000",
  58196=>"000111111",
  58197=>"111111011",
  58198=>"111000000",
  58199=>"000000000",
  58200=>"000000111",
  58201=>"101000100",
  58202=>"111111000",
  58203=>"110110111",
  58204=>"111111111",
  58205=>"111000000",
  58206=>"000101001",
  58207=>"000000000",
  58208=>"100110000",
  58209=>"111111000",
  58210=>"000100100",
  58211=>"000110111",
  58212=>"000001011",
  58213=>"010111111",
  58214=>"111111111",
  58215=>"111110110",
  58216=>"000000100",
  58217=>"111111111",
  58218=>"001000011",
  58219=>"110111111",
  58220=>"110110110",
  58221=>"001111111",
  58222=>"000000000",
  58223=>"111111111",
  58224=>"100110111",
  58225=>"000000000",
  58226=>"001001111",
  58227=>"111011111",
  58228=>"000000000",
  58229=>"110000000",
  58230=>"000010001",
  58231=>"000000011",
  58232=>"011000000",
  58233=>"000100111",
  58234=>"111001000",
  58235=>"101111111",
  58236=>"101000000",
  58237=>"111111001",
  58238=>"000111111",
  58239=>"001000000",
  58240=>"000000000",
  58241=>"000001101",
  58242=>"111111111",
  58243=>"111110110",
  58244=>"011000000",
  58245=>"111111100",
  58246=>"111011111",
  58247=>"000000000",
  58248=>"111111111",
  58249=>"000000001",
  58250=>"000000110",
  58251=>"101101101",
  58252=>"000111111",
  58253=>"010010111",
  58254=>"000111111",
  58255=>"010100100",
  58256=>"000000111",
  58257=>"111111000",
  58258=>"010110100",
  58259=>"000010011",
  58260=>"111111111",
  58261=>"000000000",
  58262=>"000000101",
  58263=>"110111111",
  58264=>"000000000",
  58265=>"001000100",
  58266=>"111111111",
  58267=>"000000000",
  58268=>"111111111",
  58269=>"111011111",
  58270=>"001100000",
  58271=>"000000000",
  58272=>"111101000",
  58273=>"110110111",
  58274=>"000010111",
  58275=>"111111111",
  58276=>"110010111",
  58277=>"111000000",
  58278=>"000111111",
  58279=>"011000000",
  58280=>"010111111",
  58281=>"000000000",
  58282=>"111000000",
  58283=>"000000111",
  58284=>"111001000",
  58285=>"101111111",
  58286=>"000111110",
  58287=>"000000000",
  58288=>"001000000",
  58289=>"000000111",
  58290=>"101001111",
  58291=>"111001000",
  58292=>"000000000",
  58293=>"101001001",
  58294=>"101101101",
  58295=>"001111111",
  58296=>"111111111",
  58297=>"111111111",
  58298=>"000000000",
  58299=>"000000000",
  58300=>"000011001",
  58301=>"110110110",
  58302=>"000000000",
  58303=>"111011000",
  58304=>"001000000",
  58305=>"111111001",
  58306=>"000000000",
  58307=>"111111111",
  58308=>"111111000",
  58309=>"011011111",
  58310=>"000000000",
  58311=>"110010111",
  58312=>"000111111",
  58313=>"111111111",
  58314=>"111111011",
  58315=>"000110000",
  58316=>"000111000",
  58317=>"011011111",
  58318=>"110000000",
  58319=>"111111100",
  58320=>"000001111",
  58321=>"111111110",
  58322=>"111111110",
  58323=>"001101111",
  58324=>"100111111",
  58325=>"101000000",
  58326=>"101101100",
  58327=>"110111111",
  58328=>"001000111",
  58329=>"111001101",
  58330=>"011010000",
  58331=>"101000100",
  58332=>"001111111",
  58333=>"100111111",
  58334=>"110111100",
  58335=>"001110110",
  58336=>"000011111",
  58337=>"111000000",
  58338=>"110000000",
  58339=>"110010011",
  58340=>"111101000",
  58341=>"111000000",
  58342=>"010010000",
  58343=>"111111111",
  58344=>"001000000",
  58345=>"110111111",
  58346=>"000000101",
  58347=>"111110000",
  58348=>"101111111",
  58349=>"111101111",
  58350=>"000000000",
  58351=>"011111111",
  58352=>"000000000",
  58353=>"000000111",
  58354=>"111111111",
  58355=>"011000000",
  58356=>"000000000",
  58357=>"111100100",
  58358=>"001111111",
  58359=>"001001101",
  58360=>"000000000",
  58361=>"111111110",
  58362=>"111111000",
  58363=>"111000000",
  58364=>"011011111",
  58365=>"111100000",
  58366=>"000000100",
  58367=>"111010000",
  58368=>"111111000",
  58369=>"011000000",
  58370=>"000000000",
  58371=>"111111111",
  58372=>"111110110",
  58373=>"001000000",
  58374=>"000111111",
  58375=>"011111111",
  58376=>"001000000",
  58377=>"111110000",
  58378=>"011010000",
  58379=>"100000001",
  58380=>"000100100",
  58381=>"111111111",
  58382=>"100110110",
  58383=>"000000000",
  58384=>"001000111",
  58385=>"000001111",
  58386=>"000000000",
  58387=>"000000000",
  58388=>"000000000",
  58389=>"111101001",
  58390=>"000000111",
  58391=>"000000110",
  58392=>"111111110",
  58393=>"011100101",
  58394=>"000000100",
  58395=>"011111000",
  58396=>"000000000",
  58397=>"111111111",
  58398=>"000000100",
  58399=>"110111111",
  58400=>"111111000",
  58401=>"000000111",
  58402=>"000100101",
  58403=>"011011001",
  58404=>"111000000",
  58405=>"000111111",
  58406=>"111010111",
  58407=>"110111101",
  58408=>"000001111",
  58409=>"000111111",
  58410=>"111100000",
  58411=>"100110111",
  58412=>"000000000",
  58413=>"100111011",
  58414=>"100110000",
  58415=>"001111111",
  58416=>"011110111",
  58417=>"000110111",
  58418=>"001001001",
  58419=>"111001000",
  58420=>"011011000",
  58421=>"111110000",
  58422=>"001001001",
  58423=>"000111111",
  58424=>"100100001",
  58425=>"010100110",
  58426=>"111111111",
  58427=>"111001011",
  58428=>"101000000",
  58429=>"011000000",
  58430=>"111100000",
  58431=>"111001100",
  58432=>"001111111",
  58433=>"110111001",
  58434=>"100110011",
  58435=>"101000100",
  58436=>"000110100",
  58437=>"011111110",
  58438=>"110000000",
  58439=>"000001000",
  58440=>"000011111",
  58441=>"111100110",
  58442=>"000011111",
  58443=>"111000000",
  58444=>"000001111",
  58445=>"000000000",
  58446=>"111001101",
  58447=>"111111111",
  58448=>"011111000",
  58449=>"111001000",
  58450=>"000000100",
  58451=>"111111100",
  58452=>"000000000",
  58453=>"000000001",
  58454=>"011000100",
  58455=>"111111000",
  58456=>"100000001",
  58457=>"111000000",
  58458=>"111011011",
  58459=>"111111110",
  58460=>"000000001",
  58461=>"000000101",
  58462=>"111000000",
  58463=>"000000111",
  58464=>"000000011",
  58465=>"000000000",
  58466=>"000000000",
  58467=>"000000000",
  58468=>"110100111",
  58469=>"111110100",
  58470=>"000000101",
  58471=>"101101111",
  58472=>"111000000",
  58473=>"110000000",
  58474=>"111000000",
  58475=>"111000000",
  58476=>"111100000",
  58477=>"000000111",
  58478=>"111111111",
  58479=>"010110111",
  58480=>"111111111",
  58481=>"111111111",
  58482=>"111000000",
  58483=>"110000000",
  58484=>"011000000",
  58485=>"000000100",
  58486=>"000000101",
  58487=>"010111000",
  58488=>"000000000",
  58489=>"000111111",
  58490=>"111111111",
  58491=>"111000000",
  58492=>"101101001",
  58493=>"111111111",
  58494=>"111111111",
  58495=>"011001000",
  58496=>"010111110",
  58497=>"101111111",
  58498=>"011001011",
  58499=>"011001000",
  58500=>"001011011",
  58501=>"100101111",
  58502=>"111001101",
  58503=>"011000000",
  58504=>"000110110",
  58505=>"000000000",
  58506=>"000000000",
  58507=>"000000000",
  58508=>"111111111",
  58509=>"111110000",
  58510=>"111111000",
  58511=>"000000000",
  58512=>"000000000",
  58513=>"010110000",
  58514=>"000000000",
  58515=>"000000000",
  58516=>"111111001",
  58517=>"101000101",
  58518=>"000111111",
  58519=>"011011001",
  58520=>"001000000",
  58521=>"001000000",
  58522=>"001000000",
  58523=>"011001101",
  58524=>"011011111",
  58525=>"001000000",
  58526=>"000000111",
  58527=>"000000010",
  58528=>"000000000",
  58529=>"000111111",
  58530=>"001001000",
  58531=>"000000111",
  58532=>"001111110",
  58533=>"111111000",
  58534=>"111101101",
  58535=>"000000100",
  58536=>"111111111",
  58537=>"000011011",
  58538=>"000000000",
  58539=>"000000100",
  58540=>"001000111",
  58541=>"100100100",
  58542=>"111101111",
  58543=>"000111111",
  58544=>"000100100",
  58545=>"111010010",
  58546=>"010010000",
  58547=>"000000000",
  58548=>"011111111",
  58549=>"000000000",
  58550=>"000111000",
  58551=>"000100111",
  58552=>"010000000",
  58553=>"100001011",
  58554=>"100000001",
  58555=>"000111111",
  58556=>"101101111",
  58557=>"110111111",
  58558=>"000000000",
  58559=>"000000010",
  58560=>"001111111",
  58561=>"010111111",
  58562=>"000000000",
  58563=>"111111111",
  58564=>"111111111",
  58565=>"111001001",
  58566=>"000000100",
  58567=>"000000000",
  58568=>"000000111",
  58569=>"111100100",
  58570=>"111111110",
  58571=>"000000111",
  58572=>"001100111",
  58573=>"000000101",
  58574=>"111111011",
  58575=>"000000000",
  58576=>"001010110",
  58577=>"011000001",
  58578=>"000000000",
  58579=>"110111111",
  58580=>"000111111",
  58581=>"110111111",
  58582=>"001001000",
  58583=>"000000011",
  58584=>"111110111",
  58585=>"111100000",
  58586=>"000100000",
  58587=>"111011111",
  58588=>"101000100",
  58589=>"001001001",
  58590=>"001000001",
  58591=>"000000000",
  58592=>"000000011",
  58593=>"110101000",
  58594=>"001000101",
  58595=>"000000011",
  58596=>"000000000",
  58597=>"010011011",
  58598=>"111000000",
  58599=>"000101111",
  58600=>"111000000",
  58601=>"011011011",
  58602=>"111110111",
  58603=>"111111111",
  58604=>"111000000",
  58605=>"111111111",
  58606=>"110111000",
  58607=>"000000000",
  58608=>"110100100",
  58609=>"000110010",
  58610=>"001001000",
  58611=>"000000110",
  58612=>"000010111",
  58613=>"100100000",
  58614=>"011011001",
  58615=>"111101000",
  58616=>"000100000",
  58617=>"000000000",
  58618=>"000000000",
  58619=>"011011010",
  58620=>"111111000",
  58621=>"110110111",
  58622=>"000000011",
  58623=>"000000000",
  58624=>"000100111",
  58625=>"111110100",
  58626=>"000000000",
  58627=>"111111110",
  58628=>"000100110",
  58629=>"110000000",
  58630=>"011100100",
  58631=>"110111111",
  58632=>"110111110",
  58633=>"111001111",
  58634=>"111111111",
  58635=>"100000000",
  58636=>"000000000",
  58637=>"011100000",
  58638=>"111111101",
  58639=>"111000000",
  58640=>"100111000",
  58641=>"001000000",
  58642=>"111111111",
  58643=>"000111111",
  58644=>"000000111",
  58645=>"111110000",
  58646=>"000111111",
  58647=>"111110000",
  58648=>"000000111",
  58649=>"111111000",
  58650=>"001101000",
  58651=>"000000000",
  58652=>"000000000",
  58653=>"111111001",
  58654=>"000000000",
  58655=>"000000000",
  58656=>"011000100",
  58657=>"111111111",
  58658=>"111110000",
  58659=>"100111111",
  58660=>"000000010",
  58661=>"000000111",
  58662=>"001111111",
  58663=>"111011011",
  58664=>"000000101",
  58665=>"111111010",
  58666=>"000111111",
  58667=>"111000000",
  58668=>"000000110",
  58669=>"000000001",
  58670=>"111011001",
  58671=>"111000001",
  58672=>"000000100",
  58673=>"011000000",
  58674=>"000000010",
  58675=>"011110110",
  58676=>"111111111",
  58677=>"011000000",
  58678=>"111111111",
  58679=>"001011111",
  58680=>"000111000",
  58681=>"000000000",
  58682=>"100111111",
  58683=>"001000000",
  58684=>"110110010",
  58685=>"111111111",
  58686=>"111111111",
  58687=>"000111000",
  58688=>"000100111",
  58689=>"111111111",
  58690=>"111110111",
  58691=>"111111111",
  58692=>"001000000",
  58693=>"111001001",
  58694=>"000000110",
  58695=>"110000000",
  58696=>"000000000",
  58697=>"000011000",
  58698=>"111000000",
  58699=>"100111111",
  58700=>"111111111",
  58701=>"000100111",
  58702=>"111111011",
  58703=>"111011000",
  58704=>"000001001",
  58705=>"000000001",
  58706=>"111000100",
  58707=>"000000001",
  58708=>"001111011",
  58709=>"000000001",
  58710=>"000000111",
  58711=>"111111100",
  58712=>"000000000",
  58713=>"111011000",
  58714=>"111100000",
  58715=>"011010000",
  58716=>"000000011",
  58717=>"000110111",
  58718=>"011000000",
  58719=>"011001111",
  58720=>"111111011",
  58721=>"000000101",
  58722=>"000000010",
  58723=>"111111111",
  58724=>"100110100",
  58725=>"000000001",
  58726=>"001000001",
  58727=>"111110000",
  58728=>"000111111",
  58729=>"111111111",
  58730=>"100111000",
  58731=>"000001111",
  58732=>"111101100",
  58733=>"000000110",
  58734=>"000001111",
  58735=>"011111011",
  58736=>"000000000",
  58737=>"000111111",
  58738=>"111100000",
  58739=>"001011111",
  58740=>"010000000",
  58741=>"000000000",
  58742=>"110110110",
  58743=>"111110100",
  58744=>"000100010",
  58745=>"010000000",
  58746=>"001111111",
  58747=>"100110110",
  58748=>"111100000",
  58749=>"001000001",
  58750=>"111111111",
  58751=>"101001000",
  58752=>"000100111",
  58753=>"101100111",
  58754=>"111111100",
  58755=>"000000000",
  58756=>"010000000",
  58757=>"000011010",
  58758=>"000000100",
  58759=>"000100101",
  58760=>"111111111",
  58761=>"000000111",
  58762=>"000000000",
  58763=>"111001000",
  58764=>"111001111",
  58765=>"100110110",
  58766=>"000000100",
  58767=>"000000100",
  58768=>"000000000",
  58769=>"111000000",
  58770=>"111111000",
  58771=>"001000100",
  58772=>"011000011",
  58773=>"001001101",
  58774=>"111111111",
  58775=>"000010100",
  58776=>"100100101",
  58777=>"000101010",
  58778=>"000000000",
  58779=>"110100101",
  58780=>"111110111",
  58781=>"000111011",
  58782=>"000000000",
  58783=>"111111000",
  58784=>"011000111",
  58785=>"111111100",
  58786=>"111111000",
  58787=>"000000111",
  58788=>"000000100",
  58789=>"111111111",
  58790=>"000000001",
  58791=>"111111000",
  58792=>"000000000",
  58793=>"000000000",
  58794=>"000000111",
  58795=>"000000110",
  58796=>"001000000",
  58797=>"000000111",
  58798=>"000000111",
  58799=>"000000000",
  58800=>"111110000",
  58801=>"111111111",
  58802=>"000000000",
  58803=>"011111111",
  58804=>"000000000",
  58805=>"111111011",
  58806=>"000011111",
  58807=>"111111101",
  58808=>"000001111",
  58809=>"101111011",
  58810=>"111111101",
  58811=>"111111111",
  58812=>"110111111",
  58813=>"000000001",
  58814=>"111111011",
  58815=>"000000000",
  58816=>"110110110",
  58817=>"000000100",
  58818=>"010111111",
  58819=>"110111111",
  58820=>"111111111",
  58821=>"001011110",
  58822=>"000111111",
  58823=>"000000110",
  58824=>"001000000",
  58825=>"000000000",
  58826=>"000001001",
  58827=>"100000111",
  58828=>"111111111",
  58829=>"111101000",
  58830=>"101101000",
  58831=>"100000100",
  58832=>"010000111",
  58833=>"111111111",
  58834=>"101101111",
  58835=>"110110111",
  58836=>"100000000",
  58837=>"000111100",
  58838=>"010111110",
  58839=>"000011011",
  58840=>"000000100",
  58841=>"000000000",
  58842=>"111100101",
  58843=>"000000000",
  58844=>"110111111",
  58845=>"111111000",
  58846=>"111001110",
  58847=>"110000000",
  58848=>"000100110",
  58849=>"100111111",
  58850=>"000000000",
  58851=>"000000111",
  58852=>"111111111",
  58853=>"111111101",
  58854=>"111111100",
  58855=>"111000000",
  58856=>"100111111",
  58857=>"111111111",
  58858=>"111111111",
  58859=>"111111000",
  58860=>"100000000",
  58861=>"000000000",
  58862=>"110000000",
  58863=>"000000000",
  58864=>"000000000",
  58865=>"111111100",
  58866=>"100111111",
  58867=>"011010000",
  58868=>"111101101",
  58869=>"000000000",
  58870=>"101101111",
  58871=>"001000100",
  58872=>"001000000",
  58873=>"001001011",
  58874=>"010000000",
  58875=>"000101111",
  58876=>"111110000",
  58877=>"110110110",
  58878=>"111111111",
  58879=>"101000000",
  58880=>"101111111",
  58881=>"011010110",
  58882=>"000111111",
  58883=>"000010011",
  58884=>"011111110",
  58885=>"111111111",
  58886=>"100000100",
  58887=>"111111000",
  58888=>"100000000",
  58889=>"111001000",
  58890=>"000000000",
  58891=>"001011111",
  58892=>"010111111",
  58893=>"000000000",
  58894=>"110110111",
  58895=>"111111111",
  58896=>"000000000",
  58897=>"101100101",
  58898=>"001000100",
  58899=>"100100000",
  58900=>"111111111",
  58901=>"000110000",
  58902=>"000100011",
  58903=>"111111001",
  58904=>"000000000",
  58905=>"011011110",
  58906=>"000000000",
  58907=>"000100110",
  58908=>"111111111",
  58909=>"101111111",
  58910=>"000000000",
  58911=>"000000000",
  58912=>"111110111",
  58913=>"100100111",
  58914=>"100100111",
  58915=>"101100110",
  58916=>"000000000",
  58917=>"110100111",
  58918=>"101100100",
  58919=>"111111000",
  58920=>"000000111",
  58921=>"000000000",
  58922=>"000000001",
  58923=>"111111111",
  58924=>"000001001",
  58925=>"111111111",
  58926=>"011111111",
  58927=>"110111111",
  58928=>"111111111",
  58929=>"011011111",
  58930=>"111111111",
  58931=>"111111000",
  58932=>"100000110",
  58933=>"000001100",
  58934=>"000011111",
  58935=>"011001000",
  58936=>"000000000",
  58937=>"001001011",
  58938=>"000000000",
  58939=>"011111000",
  58940=>"111111110",
  58941=>"111111111",
  58942=>"111111110",
  58943=>"111111111",
  58944=>"001001000",
  58945=>"000010011",
  58946=>"011111001",
  58947=>"000000000",
  58948=>"000000000",
  58949=>"111111111",
  58950=>"000110011",
  58951=>"111111111",
  58952=>"000100000",
  58953=>"011000100",
  58954=>"000010010",
  58955=>"101101111",
  58956=>"000000100",
  58957=>"000000001",
  58958=>"111111011",
  58959=>"000000000",
  58960=>"011001111",
  58961=>"110111111",
  58962=>"010011000",
  58963=>"000011111",
  58964=>"100000110",
  58965=>"111111011",
  58966=>"000100000",
  58967=>"000111111",
  58968=>"111110110",
  58969=>"000000000",
  58970=>"111111111",
  58971=>"111100000",
  58972=>"111111111",
  58973=>"000000000",
  58974=>"111111100",
  58975=>"011000110",
  58976=>"000000000",
  58977=>"111111000",
  58978=>"111111111",
  58979=>"011111111",
  58980=>"000000000",
  58981=>"111101001",
  58982=>"111111100",
  58983=>"111001001",
  58984=>"000000111",
  58985=>"110111110",
  58986=>"111100000",
  58987=>"000011111",
  58988=>"110110111",
  58989=>"101100000",
  58990=>"111001000",
  58991=>"111101001",
  58992=>"000001000",
  58993=>"000000011",
  58994=>"000000000",
  58995=>"110100000",
  58996=>"111111111",
  58997=>"001101000",
  58998=>"111111000",
  58999=>"111111111",
  59000=>"111111111",
  59001=>"000000000",
  59002=>"111111000",
  59003=>"000000100",
  59004=>"111000000",
  59005=>"100010010",
  59006=>"111111110",
  59007=>"111111110",
  59008=>"111000111",
  59009=>"000000000",
  59010=>"111011010",
  59011=>"111111110",
  59012=>"110110110",
  59013=>"011111111",
  59014=>"111111111",
  59015=>"000000100",
  59016=>"111111111",
  59017=>"000000000",
  59018=>"110111111",
  59019=>"100111001",
  59020=>"011000000",
  59021=>"111111111",
  59022=>"111011000",
  59023=>"000000000",
  59024=>"000000000",
  59025=>"100111111",
  59026=>"000000000",
  59027=>"111111111",
  59028=>"011011001",
  59029=>"111111111",
  59030=>"111111111",
  59031=>"111001111",
  59032=>"101111011",
  59033=>"011001001",
  59034=>"011111111",
  59035=>"111000000",
  59036=>"000110111",
  59037=>"101000000",
  59038=>"000000110",
  59039=>"111111000",
  59040=>"111111111",
  59041=>"000000000",
  59042=>"001001011",
  59043=>"000000000",
  59044=>"001000000",
  59045=>"000100100",
  59046=>"111111111",
  59047=>"111111001",
  59048=>"111111111",
  59049=>"111011011",
  59050=>"000000000",
  59051=>"000000000",
  59052=>"111101001",
  59053=>"111111111",
  59054=>"001111110",
  59055=>"000000111",
  59056=>"111111111",
  59057=>"000010001",
  59058=>"111111001",
  59059=>"000000000",
  59060=>"000000000",
  59061=>"001001111",
  59062=>"001001111",
  59063=>"011000000",
  59064=>"111111111",
  59065=>"000000011",
  59066=>"000000000",
  59067=>"000000000",
  59068=>"000000000",
  59069=>"001001000",
  59070=>"111001000",
  59071=>"111111111",
  59072=>"111111111",
  59073=>"000000000",
  59074=>"000111111",
  59075=>"000111111",
  59076=>"000000000",
  59077=>"111111111",
  59078=>"000000000",
  59079=>"111111110",
  59080=>"010000000",
  59081=>"000000000",
  59082=>"100100100",
  59083=>"010000001",
  59084=>"000000000",
  59085=>"001001111",
  59086=>"000000000",
  59087=>"111111001",
  59088=>"111111111",
  59089=>"101101111",
  59090=>"111111111",
  59091=>"100000000",
  59092=>"111011111",
  59093=>"111111000",
  59094=>"111001111",
  59095=>"111101110",
  59096=>"111111111",
  59097=>"001000111",
  59098=>"111111111",
  59099=>"011111111",
  59100=>"111111111",
  59101=>"000000100",
  59102=>"000001000",
  59103=>"000000000",
  59104=>"010011000",
  59105=>"011011111",
  59106=>"001010000",
  59107=>"000000011",
  59108=>"111000100",
  59109=>"101000001",
  59110=>"111111111",
  59111=>"011111111",
  59112=>"011011010",
  59113=>"111111111",
  59114=>"001000111",
  59115=>"000000000",
  59116=>"000111010",
  59117=>"101101111",
  59118=>"111110101",
  59119=>"010010111",
  59120=>"110001000",
  59121=>"000000111",
  59122=>"110000000",
  59123=>"000000000",
  59124=>"000001001",
  59125=>"100001111",
  59126=>"111110111",
  59127=>"000000001",
  59128=>"000000000",
  59129=>"000000000",
  59130=>"010111111",
  59131=>"000001001",
  59132=>"000000100",
  59133=>"000110110",
  59134=>"100100001",
  59135=>"000100111",
  59136=>"000000001",
  59137=>"110111110",
  59138=>"000000111",
  59139=>"000010111",
  59140=>"111110000",
  59141=>"111110110",
  59142=>"000000000",
  59143=>"000000000",
  59144=>"111101100",
  59145=>"000000111",
  59146=>"011101001",
  59147=>"000100100",
  59148=>"011011001",
  59149=>"011011011",
  59150=>"000000110",
  59151=>"000000000",
  59152=>"011110111",
  59153=>"000001000",
  59154=>"010000000",
  59155=>"111101101",
  59156=>"000000000",
  59157=>"111111111",
  59158=>"011110111",
  59159=>"000000000",
  59160=>"111111111",
  59161=>"111111111",
  59162=>"111111011",
  59163=>"110010001",
  59164=>"100000000",
  59165=>"000000000",
  59166=>"111111111",
  59167=>"111001000",
  59168=>"000000111",
  59169=>"001001111",
  59170=>"000100111",
  59171=>"010110111",
  59172=>"000000010",
  59173=>"111111000",
  59174=>"011111111",
  59175=>"000000001",
  59176=>"000000000",
  59177=>"000000000",
  59178=>"000000111",
  59179=>"110110000",
  59180=>"111111110",
  59181=>"101000000",
  59182=>"111111111",
  59183=>"101001000",
  59184=>"000000000",
  59185=>"000001011",
  59186=>"111111111",
  59187=>"111110000",
  59188=>"111111111",
  59189=>"111000000",
  59190=>"111111111",
  59191=>"111111111",
  59192=>"111111111",
  59193=>"111000000",
  59194=>"111100000",
  59195=>"000111011",
  59196=>"011011001",
  59197=>"000001000",
  59198=>"000001111",
  59199=>"111111111",
  59200=>"000000000",
  59201=>"000000000",
  59202=>"100111111",
  59203=>"111111111",
  59204=>"111111111",
  59205=>"000000000",
  59206=>"011000000",
  59207=>"000010010",
  59208=>"111111101",
  59209=>"111000000",
  59210=>"111000110",
  59211=>"110010000",
  59212=>"001000000",
  59213=>"101111000",
  59214=>"001000000",
  59215=>"101001001",
  59216=>"000000000",
  59217=>"000000000",
  59218=>"111000000",
  59219=>"111111100",
  59220=>"111000000",
  59221=>"001010001",
  59222=>"000011011",
  59223=>"000000000",
  59224=>"001000111",
  59225=>"111111111",
  59226=>"001011010",
  59227=>"000101111",
  59228=>"010110111",
  59229=>"111111000",
  59230=>"100000001",
  59231=>"000000000",
  59232=>"111111111",
  59233=>"000000000",
  59234=>"110011111",
  59235=>"000000000",
  59236=>"011011000",
  59237=>"001101111",
  59238=>"000000000",
  59239=>"001110111",
  59240=>"111001000",
  59241=>"000000000",
  59242=>"111111010",
  59243=>"000111111",
  59244=>"000000000",
  59245=>"000000001",
  59246=>"000001001",
  59247=>"000011000",
  59248=>"000000000",
  59249=>"111111011",
  59250=>"000111000",
  59251=>"111110111",
  59252=>"011000000",
  59253=>"100100110",
  59254=>"000000000",
  59255=>"100110000",
  59256=>"001000000",
  59257=>"000001000",
  59258=>"000000000",
  59259=>"011111110",
  59260=>"000000111",
  59261=>"010000000",
  59262=>"111000000",
  59263=>"001001001",
  59264=>"001001000",
  59265=>"000111111",
  59266=>"111111111",
  59267=>"111111111",
  59268=>"000000001",
  59269=>"000001111",
  59270=>"111110000",
  59271=>"000000000",
  59272=>"000000000",
  59273=>"000011111",
  59274=>"111101111",
  59275=>"001000111",
  59276=>"111111111",
  59277=>"101111111",
  59278=>"000001111",
  59279=>"111111111",
  59280=>"111111111",
  59281=>"000000000",
  59282=>"001000000",
  59283=>"110110110",
  59284=>"111111111",
  59285=>"000000000",
  59286=>"111101111",
  59287=>"011011111",
  59288=>"000100100",
  59289=>"000001000",
  59290=>"111111111",
  59291=>"001101111",
  59292=>"011000000",
  59293=>"111111110",
  59294=>"000000001",
  59295=>"111111100",
  59296=>"111111111",
  59297=>"100100111",
  59298=>"111110111",
  59299=>"000001111",
  59300=>"110111111",
  59301=>"010000000",
  59302=>"110011011",
  59303=>"000001000",
  59304=>"000000000",
  59305=>"110100010",
  59306=>"001001011",
  59307=>"000000000",
  59308=>"111111010",
  59309=>"000000000",
  59310=>"000000001",
  59311=>"111111110",
  59312=>"000111111",
  59313=>"111100000",
  59314=>"000000000",
  59315=>"111111111",
  59316=>"001001001",
  59317=>"110000000",
  59318=>"000000010",
  59319=>"001101000",
  59320=>"011000100",
  59321=>"001001111",
  59322=>"000000000",
  59323=>"000111101",
  59324=>"000000000",
  59325=>"111011000",
  59326=>"001000000",
  59327=>"011011011",
  59328=>"000011000",
  59329=>"111000000",
  59330=>"111111111",
  59331=>"000010010",
  59332=>"111111000",
  59333=>"111111100",
  59334=>"000000000",
  59335=>"001001001",
  59336=>"000111111",
  59337=>"100000000",
  59338=>"001111111",
  59339=>"101111111",
  59340=>"111011000",
  59341=>"111111111",
  59342=>"111111111",
  59343=>"110111111",
  59344=>"000000000",
  59345=>"000011001",
  59346=>"000111111",
  59347=>"000000001",
  59348=>"000000000",
  59349=>"001010000",
  59350=>"100100000",
  59351=>"000000000",
  59352=>"000111110",
  59353=>"000000100",
  59354=>"000000000",
  59355=>"100100101",
  59356=>"000001111",
  59357=>"001001001",
  59358=>"000000111",
  59359=>"000100000",
  59360=>"000111111",
  59361=>"001000000",
  59362=>"100100000",
  59363=>"000000111",
  59364=>"111111111",
  59365=>"111111111",
  59366=>"111010000",
  59367=>"111111101",
  59368=>"001011111",
  59369=>"000000101",
  59370=>"000000000",
  59371=>"000111111",
  59372=>"000000111",
  59373=>"110110111",
  59374=>"010111110",
  59375=>"111111111",
  59376=>"000001101",
  59377=>"111111011",
  59378=>"000000000",
  59379=>"001001000",
  59380=>"000000000",
  59381=>"000000101",
  59382=>"110111100",
  59383=>"001001000",
  59384=>"111111001",
  59385=>"111101101",
  59386=>"010000000",
  59387=>"000000000",
  59388=>"111111110",
  59389=>"000000000",
  59390=>"010111111",
  59391=>"111111111",
  59392=>"111000011",
  59393=>"111011111",
  59394=>"000000000",
  59395=>"000000000",
  59396=>"011001100",
  59397=>"011000001",
  59398=>"000001001",
  59399=>"111111111",
  59400=>"000000011",
  59401=>"000010000",
  59402=>"111111111",
  59403=>"111100101",
  59404=>"110110111",
  59405=>"111111101",
  59406=>"100111011",
  59407=>"111111000",
  59408=>"001001000",
  59409=>"000000000",
  59410=>"111101100",
  59411=>"000000000",
  59412=>"100100110",
  59413=>"111111111",
  59414=>"000100111",
  59415=>"011110111",
  59416=>"001000001",
  59417=>"000000000",
  59418=>"100000000",
  59419=>"111100101",
  59420=>"000000001",
  59421=>"100100110",
  59422=>"110110110",
  59423=>"000000000",
  59424=>"111000000",
  59425=>"100101110",
  59426=>"001101100",
  59427=>"111111111",
  59428=>"111111111",
  59429=>"011000001",
  59430=>"111111111",
  59431=>"100100100",
  59432=>"000000000",
  59433=>"000000011",
  59434=>"101001001",
  59435=>"000000000",
  59436=>"000000000",
  59437=>"111111111",
  59438=>"111111111",
  59439=>"111000000",
  59440=>"111111000",
  59441=>"000000000",
  59442=>"111111101",
  59443=>"111111111",
  59444=>"000110000",
  59445=>"010010000",
  59446=>"011001000",
  59447=>"000000000",
  59448=>"000000000",
  59449=>"000101111",
  59450=>"111111111",
  59451=>"000010000",
  59452=>"100111111",
  59453=>"101101100",
  59454=>"001100000",
  59455=>"101001000",
  59456=>"000000000",
  59457=>"000010111",
  59458=>"000101111",
  59459=>"111111111",
  59460=>"011011011",
  59461=>"010000000",
  59462=>"011011011",
  59463=>"111111111",
  59464=>"011001000",
  59465=>"000110111",
  59466=>"000000111",
  59467=>"011111110",
  59468=>"111111111",
  59469=>"000100000",
  59470=>"011000111",
  59471=>"000000000",
  59472=>"000000000",
  59473=>"111111111",
  59474=>"001001000",
  59475=>"011011110",
  59476=>"111101101",
  59477=>"000010000",
  59478=>"111110110",
  59479=>"000000000",
  59480=>"111111111",
  59481=>"001001111",
  59482=>"100100100",
  59483=>"100100000",
  59484=>"000111111",
  59485=>"111110100",
  59486=>"100000000",
  59487=>"000011111",
  59488=>"000001111",
  59489=>"101111111",
  59490=>"000001101",
  59491=>"000000000",
  59492=>"000000100",
  59493=>"000100000",
  59494=>"000000011",
  59495=>"000000000",
  59496=>"000110111",
  59497=>"000000000",
  59498=>"111111010",
  59499=>"111111111",
  59500=>"100110110",
  59501=>"000000011",
  59502=>"111001111",
  59503=>"110111000",
  59504=>"111111111",
  59505=>"000000010",
  59506=>"100101000",
  59507=>"000000000",
  59508=>"000110000",
  59509=>"011110000",
  59510=>"110110111",
  59511=>"000000111",
  59512=>"000111000",
  59513=>"111111100",
  59514=>"000000000",
  59515=>"000000000",
  59516=>"111111111",
  59517=>"111101111",
  59518=>"000010000",
  59519=>"001101101",
  59520=>"000000000",
  59521=>"111111111",
  59522=>"111111111",
  59523=>"101111000",
  59524=>"001010111",
  59525=>"000000010",
  59526=>"111111110",
  59527=>"000000000",
  59528=>"111000000",
  59529=>"001001001",
  59530=>"110100000",
  59531=>"100000000",
  59532=>"000001011",
  59533=>"111111001",
  59534=>"000100100",
  59535=>"000000000",
  59536=>"000011111",
  59537=>"000001000",
  59538=>"000000001",
  59539=>"111001001",
  59540=>"010111100",
  59541=>"000001001",
  59542=>"000000100",
  59543=>"111111111",
  59544=>"011011111",
  59545=>"000000000",
  59546=>"000000000",
  59547=>"011000000",
  59548=>"000000000",
  59549=>"000000011",
  59550=>"000001111",
  59551=>"000111111",
  59552=>"000001111",
  59553=>"011000111",
  59554=>"000000110",
  59555=>"000000000",
  59556=>"010011000",
  59557=>"000000001",
  59558=>"000000000",
  59559=>"110110000",
  59560=>"101101111",
  59561=>"011111111",
  59562=>"000000000",
  59563=>"111111111",
  59564=>"000111111",
  59565=>"111111011",
  59566=>"111111111",
  59567=>"000000000",
  59568=>"110110000",
  59569=>"001011011",
  59570=>"111110000",
  59571=>"000000000",
  59572=>"000000000",
  59573=>"110100111",
  59574=>"000101111",
  59575=>"111001001",
  59576=>"111111111",
  59577=>"111000000",
  59578=>"000000000",
  59579=>"011000100",
  59580=>"111111111",
  59581=>"110100110",
  59582=>"111111110",
  59583=>"111111111",
  59584=>"000000000",
  59585=>"011101101",
  59586=>"111000111",
  59587=>"000000000",
  59588=>"100100100",
  59589=>"000000000",
  59590=>"111111111",
  59591=>"011001111",
  59592=>"000000000",
  59593=>"101111111",
  59594=>"001001111",
  59595=>"110000100",
  59596=>"000000000",
  59597=>"010110111",
  59598=>"100000000",
  59599=>"111111111",
  59600=>"100100111",
  59601=>"111111111",
  59602=>"111111111",
  59603=>"001111111",
  59604=>"000000100",
  59605=>"111111111",
  59606=>"110010000",
  59607=>"100010111",
  59608=>"000000000",
  59609=>"111111111",
  59610=>"000000000",
  59611=>"000010111",
  59612=>"100111111",
  59613=>"100111111",
  59614=>"000000000",
  59615=>"000000100",
  59616=>"000000000",
  59617=>"000000000",
  59618=>"000000011",
  59619=>"000000100",
  59620=>"111111111",
  59621=>"001000000",
  59622=>"111111111",
  59623=>"111000100",
  59624=>"111111001",
  59625=>"010110111",
  59626=>"111111111",
  59627=>"100101111",
  59628=>"111111111",
  59629=>"000000111",
  59630=>"000000111",
  59631=>"000001011",
  59632=>"000111111",
  59633=>"000110100",
  59634=>"111100110",
  59635=>"111111111",
  59636=>"111111110",
  59637=>"000000100",
  59638=>"001011011",
  59639=>"111111111",
  59640=>"111000000",
  59641=>"000000000",
  59642=>"110110111",
  59643=>"000000111",
  59644=>"000000000",
  59645=>"000000000",
  59646=>"000111011",
  59647=>"110110110",
  59648=>"011000110",
  59649=>"001001101",
  59650=>"000000000",
  59651=>"101111111",
  59652=>"111110110",
  59653=>"110111111",
  59654=>"111100000",
  59655=>"101101111",
  59656=>"110111111",
  59657=>"111100100",
  59658=>"111111111",
  59659=>"000000111",
  59660=>"111111111",
  59661=>"111111111",
  59662=>"010000000",
  59663=>"111111111",
  59664=>"010110111",
  59665=>"011111111",
  59666=>"000000000",
  59667=>"011001111",
  59668=>"001111000",
  59669=>"000111111",
  59670=>"111011001",
  59671=>"111111111",
  59672=>"001011001",
  59673=>"000000100",
  59674=>"000000000",
  59675=>"000000100",
  59676=>"111011000",
  59677=>"000000000",
  59678=>"000000000",
  59679=>"001101111",
  59680=>"000100111",
  59681=>"111101100",
  59682=>"111111111",
  59683=>"111111111",
  59684=>"111011011",
  59685=>"111111111",
  59686=>"111111111",
  59687=>"111111000",
  59688=>"000011101",
  59689=>"101000000",
  59690=>"111000000",
  59691=>"000000000",
  59692=>"000000000",
  59693=>"011011011",
  59694=>"110000000",
  59695=>"000000000",
  59696=>"110111111",
  59697=>"000000000",
  59698=>"111101000",
  59699=>"000000001",
  59700=>"111111111",
  59701=>"000000101",
  59702=>"010010000",
  59703=>"111111111",
  59704=>"111111000",
  59705=>"110111111",
  59706=>"010000111",
  59707=>"110111111",
  59708=>"111101101",
  59709=>"000000000",
  59710=>"000000000",
  59711=>"000000000",
  59712=>"000000000",
  59713=>"000100000",
  59714=>"001100110",
  59715=>"111111111",
  59716=>"000100000",
  59717=>"110111111",
  59718=>"000000000",
  59719=>"000000001",
  59720=>"000000000",
  59721=>"000000110",
  59722=>"001000011",
  59723=>"101101111",
  59724=>"011001101",
  59725=>"111111011",
  59726=>"001100000",
  59727=>"001001001",
  59728=>"011011011",
  59729=>"000000010",
  59730=>"111111111",
  59731=>"000000000",
  59732=>"000000000",
  59733=>"011011011",
  59734=>"000000000",
  59735=>"000000000",
  59736=>"111000001",
  59737=>"011111111",
  59738=>"101101001",
  59739=>"000000000",
  59740=>"000011111",
  59741=>"000000000",
  59742=>"011111111",
  59743=>"110000000",
  59744=>"011011111",
  59745=>"111000000",
  59746=>"001001000",
  59747=>"111111111",
  59748=>"000010000",
  59749=>"011001111",
  59750=>"001000111",
  59751=>"001101110",
  59752=>"110110111",
  59753=>"111010000",
  59754=>"111000000",
  59755=>"010111000",
  59756=>"110110110",
  59757=>"011111111",
  59758=>"000000000",
  59759=>"011011111",
  59760=>"011000000",
  59761=>"110011111",
  59762=>"111111000",
  59763=>"111111011",
  59764=>"111000000",
  59765=>"011111110",
  59766=>"000110111",
  59767=>"000000000",
  59768=>"000000000",
  59769=>"110011111",
  59770=>"000000000",
  59771=>"011111111",
  59772=>"000000011",
  59773=>"000000000",
  59774=>"011001000",
  59775=>"111111011",
  59776=>"011111111",
  59777=>"000000000",
  59778=>"000000000",
  59779=>"000000000",
  59780=>"000011000",
  59781=>"000110111",
  59782=>"000000000",
  59783=>"000000000",
  59784=>"111111000",
  59785=>"111111110",
  59786=>"000000001",
  59787=>"000000010",
  59788=>"111101111",
  59789=>"100111111",
  59790=>"101111111",
  59791=>"000000000",
  59792=>"011001001",
  59793=>"111111111",
  59794=>"110000001",
  59795=>"100100100",
  59796=>"000000000",
  59797=>"000010000",
  59798=>"001000000",
  59799=>"011001011",
  59800=>"111111111",
  59801=>"010011001",
  59802=>"000000000",
  59803=>"001111110",
  59804=>"011000001",
  59805=>"000000000",
  59806=>"000000000",
  59807=>"000000000",
  59808=>"000110110",
  59809=>"000000001",
  59810=>"001000000",
  59811=>"000000000",
  59812=>"001000000",
  59813=>"000111110",
  59814=>"111100000",
  59815=>"000111111",
  59816=>"010010000",
  59817=>"110110111",
  59818=>"111111111",
  59819=>"111111001",
  59820=>"000111111",
  59821=>"100011001",
  59822=>"000000000",
  59823=>"000100101",
  59824=>"111000000",
  59825=>"100001111",
  59826=>"010011101",
  59827=>"000000000",
  59828=>"111111111",
  59829=>"000000000",
  59830=>"011010110",
  59831=>"011011000",
  59832=>"000000000",
  59833=>"000001001",
  59834=>"011000011",
  59835=>"001100100",
  59836=>"111111000",
  59837=>"000000000",
  59838=>"001000000",
  59839=>"100100101",
  59840=>"111111111",
  59841=>"000000000",
  59842=>"111111111",
  59843=>"000000000",
  59844=>"111111111",
  59845=>"000000001",
  59846=>"000000000",
  59847=>"100000000",
  59848=>"011111111",
  59849=>"111111000",
  59850=>"000000000",
  59851=>"111111011",
  59852=>"000000000",
  59853=>"110100100",
  59854=>"111101000",
  59855=>"100110001",
  59856=>"000000001",
  59857=>"001111111",
  59858=>"000100100",
  59859=>"001001011",
  59860=>"100000000",
  59861=>"100100100",
  59862=>"000000000",
  59863=>"111111111",
  59864=>"111111000",
  59865=>"000000000",
  59866=>"111101111",
  59867=>"111011001",
  59868=>"000000000",
  59869=>"111010000",
  59870=>"000000000",
  59871=>"000000000",
  59872=>"000000000",
  59873=>"111111111",
  59874=>"000000000",
  59875=>"111111010",
  59876=>"111111111",
  59877=>"000001000",
  59878=>"000000000",
  59879=>"000000100",
  59880=>"111011101",
  59881=>"011011011",
  59882=>"001101101",
  59883=>"000100101",
  59884=>"100000001",
  59885=>"101101110",
  59886=>"100100000",
  59887=>"000000000",
  59888=>"011001111",
  59889=>"111001000",
  59890=>"000101101",
  59891=>"111111001",
  59892=>"111110111",
  59893=>"110000000",
  59894=>"111111111",
  59895=>"101100000",
  59896=>"000011011",
  59897=>"011001110",
  59898=>"000001001",
  59899=>"111000000",
  59900=>"111111111",
  59901=>"010111111",
  59902=>"111111011",
  59903=>"000000000",
  59904=>"101110111",
  59905=>"110110110",
  59906=>"111111000",
  59907=>"000111111",
  59908=>"101100000",
  59909=>"000000000",
  59910=>"111001001",
  59911=>"000100111",
  59912=>"111111111",
  59913=>"000000000",
  59914=>"111000000",
  59915=>"000000000",
  59916=>"110010011",
  59917=>"010000000",
  59918=>"111111111",
  59919=>"000010010",
  59920=>"000000011",
  59921=>"111110000",
  59922=>"111000000",
  59923=>"111110000",
  59924=>"000000011",
  59925=>"000000000",
  59926=>"000100111",
  59927=>"111111111",
  59928=>"111111111",
  59929=>"000011111",
  59930=>"000000000",
  59931=>"100111111",
  59932=>"000111111",
  59933=>"001000000",
  59934=>"110000000",
  59935=>"000000001",
  59936=>"001111111",
  59937=>"000000111",
  59938=>"001101111",
  59939=>"110000000",
  59940=>"111111111",
  59941=>"000111001",
  59942=>"110000110",
  59943=>"111111000",
  59944=>"000000001",
  59945=>"000000001",
  59946=>"000000111",
  59947=>"111110111",
  59948=>"111110111",
  59949=>"000010111",
  59950=>"000000100",
  59951=>"001000000",
  59952=>"111101000",
  59953=>"000001111",
  59954=>"000110100",
  59955=>"110010111",
  59956=>"010110100",
  59957=>"110110001",
  59958=>"111011010",
  59959=>"000000111",
  59960=>"000001001",
  59961=>"011010111",
  59962=>"110111111",
  59963=>"010100111",
  59964=>"000000000",
  59965=>"111000000",
  59966=>"000111111",
  59967=>"000000110",
  59968=>"011111001",
  59969=>"000111111",
  59970=>"111110101",
  59971=>"000000111",
  59972=>"111111110",
  59973=>"111111111",
  59974=>"111100000",
  59975=>"000000111",
  59976=>"001011000",
  59977=>"111000111",
  59978=>"000101111",
  59979=>"001011001",
  59980=>"011111111",
  59981=>"111111000",
  59982=>"101000000",
  59983=>"001000000",
  59984=>"110101111",
  59985=>"000000010",
  59986=>"000000000",
  59987=>"000000110",
  59988=>"000000000",
  59989=>"110111111",
  59990=>"000010010",
  59991=>"111111000",
  59992=>"001000000",
  59993=>"111111111",
  59994=>"000000000",
  59995=>"000000110",
  59996=>"110110111",
  59997=>"111111110",
  59998=>"101100111",
  59999=>"101111110",
  60000=>"010111111",
  60001=>"011010000",
  60002=>"000001111",
  60003=>"111111111",
  60004=>"100111001",
  60005=>"000001111",
  60006=>"000110110",
  60007=>"000000000",
  60008=>"111111111",
  60009=>"000001001",
  60010=>"000110111",
  60011=>"010010000",
  60012=>"000111111",
  60013=>"111111011",
  60014=>"001000000",
  60015=>"111111111",
  60016=>"000010000",
  60017=>"000000110",
  60018=>"001001001",
  60019=>"001111111",
  60020=>"101000111",
  60021=>"111111000",
  60022=>"111000000",
  60023=>"110111101",
  60024=>"001000001",
  60025=>"001111111",
  60026=>"000000000",
  60027=>"111000000",
  60028=>"011111001",
  60029=>"110110100",
  60030=>"000000001",
  60031=>"000000000",
  60032=>"101111000",
  60033=>"000000000",
  60034=>"000000000",
  60035=>"000011111",
  60036=>"000101111",
  60037=>"111000000",
  60038=>"111100111",
  60039=>"110000000",
  60040=>"000111111",
  60041=>"000011111",
  60042=>"111101111",
  60043=>"111000000",
  60044=>"000001001",
  60045=>"000000111",
  60046=>"111111111",
  60047=>"111111000",
  60048=>"111100000",
  60049=>"100000000",
  60050=>"111111111",
  60051=>"011011011",
  60052=>"001000100",
  60053=>"000010000",
  60054=>"000000000",
  60055=>"111111111",
  60056=>"111001111",
  60057=>"000000001",
  60058=>"111000000",
  60059=>"000000000",
  60060=>"000010111",
  60061=>"000000001",
  60062=>"110111000",
  60063=>"100100010",
  60064=>"000000000",
  60065=>"100100000",
  60066=>"111111010",
  60067=>"000000111",
  60068=>"111100000",
  60069=>"000111111",
  60070=>"001001001",
  60071=>"000000000",
  60072=>"111100000",
  60073=>"101000000",
  60074=>"000000001",
  60075=>"000000110",
  60076=>"011111111",
  60077=>"000001000",
  60078=>"111111000",
  60079=>"000000111",
  60080=>"111111111",
  60081=>"000001111",
  60082=>"110111010",
  60083=>"111001000",
  60084=>"000010000",
  60085=>"000010000",
  60086=>"000011111",
  60087=>"000110111",
  60088=>"111111111",
  60089=>"111111011",
  60090=>"111110000",
  60091=>"110110100",
  60092=>"000000000",
  60093=>"010111111",
  60094=>"000000000",
  60095=>"111111111",
  60096=>"000000111",
  60097=>"111001000",
  60098=>"011000001",
  60099=>"111000000",
  60100=>"111000111",
  60101=>"001001100",
  60102=>"100100111",
  60103=>"111011000",
  60104=>"000000110",
  60105=>"111000110",
  60106=>"000000100",
  60107=>"000000000",
  60108=>"111111111",
  60109=>"110111000",
  60110=>"000000010",
  60111=>"000000000",
  60112=>"101000000",
  60113=>"000000011",
  60114=>"000000011",
  60115=>"000000000",
  60116=>"000000000",
  60117=>"111111111",
  60118=>"000100100",
  60119=>"111001111",
  60120=>"111111111",
  60121=>"111111000",
  60122=>"111111110",
  60123=>"010111111",
  60124=>"000000111",
  60125=>"110100110",
  60126=>"000011111",
  60127=>"000110111",
  60128=>"000000000",
  60129=>"000000000",
  60130=>"000000000",
  60131=>"000111111",
  60132=>"101000111",
  60133=>"000000011",
  60134=>"011000000",
  60135=>"111111101",
  60136=>"111111011",
  60137=>"001000000",
  60138=>"010000000",
  60139=>"000110111",
  60140=>"000111100",
  60141=>"000000000",
  60142=>"011000000",
  60143=>"000000010",
  60144=>"111000000",
  60145=>"001001111",
  60146=>"000000000",
  60147=>"110110000",
  60148=>"000000100",
  60149=>"111011001",
  60150=>"100111011",
  60151=>"111111111",
  60152=>"000000100",
  60153=>"111111111",
  60154=>"111110000",
  60155=>"100101111",
  60156=>"111111001",
  60157=>"100100001",
  60158=>"011000000",
  60159=>"111111000",
  60160=>"000000000",
  60161=>"000000110",
  60162=>"111110111",
  60163=>"000001111",
  60164=>"111001000",
  60165=>"001000000",
  60166=>"111111111",
  60167=>"111000110",
  60168=>"000000001",
  60169=>"000000000",
  60170=>"100000110",
  60171=>"111111010",
  60172=>"110000110",
  60173=>"000000110",
  60174=>"000000110",
  60175=>"010111100",
  60176=>"111111111",
  60177=>"000000100",
  60178=>"000000000",
  60179=>"011111111",
  60180=>"111111111",
  60181=>"111101111",
  60182=>"000000111",
  60183=>"000000000",
  60184=>"000000000",
  60185=>"000111111",
  60186=>"000000000",
  60187=>"001000000",
  60188=>"011001111",
  60189=>"110111010",
  60190=>"111101010",
  60191=>"110100100",
  60192=>"100001011",
  60193=>"000100111",
  60194=>"110111111",
  60195=>"001000000",
  60196=>"000000011",
  60197=>"100000011",
  60198=>"000110110",
  60199=>"000000111",
  60200=>"111100000",
  60201=>"111111000",
  60202=>"110000111",
  60203=>"000011111",
  60204=>"000110000",
  60205=>"000000000",
  60206=>"000000000",
  60207=>"000000000",
  60208=>"000001110",
  60209=>"111110000",
  60210=>"011010100",
  60211=>"000000111",
  60212=>"000000000",
  60213=>"000100111",
  60214=>"111001000",
  60215=>"000000001",
  60216=>"100111000",
  60217=>"111111111",
  60218=>"000000100",
  60219=>"000011101",
  60220=>"001111111",
  60221=>"010111111",
  60222=>"001001001",
  60223=>"000000010",
  60224=>"001000000",
  60225=>"111110001",
  60226=>"101000110",
  60227=>"001000000",
  60228=>"001000001",
  60229=>"001111000",
  60230=>"111010000",
  60231=>"000000111",
  60232=>"000000000",
  60233=>"110000000",
  60234=>"000000000",
  60235=>"001110111",
  60236=>"101000000",
  60237=>"001111000",
  60238=>"000000111",
  60239=>"100111011",
  60240=>"101001101",
  60241=>"011001000",
  60242=>"000001110",
  60243=>"111110111",
  60244=>"000000000",
  60245=>"001011011",
  60246=>"000001000",
  60247=>"000000001",
  60248=>"110111111",
  60249=>"011000000",
  60250=>"111000111",
  60251=>"111001001",
  60252=>"000011111",
  60253=>"111101000",
  60254=>"000000010",
  60255=>"011011000",
  60256=>"111111000",
  60257=>"111111000",
  60258=>"111101001",
  60259=>"111111111",
  60260=>"011011111",
  60261=>"111110111",
  60262=>"111000000",
  60263=>"001000001",
  60264=>"000000010",
  60265=>"110110111",
  60266=>"011000010",
  60267=>"000100100",
  60268=>"011011001",
  60269=>"001111110",
  60270=>"111111000",
  60271=>"111111101",
  60272=>"000001011",
  60273=>"001001000",
  60274=>"111000111",
  60275=>"000000001",
  60276=>"000001111",
  60277=>"101000001",
  60278=>"001000000",
  60279=>"110011101",
  60280=>"000000011",
  60281=>"111111001",
  60282=>"111111111",
  60283=>"101100100",
  60284=>"000000101",
  60285=>"111111101",
  60286=>"001000000",
  60287=>"111110111",
  60288=>"000000011",
  60289=>"111111010",
  60290=>"111111011",
  60291=>"000000000",
  60292=>"111111111",
  60293=>"110110000",
  60294=>"111001000",
  60295=>"110110110",
  60296=>"000000100",
  60297=>"011011111",
  60298=>"000010111",
  60299=>"000110111",
  60300=>"111000111",
  60301=>"111111100",
  60302=>"111111000",
  60303=>"111111001",
  60304=>"101000000",
  60305=>"000000111",
  60306=>"110110010",
  60307=>"000011010",
  60308=>"111111110",
  60309=>"000000000",
  60310=>"000000010",
  60311=>"000011111",
  60312=>"000000000",
  60313=>"100110110",
  60314=>"111100101",
  60315=>"100010111",
  60316=>"000110111",
  60317=>"100000100",
  60318=>"111111000",
  60319=>"000000000",
  60320=>"111111000",
  60321=>"001000000",
  60322=>"000000111",
  60323=>"111010100",
  60324=>"111111001",
  60325=>"001001001",
  60326=>"111100000",
  60327=>"001001000",
  60328=>"000001111",
  60329=>"111111111",
  60330=>"010111010",
  60331=>"101000000",
  60332=>"111111010",
  60333=>"111111111",
  60334=>"011111111",
  60335=>"111111111",
  60336=>"110111110",
  60337=>"111111001",
  60338=>"000000111",
  60339=>"111111000",
  60340=>"111111111",
  60341=>"111111000",
  60342=>"000000001",
  60343=>"100000000",
  60344=>"000111111",
  60345=>"000011111",
  60346=>"010000000",
  60347=>"111000000",
  60348=>"000000000",
  60349=>"111100110",
  60350=>"000000100",
  60351=>"001100111",
  60352=>"000111111",
  60353=>"000000000",
  60354=>"000111010",
  60355=>"011111000",
  60356=>"111111111",
  60357=>"111011000",
  60358=>"001010010",
  60359=>"000000000",
  60360=>"000011010",
  60361=>"000000101",
  60362=>"111111001",
  60363=>"100100111",
  60364=>"000000011",
  60365=>"000000010",
  60366=>"111101011",
  60367=>"000000001",
  60368=>"001001000",
  60369=>"010111000",
  60370=>"000000000",
  60371=>"111010111",
  60372=>"011111011",
  60373=>"000000000",
  60374=>"111111000",
  60375=>"110100110",
  60376=>"000000111",
  60377=>"111111000",
  60378=>"000000000",
  60379=>"000010111",
  60380=>"111111110",
  60381=>"111111111",
  60382=>"101011000",
  60383=>"000000111",
  60384=>"001111000",
  60385=>"101000000",
  60386=>"101100110",
  60387=>"100100110",
  60388=>"111000000",
  60389=>"100111100",
  60390=>"000110110",
  60391=>"111110000",
  60392=>"111101010",
  60393=>"000000000",
  60394=>"000000111",
  60395=>"100000100",
  60396=>"000000001",
  60397=>"000000001",
  60398=>"111111000",
  60399=>"010000000",
  60400=>"000111111",
  60401=>"000000000",
  60402=>"111000000",
  60403=>"010111011",
  60404=>"010000000",
  60405=>"000000000",
  60406=>"000000000",
  60407=>"110001000",
  60408=>"000111111",
  60409=>"011000110",
  60410=>"111000000",
  60411=>"000000111",
  60412=>"111000000",
  60413=>"111111110",
  60414=>"000001011",
  60415=>"000111111",
  60416=>"000000000",
  60417=>"111111111",
  60418=>"000000000",
  60419=>"010000000",
  60420=>"111111011",
  60421=>"110000000",
  60422=>"111111101",
  60423=>"000000000",
  60424=>"000101001",
  60425=>"110000000",
  60426=>"001000000",
  60427=>"000000011",
  60428=>"111111001",
  60429=>"000000010",
  60430=>"000100100",
  60431=>"111111111",
  60432=>"111000111",
  60433=>"111111111",
  60434=>"111111010",
  60435=>"000000000",
  60436=>"111111111",
  60437=>"000001111",
  60438=>"000000000",
  60439=>"001001001",
  60440=>"000001001",
  60441=>"011111001",
  60442=>"001011111",
  60443=>"111111111",
  60444=>"100000000",
  60445=>"000011111",
  60446=>"000000000",
  60447=>"000001111",
  60448=>"000000000",
  60449=>"101000000",
  60450=>"011111111",
  60451=>"111111111",
  60452=>"000000100",
  60453=>"011110111",
  60454=>"111111111",
  60455=>"100100000",
  60456=>"111111111",
  60457=>"001001101",
  60458=>"000000101",
  60459=>"110110110",
  60460=>"001000111",
  60461=>"011011100",
  60462=>"111111111",
  60463=>"111111000",
  60464=>"000010110",
  60465=>"000000111",
  60466=>"100111100",
  60467=>"111111111",
  60468=>"000111110",
  60469=>"100110010",
  60470=>"000001000",
  60471=>"110100110",
  60472=>"000000000",
  60473=>"111000000",
  60474=>"111111111",
  60475=>"000000000",
  60476=>"111111111",
  60477=>"000011011",
  60478=>"110111011",
  60479=>"000000000",
  60480=>"001000011",
  60481=>"111001100",
  60482=>"111001001",
  60483=>"000000000",
  60484=>"111000011",
  60485=>"100001111",
  60486=>"110010010",
  60487=>"111111111",
  60488=>"111110110",
  60489=>"110000000",
  60490=>"000000001",
  60491=>"111011011",
  60492=>"100110111",
  60493=>"000000111",
  60494=>"111111111",
  60495=>"110111111",
  60496=>"111111111",
  60497=>"000000000",
  60498=>"000000000",
  60499=>"110110010",
  60500=>"000001001",
  60501=>"000111111",
  60502=>"110110000",
  60503=>"000010111",
  60504=>"000000110",
  60505=>"110010010",
  60506=>"100000000",
  60507=>"011000000",
  60508=>"000001000",
  60509=>"010111111",
  60510=>"111111111",
  60511=>"111011000",
  60512=>"111011111",
  60513=>"000001000",
  60514=>"111000000",
  60515=>"000000000",
  60516=>"101101011",
  60517=>"110000101",
  60518=>"111000000",
  60519=>"000000001",
  60520=>"000000000",
  60521=>"000010010",
  60522=>"011011011",
  60523=>"111111111",
  60524=>"000000000",
  60525=>"111111001",
  60526=>"100100100",
  60527=>"110111111",
  60528=>"100110100",
  60529=>"111111011",
  60530=>"100100100",
  60531=>"000000000",
  60532=>"111000001",
  60533=>"000000000",
  60534=>"111010000",
  60535=>"000000001",
  60536=>"111100110",
  60537=>"000001111",
  60538=>"110110111",
  60539=>"111111111",
  60540=>"100000000",
  60541=>"111011001",
  60542=>"000000000",
  60543=>"000000000",
  60544=>"111111110",
  60545=>"111110000",
  60546=>"111111111",
  60547=>"111101111",
  60548=>"111111111",
  60549=>"110110110",
  60550=>"111111111",
  60551=>"000000000",
  60552=>"000000000",
  60553=>"110000001",
  60554=>"000000000",
  60555=>"000000111",
  60556=>"111101011",
  60557=>"000000110",
  60558=>"000001011",
  60559=>"011110110",
  60560=>"000000000",
  60561=>"000000001",
  60562=>"110100101",
  60563=>"111111001",
  60564=>"000000000",
  60565=>"000000001",
  60566=>"000000000",
  60567=>"000000000",
  60568=>"001001101",
  60569=>"000011111",
  60570=>"111110110",
  60571=>"000000000",
  60572=>"111111111",
  60573=>"000001001",
  60574=>"000001111",
  60575=>"111111111",
  60576=>"111111110",
  60577=>"110110111",
  60578=>"111110110",
  60579=>"000000000",
  60580=>"011110000",
  60581=>"101111101",
  60582=>"100000000",
  60583=>"011011000",
  60584=>"010111011",
  60585=>"000000000",
  60586=>"100100100",
  60587=>"000000000",
  60588=>"111011011",
  60589=>"110110110",
  60590=>"000010000",
  60591=>"000011001",
  60592=>"111111101",
  60593=>"101101001",
  60594=>"111000000",
  60595=>"000000000",
  60596=>"111111100",
  60597=>"110111111",
  60598=>"000000000",
  60599=>"111000000",
  60600=>"001111111",
  60601=>"101000000",
  60602=>"000000000",
  60603=>"010010011",
  60604=>"000000111",
  60605=>"000000001",
  60606=>"000110010",
  60607=>"011000000",
  60608=>"100000000",
  60609=>"111111111",
  60610=>"011001000",
  60611=>"000000001",
  60612=>"111010000",
  60613=>"101111000",
  60614=>"000000110",
  60615=>"000000000",
  60616=>"111111111",
  60617=>"111111111",
  60618=>"000000000",
  60619=>"111111111",
  60620=>"000110110",
  60621=>"111111111",
  60622=>"101001001",
  60623=>"000000001",
  60624=>"010011000",
  60625=>"100000000",
  60626=>"010110000",
  60627=>"001001111",
  60628=>"111010111",
  60629=>"010011000",
  60630=>"000111111",
  60631=>"101001001",
  60632=>"000000001",
  60633=>"000000000",
  60634=>"000000111",
  60635=>"000100101",
  60636=>"000000000",
  60637=>"000010111",
  60638=>"001111111",
  60639=>"111111111",
  60640=>"111111110",
  60641=>"111100110",
  60642=>"010111110",
  60643=>"000110111",
  60644=>"011111111",
  60645=>"110111111",
  60646=>"001000100",
  60647=>"111111001",
  60648=>"111111111",
  60649=>"001000001",
  60650=>"111111111",
  60651=>"111111111",
  60652=>"000111111",
  60653=>"111111000",
  60654=>"000000111",
  60655=>"000111111",
  60656=>"101111111",
  60657=>"111111111",
  60658=>"111111111",
  60659=>"111111111",
  60660=>"111110000",
  60661=>"110000000",
  60662=>"001001011",
  60663=>"000000000",
  60664=>"000000000",
  60665=>"111110101",
  60666=>"000111111",
  60667=>"000100100",
  60668=>"110111111",
  60669=>"111111011",
  60670=>"001011111",
  60671=>"001000000",
  60672=>"001011011",
  60673=>"000000000",
  60674=>"000001000",
  60675=>"111111111",
  60676=>"111111000",
  60677=>"001001001",
  60678=>"111110000",
  60679=>"111110001",
  60680=>"111111110",
  60681=>"000000000",
  60682=>"110000111",
  60683=>"111011001",
  60684=>"000000110",
  60685=>"000110111",
  60686=>"111111111",
  60687=>"000110111",
  60688=>"000100101",
  60689=>"000110000",
  60690=>"111011011",
  60691=>"100111111",
  60692=>"000000001",
  60693=>"000000000",
  60694=>"100000000",
  60695=>"000000000",
  60696=>"111111111",
  60697=>"000000111",
  60698=>"100111001",
  60699=>"011010000",
  60700=>"111011001",
  60701=>"111111111",
  60702=>"000000000",
  60703=>"000000000",
  60704=>"110111000",
  60705=>"000000000",
  60706=>"100100111",
  60707=>"000000000",
  60708=>"110110110",
  60709=>"111101000",
  60710=>"000000000",
  60711=>"100000001",
  60712=>"111111111",
  60713=>"111111111",
  60714=>"000110110",
  60715=>"110111010",
  60716=>"000000000",
  60717=>"000000000",
  60718=>"000000000",
  60719=>"001001000",
  60720=>"100000000",
  60721=>"001000000",
  60722=>"100110110",
  60723=>"000000000",
  60724=>"000000000",
  60725=>"110100000",
  60726=>"000111111",
  60727=>"111000000",
  60728=>"001000000",
  60729=>"111100100",
  60730=>"000000111",
  60731=>"101100100",
  60732=>"000111111",
  60733=>"111010000",
  60734=>"010000000",
  60735=>"011001001",
  60736=>"111110110",
  60737=>"111111111",
  60738=>"000000000",
  60739=>"111111111",
  60740=>"000000010",
  60741=>"111100111",
  60742=>"111111000",
  60743=>"111100100",
  60744=>"000000000",
  60745=>"111111111",
  60746=>"000100110",
  60747=>"111111001",
  60748=>"000000000",
  60749=>"001111111",
  60750=>"000000000",
  60751=>"001001001",
  60752=>"000000001",
  60753=>"000000000",
  60754=>"111111111",
  60755=>"011001011",
  60756=>"001000000",
  60757=>"111101101",
  60758=>"000000110",
  60759=>"110110100",
  60760=>"111111111",
  60761=>"111111111",
  60762=>"000001111",
  60763=>"110100000",
  60764=>"111100100",
  60765=>"000000000",
  60766=>"111111111",
  60767=>"100000000",
  60768=>"000011111",
  60769=>"000000111",
  60770=>"000000000",
  60771=>"100100111",
  60772=>"001001111",
  60773=>"001110000",
  60774=>"000000000",
  60775=>"011011001",
  60776=>"110110110",
  60777=>"111111010",
  60778=>"100000111",
  60779=>"111111111",
  60780=>"111111011",
  60781=>"111111111",
  60782=>"111111111",
  60783=>"000000000",
  60784=>"111010000",
  60785=>"000000101",
  60786=>"000000000",
  60787=>"111111111",
  60788=>"000000001",
  60789=>"000000000",
  60790=>"000000010",
  60791=>"000000000",
  60792=>"000000111",
  60793=>"110111111",
  60794=>"111011000",
  60795=>"000011111",
  60796=>"010110110",
  60797=>"000000000",
  60798=>"000000011",
  60799=>"000000000",
  60800=>"001001011",
  60801=>"000111101",
  60802=>"110110111",
  60803=>"000000000",
  60804=>"000111111",
  60805=>"000000000",
  60806=>"000000000",
  60807=>"000001001",
  60808=>"100000000",
  60809=>"000000000",
  60810=>"001000000",
  60811=>"000000000",
  60812=>"111111111",
  60813=>"110110110",
  60814=>"000011010",
  60815=>"111111111",
  60816=>"000000000",
  60817=>"011011011",
  60818=>"000011011",
  60819=>"000011111",
  60820=>"111111111",
  60821=>"000001001",
  60822=>"000000000",
  60823=>"110010000",
  60824=>"111111111",
  60825=>"110111111",
  60826=>"000000000",
  60827=>"011111111",
  60828=>"111100111",
  60829=>"000000000",
  60830=>"000111111",
  60831=>"100000000",
  60832=>"000000100",
  60833=>"010110110",
  60834=>"111111101",
  60835=>"000000000",
  60836=>"100100111",
  60837=>"000000000",
  60838=>"000111000",
  60839=>"000111111",
  60840=>"100000000",
  60841=>"111100100",
  60842=>"110110111",
  60843=>"000010110",
  60844=>"111100000",
  60845=>"000000100",
  60846=>"000000111",
  60847=>"111011000",
  60848=>"111100100",
  60849=>"111001011",
  60850=>"000000000",
  60851=>"000000111",
  60852=>"001001011",
  60853=>"000100000",
  60854=>"101111111",
  60855=>"111110001",
  60856=>"011011111",
  60857=>"111111111",
  60858=>"110000000",
  60859=>"111111111",
  60860=>"111111111",
  60861=>"000000000",
  60862=>"111111111",
  60863=>"010010010",
  60864=>"000000000",
  60865=>"000000000",
  60866=>"000000000",
  60867=>"000000000",
  60868=>"000000000",
  60869=>"000000010",
  60870=>"010110000",
  60871=>"000000100",
  60872=>"000010000",
  60873=>"011000000",
  60874=>"110111111",
  60875=>"111111111",
  60876=>"111110000",
  60877=>"000000111",
  60878=>"000000000",
  60879=>"000000100",
  60880=>"110111110",
  60881=>"001001001",
  60882=>"000000000",
  60883=>"111111111",
  60884=>"000111111",
  60885=>"000110110",
  60886=>"011011000",
  60887=>"100100100",
  60888=>"100100001",
  60889=>"111110111",
  60890=>"111110000",
  60891=>"110000000",
  60892=>"111111111",
  60893=>"111111111",
  60894=>"000000000",
  60895=>"001001111",
  60896=>"111000100",
  60897=>"111110110",
  60898=>"111111110",
  60899=>"111101111",
  60900=>"100100110",
  60901=>"111111111",
  60902=>"000000000",
  60903=>"000000000",
  60904=>"101001001",
  60905=>"000000000",
  60906=>"111111011",
  60907=>"111111111",
  60908=>"110100100",
  60909=>"111011000",
  60910=>"001000111",
  60911=>"111110000",
  60912=>"000011000",
  60913=>"111111111",
  60914=>"000100111",
  60915=>"000000000",
  60916=>"000000000",
  60917=>"000001001",
  60918=>"000000000",
  60919=>"000000000",
  60920=>"000110111",
  60921=>"000010010",
  60922=>"111111000",
  60923=>"100100000",
  60924=>"111100000",
  60925=>"001110111",
  60926=>"000000001",
  60927=>"111111111",
  60928=>"001101000",
  60929=>"111011000",
  60930=>"000000000",
  60931=>"000000011",
  60932=>"111001101",
  60933=>"111101000",
  60934=>"001000000",
  60935=>"111111111",
  60936=>"000000000",
  60937=>"110110111",
  60938=>"000100111",
  60939=>"101111100",
  60940=>"100000010",
  60941=>"000110110",
  60942=>"000111111",
  60943=>"100000011",
  60944=>"000000000",
  60945=>"100001111",
  60946=>"111111101",
  60947=>"111111100",
  60948=>"000000000",
  60949=>"111111111",
  60950=>"111111111",
  60951=>"111100111",
  60952=>"000000000",
  60953=>"111001001",
  60954=>"110010011",
  60955=>"000000000",
  60956=>"000000000",
  60957=>"100111111",
  60958=>"011000000",
  60959=>"111110000",
  60960=>"000111111",
  60961=>"000001000",
  60962=>"001111111",
  60963=>"100111111",
  60964=>"011001000",
  60965=>"000001000",
  60966=>"000000111",
  60967=>"001001111",
  60968=>"000111110",
  60969=>"000000111",
  60970=>"111111010",
  60971=>"010011111",
  60972=>"000000000",
  60973=>"011111000",
  60974=>"001001001",
  60975=>"110100000",
  60976=>"011000000",
  60977=>"111001111",
  60978=>"101111111",
  60979=>"000000100",
  60980=>"111101111",
  60981=>"101000000",
  60982=>"000111111",
  60983=>"111111111",
  60984=>"000110000",
  60985=>"000000110",
  60986=>"111111011",
  60987=>"000000000",
  60988=>"000000111",
  60989=>"000011111",
  60990=>"000000000",
  60991=>"001001000",
  60992=>"000000111",
  60993=>"011111111",
  60994=>"011011111",
  60995=>"000100110",
  60996=>"000010100",
  60997=>"011000000",
  60998=>"010111110",
  60999=>"100100111",
  61000=>"111100001",
  61001=>"110110111",
  61002=>"000111111",
  61003=>"000000000",
  61004=>"110111100",
  61005=>"111000000",
  61006=>"100000000",
  61007=>"011111111",
  61008=>"000101110",
  61009=>"100110111",
  61010=>"010111110",
  61011=>"001000011",
  61012=>"101100111",
  61013=>"000000110",
  61014=>"000000011",
  61015=>"111000011",
  61016=>"000000000",
  61017=>"000000111",
  61018=>"000000100",
  61019=>"100110100",
  61020=>"000000000",
  61021=>"000000000",
  61022=>"111111100",
  61023=>"100000001",
  61024=>"100000000",
  61025=>"110110110",
  61026=>"111111111",
  61027=>"100100111",
  61028=>"111111111",
  61029=>"000000011",
  61030=>"111111011",
  61031=>"110100100",
  61032=>"000000110",
  61033=>"111110000",
  61034=>"000000000",
  61035=>"111000000",
  61036=>"000100001",
  61037=>"111111111",
  61038=>"100111000",
  61039=>"000000000",
  61040=>"110111110",
  61041=>"000010111",
  61042=>"101001111",
  61043=>"110110110",
  61044=>"011111111",
  61045=>"010000000",
  61046=>"001000111",
  61047=>"111111111",
  61048=>"110111111",
  61049=>"100000000",
  61050=>"110000110",
  61051=>"000010110",
  61052=>"000001000",
  61053=>"000011111",
  61054=>"100000000",
  61055=>"111111111",
  61056=>"000000000",
  61057=>"011111111",
  61058=>"110110000",
  61059=>"000000000",
  61060=>"000000000",
  61061=>"110100111",
  61062=>"000111111",
  61063=>"111100000",
  61064=>"000000000",
  61065=>"000000000",
  61066=>"111111111",
  61067=>"001111111",
  61068=>"101111000",
  61069=>"000001111",
  61070=>"001001111",
  61071=>"111111100",
  61072=>"000000000",
  61073=>"111011001",
  61074=>"000111111",
  61075=>"000000000",
  61076=>"001000000",
  61077=>"111000000",
  61078=>"000000000",
  61079=>"100111000",
  61080=>"000111100",
  61081=>"000000000",
  61082=>"000000100",
  61083=>"111100000",
  61084=>"000111111",
  61085=>"000111101",
  61086=>"111011110",
  61087=>"000000000",
  61088=>"111111110",
  61089=>"000000000",
  61090=>"011011111",
  61091=>"111111111",
  61092=>"000000100",
  61093=>"011000010",
  61094=>"000000111",
  61095=>"100100101",
  61096=>"000111111",
  61097=>"000101101",
  61098=>"111111111",
  61099=>"111111000",
  61100=>"000000001",
  61101=>"000100000",
  61102=>"101000111",
  61103=>"110111111",
  61104=>"000111000",
  61105=>"111000001",
  61106=>"110110111",
  61107=>"111000000",
  61108=>"110000111",
  61109=>"100111111",
  61110=>"111000000",
  61111=>"101000111",
  61112=>"101111111",
  61113=>"000000000",
  61114=>"110000111",
  61115=>"100001111",
  61116=>"000111111",
  61117=>"001111111",
  61118=>"100111110",
  61119=>"000001001",
  61120=>"111111111",
  61121=>"111110100",
  61122=>"001000000",
  61123=>"000000100",
  61124=>"111111000",
  61125=>"000000100",
  61126=>"110000111",
  61127=>"000001111",
  61128=>"100111111",
  61129=>"111111110",
  61130=>"100100101",
  61131=>"111101111",
  61132=>"000111111",
  61133=>"101101111",
  61134=>"000000000",
  61135=>"000100111",
  61136=>"000000000",
  61137=>"111111000",
  61138=>"111010000",
  61139=>"000000000",
  61140=>"100100111",
  61141=>"000001000",
  61142=>"000000010",
  61143=>"000001001",
  61144=>"110000100",
  61145=>"100111000",
  61146=>"010000000",
  61147=>"000111111",
  61148=>"000001000",
  61149=>"000000000",
  61150=>"111000000",
  61151=>"111001001",
  61152=>"000000000",
  61153=>"000110000",
  61154=>"110111000",
  61155=>"111111100",
  61156=>"111010111",
  61157=>"101111111",
  61158=>"110111111",
  61159=>"111111111",
  61160=>"001111011",
  61161=>"010100111",
  61162=>"111111111",
  61163=>"000000000",
  61164=>"000000000",
  61165=>"111111011",
  61166=>"111000011",
  61167=>"111100000",
  61168=>"101100111",
  61169=>"111000000",
  61170=>"110111111",
  61171=>"000001111",
  61172=>"111111100",
  61173=>"000000100",
  61174=>"000100000",
  61175=>"110000100",
  61176=>"001000000",
  61177=>"110001111",
  61178=>"000111111",
  61179=>"000000001",
  61180=>"111111011",
  61181=>"111111101",
  61182=>"001001001",
  61183=>"011011000",
  61184=>"100111111",
  61185=>"110110110",
  61186=>"111111000",
  61187=>"101111101",
  61188=>"110111111",
  61189=>"000011000",
  61190=>"010111011",
  61191=>"001011011",
  61192=>"000001111",
  61193=>"000000000",
  61194=>"000000000",
  61195=>"001000000",
  61196=>"010110110",
  61197=>"000000100",
  61198=>"000000000",
  61199=>"000001001",
  61200=>"011000000",
  61201=>"000000000",
  61202=>"111011011",
  61203=>"111111000",
  61204=>"111111110",
  61205=>"000000000",
  61206=>"110001001",
  61207=>"111111111",
  61208=>"111111111",
  61209=>"111000000",
  61210=>"010110000",
  61211=>"111111011",
  61212=>"000000100",
  61213=>"001000000",
  61214=>"000000111",
  61215=>"111100000",
  61216=>"000011001",
  61217=>"011011000",
  61218=>"111111111",
  61219=>"111111111",
  61220=>"000011000",
  61221=>"000000000",
  61222=>"001101111",
  61223=>"000010001",
  61224=>"111000000",
  61225=>"000000101",
  61226=>"000000000",
  61227=>"000000010",
  61228=>"101001101",
  61229=>"000000101",
  61230=>"000000000",
  61231=>"000000111",
  61232=>"001001111",
  61233=>"111111001",
  61234=>"000011111",
  61235=>"110000000",
  61236=>"000111000",
  61237=>"000001111",
  61238=>"111100000",
  61239=>"100000000",
  61240=>"000000010",
  61241=>"000100110",
  61242=>"111000001",
  61243=>"001011011",
  61244=>"000000111",
  61245=>"100100111",
  61246=>"111111111",
  61247=>"111111111",
  61248=>"000001000",
  61249=>"100111110",
  61250=>"000000000",
  61251=>"000000000",
  61252=>"101111111",
  61253=>"000111011",
  61254=>"100100110",
  61255=>"111111111",
  61256=>"000000011",
  61257=>"010000000",
  61258=>"001000000",
  61259=>"111111111",
  61260=>"111111000",
  61261=>"010000000",
  61262=>"000111010",
  61263=>"001001001",
  61264=>"101101110",
  61265=>"011011010",
  61266=>"101000111",
  61267=>"100000111",
  61268=>"111100111",
  61269=>"111111111",
  61270=>"101000000",
  61271=>"110110111",
  61272=>"000000000",
  61273=>"110110000",
  61274=>"101111111",
  61275=>"000110000",
  61276=>"111111111",
  61277=>"001001001",
  61278=>"110111111",
  61279=>"111111111",
  61280=>"011111111",
  61281=>"111111111",
  61282=>"100000000",
  61283=>"100000000",
  61284=>"000000000",
  61285=>"000001011",
  61286=>"000000001",
  61287=>"000000000",
  61288=>"111111111",
  61289=>"000111000",
  61290=>"000000111",
  61291=>"010010110",
  61292=>"011111010",
  61293=>"110011111",
  61294=>"001001001",
  61295=>"111111110",
  61296=>"111111101",
  61297=>"111011111",
  61298=>"000100100",
  61299=>"101001001",
  61300=>"111111111",
  61301=>"111011000",
  61302=>"011111100",
  61303=>"000000000",
  61304=>"000000100",
  61305=>"000000000",
  61306=>"000000111",
  61307=>"111101001",
  61308=>"011110100",
  61309=>"000111111",
  61310=>"000000000",
  61311=>"111111000",
  61312=>"000010000",
  61313=>"011010000",
  61314=>"110000000",
  61315=>"000000000",
  61316=>"000000000",
  61317=>"000100000",
  61318=>"111111111",
  61319=>"111111111",
  61320=>"010110000",
  61321=>"110110111",
  61322=>"000000000",
  61323=>"100101000",
  61324=>"000100101",
  61325=>"110111011",
  61326=>"001111000",
  61327=>"000000111",
  61328=>"111111111",
  61329=>"111111110",
  61330=>"000111111",
  61331=>"000000000",
  61332=>"000000000",
  61333=>"011000001",
  61334=>"111101100",
  61335=>"100000100",
  61336=>"011000000",
  61337=>"010111110",
  61338=>"000000111",
  61339=>"001001001",
  61340=>"000000101",
  61341=>"000000000",
  61342=>"111000111",
  61343=>"111111010",
  61344=>"011110111",
  61345=>"111011011",
  61346=>"100111111",
  61347=>"000010010",
  61348=>"000111110",
  61349=>"011111011",
  61350=>"000000000",
  61351=>"100000110",
  61352=>"111111111",
  61353=>"000000101",
  61354=>"111111100",
  61355=>"101101001",
  61356=>"000110111",
  61357=>"111111010",
  61358=>"000001111",
  61359=>"011000111",
  61360=>"000000000",
  61361=>"011000000",
  61362=>"111111100",
  61363=>"000000000",
  61364=>"000100000",
  61365=>"000001101",
  61366=>"100110000",
  61367=>"100000000",
  61368=>"000000000",
  61369=>"110110011",
  61370=>"111111110",
  61371=>"111111000",
  61372=>"011110111",
  61373=>"000111111",
  61374=>"000010111",
  61375=>"100110110",
  61376=>"000000000",
  61377=>"110110010",
  61378=>"100100110",
  61379=>"111111001",
  61380=>"100110000",
  61381=>"101100001",
  61382=>"100000111",
  61383=>"111110000",
  61384=>"000000000",
  61385=>"001001001",
  61386=>"000110100",
  61387=>"000111111",
  61388=>"000000000",
  61389=>"100000000",
  61390=>"110110001",
  61391=>"000000000",
  61392=>"001001111",
  61393=>"100000000",
  61394=>"100010000",
  61395=>"111111111",
  61396=>"000010000",
  61397=>"111000000",
  61398=>"000010110",
  61399=>"000000101",
  61400=>"000100011",
  61401=>"000000110",
  61402=>"101100000",
  61403=>"100100100",
  61404=>"111101101",
  61405=>"001011011",
  61406=>"100000000",
  61407=>"110100011",
  61408=>"111111111",
  61409=>"001111111",
  61410=>"010000111",
  61411=>"000000000",
  61412=>"011111111",
  61413=>"000000010",
  61414=>"011011000",
  61415=>"111100000",
  61416=>"001111101",
  61417=>"101111111",
  61418=>"100100101",
  61419=>"111111100",
  61420=>"000000000",
  61421=>"111100011",
  61422=>"101111110",
  61423=>"100111111",
  61424=>"100000100",
  61425=>"111001000",
  61426=>"000000000",
  61427=>"000000111",
  61428=>"000111001",
  61429=>"111111010",
  61430=>"111111111",
  61431=>"111111001",
  61432=>"110110110",
  61433=>"001101111",
  61434=>"111000001",
  61435=>"100100110",
  61436=>"110100000",
  61437=>"001000000",
  61438=>"000111111",
  61439=>"001111001",
  61440=>"000000000",
  61441=>"000001111",
  61442=>"000111111",
  61443=>"000111111",
  61444=>"100000100",
  61445=>"001111111",
  61446=>"111111000",
  61447=>"100110111",
  61448=>"111111010",
  61449=>"111111111",
  61450=>"111011011",
  61451=>"100000000",
  61452=>"100111111",
  61453=>"000000011",
  61454=>"110111111",
  61455=>"100101111",
  61456=>"110110111",
  61457=>"110111111",
  61458=>"000011110",
  61459=>"000101101",
  61460=>"111111111",
  61461=>"111101111",
  61462=>"111011011",
  61463=>"011001110",
  61464=>"000000100",
  61465=>"000000000",
  61466=>"111111111",
  61467=>"110100111",
  61468=>"111010000",
  61469=>"111000000",
  61470=>"000001001",
  61471=>"000000000",
  61472=>"111111010",
  61473=>"101111000",
  61474=>"111111111",
  61475=>"010010000",
  61476=>"001111111",
  61477=>"000110111",
  61478=>"111101110",
  61479=>"000000000",
  61480=>"000000000",
  61481=>"000100101",
  61482=>"000000000",
  61483=>"000000110",
  61484=>"110111111",
  61485=>"001101100",
  61486=>"111100000",
  61487=>"111111000",
  61488=>"110111111",
  61489=>"000000000",
  61490=>"000000000",
  61491=>"000000000",
  61492=>"000101000",
  61493=>"110111110",
  61494=>"111111111",
  61495=>"000000010",
  61496=>"111111111",
  61497=>"100100000",
  61498=>"111101000",
  61499=>"001000111",
  61500=>"111111010",
  61501=>"001011010",
  61502=>"000000000",
  61503=>"100110111",
  61504=>"000000000",
  61505=>"000000000",
  61506=>"111111110",
  61507=>"110111011",
  61508=>"000000000",
  61509=>"111111111",
  61510=>"000000000",
  61511=>"111111111",
  61512=>"011011011",
  61513=>"011111111",
  61514=>"000001000",
  61515=>"111000000",
  61516=>"000000000",
  61517=>"110110001",
  61518=>"111111111",
  61519=>"100111111",
  61520=>"000000000",
  61521=>"000000000",
  61522=>"110111111",
  61523=>"000001111",
  61524=>"000000000",
  61525=>"000111111",
  61526=>"111111111",
  61527=>"111111111",
  61528=>"000000000",
  61529=>"010000000",
  61530=>"000000000",
  61531=>"000000001",
  61532=>"111000111",
  61533=>"000111111",
  61534=>"111111111",
  61535=>"000011111",
  61536=>"000000000",
  61537=>"111111111",
  61538=>"111111111",
  61539=>"000000100",
  61540=>"001111101",
  61541=>"000000001",
  61542=>"001101001",
  61543=>"000011000",
  61544=>"000000000",
  61545=>"111111111",
  61546=>"111111111",
  61547=>"111111111",
  61548=>"000000000",
  61549=>"110000000",
  61550=>"111000000",
  61551=>"011111111",
  61552=>"100111111",
  61553=>"001111111",
  61554=>"011111000",
  61555=>"000111100",
  61556=>"111111011",
  61557=>"000000010",
  61558=>"111111111",
  61559=>"111111111",
  61560=>"000000000",
  61561=>"000000000",
  61562=>"010001000",
  61563=>"000000000",
  61564=>"100000000",
  61565=>"011011000",
  61566=>"111111000",
  61567=>"011001001",
  61568=>"000000000",
  61569=>"011000011",
  61570=>"111101000",
  61571=>"000000000",
  61572=>"100111111",
  61573=>"000000000",
  61574=>"111111110",
  61575=>"111111110",
  61576=>"111111111",
  61577=>"111111111",
  61578=>"000000000",
  61579=>"000000010",
  61580=>"011111110",
  61581=>"111111000",
  61582=>"000010111",
  61583=>"111111000",
  61584=>"000000000",
  61585=>"000000000",
  61586=>"000000111",
  61587=>"111111111",
  61588=>"110111000",
  61589=>"000000000",
  61590=>"111011001",
  61591=>"111100000",
  61592=>"111110111",
  61593=>"101111111",
  61594=>"000111111",
  61595=>"000000000",
  61596=>"111110111",
  61597=>"000000001",
  61598=>"000000000",
  61599=>"001001101",
  61600=>"111001111",
  61601=>"111111010",
  61602=>"001001011",
  61603=>"111111111",
  61604=>"101101000",
  61605=>"111111111",
  61606=>"000110110",
  61607=>"010110000",
  61608=>"000010000",
  61609=>"111111111",
  61610=>"101000111",
  61611=>"011000000",
  61612=>"111110110",
  61613=>"000100000",
  61614=>"000000000",
  61615=>"000001000",
  61616=>"001111001",
  61617=>"000001011",
  61618=>"111111100",
  61619=>"011111000",
  61620=>"011001000",
  61621=>"001001111",
  61622=>"110000000",
  61623=>"111111111",
  61624=>"000000000",
  61625=>"111111000",
  61626=>"111111011",
  61627=>"110010010",
  61628=>"000000111",
  61629=>"000000001",
  61630=>"000000000",
  61631=>"110000001",
  61632=>"110110111",
  61633=>"110010000",
  61634=>"111011001",
  61635=>"000000000",
  61636=>"000110000",
  61637=>"111000010",
  61638=>"010010111",
  61639=>"000001011",
  61640=>"000000000",
  61641=>"000111111",
  61642=>"000011011",
  61643=>"001001111",
  61644=>"000110110",
  61645=>"110110111",
  61646=>"000000111",
  61647=>"111010000",
  61648=>"000111111",
  61649=>"000101000",
  61650=>"000001111",
  61651=>"000000111",
  61652=>"101111001",
  61653=>"100110100",
  61654=>"010011010",
  61655=>"001001000",
  61656=>"111111111",
  61657=>"000000000",
  61658=>"111111000",
  61659=>"111111111",
  61660=>"101000000",
  61661=>"010001000",
  61662=>"000110100",
  61663=>"011000000",
  61664=>"000000000",
  61665=>"101111111",
  61666=>"111000000",
  61667=>"001000001",
  61668=>"000000000",
  61669=>"110000100",
  61670=>"001000000",
  61671=>"011010000",
  61672=>"000000000",
  61673=>"000000000",
  61674=>"000010111",
  61675=>"111101111",
  61676=>"111111111",
  61677=>"001000001",
  61678=>"000101111",
  61679=>"111011011",
  61680=>"111110000",
  61681=>"000010010",
  61682=>"000011111",
  61683=>"011111001",
  61684=>"111111001",
  61685=>"000011111",
  61686=>"111101000",
  61687=>"111110000",
  61688=>"000000000",
  61689=>"100110110",
  61690=>"111111111",
  61691=>"110111111",
  61692=>"000000000",
  61693=>"000110011",
  61694=>"111111000",
  61695=>"010010000",
  61696=>"000010011",
  61697=>"010010010",
  61698=>"000011001",
  61699=>"100111100",
  61700=>"000000000",
  61701=>"111111111",
  61702=>"110000000",
  61703=>"111111100",
  61704=>"111111111",
  61705=>"000100000",
  61706=>"111000110",
  61707=>"000000000",
  61708=>"000000000",
  61709=>"111000000",
  61710=>"111110110",
  61711=>"000000000",
  61712=>"100111111",
  61713=>"111111111",
  61714=>"111111010",
  61715=>"100110111",
  61716=>"111100000",
  61717=>"111111111",
  61718=>"000000000",
  61719=>"110110000",
  61720=>"000000000",
  61721=>"000011000",
  61722=>"101111001",
  61723=>"011000110",
  61724=>"100000000",
  61725=>"001000111",
  61726=>"001001000",
  61727=>"111101101",
  61728=>"000000000",
  61729=>"111111111",
  61730=>"111000000",
  61731=>"111011111",
  61732=>"000000001",
  61733=>"001001111",
  61734=>"001001000",
  61735=>"111001101",
  61736=>"000000000",
  61737=>"001000000",
  61738=>"000111111",
  61739=>"000000000",
  61740=>"101001000",
  61741=>"110100000",
  61742=>"000111001",
  61743=>"000000000",
  61744=>"000000010",
  61745=>"111111111",
  61746=>"011111111",
  61747=>"111111111",
  61748=>"111111111",
  61749=>"000000000",
  61750=>"100000000",
  61751=>"000111111",
  61752=>"000000000",
  61753=>"011000000",
  61754=>"011111011",
  61755=>"100000000",
  61756=>"011011000",
  61757=>"000111111",
  61758=>"110111111",
  61759=>"101000000",
  61760=>"000111111",
  61761=>"111111011",
  61762=>"000010111",
  61763=>"000000000",
  61764=>"000111111",
  61765=>"000110111",
  61766=>"000011001",
  61767=>"011000000",
  61768=>"000000000",
  61769=>"111111111",
  61770=>"111010011",
  61771=>"110100100",
  61772=>"000011001",
  61773=>"111111111",
  61774=>"110000000",
  61775=>"110110110",
  61776=>"000000000",
  61777=>"111110110",
  61778=>"111101000",
  61779=>"001111111",
  61780=>"000010010",
  61781=>"111111000",
  61782=>"000000101",
  61783=>"111111111",
  61784=>"000001100",
  61785=>"111111110",
  61786=>"111111111",
  61787=>"111111111",
  61788=>"011001000",
  61789=>"000000000",
  61790=>"111011000",
  61791=>"111111111",
  61792=>"111111111",
  61793=>"000000011",
  61794=>"000010010",
  61795=>"000000011",
  61796=>"000000100",
  61797=>"011001001",
  61798=>"111011111",
  61799=>"111010110",
  61800=>"000110010",
  61801=>"111111111",
  61802=>"101001000",
  61803=>"000111111",
  61804=>"110111111",
  61805=>"111111011",
  61806=>"000000000",
  61807=>"000110110",
  61808=>"001011111",
  61809=>"111111111",
  61810=>"100100101",
  61811=>"000111111",
  61812=>"111111111",
  61813=>"110110110",
  61814=>"000000000",
  61815=>"111111111",
  61816=>"000000000",
  61817=>"000110111",
  61818=>"000000001",
  61819=>"000000000",
  61820=>"111111111",
  61821=>"100100100",
  61822=>"000011110",
  61823=>"011110000",
  61824=>"110110010",
  61825=>"101110000",
  61826=>"111111111",
  61827=>"000000100",
  61828=>"000011111",
  61829=>"110010111",
  61830=>"000000010",
  61831=>"111100111",
  61832=>"000000000",
  61833=>"110111011",
  61834=>"000000000",
  61835=>"000000111",
  61836=>"111111111",
  61837=>"000110111",
  61838=>"010010110",
  61839=>"000000000",
  61840=>"111111100",
  61841=>"000101111",
  61842=>"111111111",
  61843=>"100111100",
  61844=>"111111111",
  61845=>"000000000",
  61846=>"000011000",
  61847=>"000100000",
  61848=>"111111101",
  61849=>"000000111",
  61850=>"111111111",
  61851=>"000000000",
  61852=>"111111001",
  61853=>"010111011",
  61854=>"110111111",
  61855=>"101000000",
  61856=>"000000000",
  61857=>"111000000",
  61858=>"000000000",
  61859=>"111111111",
  61860=>"000000000",
  61861=>"111111000",
  61862=>"111111100",
  61863=>"110111111",
  61864=>"000000000",
  61865=>"101111111",
  61866=>"011111011",
  61867=>"001000001",
  61868=>"000111000",
  61869=>"000000111",
  61870=>"100000000",
  61871=>"111010000",
  61872=>"111000111",
  61873=>"111111111",
  61874=>"001001111",
  61875=>"111011001",
  61876=>"111111011",
  61877=>"111111111",
  61878=>"111111010",
  61879=>"000100100",
  61880=>"111111000",
  61881=>"111111111",
  61882=>"111111111",
  61883=>"010010011",
  61884=>"001101111",
  61885=>"111111000",
  61886=>"000000000",
  61887=>"000000000",
  61888=>"000000000",
  61889=>"111001001",
  61890=>"000000000",
  61891=>"000000111",
  61892=>"111001000",
  61893=>"110000000",
  61894=>"000000000",
  61895=>"000111111",
  61896=>"111111111",
  61897=>"110110110",
  61898=>"111100000",
  61899=>"111111111",
  61900=>"111101111",
  61901=>"000101001",
  61902=>"000111100",
  61903=>"010000000",
  61904=>"000000111",
  61905=>"000000001",
  61906=>"001001001",
  61907=>"100100000",
  61908=>"000110110",
  61909=>"000000000",
  61910=>"000011010",
  61911=>"000001000",
  61912=>"111111110",
  61913=>"000000001",
  61914=>"000001111",
  61915=>"111111100",
  61916=>"111011111",
  61917=>"001000110",
  61918=>"011000000",
  61919=>"001001011",
  61920=>"111111111",
  61921=>"010000000",
  61922=>"000000000",
  61923=>"001011011",
  61924=>"111111000",
  61925=>"000000000",
  61926=>"000100100",
  61927=>"111111111",
  61928=>"001000011",
  61929=>"111011011",
  61930=>"010110000",
  61931=>"000111111",
  61932=>"000000111",
  61933=>"000000000",
  61934=>"111101001",
  61935=>"010000000",
  61936=>"110000000",
  61937=>"010110111",
  61938=>"001011111",
  61939=>"000000001",
  61940=>"000111111",
  61941=>"001011011",
  61942=>"000110000",
  61943=>"001000010",
  61944=>"000000000",
  61945=>"000000000",
  61946=>"111111010",
  61947=>"000000000",
  61948=>"000000010",
  61949=>"001000000",
  61950=>"111111111",
  61951=>"000000000",
  61952=>"001001001",
  61953=>"111111001",
  61954=>"111111111",
  61955=>"000000000",
  61956=>"111101111",
  61957=>"011011111",
  61958=>"000000000",
  61959=>"111111111",
  61960=>"111100110",
  61961=>"000000111",
  61962=>"111111111",
  61963=>"000001001",
  61964=>"000100100",
  61965=>"000000000",
  61966=>"111111111",
  61967=>"100100000",
  61968=>"111010000",
  61969=>"000000000",
  61970=>"011111000",
  61971=>"000000011",
  61972=>"111111111",
  61973=>"000000011",
  61974=>"110111101",
  61975=>"111111111",
  61976=>"001101101",
  61977=>"111111111",
  61978=>"111011000",
  61979=>"100100100",
  61980=>"110110111",
  61981=>"101101111",
  61982=>"010000000",
  61983=>"000011111",
  61984=>"000000000",
  61985=>"001001110",
  61986=>"111111111",
  61987=>"101111111",
  61988=>"010111111",
  61989=>"000000000",
  61990=>"000000000",
  61991=>"111111111",
  61992=>"111100101",
  61993=>"000000000",
  61994=>"111111111",
  61995=>"100111111",
  61996=>"111111111",
  61997=>"000100111",
  61998=>"011011111",
  61999=>"000000111",
  62000=>"000000000",
  62001=>"000000000",
  62002=>"111111111",
  62003=>"110000110",
  62004=>"000111111",
  62005=>"000100100",
  62006=>"100000000",
  62007=>"110110101",
  62008=>"001011111",
  62009=>"111111111",
  62010=>"000000000",
  62011=>"110111111",
  62012=>"011011111",
  62013=>"111100000",
  62014=>"001011011",
  62015=>"111111111",
  62016=>"000000000",
  62017=>"111111111",
  62018=>"000000110",
  62019=>"111111111",
  62020=>"100100000",
  62021=>"100000110",
  62022=>"000000000",
  62023=>"000000000",
  62024=>"100110111",
  62025=>"000000000",
  62026=>"111011001",
  62027=>"001000000",
  62028=>"000000000",
  62029=>"000000110",
  62030=>"101001000",
  62031=>"001111111",
  62032=>"111111111",
  62033=>"011011011",
  62034=>"011000000",
  62035=>"111111111",
  62036=>"011111111",
  62037=>"000100111",
  62038=>"100100111",
  62039=>"000000000",
  62040=>"111001110",
  62041=>"000000000",
  62042=>"000000000",
  62043=>"000011111",
  62044=>"101111001",
  62045=>"111111111",
  62046=>"100111111",
  62047=>"000100100",
  62048=>"000100011",
  62049=>"011000100",
  62050=>"000000000",
  62051=>"111011000",
  62052=>"001001011",
  62053=>"001000110",
  62054=>"000000000",
  62055=>"000000010",
  62056=>"110100000",
  62057=>"110111000",
  62058=>"110010000",
  62059=>"111111010",
  62060=>"001100111",
  62061=>"000000010",
  62062=>"111111110",
  62063=>"001000000",
  62064=>"010010010",
  62065=>"000110110",
  62066=>"000000000",
  62067=>"000000011",
  62068=>"000001001",
  62069=>"000110000",
  62070=>"111111111",
  62071=>"111111111",
  62072=>"000000000",
  62073=>"100000100",
  62074=>"000001001",
  62075=>"000000000",
  62076=>"110000110",
  62077=>"000000000",
  62078=>"110110110",
  62079=>"000000000",
  62080=>"111111111",
  62081=>"101100111",
  62082=>"111111111",
  62083=>"011000011",
  62084=>"000100111",
  62085=>"000000000",
  62086=>"010000000",
  62087=>"111111001",
  62088=>"001000011",
  62089=>"000000011",
  62090=>"111000000",
  62091=>"111010011",
  62092=>"110110111",
  62093=>"000100101",
  62094=>"111111000",
  62095=>"111110111",
  62096=>"000000000",
  62097=>"011011001",
  62098=>"001010100",
  62099=>"111111111",
  62100=>"101111010",
  62101=>"110111111",
  62102=>"100100100",
  62103=>"000100111",
  62104=>"100000000",
  62105=>"110110100",
  62106=>"111111111",
  62107=>"000000110",
  62108=>"110010000",
  62109=>"100000000",
  62110=>"000000000",
  62111=>"110111111",
  62112=>"101111111",
  62113=>"110110101",
  62114=>"000000000",
  62115=>"111101110",
  62116=>"000000000",
  62117=>"000100111",
  62118=>"111000000",
  62119=>"001000001",
  62120=>"111111110",
  62121=>"000111111",
  62122=>"111111011",
  62123=>"111111111",
  62124=>"111010111",
  62125=>"110110111",
  62126=>"000000000",
  62127=>"000000000",
  62128=>"000000000",
  62129=>"011000111",
  62130=>"110111000",
  62131=>"000000110",
  62132=>"000000001",
  62133=>"110110110",
  62134=>"000000000",
  62135=>"011011000",
  62136=>"111000000",
  62137=>"000000011",
  62138=>"100100100",
  62139=>"110110100",
  62140=>"111111111",
  62141=>"000000000",
  62142=>"000000110",
  62143=>"111111111",
  62144=>"111111101",
  62145=>"011001000",
  62146=>"000000001",
  62147=>"111010000",
  62148=>"000000000",
  62149=>"001100000",
  62150=>"000000000",
  62151=>"000001000",
  62152=>"000111110",
  62153=>"001000100",
  62154=>"100100000",
  62155=>"000000000",
  62156=>"100100000",
  62157=>"111111111",
  62158=>"111111111",
  62159=>"000100111",
  62160=>"000000001",
  62161=>"100110000",
  62162=>"000000000",
  62163=>"001001101",
  62164=>"010110111",
  62165=>"111111011",
  62166=>"111111111",
  62167=>"110010000",
  62168=>"111000000",
  62169=>"000000000",
  62170=>"101001101",
  62171=>"000000111",
  62172=>"000000000",
  62173=>"110111111",
  62174=>"000000000",
  62175=>"111111111",
  62176=>"001000000",
  62177=>"001111111",
  62178=>"111111111",
  62179=>"110111110",
  62180=>"111000111",
  62181=>"111110100",
  62182=>"000000000",
  62183=>"000011111",
  62184=>"100111111",
  62185=>"010000000",
  62186=>"000000000",
  62187=>"111111111",
  62188=>"111111010",
  62189=>"111111111",
  62190=>"001000101",
  62191=>"000111000",
  62192=>"000000011",
  62193=>"000100100",
  62194=>"111111111",
  62195=>"110111000",
  62196=>"000100100",
  62197=>"010000010",
  62198=>"111111111",
  62199=>"000100000",
  62200=>"000000001",
  62201=>"111111011",
  62202=>"110111111",
  62203=>"011000000",
  62204=>"100110111",
  62205=>"001001000",
  62206=>"101000000",
  62207=>"000000000",
  62208=>"001000110",
  62209=>"011111111",
  62210=>"111100000",
  62211=>"000000111",
  62212=>"011111111",
  62213=>"000000000",
  62214=>"000000000",
  62215=>"000110110",
  62216=>"001001000",
  62217=>"101001111",
  62218=>"111111111",
  62219=>"111110111",
  62220=>"011001000",
  62221=>"000110110",
  62222=>"100111111",
  62223=>"000000000",
  62224=>"111111001",
  62225=>"000000000",
  62226=>"111111111",
  62227=>"111111111",
  62228=>"000000000",
  62229=>"111111111",
  62230=>"011011011",
  62231=>"000000111",
  62232=>"110110100",
  62233=>"000000000",
  62234=>"000000000",
  62235=>"100000000",
  62236=>"001001111",
  62237=>"111110000",
  62238=>"000000000",
  62239=>"111111111",
  62240=>"000000000",
  62241=>"111111111",
  62242=>"111111111",
  62243=>"000000000",
  62244=>"011011000",
  62245=>"001000000",
  62246=>"010110110",
  62247=>"000000000",
  62248=>"000000100",
  62249=>"001111111",
  62250=>"000100111",
  62251=>"000000000",
  62252=>"000000000",
  62253=>"111000000",
  62254=>"111000000",
  62255=>"010010000",
  62256=>"001000000",
  62257=>"000000000",
  62258=>"111111111",
  62259=>"000000000",
  62260=>"111111111",
  62261=>"111111110",
  62262=>"111111111",
  62263=>"100000000",
  62264=>"000000000",
  62265=>"000101111",
  62266=>"111111111",
  62267=>"000110111",
  62268=>"110111111",
  62269=>"100100000",
  62270=>"101100111",
  62271=>"111111000",
  62272=>"000000000",
  62273=>"000000000",
  62274=>"000100000",
  62275=>"000000000",
  62276=>"000000000",
  62277=>"111111110",
  62278=>"111111011",
  62279=>"111111000",
  62280=>"000000000",
  62281=>"111100000",
  62282=>"111111111",
  62283=>"000000000",
  62284=>"000000000",
  62285=>"101001000",
  62286=>"010000000",
  62287=>"111101101",
  62288=>"000000010",
  62289=>"111111000",
  62290=>"000000000",
  62291=>"111111000",
  62292=>"000101000",
  62293=>"011011011",
  62294=>"111111000",
  62295=>"001000000",
  62296=>"110111111",
  62297=>"001101101",
  62298=>"101111111",
  62299=>"101011000",
  62300=>"000000110",
  62301=>"111111111",
  62302=>"000000000",
  62303=>"110111111",
  62304=>"000000000",
  62305=>"000000000",
  62306=>"000000001",
  62307=>"000000111",
  62308=>"100100000",
  62309=>"111111111",
  62310=>"111111101",
  62311=>"111111111",
  62312=>"000000001",
  62313=>"010010110",
  62314=>"111000000",
  62315=>"111001001",
  62316=>"011111111",
  62317=>"110110111",
  62318=>"000000100",
  62319=>"000000000",
  62320=>"000000000",
  62321=>"111111111",
  62322=>"111111000",
  62323=>"001011011",
  62324=>"111000000",
  62325=>"111000000",
  62326=>"111010000",
  62327=>"111011000",
  62328=>"011000000",
  62329=>"000000000",
  62330=>"111111011",
  62331=>"000100011",
  62332=>"000111111",
  62333=>"111111000",
  62334=>"111110000",
  62335=>"111000101",
  62336=>"111100100",
  62337=>"000000000",
  62338=>"000001011",
  62339=>"111000000",
  62340=>"000101000",
  62341=>"000000000",
  62342=>"000000000",
  62343=>"111111111",
  62344=>"111110010",
  62345=>"111111111",
  62346=>"111111101",
  62347=>"000000000",
  62348=>"111101111",
  62349=>"110110111",
  62350=>"000000111",
  62351=>"000000000",
  62352=>"000000000",
  62353=>"000001110",
  62354=>"101101000",
  62355=>"111111111",
  62356=>"100111100",
  62357=>"011011010",
  62358=>"101101011",
  62359=>"000001101",
  62360=>"000000001",
  62361=>"001001111",
  62362=>"000000000",
  62363=>"111111111",
  62364=>"111111011",
  62365=>"000000000",
  62366=>"000000000",
  62367=>"000000000",
  62368=>"000000010",
  62369=>"000000000",
  62370=>"111111111",
  62371=>"100101000",
  62372=>"100101111",
  62373=>"111111010",
  62374=>"111111111",
  62375=>"111111111",
  62376=>"110111111",
  62377=>"011111111",
  62378=>"110100000",
  62379=>"000000000",
  62380=>"000000000",
  62381=>"110111110",
  62382=>"000000000",
  62383=>"110100110",
  62384=>"000000000",
  62385=>"000101000",
  62386=>"111111100",
  62387=>"000010000",
  62388=>"111111111",
  62389=>"011011011",
  62390=>"100101100",
  62391=>"000001000",
  62392=>"000110111",
  62393=>"111111111",
  62394=>"000000000",
  62395=>"111110111",
  62396=>"000000010",
  62397=>"000000100",
  62398=>"000000111",
  62399=>"000010011",
  62400=>"110100000",
  62401=>"011000000",
  62402=>"101000000",
  62403=>"111110111",
  62404=>"111111100",
  62405=>"110110111",
  62406=>"000000000",
  62407=>"000000000",
  62408=>"011001000",
  62409=>"000000000",
  62410=>"000000000",
  62411=>"000110111",
  62412=>"111001000",
  62413=>"100111000",
  62414=>"000000000",
  62415=>"110111111",
  62416=>"000000000",
  62417=>"010000100",
  62418=>"111111111",
  62419=>"111101111",
  62420=>"000000011",
  62421=>"111111111",
  62422=>"001000111",
  62423=>"001010010",
  62424=>"011001011",
  62425=>"000100000",
  62426=>"111111111",
  62427=>"111111101",
  62428=>"010001001",
  62429=>"010110110",
  62430=>"011000000",
  62431=>"111111111",
  62432=>"111111010",
  62433=>"011011000",
  62434=>"000000111",
  62435=>"000100101",
  62436=>"000000000",
  62437=>"111111111",
  62438=>"100111011",
  62439=>"101101111",
  62440=>"011111011",
  62441=>"000110100",
  62442=>"000000000",
  62443=>"000110110",
  62444=>"000000000",
  62445=>"000000111",
  62446=>"110111111",
  62447=>"000100100",
  62448=>"111111111",
  62449=>"000111111",
  62450=>"111100111",
  62451=>"000000000",
  62452=>"000000000",
  62453=>"000110110",
  62454=>"011011001",
  62455=>"001000011",
  62456=>"000000000",
  62457=>"111000110",
  62458=>"010011011",
  62459=>"111111111",
  62460=>"111111011",
  62461=>"100110111",
  62462=>"000000000",
  62463=>"000100111",
  62464=>"111111111",
  62465=>"000000000",
  62466=>"111111111",
  62467=>"000000001",
  62468=>"100100111",
  62469=>"111111011",
  62470=>"111000000",
  62471=>"111111100",
  62472=>"000000000",
  62473=>"000100110",
  62474=>"000000001",
  62475=>"000000000",
  62476=>"000000000",
  62477=>"011001000",
  62478=>"011010000",
  62479=>"011111111",
  62480=>"111111000",
  62481=>"000101111",
  62482=>"111000000",
  62483=>"111111111",
  62484=>"000000000",
  62485=>"001000100",
  62486=>"001101101",
  62487=>"000000000",
  62488=>"100110110",
  62489=>"101000001",
  62490=>"111111111",
  62491=>"100110000",
  62492=>"001100111",
  62493=>"111110000",
  62494=>"000000000",
  62495=>"001001111",
  62496=>"001111101",
  62497=>"000000000",
  62498=>"011111000",
  62499=>"010000011",
  62500=>"111111111",
  62501=>"111111111",
  62502=>"000001011",
  62503=>"101101111",
  62504=>"011111111",
  62505=>"000000000",
  62506=>"000000111",
  62507=>"111111111",
  62508=>"000000000",
  62509=>"000011011",
  62510=>"000000000",
  62511=>"111111111",
  62512=>"000000000",
  62513=>"101000000",
  62514=>"111111111",
  62515=>"101110111",
  62516=>"111111111",
  62517=>"110110101",
  62518=>"100111111",
  62519=>"100000000",
  62520=>"011011011",
  62521=>"111111111",
  62522=>"111111000",
  62523=>"110011001",
  62524=>"111001001",
  62525=>"111111000",
  62526=>"000000000",
  62527=>"111111010",
  62528=>"001000000",
  62529=>"010010011",
  62530=>"101111111",
  62531=>"111101100",
  62532=>"111100000",
  62533=>"101000001",
  62534=>"111111011",
  62535=>"111111111",
  62536=>"000000000",
  62537=>"000000000",
  62538=>"101111111",
  62539=>"111101000",
  62540=>"011111101",
  62541=>"001000101",
  62542=>"111111011",
  62543=>"000111111",
  62544=>"011111010",
  62545=>"111111111",
  62546=>"000000000",
  62547=>"010000011",
  62548=>"111101111",
  62549=>"000000111",
  62550=>"101100101",
  62551=>"100100000",
  62552=>"000000011",
  62553=>"111111111",
  62554=>"001100000",
  62555=>"000110110",
  62556=>"000100000",
  62557=>"111111111",
  62558=>"001001111",
  62559=>"111111111",
  62560=>"000100000",
  62561=>"000000000",
  62562=>"000000000",
  62563=>"000000000",
  62564=>"000000000",
  62565=>"100101111",
  62566=>"011110111",
  62567=>"110010000",
  62568=>"000000000",
  62569=>"101111111",
  62570=>"000000000",
  62571=>"000000000",
  62572=>"111111101",
  62573=>"111111111",
  62574=>"000000111",
  62575=>"010000000",
  62576=>"111011010",
  62577=>"000000111",
  62578=>"011011000",
  62579=>"111111000",
  62580=>"100000000",
  62581=>"110100000",
  62582=>"000111111",
  62583=>"001000000",
  62584=>"000100100",
  62585=>"000001111",
  62586=>"111111111",
  62587=>"111111000",
  62588=>"110110110",
  62589=>"000000000",
  62590=>"111111111",
  62591=>"111101011",
  62592=>"111111110",
  62593=>"000000000",
  62594=>"111010110",
  62595=>"011011111",
  62596=>"101111011",
  62597=>"000000000",
  62598=>"011111000",
  62599=>"001111111",
  62600=>"000000000",
  62601=>"000000000",
  62602=>"000000000",
  62603=>"011100101",
  62604=>"000000000",
  62605=>"000000111",
  62606=>"111010111",
  62607=>"001000000",
  62608=>"111001000",
  62609=>"100100000",
  62610=>"001001111",
  62611=>"000001000",
  62612=>"100111101",
  62613=>"111110011",
  62614=>"111001111",
  62615=>"110110110",
  62616=>"000000000",
  62617=>"111111111",
  62618=>"000000011",
  62619=>"000000000",
  62620=>"100100000",
  62621=>"000000000",
  62622=>"000100100",
  62623=>"000000000",
  62624=>"101011111",
  62625=>"011001000",
  62626=>"111000000",
  62627=>"101111111",
  62628=>"000001101",
  62629=>"101000001",
  62630=>"111111011",
  62631=>"011011111",
  62632=>"000000000",
  62633=>"111111111",
  62634=>"000010000",
  62635=>"111111111",
  62636=>"001101101",
  62637=>"000000110",
  62638=>"101011011",
  62639=>"111111111",
  62640=>"111111011",
  62641=>"111011011",
  62642=>"000000000",
  62643=>"011111000",
  62644=>"000000000",
  62645=>"111110000",
  62646=>"001001000",
  62647=>"000000000",
  62648=>"000000000",
  62649=>"111110111",
  62650=>"101000001",
  62651=>"000000000",
  62652=>"111111111",
  62653=>"111111111",
  62654=>"111110111",
  62655=>"000000000",
  62656=>"111111111",
  62657=>"000000000",
  62658=>"001111101",
  62659=>"100100101",
  62660=>"000000000",
  62661=>"000010000",
  62662=>"000101101",
  62663=>"000000010",
  62664=>"111111000",
  62665=>"100000111",
  62666=>"000000000",
  62667=>"111111111",
  62668=>"101001011",
  62669=>"011000001",
  62670=>"000111111",
  62671=>"111001111",
  62672=>"011111000",
  62673=>"111111000",
  62674=>"011011000",
  62675=>"000000010",
  62676=>"000000000",
  62677=>"111111111",
  62678=>"010011011",
  62679=>"000011000",
  62680=>"000010011",
  62681=>"001000101",
  62682=>"000000001",
  62683=>"011001001",
  62684=>"000111111",
  62685=>"101000111",
  62686=>"111111111",
  62687=>"111111101",
  62688=>"000000000",
  62689=>"000010010",
  62690=>"111111001",
  62691=>"100111111",
  62692=>"111101111",
  62693=>"001110110",
  62694=>"111111111",
  62695=>"001111111",
  62696=>"000000111",
  62697=>"001101000",
  62698=>"000000000",
  62699=>"111001101",
  62700=>"111111100",
  62701=>"000010010",
  62702=>"000001111",
  62703=>"000000000",
  62704=>"000000000",
  62705=>"000000001",
  62706=>"000000000",
  62707=>"011001000",
  62708=>"000000000",
  62709=>"110111111",
  62710=>"100101011",
  62711=>"000000000",
  62712=>"111111100",
  62713=>"011111111",
  62714=>"111111111",
  62715=>"010111111",
  62716=>"000100100",
  62717=>"100100100",
  62718=>"101000000",
  62719=>"111111111",
  62720=>"000000000",
  62721=>"011011011",
  62722=>"000000000",
  62723=>"110111111",
  62724=>"000000000",
  62725=>"000000000",
  62726=>"110000100",
  62727=>"110111000",
  62728=>"001000010",
  62729=>"111111110",
  62730=>"111010110",
  62731=>"000000001",
  62732=>"000100100",
  62733=>"011000000",
  62734=>"101101111",
  62735=>"000100111",
  62736=>"000001101",
  62737=>"111111000",
  62738=>"111011001",
  62739=>"111111111",
  62740=>"000000000",
  62741=>"111111110",
  62742=>"111111110",
  62743=>"111111111",
  62744=>"111101011",
  62745=>"110101001",
  62746=>"000000001",
  62747=>"111111111",
  62748=>"000000000",
  62749=>"011111111",
  62750=>"000011000",
  62751=>"001111001",
  62752=>"110111011",
  62753=>"001111111",
  62754=>"111110111",
  62755=>"111111011",
  62756=>"011000000",
  62757=>"111110000",
  62758=>"000000000",
  62759=>"111111111",
  62760=>"000000000",
  62761=>"011111111",
  62762=>"001011111",
  62763=>"100101111",
  62764=>"111000000",
  62765=>"000000000",
  62766=>"000000000",
  62767=>"000000000",
  62768=>"100000000",
  62769=>"000000000",
  62770=>"000011000",
  62771=>"000111111",
  62772=>"010110110",
  62773=>"111001101",
  62774=>"000000000",
  62775=>"110110110",
  62776=>"100100101",
  62777=>"100000000",
  62778=>"111101111",
  62779=>"000000111",
  62780=>"001001011",
  62781=>"001001011",
  62782=>"000000000",
  62783=>"100000111",
  62784=>"111011000",
  62785=>"000000000",
  62786=>"000110110",
  62787=>"000000000",
  62788=>"000000000",
  62789=>"101100100",
  62790=>"100000111",
  62791=>"111000000",
  62792=>"111111111",
  62793=>"000000000",
  62794=>"000000000",
  62795=>"111111100",
  62796=>"100000000",
  62797=>"000000000",
  62798=>"111111111",
  62799=>"000100100",
  62800=>"011111111",
  62801=>"000001001",
  62802=>"000000000",
  62803=>"111111111",
  62804=>"111101101",
  62805=>"001001001",
  62806=>"000111111",
  62807=>"111111111",
  62808=>"111111111",
  62809=>"010111111",
  62810=>"111110000",
  62811=>"111111111",
  62812=>"000000000",
  62813=>"111111111",
  62814=>"000110000",
  62815=>"000000011",
  62816=>"000000000",
  62817=>"011111111",
  62818=>"000000000",
  62819=>"111111111",
  62820=>"001001001",
  62821=>"000111111",
  62822=>"000000100",
  62823=>"111111111",
  62824=>"100111011",
  62825=>"111111011",
  62826=>"100000000",
  62827=>"001101111",
  62828=>"011111110",
  62829=>"101111100",
  62830=>"000000000",
  62831=>"011011000",
  62832=>"010000000",
  62833=>"111111111",
  62834=>"000100111",
  62835=>"000101100",
  62836=>"111111001",
  62837=>"000000000",
  62838=>"000000011",
  62839=>"010010011",
  62840=>"111111111",
  62841=>"000000000",
  62842=>"001000000",
  62843=>"000001000",
  62844=>"111010010",
  62845=>"111101111",
  62846=>"111111101",
  62847=>"111111100",
  62848=>"000000000",
  62849=>"111011111",
  62850=>"000000000",
  62851=>"000000000",
  62852=>"101000001",
  62853=>"000010010",
  62854=>"110111111",
  62855=>"111111111",
  62856=>"110110000",
  62857=>"000000100",
  62858=>"010010111",
  62859=>"000000110",
  62860=>"111111111",
  62861=>"110111110",
  62862=>"111111111",
  62863=>"000000000",
  62864=>"000000000",
  62865=>"000000000",
  62866=>"111011111",
  62867=>"000000100",
  62868=>"111111111",
  62869=>"000000000",
  62870=>"000000000",
  62871=>"100001111",
  62872=>"001000000",
  62873=>"111111111",
  62874=>"111111111",
  62875=>"000100111",
  62876=>"000000000",
  62877=>"000000000",
  62878=>"011001111",
  62879=>"111111111",
  62880=>"111101111",
  62881=>"110111111",
  62882=>"111111111",
  62883=>"000000011",
  62884=>"111011010",
  62885=>"100010000",
  62886=>"000000000",
  62887=>"000001111",
  62888=>"000011010",
  62889=>"100110100",
  62890=>"011111110",
  62891=>"001011000",
  62892=>"000000000",
  62893=>"000000000",
  62894=>"101001011",
  62895=>"101001000",
  62896=>"011110100",
  62897=>"111111111",
  62898=>"000000000",
  62899=>"000000000",
  62900=>"000000000",
  62901=>"111000000",
  62902=>"111111001",
  62903=>"000010000",
  62904=>"001000111",
  62905=>"000000100",
  62906=>"000111101",
  62907=>"111000011",
  62908=>"101111111",
  62909=>"000110100",
  62910=>"000101111",
  62911=>"010110110",
  62912=>"000100100",
  62913=>"000000000",
  62914=>"101111110",
  62915=>"111111011",
  62916=>"000000100",
  62917=>"100100100",
  62918=>"101001110",
  62919=>"000100100",
  62920=>"001000000",
  62921=>"111111111",
  62922=>"111101111",
  62923=>"111111000",
  62924=>"101101000",
  62925=>"111000000",
  62926=>"000000000",
  62927=>"001000000",
  62928=>"000011001",
  62929=>"000000100",
  62930=>"000001111",
  62931=>"111111111",
  62932=>"111111001",
  62933=>"000000001",
  62934=>"011011000",
  62935=>"110011000",
  62936=>"100100001",
  62937=>"111111111",
  62938=>"000000100",
  62939=>"111111111",
  62940=>"000000110",
  62941=>"000000000",
  62942=>"000000000",
  62943=>"001001011",
  62944=>"110100100",
  62945=>"111001000",
  62946=>"000000100",
  62947=>"000000110",
  62948=>"111111111",
  62949=>"100111111",
  62950=>"000001000",
  62951=>"010100111",
  62952=>"000000111",
  62953=>"000100000",
  62954=>"000001001",
  62955=>"000010111",
  62956=>"000111000",
  62957=>"111101101",
  62958=>"000111111",
  62959=>"110111111",
  62960=>"000000000",
  62961=>"000000000",
  62962=>"011011111",
  62963=>"000100100",
  62964=>"111110110",
  62965=>"111000000",
  62966=>"000000111",
  62967=>"011011111",
  62968=>"000010000",
  62969=>"100111111",
  62970=>"000000000",
  62971=>"111011110",
  62972=>"110100000",
  62973=>"011011111",
  62974=>"011001111",
  62975=>"111001101",
  62976=>"011011000",
  62977=>"111010000",
  62978=>"000000000",
  62979=>"100000101",
  62980=>"011001111",
  62981=>"111010010",
  62982=>"111111111",
  62983=>"000000000",
  62984=>"001000001",
  62985=>"111111100",
  62986=>"001000000",
  62987=>"010111000",
  62988=>"011001001",
  62989=>"000000000",
  62990=>"001001111",
  62991=>"111111111",
  62992=>"111110100",
  62993=>"111111111",
  62994=>"001111111",
  62995=>"100000100",
  62996=>"000010000",
  62997=>"010010000",
  62998=>"000000101",
  62999=>"011111110",
  63000=>"111011000",
  63001=>"111111011",
  63002=>"000000011",
  63003=>"011001000",
  63004=>"111000000",
  63005=>"000000000",
  63006=>"111111111",
  63007=>"000000100",
  63008=>"111110111",
  63009=>"111111111",
  63010=>"001001001",
  63011=>"000110100",
  63012=>"011111111",
  63013=>"011000001",
  63014=>"000000000",
  63015=>"000100100",
  63016=>"111101001",
  63017=>"111010000",
  63018=>"111111111",
  63019=>"000000000",
  63020=>"011111101",
  63021=>"011111111",
  63022=>"000000000",
  63023=>"111110010",
  63024=>"110000011",
  63025=>"111111111",
  63026=>"101110111",
  63027=>"001001001",
  63028=>"000000000",
  63029=>"111001111",
  63030=>"001001000",
  63031=>"000000000",
  63032=>"111111111",
  63033=>"111100111",
  63034=>"000000001",
  63035=>"110000000",
  63036=>"000000000",
  63037=>"001001101",
  63038=>"000000011",
  63039=>"000000000",
  63040=>"111111111",
  63041=>"000100001",
  63042=>"110111001",
  63043=>"000000111",
  63044=>"001001011",
  63045=>"000000000",
  63046=>"010111010",
  63047=>"111111111",
  63048=>"100100100",
  63049=>"111101111",
  63050=>"000000000",
  63051=>"110111111",
  63052=>"000111111",
  63053=>"000010000",
  63054=>"111000000",
  63055=>"000001000",
  63056=>"010011111",
  63057=>"110010111",
  63058=>"111000110",
  63059=>"111110110",
  63060=>"000000000",
  63061=>"110110110",
  63062=>"111000000",
  63063=>"000000100",
  63064=>"111111111",
  63065=>"000000000",
  63066=>"101101001",
  63067=>"001111101",
  63068=>"111111111",
  63069=>"000010000",
  63070=>"111001000",
  63071=>"000111010",
  63072=>"000001111",
  63073=>"110000101",
  63074=>"011010000",
  63075=>"111000101",
  63076=>"000000111",
  63077=>"111111001",
  63078=>"111111111",
  63079=>"000000000",
  63080=>"000000010",
  63081=>"111011000",
  63082=>"001111111",
  63083=>"111110110",
  63084=>"000001001",
  63085=>"111010000",
  63086=>"000000000",
  63087=>"111011111",
  63088=>"001001011",
  63089=>"111111111",
  63090=>"100100100",
  63091=>"110000011",
  63092=>"111000000",
  63093=>"000110110",
  63094=>"111111111",
  63095=>"000110111",
  63096=>"000000110",
  63097=>"111111000",
  63098=>"000110111",
  63099=>"000000000",
  63100=>"000011011",
  63101=>"000000000",
  63102=>"000110110",
  63103=>"010111111",
  63104=>"000000000",
  63105=>"000000011",
  63106=>"000111111",
  63107=>"100111111",
  63108=>"000000000",
  63109=>"000000000",
  63110=>"001011111",
  63111=>"111111111",
  63112=>"100110111",
  63113=>"111111001",
  63114=>"111100100",
  63115=>"001000000",
  63116=>"111111000",
  63117=>"111111111",
  63118=>"000011000",
  63119=>"111111111",
  63120=>"110111111",
  63121=>"011000000",
  63122=>"001101010",
  63123=>"111111111",
  63124=>"001111110",
  63125=>"111111100",
  63126=>"000000001",
  63127=>"111111011",
  63128=>"111111001",
  63129=>"111111000",
  63130=>"111111111",
  63131=>"111001111",
  63132=>"111000011",
  63133=>"010010000",
  63134=>"111111000",
  63135=>"010111110",
  63136=>"000000000",
  63137=>"110000000",
  63138=>"000000000",
  63139=>"101000101",
  63140=>"111010110",
  63141=>"000110000",
  63142=>"000000000",
  63143=>"110110110",
  63144=>"111111111",
  63145=>"001001001",
  63146=>"000000000",
  63147=>"000000111",
  63148=>"111111111",
  63149=>"000001000",
  63150=>"111110110",
  63151=>"000000110",
  63152=>"000000100",
  63153=>"010000100",
  63154=>"000000111",
  63155=>"111000111",
  63156=>"111010010",
  63157=>"111011111",
  63158=>"111000000",
  63159=>"111111111",
  63160=>"011111111",
  63161=>"000111101",
  63162=>"111110111",
  63163=>"000000111",
  63164=>"111010010",
  63165=>"111111111",
  63166=>"000000000",
  63167=>"010000000",
  63168=>"000101111",
  63169=>"011111111",
  63170=>"110110110",
  63171=>"000010000",
  63172=>"111111111",
  63173=>"111111111",
  63174=>"111000000",
  63175=>"000000000",
  63176=>"000000011",
  63177=>"111111000",
  63178=>"111111100",
  63179=>"111111111",
  63180=>"000110111",
  63181=>"000110010",
  63182=>"011000000",
  63183=>"111111111",
  63184=>"111000000",
  63185=>"111000000",
  63186=>"111000111",
  63187=>"001111111",
  63188=>"111111111",
  63189=>"100000111",
  63190=>"011000000",
  63191=>"000110000",
  63192=>"111111111",
  63193=>"110100000",
  63194=>"111111111",
  63195=>"000001011",
  63196=>"000000000",
  63197=>"000111000",
  63198=>"001000010",
  63199=>"111010000",
  63200=>"001111000",
  63201=>"000000000",
  63202=>"000000000",
  63203=>"111111111",
  63204=>"011000000",
  63205=>"000010000",
  63206=>"000000101",
  63207=>"000000000",
  63208=>"111000100",
  63209=>"111110111",
  63210=>"000001111",
  63211=>"000000000",
  63212=>"111111111",
  63213=>"000000110",
  63214=>"111000010",
  63215=>"000000000",
  63216=>"111111111",
  63217=>"111111111",
  63218=>"111111111",
  63219=>"010111101",
  63220=>"111111111",
  63221=>"011000001",
  63222=>"001001000",
  63223=>"000000000",
  63224=>"111111111",
  63225=>"111011011",
  63226=>"010010000",
  63227=>"000000000",
  63228=>"000110100",
  63229=>"111111011",
  63230=>"111110110",
  63231=>"001111111",
  63232=>"101000111",
  63233=>"111111111",
  63234=>"101000000",
  63235=>"001001111",
  63236=>"000000111",
  63237=>"000000101",
  63238=>"000000000",
  63239=>"011111111",
  63240=>"000010010",
  63241=>"000000000",
  63242=>"000001000",
  63243=>"011011111",
  63244=>"000000101",
  63245=>"000000000",
  63246=>"111111111",
  63247=>"000100100",
  63248=>"011011111",
  63249=>"000000000",
  63250=>"110001001",
  63251=>"101111111",
  63252=>"000000101",
  63253=>"000111111",
  63254=>"000000100",
  63255=>"111111111",
  63256=>"111111001",
  63257=>"111000111",
  63258=>"110111111",
  63259=>"111111111",
  63260=>"001011001",
  63261=>"101101101",
  63262=>"011010111",
  63263=>"000000100",
  63264=>"011000000",
  63265=>"000000000",
  63266=>"111111110",
  63267=>"000000110",
  63268=>"111111111",
  63269=>"111111111",
  63270=>"000000111",
  63271=>"110110111",
  63272=>"000000000",
  63273=>"100111111",
  63274=>"000000000",
  63275=>"000111011",
  63276=>"000100100",
  63277=>"000100100",
  63278=>"000111111",
  63279=>"110000000",
  63280=>"111111111",
  63281=>"000000010",
  63282=>"011001000",
  63283=>"110000000",
  63284=>"000000011",
  63285=>"011111010",
  63286=>"000000010",
  63287=>"011011011",
  63288=>"000000111",
  63289=>"001111111",
  63290=>"111011000",
  63291=>"111101101",
  63292=>"111111111",
  63293=>"110110000",
  63294=>"111111111",
  63295=>"000000000",
  63296=>"111110100",
  63297=>"111111111",
  63298=>"011010111",
  63299=>"000010000",
  63300=>"000000100",
  63301=>"000000010",
  63302=>"000011111",
  63303=>"100100101",
  63304=>"111111111",
  63305=>"010000000",
  63306=>"111111111",
  63307=>"011111111",
  63308=>"100000000",
  63309=>"000010011",
  63310=>"110100100",
  63311=>"000001001",
  63312=>"001001011",
  63313=>"000101000",
  63314=>"111111111",
  63315=>"111110111",
  63316=>"111100110",
  63317=>"000110000",
  63318=>"111110111",
  63319=>"111111010",
  63320=>"111111111",
  63321=>"000000001",
  63322=>"001001111",
  63323=>"111010110",
  63324=>"000000000",
  63325=>"000000000",
  63326=>"111111111",
  63327=>"110000000",
  63328=>"111111111",
  63329=>"101000001",
  63330=>"111111101",
  63331=>"001011001",
  63332=>"100010001",
  63333=>"000011001",
  63334=>"000001001",
  63335=>"011011000",
  63336=>"100111101",
  63337=>"000000000",
  63338=>"110111111",
  63339=>"111111111",
  63340=>"011111011",
  63341=>"110100011",
  63342=>"000000000",
  63343=>"111111111",
  63344=>"111111111",
  63345=>"111111111",
  63346=>"000000000",
  63347=>"110100100",
  63348=>"110111111",
  63349=>"111111111",
  63350=>"111100000",
  63351=>"000000110",
  63352=>"000111111",
  63353=>"000100101",
  63354=>"000000101",
  63355=>"110011111",
  63356=>"010000010",
  63357=>"000000011",
  63358=>"010111111",
  63359=>"111111000",
  63360=>"011111111",
  63361=>"111111000",
  63362=>"110110100",
  63363=>"000000000",
  63364=>"111111011",
  63365=>"000000010",
  63366=>"000000100",
  63367=>"110111011",
  63368=>"111111111",
  63369=>"100100100",
  63370=>"111011000",
  63371=>"010000000",
  63372=>"101011001",
  63373=>"000000000",
  63374=>"000100111",
  63375=>"111111111",
  63376=>"100000000",
  63377=>"000000000",
  63378=>"000000001",
  63379=>"111111111",
  63380=>"000000011",
  63381=>"111111111",
  63382=>"111111111",
  63383=>"000011111",
  63384=>"100000000",
  63385=>"111101011",
  63386=>"000000010",
  63387=>"001111111",
  63388=>"000111111",
  63389=>"111111111",
  63390=>"000000111",
  63391=>"111111111",
  63392=>"011111000",
  63393=>"110000100",
  63394=>"000111111",
  63395=>"111110010",
  63396=>"000000010",
  63397=>"001000000",
  63398=>"000000111",
  63399=>"001111000",
  63400=>"111111111",
  63401=>"000000000",
  63402=>"111101101",
  63403=>"111000000",
  63404=>"110111000",
  63405=>"000010010",
  63406=>"100000000",
  63407=>"001100111",
  63408=>"000000000",
  63409=>"000100000",
  63410=>"000000111",
  63411=>"000000000",
  63412=>"000001001",
  63413=>"010010100",
  63414=>"011000111",
  63415=>"100100000",
  63416=>"001011000",
  63417=>"111000100",
  63418=>"100000011",
  63419=>"000000001",
  63420=>"111111010",
  63421=>"000010000",
  63422=>"111000000",
  63423=>"100100100",
  63424=>"000100100",
  63425=>"000000000",
  63426=>"000000000",
  63427=>"000000000",
  63428=>"101100110",
  63429=>"001001111",
  63430=>"100100111",
  63431=>"111111100",
  63432=>"111111110",
  63433=>"011011110",
  63434=>"111111111",
  63435=>"010011111",
  63436=>"100100111",
  63437=>"000000000",
  63438=>"111001000",
  63439=>"111100111",
  63440=>"101001101",
  63441=>"001110100",
  63442=>"111011001",
  63443=>"000000011",
  63444=>"110000000",
  63445=>"111110001",
  63446=>"110110110",
  63447=>"100000100",
  63448=>"000001101",
  63449=>"111110100",
  63450=>"000000000",
  63451=>"111000110",
  63452=>"111111111",
  63453=>"111111111",
  63454=>"111000111",
  63455=>"111110110",
  63456=>"000111111",
  63457=>"001101110",
  63458=>"111000001",
  63459=>"000000000",
  63460=>"101000000",
  63461=>"000010011",
  63462=>"110010001",
  63463=>"010000000",
  63464=>"001001001",
  63465=>"100001001",
  63466=>"000000000",
  63467=>"101110100",
  63468=>"111000101",
  63469=>"000000000",
  63470=>"001000000",
  63471=>"000000000",
  63472=>"111111111",
  63473=>"111111111",
  63474=>"111111100",
  63475=>"111111111",
  63476=>"110100111",
  63477=>"001000001",
  63478=>"000000001",
  63479=>"011011010",
  63480=>"000000000",
  63481=>"011001001",
  63482=>"111111110",
  63483=>"000000000",
  63484=>"111111111",
  63485=>"000000000",
  63486=>"000111000",
  63487=>"000000001",
  63488=>"111111111",
  63489=>"001011000",
  63490=>"111111011",
  63491=>"000000000",
  63492=>"111010100",
  63493=>"000000000",
  63494=>"000000000",
  63495=>"111111111",
  63496=>"111111111",
  63497=>"000000111",
  63498=>"011111111",
  63499=>"000101101",
  63500=>"111111111",
  63501=>"101101101",
  63502=>"100000000",
  63503=>"000100000",
  63504=>"111111001",
  63505=>"000000000",
  63506=>"011111111",
  63507=>"010010000",
  63508=>"011000000",
  63509=>"000000110",
  63510=>"101111101",
  63511=>"100111111",
  63512=>"110110111",
  63513=>"111111101",
  63514=>"101000001",
  63515=>"110111000",
  63516=>"001011111",
  63517=>"000111111",
  63518=>"111111111",
  63519=>"000000111",
  63520=>"000001001",
  63521=>"110000111",
  63522=>"000000000",
  63523=>"111111001",
  63524=>"010011000",
  63525=>"000011111",
  63526=>"000000000",
  63527=>"000000000",
  63528=>"111111000",
  63529=>"000000000",
  63530=>"000000000",
  63531=>"110100000",
  63532=>"000000000",
  63533=>"111111100",
  63534=>"000000000",
  63535=>"111111000",
  63536=>"000000111",
  63537=>"001001001",
  63538=>"001011000",
  63539=>"000000000",
  63540=>"111111110",
  63541=>"000011011",
  63542=>"011111111",
  63543=>"000000000",
  63544=>"110110111",
  63545=>"111111010",
  63546=>"000000000",
  63547=>"001111111",
  63548=>"000000111",
  63549=>"011111000",
  63550=>"001011000",
  63551=>"000000000",
  63552=>"000110111",
  63553=>"010000110",
  63554=>"111111111",
  63555=>"101110110",
  63556=>"100111111",
  63557=>"000000001",
  63558=>"000011111",
  63559=>"111100000",
  63560=>"001000000",
  63561=>"000000001",
  63562=>"111111011",
  63563=>"000101100",
  63564=>"111111000",
  63565=>"011011001",
  63566=>"011111001",
  63567=>"000000000",
  63568=>"000110110",
  63569=>"000000111",
  63570=>"000100110",
  63571=>"001001000",
  63572=>"000000000",
  63573=>"000000111",
  63574=>"101111111",
  63575=>"101111111",
  63576=>"111111100",
  63577=>"000000000",
  63578=>"001101111",
  63579=>"000001001",
  63580=>"111111111",
  63581=>"000000000",
  63582=>"110100000",
  63583=>"001000110",
  63584=>"000111111",
  63585=>"000000111",
  63586=>"000000000",
  63587=>"000000111",
  63588=>"010000000",
  63589=>"000000110",
  63590=>"111111111",
  63591=>"000000000",
  63592=>"000000000",
  63593=>"010010111",
  63594=>"000000111",
  63595=>"101000000",
  63596=>"100100000",
  63597=>"111111110",
  63598=>"111111111",
  63599=>"000000111",
  63600=>"001110111",
  63601=>"000000000",
  63602=>"001001101",
  63603=>"100000001",
  63604=>"000100100",
  63605=>"100010000",
  63606=>"111111111",
  63607=>"000000000",
  63608=>"111100111",
  63609=>"111111101",
  63610=>"000000000",
  63611=>"011011101",
  63612=>"000001000",
  63613=>"001001000",
  63614=>"111111111",
  63615=>"001000000",
  63616=>"000000001",
  63617=>"000001000",
  63618=>"000000101",
  63619=>"011011011",
  63620=>"000000000",
  63621=>"000001111",
  63622=>"111111111",
  63623=>"111111111",
  63624=>"111110100",
  63625=>"001001111",
  63626=>"111111111",
  63627=>"011000001",
  63628=>"100000000",
  63629=>"000000000",
  63630=>"101111101",
  63631=>"110000110",
  63632=>"101001001",
  63633=>"000000000",
  63634=>"011111011",
  63635=>"110111111",
  63636=>"000000111",
  63637=>"000111110",
  63638=>"000000000",
  63639=>"000000001",
  63640=>"001001111",
  63641=>"101111000",
  63642=>"111111000",
  63643=>"000000000",
  63644=>"000011000",
  63645=>"000000000",
  63646=>"111111000",
  63647=>"001000000",
  63648=>"000110111",
  63649=>"000110010",
  63650=>"000000110",
  63651=>"111111100",
  63652=>"111000000",
  63653=>"100100100",
  63654=>"111000000",
  63655=>"110000000",
  63656=>"111111111",
  63657=>"000000000",
  63658=>"111111111",
  63659=>"000101100",
  63660=>"111001000",
  63661=>"011011001",
  63662=>"111111000",
  63663=>"000000001",
  63664=>"110110000",
  63665=>"100111001",
  63666=>"111111000",
  63667=>"111100001",
  63668=>"000000000",
  63669=>"000001000",
  63670=>"000000000",
  63671=>"010000110",
  63672=>"110100000",
  63673=>"001000111",
  63674=>"111111101",
  63675=>"101111001",
  63676=>"000000000",
  63677=>"000000000",
  63678=>"111111111",
  63679=>"111111111",
  63680=>"000011011",
  63681=>"110110000",
  63682=>"111111111",
  63683=>"111111111",
  63684=>"000000000",
  63685=>"000000000",
  63686=>"111000000",
  63687=>"001000110",
  63688=>"111111000",
  63689=>"000000000",
  63690=>"001000000",
  63691=>"100000111",
  63692=>"000000111",
  63693=>"101101000",
  63694=>"111111111",
  63695=>"001100111",
  63696=>"111100000",
  63697=>"111111111",
  63698=>"111101101",
  63699=>"110111111",
  63700=>"000100100",
  63701=>"100001011",
  63702=>"111111111",
  63703=>"000000000",
  63704=>"101000110",
  63705=>"111111111",
  63706=>"000000111",
  63707=>"111111111",
  63708=>"000111100",
  63709=>"001000101",
  63710=>"000000000",
  63711=>"101011100",
  63712=>"000000000",
  63713=>"110010010",
  63714=>"111111110",
  63715=>"011011011",
  63716=>"111111111",
  63717=>"000000100",
  63718=>"000000000",
  63719=>"111111111",
  63720=>"111000111",
  63721=>"000000001",
  63722=>"111111111",
  63723=>"100011100",
  63724=>"111111111",
  63725=>"111111111",
  63726=>"111101000",
  63727=>"000011001",
  63728=>"111111111",
  63729=>"001001111",
  63730=>"100000100",
  63731=>"011111000",
  63732=>"011000000",
  63733=>"000110011",
  63734=>"100100111",
  63735=>"100110111",
  63736=>"101100111",
  63737=>"111111111",
  63738=>"000000000",
  63739=>"000000000",
  63740=>"111111111",
  63741=>"110111011",
  63742=>"111111001",
  63743=>"000000000",
  63744=>"001001000",
  63745=>"101101101",
  63746=>"110110111",
  63747=>"001001111",
  63748=>"000000000",
  63749=>"111100000",
  63750=>"000000000",
  63751=>"000000100",
  63752=>"111111000",
  63753=>"111111111",
  63754=>"000000000",
  63755=>"111000000",
  63756=>"111111111",
  63757=>"000100100",
  63758=>"100110110",
  63759=>"000000000",
  63760=>"000000100",
  63761=>"100111111",
  63762=>"000000000",
  63763=>"001001000",
  63764=>"111111001",
  63765=>"111111111",
  63766=>"100000000",
  63767=>"001101100",
  63768=>"111111111",
  63769=>"111111001",
  63770=>"000000000",
  63771=>"110110111",
  63772=>"111101000",
  63773=>"110000010",
  63774=>"000100111",
  63775=>"011110111",
  63776=>"111111110",
  63777=>"000000000",
  63778=>"000111010",
  63779=>"111111000",
  63780=>"010000000",
  63781=>"111111111",
  63782=>"001101110",
  63783=>"111111111",
  63784=>"111101101",
  63785=>"000000000",
  63786=>"111111001",
  63787=>"111111111",
  63788=>"000000100",
  63789=>"111111111",
  63790=>"100000010",
  63791=>"000000000",
  63792=>"100000000",
  63793=>"111111110",
  63794=>"000000011",
  63795=>"100001011",
  63796=>"000000001",
  63797=>"101111110",
  63798=>"000000111",
  63799=>"000000000",
  63800=>"000000000",
  63801=>"111001000",
  63802=>"100000101",
  63803=>"000000000",
  63804=>"111111111",
  63805=>"101111111",
  63806=>"100101101",
  63807=>"111001111",
  63808=>"111111111",
  63809=>"111111111",
  63810=>"111111010",
  63811=>"111111111",
  63812=>"011011011",
  63813=>"000110111",
  63814=>"000000000",
  63815=>"111111011",
  63816=>"000000000",
  63817=>"000000000",
  63818=>"001110000",
  63819=>"100110100",
  63820=>"111111111",
  63821=>"100111110",
  63822=>"011111110",
  63823=>"110000000",
  63824=>"001101111",
  63825=>"000000000",
  63826=>"001011000",
  63827=>"000000000",
  63828=>"111100000",
  63829=>"001001011",
  63830=>"110000000",
  63831=>"111111111",
  63832=>"111111111",
  63833=>"000011011",
  63834=>"111000000",
  63835=>"101100000",
  63836=>"000000000",
  63837=>"000000000",
  63838=>"110110010",
  63839=>"111111001",
  63840=>"000000000",
  63841=>"111111111",
  63842=>"111110000",
  63843=>"111111111",
  63844=>"101101001",
  63845=>"101111111",
  63846=>"110111111",
  63847=>"001011111",
  63848=>"110111011",
  63849=>"111000000",
  63850=>"111111100",
  63851=>"111111111",
  63852=>"111110100",
  63853=>"011001000",
  63854=>"000000111",
  63855=>"111100100",
  63856=>"000000000",
  63857=>"000000001",
  63858=>"000001110",
  63859=>"100100101",
  63860=>"000001011",
  63861=>"101000000",
  63862=>"001011001",
  63863=>"101111000",
  63864=>"000000100",
  63865=>"000000001",
  63866=>"000111111",
  63867=>"000111001",
  63868=>"000000000",
  63869=>"111111000",
  63870=>"000001111",
  63871=>"111111111",
  63872=>"000000001",
  63873=>"000000000",
  63874=>"001001010",
  63875=>"000000000",
  63876=>"000000111",
  63877=>"000000000",
  63878=>"011111011",
  63879=>"001111010",
  63880=>"000000000",
  63881=>"111100000",
  63882=>"000000000",
  63883=>"111111010",
  63884=>"101000111",
  63885=>"100100111",
  63886=>"110000000",
  63887=>"111111111",
  63888=>"000000000",
  63889=>"011011000",
  63890=>"000000000",
  63891=>"111111110",
  63892=>"000000000",
  63893=>"010100000",
  63894=>"011111111",
  63895=>"001011001",
  63896=>"000001111",
  63897=>"011000001",
  63898=>"000000000",
  63899=>"000000001",
  63900=>"000000001",
  63901=>"001000000",
  63902=>"111101101",
  63903=>"100111111",
  63904=>"000011000",
  63905=>"111001101",
  63906=>"011111000",
  63907=>"001000000",
  63908=>"000000111",
  63909=>"111111111",
  63910=>"000000001",
  63911=>"000000101",
  63912=>"110100110",
  63913=>"101000000",
  63914=>"111111111",
  63915=>"111111111",
  63916=>"011000000",
  63917=>"111111111",
  63918=>"011111010",
  63919=>"111111100",
  63920=>"000000000",
  63921=>"001000000",
  63922=>"111011111",
  63923=>"111111111",
  63924=>"000000000",
  63925=>"111100000",
  63926=>"111111111",
  63927=>"110100000",
  63928=>"101001111",
  63929=>"111111110",
  63930=>"110110010",
  63931=>"000000000",
  63932=>"000000100",
  63933=>"000000000",
  63934=>"000000000",
  63935=>"111111111",
  63936=>"111111001",
  63937=>"111111111",
  63938=>"111111111",
  63939=>"000000000",
  63940=>"111110000",
  63941=>"011000101",
  63942=>"000000000",
  63943=>"111111100",
  63944=>"001111101",
  63945=>"101000000",
  63946=>"001001111",
  63947=>"111011010",
  63948=>"100111111",
  63949=>"111111000",
  63950=>"001000000",
  63951=>"101111000",
  63952=>"111111111",
  63953=>"111010100",
  63954=>"111111111",
  63955=>"110111111",
  63956=>"110110111",
  63957=>"111111000",
  63958=>"111001011",
  63959=>"100100100",
  63960=>"110111001",
  63961=>"000000000",
  63962=>"000010000",
  63963=>"000000000",
  63964=>"000011011",
  63965=>"000000000",
  63966=>"111110000",
  63967=>"001101101",
  63968=>"101100000",
  63969=>"000110110",
  63970=>"000110010",
  63971=>"010010001",
  63972=>"111111000",
  63973=>"001000000",
  63974=>"100100001",
  63975=>"000000000",
  63976=>"001000001",
  63977=>"111111011",
  63978=>"000011000",
  63979=>"101000101",
  63980=>"000000000",
  63981=>"100100100",
  63982=>"000000111",
  63983=>"111111111",
  63984=>"000000000",
  63985=>"000000111",
  63986=>"010100111",
  63987=>"011000000",
  63988=>"111111111",
  63989=>"111111111",
  63990=>"000000111",
  63991=>"000101111",
  63992=>"111111000",
  63993=>"101100111",
  63994=>"110110110",
  63995=>"111111011",
  63996=>"000000000",
  63997=>"000110111",
  63998=>"001000000",
  63999=>"001000001",
  64000=>"110111111",
  64001=>"010110000",
  64002=>"000010011",
  64003=>"000100100",
  64004=>"110110111",
  64005=>"100000000",
  64006=>"111111111",
  64007=>"000000000",
  64008=>"100000000",
  64009=>"111011001",
  64010=>"001000000",
  64011=>"111111100",
  64012=>"000000000",
  64013=>"000110100",
  64014=>"001001011",
  64015=>"011111111",
  64016=>"100100111",
  64017=>"000111111",
  64018=>"000000000",
  64019=>"101111111",
  64020=>"010010010",
  64021=>"000000000",
  64022=>"110110000",
  64023=>"010110100",
  64024=>"100111111",
  64025=>"100100100",
  64026=>"110111000",
  64027=>"111011011",
  64028=>"001011111",
  64029=>"111000000",
  64030=>"111111111",
  64031=>"000000100",
  64032=>"111111011",
  64033=>"111111111",
  64034=>"111100100",
  64035=>"100111111",
  64036=>"000000000",
  64037=>"001000000",
  64038=>"111110100",
  64039=>"100000000",
  64040=>"100000100",
  64041=>"011000000",
  64042=>"001001111",
  64043=>"111111000",
  64044=>"000000001",
  64045=>"000000111",
  64046=>"101001111",
  64047=>"111111111",
  64048=>"111111111",
  64049=>"001001011",
  64050=>"000000000",
  64051=>"001011011",
  64052=>"101101111",
  64053=>"011111111",
  64054=>"110101111",
  64055=>"000001000",
  64056=>"000011001",
  64057=>"000000000",
  64058=>"100000100",
  64059=>"111010000",
  64060=>"000000001",
  64061=>"000110111",
  64062=>"111101101",
  64063=>"111111111",
  64064=>"110011111",
  64065=>"000000110",
  64066=>"111111101",
  64067=>"110111100",
  64068=>"100000101",
  64069=>"111111111",
  64070=>"000000010",
  64071=>"110110111",
  64072=>"000001111",
  64073=>"111111000",
  64074=>"011011011",
  64075=>"111111100",
  64076=>"001000100",
  64077=>"100100100",
  64078=>"111011001",
  64079=>"001001001",
  64080=>"000100111",
  64081=>"100101111",
  64082=>"000000000",
  64083=>"100110110",
  64084=>"000000111",
  64085=>"000100110",
  64086=>"011011011",
  64087=>"000000000",
  64088=>"110111100",
  64089=>"111111100",
  64090=>"111111111",
  64091=>"110110000",
  64092=>"000011010",
  64093=>"111101000",
  64094=>"000000000",
  64095=>"111111110",
  64096=>"111111111",
  64097=>"000010000",
  64098=>"111111111",
  64099=>"001011111",
  64100=>"110110110",
  64101=>"111111111",
  64102=>"111111001",
  64103=>"111111111",
  64104=>"000000000",
  64105=>"111000000",
  64106=>"001001011",
  64107=>"111111000",
  64108=>"110110110",
  64109=>"011000000",
  64110=>"111111000",
  64111=>"101000000",
  64112=>"000001001",
  64113=>"011111111",
  64114=>"111111011",
  64115=>"010000000",
  64116=>"111011111",
  64117=>"110111111",
  64118=>"111111111",
  64119=>"000000000",
  64120=>"111110010",
  64121=>"110000001",
  64122=>"000000100",
  64123=>"111111111",
  64124=>"000000101",
  64125=>"101100100",
  64126=>"000000000",
  64127=>"000000000",
  64128=>"000000100",
  64129=>"111111000",
  64130=>"011001000",
  64131=>"000000000",
  64132=>"100100111",
  64133=>"000000011",
  64134=>"110000000",
  64135=>"111111000",
  64136=>"100110000",
  64137=>"000000000",
  64138=>"111111010",
  64139=>"110010000",
  64140=>"011000000",
  64141=>"111001000",
  64142=>"000001111",
  64143=>"000000000",
  64144=>"111111111",
  64145=>"111111111",
  64146=>"110000000",
  64147=>"100110110",
  64148=>"000001000",
  64149=>"111000000",
  64150=>"000000000",
  64151=>"111110000",
  64152=>"000100111",
  64153=>"000000000",
  64154=>"000000000",
  64155=>"010011011",
  64156=>"000111110",
  64157=>"110110011",
  64158=>"111111111",
  64159=>"000000000",
  64160=>"111000000",
  64161=>"101001011",
  64162=>"000000000",
  64163=>"101111111",
  64164=>"110100100",
  64165=>"000000000",
  64166=>"110111111",
  64167=>"110100000",
  64168=>"111001000",
  64169=>"111111111",
  64170=>"001000000",
  64171=>"111100000",
  64172=>"111111111",
  64173=>"100001000",
  64174=>"100100101",
  64175=>"011111111",
  64176=>"111010111",
  64177=>"000000000",
  64178=>"000000000",
  64179=>"111100000",
  64180=>"000000000",
  64181=>"110000111",
  64182=>"001111111",
  64183=>"000001111",
  64184=>"110000000",
  64185=>"110110111",
  64186=>"011111111",
  64187=>"111101101",
  64188=>"000011111",
  64189=>"110000000",
  64190=>"111000000",
  64191=>"111001001",
  64192=>"000000000",
  64193=>"110111111",
  64194=>"101011010",
  64195=>"100100111",
  64196=>"000100111",
  64197=>"000000111",
  64198=>"111111111",
  64199=>"000000000",
  64200=>"110110000",
  64201=>"111111111",
  64202=>"000001001",
  64203=>"000000000",
  64204=>"000000000",
  64205=>"001111111",
  64206=>"000000001",
  64207=>"111111010",
  64208=>"110111111",
  64209=>"111110000",
  64210=>"111111000",
  64211=>"000000000",
  64212=>"111000000",
  64213=>"111011111",
  64214=>"111111111",
  64215=>"110111111",
  64216=>"100000001",
  64217=>"001111111",
  64218=>"111111010",
  64219=>"111000000",
  64220=>"111111111",
  64221=>"110100101",
  64222=>"000100110",
  64223=>"110100000",
  64224=>"111011011",
  64225=>"000010011",
  64226=>"000000000",
  64227=>"000000000",
  64228=>"100111111",
  64229=>"000001001",
  64230=>"000001000",
  64231=>"111111101",
  64232=>"111111111",
  64233=>"000001001",
  64234=>"001001111",
  64235=>"111001111",
  64236=>"000000000",
  64237=>"111111111",
  64238=>"111111110",
  64239=>"111111111",
  64240=>"000001011",
  64241=>"011000101",
  64242=>"000000000",
  64243=>"111111010",
  64244=>"000000000",
  64245=>"110110100",
  64246=>"011010000",
  64247=>"111001000",
  64248=>"000001011",
  64249=>"011111111",
  64250=>"000000111",
  64251=>"000100100",
  64252=>"001011111",
  64253=>"110110111",
  64254=>"001000000",
  64255=>"000000001",
  64256=>"111110000",
  64257=>"000000000",
  64258=>"000000111",
  64259=>"111111001",
  64260=>"000000100",
  64261=>"000000100",
  64262=>"000101111",
  64263=>"011101111",
  64264=>"000000000",
  64265=>"100100100",
  64266=>"111111100",
  64267=>"000010110",
  64268=>"110000100",
  64269=>"111000000",
  64270=>"111111111",
  64271=>"111000000",
  64272=>"000000000",
  64273=>"100110100",
  64274=>"000000000",
  64275=>"000000000",
  64276=>"001001111",
  64277=>"000000000",
  64278=>"000000000",
  64279=>"111111011",
  64280=>"111111111",
  64281=>"000000000",
  64282=>"101001000",
  64283=>"011111111",
  64284=>"110000000",
  64285=>"000000000",
  64286=>"110111111",
  64287=>"100000000",
  64288=>"011001100",
  64289=>"000000000",
  64290=>"011011011",
  64291=>"111111111",
  64292=>"000011011",
  64293=>"110000000",
  64294=>"100000000",
  64295=>"011011001",
  64296=>"111111111",
  64297=>"111000000",
  64298=>"111011111",
  64299=>"000000000",
  64300=>"000000000",
  64301=>"100100100",
  64302=>"000000000",
  64303=>"001000000",
  64304=>"000000000",
  64305=>"000100110",
  64306=>"111111111",
  64307=>"001111111",
  64308=>"000000000",
  64309=>"000000011",
  64310=>"100100000",
  64311=>"000000000",
  64312=>"010000000",
  64313=>"000000111",
  64314=>"111111110",
  64315=>"000000000",
  64316=>"000000000",
  64317=>"111101111",
  64318=>"000000000",
  64319=>"001011111",
  64320=>"000000000",
  64321=>"111111111",
  64322=>"100000000",
  64323=>"111111111",
  64324=>"000110111",
  64325=>"100110100",
  64326=>"010000001",
  64327=>"000000000",
  64328=>"000000111",
  64329=>"111011010",
  64330=>"111111111",
  64331=>"100100100",
  64332=>"110100000",
  64333=>"000000111",
  64334=>"001111000",
  64335=>"110111111",
  64336=>"011011111",
  64337=>"000000111",
  64338=>"011000001",
  64339=>"000000110",
  64340=>"000000000",
  64341=>"111111111",
  64342=>"111101000",
  64343=>"111001000",
  64344=>"101111111",
  64345=>"110000000",
  64346=>"000000011",
  64347=>"000000111",
  64348=>"111111011",
  64349=>"111111111",
  64350=>"000011011",
  64351=>"001001000",
  64352=>"000000000",
  64353=>"111111111",
  64354=>"111111010",
  64355=>"111111011",
  64356=>"111111111",
  64357=>"100111111",
  64358=>"000000000",
  64359=>"110100100",
  64360=>"001001001",
  64361=>"111110000",
  64362=>"000000000",
  64363=>"000000011",
  64364=>"000100000",
  64365=>"111000111",
  64366=>"000000000",
  64367=>"011011011",
  64368=>"111111111",
  64369=>"001000000",
  64370=>"001011000",
  64371=>"000000000",
  64372=>"111111001",
  64373=>"000011111",
  64374=>"000000000",
  64375=>"010000000",
  64376=>"001001000",
  64377=>"000110100",
  64378=>"111100000",
  64379=>"100101100",
  64380=>"111011010",
  64381=>"001001011",
  64382=>"111111111",
  64383=>"111000000",
  64384=>"100000000",
  64385=>"100111011",
  64386=>"111111111",
  64387=>"000000000",
  64388=>"111100000",
  64389=>"100111101",
  64390=>"011011011",
  64391=>"111111001",
  64392=>"000001001",
  64393=>"111100000",
  64394=>"000000100",
  64395=>"111000000",
  64396=>"111111111",
  64397=>"001111111",
  64398=>"000000000",
  64399=>"000000000",
  64400=>"000110110",
  64401=>"111101100",
  64402=>"111110100",
  64403=>"000000000",
  64404=>"111000000",
  64405=>"001000000",
  64406=>"100100000",
  64407=>"100100110",
  64408=>"000000000",
  64409=>"111111111",
  64410=>"010110111",
  64411=>"000100111",
  64412=>"111111111",
  64413=>"111111111",
  64414=>"111111111",
  64415=>"000000000",
  64416=>"111111110",
  64417=>"111111101",
  64418=>"000000000",
  64419=>"110111110",
  64420=>"000000111",
  64421=>"000100110",
  64422=>"000000100",
  64423=>"110110111",
  64424=>"111110111",
  64425=>"001001001",
  64426=>"111001111",
  64427=>"111000011",
  64428=>"011111111",
  64429=>"001011001",
  64430=>"111111010",
  64431=>"111100111",
  64432=>"000000010",
  64433=>"111111000",
  64434=>"000000000",
  64435=>"111111111",
  64436=>"110000000",
  64437=>"111111111",
  64438=>"111111111",
  64439=>"001000001",
  64440=>"010100000",
  64441=>"000000000",
  64442=>"111101000",
  64443=>"111111111",
  64444=>"000111111",
  64445=>"111111001",
  64446=>"000000001",
  64447=>"110001011",
  64448=>"100111111",
  64449=>"000000011",
  64450=>"000000000",
  64451=>"111000000",
  64452=>"000000100",
  64453=>"100110111",
  64454=>"111110000",
  64455=>"000100110",
  64456=>"000100000",
  64457=>"111111110",
  64458=>"111111100",
  64459=>"110111111",
  64460=>"110000111",
  64461=>"000000000",
  64462=>"111111000",
  64463=>"110000000",
  64464=>"000000000",
  64465=>"000100100",
  64466=>"000001101",
  64467=>"000000111",
  64468=>"111111111",
  64469=>"100100110",
  64470=>"100110111",
  64471=>"000000110",
  64472=>"111111011",
  64473=>"101000111",
  64474=>"110101000",
  64475=>"011011011",
  64476=>"111111111",
  64477=>"111111111",
  64478=>"111111010",
  64479=>"010000000",
  64480=>"000111111",
  64481=>"000000000",
  64482=>"011000000",
  64483=>"000001011",
  64484=>"000111111",
  64485=>"000101111",
  64486=>"111000000",
  64487=>"000110000",
  64488=>"000100000",
  64489=>"001110111",
  64490=>"000000000",
  64491=>"000000000",
  64492=>"000000000",
  64493=>"000000001",
  64494=>"000000000",
  64495=>"000000100",
  64496=>"011011001",
  64497=>"111111111",
  64498=>"000000111",
  64499=>"111000000",
  64500=>"000000000",
  64501=>"111111101",
  64502=>"111111111",
  64503=>"101111001",
  64504=>"111111001",
  64505=>"000100100",
  64506=>"000111011",
  64507=>"111111011",
  64508=>"000000001",
  64509=>"100100100",
  64510=>"000000000",
  64511=>"001000000",
  64512=>"111111011",
  64513=>"000000111",
  64514=>"111110110",
  64515=>"001000000",
  64516=>"111011010",
  64517=>"000010011",
  64518=>"111111111",
  64519=>"110111111",
  64520=>"111111111",
  64521=>"111111000",
  64522=>"001000011",
  64523=>"011000111",
  64524=>"001000000",
  64525=>"111001011",
  64526=>"000000000",
  64527=>"111111111",
  64528=>"111111001",
  64529=>"111011111",
  64530=>"111001000",
  64531=>"000100000",
  64532=>"010111111",
  64533=>"111111000",
  64534=>"111111001",
  64535=>"011011001",
  64536=>"000110110",
  64537=>"101001000",
  64538=>"000000000",
  64539=>"000100110",
  64540=>"000000111",
  64541=>"111110111",
  64542=>"110111111",
  64543=>"001111111",
  64544=>"000000111",
  64545=>"111000011",
  64546=>"000100111",
  64547=>"111111111",
  64548=>"010110010",
  64549=>"010111111",
  64550=>"011111111",
  64551=>"000000000",
  64552=>"111111000",
  64553=>"000000000",
  64554=>"000000110",
  64555=>"000010111",
  64556=>"000111111",
  64557=>"111110000",
  64558=>"000000111",
  64559=>"000000000",
  64560=>"110000000",
  64561=>"000000000",
  64562=>"001111000",
  64563=>"111000000",
  64564=>"011001001",
  64565=>"111001011",
  64566=>"111000000",
  64567=>"110111000",
  64568=>"000111110",
  64569=>"110100000",
  64570=>"000000111",
  64571=>"000000111",
  64572=>"111110000",
  64573=>"000100111",
  64574=>"110110110",
  64575=>"101000001",
  64576=>"111110111",
  64577=>"000011111",
  64578=>"000110111",
  64579=>"000000000",
  64580=>"000000000",
  64581=>"111111000",
  64582=>"000000000",
  64583=>"011000000",
  64584=>"001001000",
  64585=>"000000110",
  64586=>"000110111",
  64587=>"000000110",
  64588=>"000000001",
  64589=>"101000111",
  64590=>"110100100",
  64591=>"000001000",
  64592=>"111000000",
  64593=>"111110000",
  64594=>"111000000",
  64595=>"110000000",
  64596=>"111000000",
  64597=>"000111111",
  64598=>"000000000",
  64599=>"000000111",
  64600=>"000000000",
  64601=>"000000000",
  64602=>"111111011",
  64603=>"000001111",
  64604=>"110111111",
  64605=>"000111111",
  64606=>"001111111",
  64607=>"001001000",
  64608=>"111011110",
  64609=>"111110010",
  64610=>"111111111",
  64611=>"111111000",
  64612=>"000010011",
  64613=>"100111111",
  64614=>"111010000",
  64615=>"000000000",
  64616=>"111111111",
  64617=>"000000000",
  64618=>"010000000",
  64619=>"000000000",
  64620=>"110110110",
  64621=>"000101101",
  64622=>"111110100",
  64623=>"000000000",
  64624=>"000010111",
  64625=>"100000000",
  64626=>"111001011",
  64627=>"111111000",
  64628=>"101000000",
  64629=>"100111100",
  64630=>"010000000",
  64631=>"000000000",
  64632=>"000000000",
  64633=>"000000111",
  64634=>"001001000",
  64635=>"111000000",
  64636=>"111101110",
  64637=>"111111001",
  64638=>"001000000",
  64639=>"000000000",
  64640=>"111011000",
  64641=>"110111111",
  64642=>"000000111",
  64643=>"000101001",
  64644=>"001011111",
  64645=>"111111111",
  64646=>"000000000",
  64647=>"100000001",
  64648=>"011111111",
  64649=>"000100000",
  64650=>"111011000",
  64651=>"011111111",
  64652=>"000111111",
  64653=>"111111111",
  64654=>"111111111",
  64655=>"001001111",
  64656=>"010111111",
  64657=>"111111111",
  64658=>"100111111",
  64659=>"000000000",
  64660=>"111111000",
  64661=>"100101001",
  64662=>"000111111",
  64663=>"111111111",
  64664=>"111001001",
  64665=>"000110111",
  64666=>"111111111",
  64667=>"000000111",
  64668=>"000010111",
  64669=>"110000011",
  64670=>"000000111",
  64671=>"001000100",
  64672=>"101010111",
  64673=>"000000110",
  64674=>"000000000",
  64675=>"000100110",
  64676=>"111011000",
  64677=>"111000000",
  64678=>"011111011",
  64679=>"111011001",
  64680=>"011111111",
  64681=>"000000111",
  64682=>"111111111",
  64683=>"111010000",
  64684=>"000000000",
  64685=>"110111110",
  64686=>"110010111",
  64687=>"011111111",
  64688=>"000000111",
  64689=>"100000001",
  64690=>"011111010",
  64691=>"111110110",
  64692=>"000111111",
  64693=>"101000010",
  64694=>"111111111",
  64695=>"000000111",
  64696=>"000111111",
  64697=>"111011011",
  64698=>"001000111",
  64699=>"000001011",
  64700=>"000000000",
  64701=>"110000000",
  64702=>"111111111",
  64703=>"000000000",
  64704=>"000110000",
  64705=>"000101111",
  64706=>"111000000",
  64707=>"101111111",
  64708=>"000000111",
  64709=>"001111111",
  64710=>"000100000",
  64711=>"111000000",
  64712=>"110111111",
  64713=>"000000000",
  64714=>"101000000",
  64715=>"000000000",
  64716=>"000101111",
  64717=>"111001000",
  64718=>"000011111",
  64719=>"000100100",
  64720=>"001010111",
  64721=>"001000111",
  64722=>"100111111",
  64723=>"000100111",
  64724=>"111111000",
  64725=>"100100011",
  64726=>"100000000",
  64727=>"111000100",
  64728=>"100111001",
  64729=>"110111111",
  64730=>"000000010",
  64731=>"111111111",
  64732=>"100000111",
  64733=>"101111111",
  64734=>"111000000",
  64735=>"100000000",
  64736=>"000111011",
  64737=>"000000000",
  64738=>"111111000",
  64739=>"000000000",
  64740=>"110101000",
  64741=>"011111111",
  64742=>"000111111",
  64743=>"010111010",
  64744=>"000100111",
  64745=>"000000000",
  64746=>"111111100",
  64747=>"101000111",
  64748=>"111001001",
  64749=>"111001000",
  64750=>"110000010",
  64751=>"000000000",
  64752=>"000000000",
  64753=>"001000000",
  64754=>"000001000",
  64755=>"000000000",
  64756=>"000000011",
  64757=>"100100000",
  64758=>"111011000",
  64759=>"000000000",
  64760=>"110110111",
  64761=>"111111111",
  64762=>"001000010",
  64763=>"011000110",
  64764=>"110100000",
  64765=>"000000100",
  64766=>"111111000",
  64767=>"111000000",
  64768=>"000000000",
  64769=>"000101111",
  64770=>"111000000",
  64771=>"111111111",
  64772=>"000000000",
  64773=>"010000000",
  64774=>"111111000",
  64775=>"100000111",
  64776=>"111011001",
  64777=>"101100111",
  64778=>"001100111",
  64779=>"000000111",
  64780=>"111001000",
  64781=>"000000111",
  64782=>"011111111",
  64783=>"000000111",
  64784=>"111100000",
  64785=>"111001000",
  64786=>"110111110",
  64787=>"000110110",
  64788=>"001000000",
  64789=>"011000000",
  64790=>"000000000",
  64791=>"111000111",
  64792=>"111111001",
  64793=>"111011000",
  64794=>"000000000",
  64795=>"001000000",
  64796=>"100000010",
  64797=>"111011000",
  64798=>"111111111",
  64799=>"111111101",
  64800=>"000010011",
  64801=>"000110111",
  64802=>"010000000",
  64803=>"000000001",
  64804=>"100110111",
  64805=>"111111001",
  64806=>"100100111",
  64807=>"000000010",
  64808=>"101111111",
  64809=>"001000000",
  64810=>"000000000",
  64811=>"000000011",
  64812=>"000001111",
  64813=>"010010110",
  64814=>"000000111",
  64815=>"000000111",
  64816=>"111000000",
  64817=>"000001000",
  64818=>"000000111",
  64819=>"000000000",
  64820=>"111111110",
  64821=>"000000000",
  64822=>"101000001",
  64823=>"111100000",
  64824=>"000110000",
  64825=>"000000000",
  64826=>"100100111",
  64827=>"111111000",
  64828=>"110111000",
  64829=>"111111111",
  64830=>"011010110",
  64831=>"111000000",
  64832=>"000000001",
  64833=>"111111111",
  64834=>"100000000",
  64835=>"000000101",
  64836=>"000000001",
  64837=>"000000101",
  64838=>"101111111",
  64839=>"000000011",
  64840=>"000000001",
  64841=>"000001111",
  64842=>"000000110",
  64843=>"010000111",
  64844=>"110000001",
  64845=>"000110110",
  64846=>"000000110",
  64847=>"111111000",
  64848=>"001000000",
  64849=>"001000000",
  64850=>"000000000",
  64851=>"000111111",
  64852=>"000000000",
  64853=>"001001001",
  64854=>"001111111",
  64855=>"100000110",
  64856=>"101000111",
  64857=>"111111101",
  64858=>"010110111",
  64859=>"111111111",
  64860=>"000101111",
  64861=>"011001011",
  64862=>"111110100",
  64863=>"000000000",
  64864=>"000010011",
  64865=>"110111111",
  64866=>"111111011",
  64867=>"101001111",
  64868=>"100000110",
  64869=>"111110000",
  64870=>"100111111",
  64871=>"111111011",
  64872=>"000001111",
  64873=>"110000000",
  64874=>"000000001",
  64875=>"000000110",
  64876=>"111111111",
  64877=>"000010111",
  64878=>"000000010",
  64879=>"000000001",
  64880=>"111000111",
  64881=>"000010000",
  64882=>"110010111",
  64883=>"100111011",
  64884=>"011010000",
  64885=>"111111001",
  64886=>"110100000",
  64887=>"001000000",
  64888=>"000000000",
  64889=>"000111011",
  64890=>"111000000",
  64891=>"100100000",
  64892=>"111001111",
  64893=>"010111111",
  64894=>"111111010",
  64895=>"001001111",
  64896=>"000000000",
  64897=>"110111111",
  64898=>"111001001",
  64899=>"000000000",
  64900=>"000000111",
  64901=>"001000000",
  64902=>"000110010",
  64903=>"000000110",
  64904=>"111010000",
  64905=>"101101100",
  64906=>"000100111",
  64907=>"000000111",
  64908=>"111111111",
  64909=>"110100101",
  64910=>"000000000",
  64911=>"000000111",
  64912=>"111000000",
  64913=>"111111011",
  64914=>"111111000",
  64915=>"000111000",
  64916=>"000111110",
  64917=>"000000000",
  64918=>"010000000",
  64919=>"101000000",
  64920=>"000000000",
  64921=>"000000100",
  64922=>"000000000",
  64923=>"111111111",
  64924=>"111000000",
  64925=>"110000110",
  64926=>"111100100",
  64927=>"010000000",
  64928=>"001001001",
  64929=>"011011000",
  64930=>"110000011",
  64931=>"111001000",
  64932=>"000000101",
  64933=>"000110111",
  64934=>"000000100",
  64935=>"111111111",
  64936=>"000011110",
  64937=>"010111111",
  64938=>"100000000",
  64939=>"011001000",
  64940=>"111001000",
  64941=>"100000100",
  64942=>"000000000",
  64943=>"111111110",
  64944=>"000000101",
  64945=>"000000100",
  64946=>"000000000",
  64947=>"100100000",
  64948=>"110110100",
  64949=>"000000000",
  64950=>"111000111",
  64951=>"111000000",
  64952=>"000000000",
  64953=>"111111111",
  64954=>"110000000",
  64955=>"111001111",
  64956=>"000000000",
  64957=>"000000000",
  64958=>"000000000",
  64959=>"000100100",
  64960=>"000010111",
  64961=>"000000000",
  64962=>"111111111",
  64963=>"111001000",
  64964=>"000000110",
  64965=>"100111000",
  64966=>"100000010",
  64967=>"101000000",
  64968=>"000000000",
  64969=>"101100000",
  64970=>"110000001",
  64971=>"000000000",
  64972=>"000001001",
  64973=>"010111010",
  64974=>"110010000",
  64975=>"000110111",
  64976=>"010010111",
  64977=>"010111111",
  64978=>"111111111",
  64979=>"111111001",
  64980=>"001000100",
  64981=>"000101100",
  64982=>"100000000",
  64983=>"011011000",
  64984=>"000001000",
  64985=>"100000100",
  64986=>"000000000",
  64987=>"110100000",
  64988=>"000111011",
  64989=>"111101111",
  64990=>"000000011",
  64991=>"000001001",
  64992=>"001000000",
  64993=>"000111101",
  64994=>"000000000",
  64995=>"010111111",
  64996=>"000010111",
  64997=>"111000000",
  64998=>"111111000",
  64999=>"111000001",
  65000=>"110010000",
  65001=>"111000000",
  65002=>"100000000",
  65003=>"100110111",
  65004=>"011010111",
  65005=>"111011001",
  65006=>"010010000",
  65007=>"111000000",
  65008=>"001100100",
  65009=>"101100110",
  65010=>"011011111",
  65011=>"000001111",
  65012=>"001000000",
  65013=>"111101001",
  65014=>"111110000",
  65015=>"100000000",
  65016=>"001111111",
  65017=>"000000011",
  65018=>"011000000",
  65019=>"110111000",
  65020=>"000000111",
  65021=>"111111001",
  65022=>"101110100",
  65023=>"111000000",
  65024=>"001111111",
  65025=>"111111111",
  65026=>"101000000",
  65027=>"000000010",
  65028=>"010000001",
  65029=>"101001111",
  65030=>"000110010",
  65031=>"101000101",
  65032=>"111111100",
  65033=>"000000111",
  65034=>"000000000",
  65035=>"111000000",
  65036=>"000111110",
  65037=>"011001000",
  65038=>"101000100",
  65039=>"111111111",
  65040=>"000011110",
  65041=>"000111111",
  65042=>"000111111",
  65043=>"000000000",
  65044=>"101000000",
  65045=>"111011000",
  65046=>"010000000",
  65047=>"111011011",
  65048=>"110110110",
  65049=>"111101000",
  65050=>"111011111",
  65051=>"111000000",
  65052=>"110000100",
  65053=>"000100100",
  65054=>"111111100",
  65055=>"000000111",
  65056=>"110000101",
  65057=>"010000110",
  65058=>"000000110",
  65059=>"011000000",
  65060=>"000010011",
  65061=>"000111111",
  65062=>"111101000",
  65063=>"111111111",
  65064=>"111100100",
  65065=>"101000000",
  65066=>"000000010",
  65067=>"111001111",
  65068=>"101100000",
  65069=>"100100000",
  65070=>"111111111",
  65071=>"000111111",
  65072=>"000011111",
  65073=>"000000000",
  65074=>"000001000",
  65075=>"000000001",
  65076=>"000000000",
  65077=>"000111110",
  65078=>"000000110",
  65079=>"000000000",
  65080=>"000000111",
  65081=>"011111100",
  65082=>"111100000",
  65083=>"110000000",
  65084=>"000000000",
  65085=>"010001000",
  65086=>"000011111",
  65087=>"001001000",
  65088=>"111000111",
  65089=>"110110100",
  65090=>"111111100",
  65091=>"011000100",
  65092=>"000000100",
  65093=>"111100000",
  65094=>"111100111",
  65095=>"111111111",
  65096=>"101100000",
  65097=>"001000111",
  65098=>"000000000",
  65099=>"000000111",
  65100=>"001100110",
  65101=>"000011111",
  65102=>"111000000",
  65103=>"000000111",
  65104=>"111011000",
  65105=>"000111111",
  65106=>"000000010",
  65107=>"011011011",
  65108=>"000011111",
  65109=>"000000111",
  65110=>"001011111",
  65111=>"111000000",
  65112=>"000001111",
  65113=>"111000101",
  65114=>"111110111",
  65115=>"110110000",
  65116=>"000000111",
  65117=>"111000010",
  65118=>"111111111",
  65119=>"000000011",
  65120=>"000110111",
  65121=>"101011010",
  65122=>"111111110",
  65123=>"111111000",
  65124=>"000000000",
  65125=>"000000001",
  65126=>"000010111",
  65127=>"000000010",
  65128=>"100110111",
  65129=>"000000111",
  65130=>"111101000",
  65131=>"111011111",
  65132=>"110111111",
  65133=>"000010000",
  65134=>"001000111",
  65135=>"100111111",
  65136=>"100100000",
  65137=>"110100100",
  65138=>"000000000",
  65139=>"001000000",
  65140=>"100111011",
  65141=>"111111111",
  65142=>"000011111",
  65143=>"000000000",
  65144=>"000000001",
  65145=>"000000000",
  65146=>"110110110",
  65147=>"000000000",
  65148=>"110111111",
  65149=>"110010000",
  65150=>"111111111",
  65151=>"010001000",
  65152=>"111110000",
  65153=>"110111111",
  65154=>"111111000",
  65155=>"111101111",
  65156=>"000010111",
  65157=>"000000111",
  65158=>"111111100",
  65159=>"111111111",
  65160=>"111001010",
  65161=>"111000000",
  65162=>"110110111",
  65163=>"100100111",
  65164=>"001000111",
  65165=>"000000101",
  65166=>"000000000",
  65167=>"000000000",
  65168=>"000111111",
  65169=>"000011111",
  65170=>"101000101",
  65171=>"110110000",
  65172=>"110100100",
  65173=>"000000011",
  65174=>"111111100",
  65175=>"111100000",
  65176=>"101111111",
  65177=>"111111111",
  65178=>"000000000",
  65179=>"001010110",
  65180=>"011000000",
  65181=>"000000000",
  65182=>"011111111",
  65183=>"101100000",
  65184=>"000000000",
  65185=>"111011000",
  65186=>"000011111",
  65187=>"011000100",
  65188=>"000000001",
  65189=>"111000000",
  65190=>"111111111",
  65191=>"000100111",
  65192=>"111011001",
  65193=>"000000000",
  65194=>"111000000",
  65195=>"000000000",
  65196=>"111111000",
  65197=>"000000110",
  65198=>"010110111",
  65199=>"101100100",
  65200=>"000000010",
  65201=>"110110110",
  65202=>"111111111",
  65203=>"000000000",
  65204=>"011001100",
  65205=>"011111111",
  65206=>"111111111",
  65207=>"000000111",
  65208=>"011000000",
  65209=>"000001000",
  65210=>"000000100",
  65211=>"111111111",
  65212=>"111000000",
  65213=>"111010000",
  65214=>"000000000",
  65215=>"110111000",
  65216=>"000000000",
  65217=>"000000000",
  65218=>"010111010",
  65219=>"000000111",
  65220=>"111111000",
  65221=>"000101111",
  65222=>"110111001",
  65223=>"011001011",
  65224=>"011111011",
  65225=>"000000000",
  65226=>"010000000",
  65227=>"000111000",
  65228=>"000000000",
  65229=>"110111000",
  65230=>"111111111",
  65231=>"111000110",
  65232=>"110000000",
  65233=>"000100000",
  65234=>"110111111",
  65235=>"000000000",
  65236=>"011111110",
  65237=>"111111110",
  65238=>"000000000",
  65239=>"111111111",
  65240=>"000001001",
  65241=>"000000000",
  65242=>"111111111",
  65243=>"111111111",
  65244=>"000100100",
  65245=>"111111111",
  65246=>"000000000",
  65247=>"000011011",
  65248=>"001101111",
  65249=>"001000011",
  65250=>"110111111",
  65251=>"111001001",
  65252=>"000111111",
  65253=>"111111101",
  65254=>"000000000",
  65255=>"110100111",
  65256=>"001010111",
  65257=>"110100000",
  65258=>"000110110",
  65259=>"001000000",
  65260=>"000100111",
  65261=>"000000000",
  65262=>"001111111",
  65263=>"000000000",
  65264=>"110111011",
  65265=>"111111000",
  65266=>"111111011",
  65267=>"000001111",
  65268=>"101000111",
  65269=>"100111111",
  65270=>"001000000",
  65271=>"000000100",
  65272=>"100000000",
  65273=>"111111111",
  65274=>"001111111",
  65275=>"000000000",
  65276=>"001111111",
  65277=>"001000000",
  65278=>"110111111",
  65279=>"110110110",
  65280=>"000111111",
  65281=>"110100100",
  65282=>"000001111",
  65283=>"000000111",
  65284=>"000000000",
  65285=>"000110000",
  65286=>"111111001",
  65287=>"001010110",
  65288=>"000000000",
  65289=>"110111110",
  65290=>"111000000",
  65291=>"000011111",
  65292=>"111111111",
  65293=>"000000111",
  65294=>"000000111",
  65295=>"111100000",
  65296=>"000110010",
  65297=>"000000010",
  65298=>"111111110",
  65299=>"000000000",
  65300=>"100000000",
  65301=>"000000000",
  65302=>"001100100",
  65303=>"000000000",
  65304=>"000111110",
  65305=>"111000000",
  65306=>"101101000",
  65307=>"000000000",
  65308=>"111111111",
  65309=>"111111111",
  65310=>"000000000",
  65311=>"000000111",
  65312=>"000100111",
  65313=>"000000110",
  65314=>"101111111",
  65315=>"111110000",
  65316=>"111010000",
  65317=>"001000000",
  65318=>"111111111",
  65319=>"000000000",
  65320=>"000000000",
  65321=>"000000000",
  65322=>"000011100",
  65323=>"101000100",
  65324=>"100000000",
  65325=>"000111101",
  65326=>"000000100",
  65327=>"000000110",
  65328=>"000000000",
  65329=>"000111111",
  65330=>"111111000",
  65331=>"111111010",
  65332=>"011000000",
  65333=>"000000111",
  65334=>"100000000",
  65335=>"111000111",
  65336=>"111111111",
  65337=>"111000000",
  65338=>"001000000",
  65339=>"100000000",
  65340=>"111001000",
  65341=>"111111111",
  65342=>"000011011",
  65343=>"000110111",
  65344=>"101111100",
  65345=>"100100110",
  65346=>"011011000",
  65347=>"001011111",
  65348=>"110010111",
  65349=>"111110000",
  65350=>"000000000",
  65351=>"011111110",
  65352=>"101000001",
  65353=>"000000110",
  65354=>"000111100",
  65355=>"011001000",
  65356=>"000000000",
  65357=>"100111001",
  65358=>"111111111",
  65359=>"000011001",
  65360=>"010011001",
  65361=>"111111101",
  65362=>"111000000",
  65363=>"000000111",
  65364=>"000000000",
  65365=>"001011111",
  65366=>"001001111",
  65367=>"111111000",
  65368=>"000001000",
  65369=>"111000000",
  65370=>"001100000",
  65371=>"000000100",
  65372=>"000000100",
  65373=>"010000000",
  65374=>"000000000",
  65375=>"011111110",
  65376=>"000000000",
  65377=>"111111000",
  65378=>"000111100",
  65379=>"000000000",
  65380=>"100110011",
  65381=>"011001001",
  65382=>"000000000",
  65383=>"000000000",
  65384=>"100110000",
  65385=>"000000010",
  65386=>"110000000",
  65387=>"111011001",
  65388=>"100110111",
  65389=>"000000000",
  65390=>"100110100",
  65391=>"111110111",
  65392=>"111001000",
  65393=>"111100111",
  65394=>"000000000",
  65395=>"111111111",
  65396=>"000111000",
  65397=>"000000000",
  65398=>"111110101",
  65399=>"000001001",
  65400=>"000000000",
  65401=>"111111111",
  65402=>"111010001",
  65403=>"110010000",
  65404=>"111111011",
  65405=>"011011010",
  65406=>"110000000",
  65407=>"100000000",
  65408=>"110000000",
  65409=>"001001000",
  65410=>"101101000",
  65411=>"000000000",
  65412=>"111101000",
  65413=>"001011111",
  65414=>"000011000",
  65415=>"111000000",
  65416=>"000000000",
  65417=>"000001000",
  65418=>"000000100",
  65419=>"011001001",
  65420=>"000111111",
  65421=>"001111111",
  65422=>"000000001",
  65423=>"010010000",
  65424=>"000000000",
  65425=>"000111111",
  65426=>"000000000",
  65427=>"110010000",
  65428=>"111111111",
  65429=>"000000000",
  65430=>"000111111",
  65431=>"010111111",
  65432=>"000011111",
  65433=>"111111111",
  65434=>"110000000",
  65435=>"000000000",
  65436=>"111111111",
  65437=>"011111111",
  65438=>"000000111",
  65439=>"000000000",
  65440=>"111111111",
  65441=>"110100101",
  65442=>"100101111",
  65443=>"110100110",
  65444=>"101100100",
  65445=>"111000000",
  65446=>"000110100",
  65447=>"011011011",
  65448=>"000000000",
  65449=>"111111001",
  65450=>"000000000",
  65451=>"000111111",
  65452=>"110010000",
  65453=>"110001001",
  65454=>"111000001",
  65455=>"111011111",
  65456=>"000111111",
  65457=>"000000000",
  65458=>"000011011",
  65459=>"000000000",
  65460=>"001111111",
  65461=>"001001000",
  65462=>"011010111",
  65463=>"111111110",
  65464=>"111110000",
  65465=>"010110111",
  65466=>"000100111",
  65467=>"000000100",
  65468=>"111001111",
  65469=>"001001000",
  65470=>"111111101",
  65471=>"000110110",
  65472=>"111111000",
  65473=>"001111111",
  65474=>"000000000",
  65475=>"110100000",
  65476=>"011111111",
  65477=>"001001110",
  65478=>"011000000",
  65479=>"000100111",
  65480=>"110100111",
  65481=>"000111111",
  65482=>"000000001",
  65483=>"111111010",
  65484=>"111110110",
  65485=>"110111111",
  65486=>"000000000",
  65487=>"011000000",
  65488=>"000000000",
  65489=>"001001011",
  65490=>"000000110",
  65491=>"000000000",
  65492=>"000111111",
  65493=>"111111111",
  65494=>"000100111",
  65495=>"000100100",
  65496=>"101101100",
  65497=>"111111111",
  65498=>"111111010",
  65499=>"101111111",
  65500=>"000000000",
  65501=>"000001111",
  65502=>"111000000",
  65503=>"110110111",
  65504=>"001111111",
  65505=>"000000000",
  65506=>"000011111",
  65507=>"001001111",
  65508=>"111001000",
  65509=>"111111110",
  65510=>"111111111",
  65511=>"111111010",
  65512=>"000010110",
  65513=>"010000111",
  65514=>"000111111",
  65515=>"111111000",
  65516=>"111111111",
  65517=>"000001111",
  65518=>"000000100",
  65519=>"000000001",
  65520=>"000111111",
  65521=>"000011111",
  65522=>"111111000",
  65523=>"010000000",
  65524=>"111111111",
  65525=>"000110110",
  65526=>"000000000",
  65527=>"101000100",
  65528=>"010000000",
  65529=>"111011001",
  65530=>"000111111",
  65531=>"111111000",
  65532=>"000110111",
  65533=>"000000000",
  65534=>"100111111",
  65535=>"001000011");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;