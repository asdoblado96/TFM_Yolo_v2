LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L7_3_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(7) - 1 DOWNTO 0));
END L7_3_WROM;

ARCHITECTURE RTL OF L7_3_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"110111111",
  1=>"000000000",
  2=>"000000111",
  3=>"000000000",
  4=>"000000000",
  5=>"001001000",
  6=>"000000111",
  7=>"111111111",
  8=>"000000111",
  9=>"101111111",
  10=>"111111100",
  11=>"100111111",
  12=>"000000100",
  13=>"000000000",
  14=>"100100100",
  15=>"000000000",
  16=>"000111111",
  17=>"000011111",
  18=>"000000000",
  19=>"111111000",
  20=>"000000110",
  21=>"111111111",
  22=>"000001101",
  23=>"100111111",
  24=>"111111111",
  25=>"110011001",
  26=>"111000000",
  27=>"000000111",
  28=>"111111111",
  29=>"000000010",
  30=>"100000000",
  31=>"010010010",
  32=>"101101111",
  33=>"111001111",
  34=>"000001111",
  35=>"111001000",
  36=>"001011000",
  37=>"111000000",
  38=>"111111101",
  39=>"000000000",
  40=>"111000000",
  41=>"000001011",
  42=>"000000000",
  43=>"111111010",
  44=>"111111111",
  45=>"000000000",
  46=>"110111111",
  47=>"111101001",
  48=>"111111111",
  49=>"000000000",
  50=>"111000000",
  51=>"100110111",
  52=>"110000100",
  53=>"000100111",
  54=>"000000000",
  55=>"000000001",
  56=>"000000111",
  57=>"001000000",
  58=>"101100110",
  59=>"111100101",
  60=>"011111111",
  61=>"111100000",
  62=>"011111111",
  63=>"111000000",
  64=>"000000111",
  65=>"010110110",
  66=>"110111000",
  67=>"111111111",
  68=>"100100100",
  69=>"001000000",
  70=>"100111111",
  71=>"111111111",
  72=>"000011011",
  73=>"111111111",
  74=>"111111111",
  75=>"101111111",
  76=>"100111111",
  77=>"011000000",
  78=>"000000100",
  79=>"111111011",
  80=>"000000000",
  81=>"000000101",
  82=>"111111111",
  83=>"000000011",
  84=>"000000000",
  85=>"101100000",
  86=>"001000000",
  87=>"000000101",
  88=>"011001101",
  89=>"101001000",
  90=>"000000111",
  91=>"010011011",
  92=>"000000000",
  93=>"111001000",
  94=>"000001011",
  95=>"111111000",
  96=>"000111111",
  97=>"000001001",
  98=>"000111111",
  99=>"000111111",
  100=>"101111000",
  101=>"000101111",
  102=>"111000000",
  103=>"000000000",
  104=>"000000111",
  105=>"000000000",
  106=>"101000111",
  107=>"111001000",
  108=>"110110111",
  109=>"111111111",
  110=>"011111111",
  111=>"111111000",
  112=>"111001000",
  113=>"000000110",
  114=>"000110111",
  115=>"000000111",
  116=>"000000000",
  117=>"000100111",
  118=>"000000001",
  119=>"111111011",
  120=>"001111111",
  121=>"111111111",
  122=>"000100000",
  123=>"101111000",
  124=>"110110110",
  125=>"101000000",
  126=>"000000000",
  127=>"011011111",
  128=>"011001100",
  129=>"000000110",
  130=>"000111111",
  131=>"101100000",
  132=>"011011011",
  133=>"001000000",
  134=>"110110000",
  135=>"000000000",
  136=>"000001111",
  137=>"000000000",
  138=>"000000011",
  139=>"111111111",
  140=>"000000000",
  141=>"111111000",
  142=>"111111111",
  143=>"101100000",
  144=>"010000000",
  145=>"111000000",
  146=>"000100111",
  147=>"000111111",
  148=>"000000111",
  149=>"111111000",
  150=>"111111011",
  151=>"000000111",
  152=>"000000110",
  153=>"000000000",
  154=>"000101111",
  155=>"110111111",
  156=>"111000000",
  157=>"000111111",
  158=>"000000000",
  159=>"100000111",
  160=>"001000000",
  161=>"000001001",
  162=>"000011001",
  163=>"001011000",
  164=>"000000001",
  165=>"111110111",
  166=>"111111111",
  167=>"000001001",
  168=>"111111000",
  169=>"001001001",
  170=>"000011111",
  171=>"110111011",
  172=>"101111111",
  173=>"000110111",
  174=>"000001011",
  175=>"111111111",
  176=>"000011000",
  177=>"001111110",
  178=>"111111111",
  179=>"000000111",
  180=>"000000000",
  181=>"111111000",
  182=>"000001000",
  183=>"000011111",
  184=>"111111001",
  185=>"111000101",
  186=>"000000000",
  187=>"011010000",
  188=>"000000000",
  189=>"000000000",
  190=>"101111101",
  191=>"101101000",
  192=>"111111111",
  193=>"000000111",
  194=>"111111100",
  195=>"010000000",
  196=>"000100111",
  197=>"111111001",
  198=>"001001101",
  199=>"111011000",
  200=>"001011111",
  201=>"111111111",
  202=>"000000000",
  203=>"000000000",
  204=>"011011011",
  205=>"111111111",
  206=>"110110110",
  207=>"000010000",
  208=>"000000000",
  209=>"000000000",
  210=>"111001111",
  211=>"111111110",
  212=>"000001000",
  213=>"110111111",
  214=>"000000000",
  215=>"000010110",
  216=>"000000010",
  217=>"001001001",
  218=>"000000000",
  219=>"100111111",
  220=>"111111000",
  221=>"000011000",
  222=>"000000000",
  223=>"000001110",
  224=>"001000100",
  225=>"100110010",
  226=>"010010011",
  227=>"110000111",
  228=>"000000000",
  229=>"000100111",
  230=>"111111111",
  231=>"000111111",
  232=>"111100000",
  233=>"111001001",
  234=>"011011101",
  235=>"000000101",
  236=>"000111000",
  237=>"000000111",
  238=>"111010010",
  239=>"011111000",
  240=>"111111110",
  241=>"000111111",
  242=>"000000010",
  243=>"000000000",
  244=>"000001011",
  245=>"111111000",
  246=>"000001001",
  247=>"110110110",
  248=>"111111001",
  249=>"111111000",
  250=>"111000000",
  251=>"000000000",
  252=>"001001001",
  253=>"000001011",
  254=>"101111011",
  255=>"000000000",
  256=>"111001001",
  257=>"110110110",
  258=>"011011100",
  259=>"000011111",
  260=>"111111111",
  261=>"000000001",
  262=>"111110111",
  263=>"000000000",
  264=>"111111111",
  265=>"000011111",
  266=>"011011011",
  267=>"111111111",
  268=>"000101111",
  269=>"100000000",
  270=>"010111111",
  271=>"000000100",
  272=>"111111000",
  273=>"000000000",
  274=>"100000000",
  275=>"110111111",
  276=>"001001000",
  277=>"111111111",
  278=>"001000000",
  279=>"111010010",
  280=>"111111001",
  281=>"111111111",
  282=>"101000111",
  283=>"000000001",
  284=>"111111111",
  285=>"000011111",
  286=>"011000000",
  287=>"010000110",
  288=>"100101000",
  289=>"110111011",
  290=>"000000111",
  291=>"101001000",
  292=>"111110111",
  293=>"111111111",
  294=>"111110000",
  295=>"111111000",
  296=>"110111111",
  297=>"000100000",
  298=>"000111111",
  299=>"000000000",
  300=>"000000000",
  301=>"001101101",
  302=>"111000000",
  303=>"000011011",
  304=>"000000111",
  305=>"001111111",
  306=>"100110100",
  307=>"111011011",
  308=>"000000110",
  309=>"111111111",
  310=>"000000011",
  311=>"000000111",
  312=>"100000111",
  313=>"100000000",
  314=>"000000000",
  315=>"110111010",
  316=>"111111111",
  317=>"111111010",
  318=>"111011000",
  319=>"010001000",
  320=>"010111000",
  321=>"111111101",
  322=>"111111000",
  323=>"000010000",
  324=>"111111100",
  325=>"000111111",
  326=>"111111000",
  327=>"000000000",
  328=>"000000000",
  329=>"000000000",
  330=>"001011111",
  331=>"100000001",
  332=>"000000110",
  333=>"000100111",
  334=>"111111000",
  335=>"111111111",
  336=>"111001000",
  337=>"010000000",
  338=>"101111111",
  339=>"000111111",
  340=>"000000000",
  341=>"001011011",
  342=>"000000000",
  343=>"101000000",
  344=>"111111111",
  345=>"000000000",
  346=>"101101000",
  347=>"000001000",
  348=>"000000000",
  349=>"111111111",
  350=>"001101111",
  351=>"110000000",
  352=>"111001000",
  353=>"111000000",
  354=>"011000000",
  355=>"000000000",
  356=>"000100100",
  357=>"000000000",
  358=>"011111110",
  359=>"111111110",
  360=>"100000000",
  361=>"000010111",
  362=>"111111111",
  363=>"111111111",
  364=>"100110000",
  365=>"000000000",
  366=>"010111011",
  367=>"111111111",
  368=>"000000000",
  369=>"000110010",
  370=>"000000011",
  371=>"001001111",
  372=>"000111111",
  373=>"111111111",
  374=>"010000111",
  375=>"000000000",
  376=>"011000000",
  377=>"111111111",
  378=>"111111111",
  379=>"000000111",
  380=>"000000011",
  381=>"111111011",
  382=>"000000000",
  383=>"111010001",
  384=>"110110100",
  385=>"111111011",
  386=>"001000000",
  387=>"111110000",
  388=>"100000010",
  389=>"001111000",
  390=>"001101111",
  391=>"111111000",
  392=>"000000111",
  393=>"111000000",
  394=>"111111011",
  395=>"010000111",
  396=>"111111111",
  397=>"000110111",
  398=>"000000011",
  399=>"001001000",
  400=>"010100000",
  401=>"111111101",
  402=>"011011000",
  403=>"110010110",
  404=>"000000000",
  405=>"000000000",
  406=>"000001111",
  407=>"011011111",
  408=>"000000110",
  409=>"000011111",
  410=>"101000000",
  411=>"011111110",
  412=>"000001101",
  413=>"111011000",
  414=>"111111111",
  415=>"000001111",
  416=>"000000010",
  417=>"000111111",
  418=>"000001111",
  419=>"110111111",
  420=>"001011000",
  421=>"000011000",
  422=>"001001111",
  423=>"111111110",
  424=>"111110000",
  425=>"011100100",
  426=>"111111111",
  427=>"011111000",
  428=>"001000000",
  429=>"001011111",
  430=>"000101111",
  431=>"111100000",
  432=>"111111111",
  433=>"000111111",
  434=>"111000000",
  435=>"001100001",
  436=>"111111000",
  437=>"010100000",
  438=>"000111111",
  439=>"111000000",
  440=>"000000000",
  441=>"100110110",
  442=>"000000000",
  443=>"000000010",
  444=>"000000000",
  445=>"101100111",
  446=>"001000111",
  447=>"010010000",
  448=>"111111000",
  449=>"111101001",
  450=>"111111111",
  451=>"000111000",
  452=>"100111111",
  453=>"000101111",
  454=>"000000000",
  455=>"000010111",
  456=>"000000000",
  457=>"110000000",
  458=>"001001111",
  459=>"111011111",
  460=>"010100100",
  461=>"111111111",
  462=>"100001001",
  463=>"111111001",
  464=>"000000000",
  465=>"111000000",
  466=>"000000101",
  467=>"111000000",
  468=>"101111111",
  469=>"100100111",
  470=>"000000000",
  471=>"000000000",
  472=>"000000010",
  473=>"101000000",
  474=>"111000000",
  475=>"010010111",
  476=>"100100101",
  477=>"111111000",
  478=>"000000100",
  479=>"001000001",
  480=>"111111111",
  481=>"000000001",
  482=>"010111111",
  483=>"011000000",
  484=>"000001000",
  485=>"111111111",
  486=>"000101111",
  487=>"000000000",
  488=>"101111111",
  489=>"111011000",
  490=>"011011111",
  491=>"000011110",
  492=>"111111111",
  493=>"000000000",
  494=>"000101111",
  495=>"111100111",
  496=>"000000000",
  497=>"111111111",
  498=>"010000100",
  499=>"110111100",
  500=>"000000111",
  501=>"100001011",
  502=>"111111111",
  503=>"000000001",
  504=>"111111111",
  505=>"000000000",
  506=>"111111101",
  507=>"000000000",
  508=>"000110111",
  509=>"110111000",
  510=>"000000000",
  511=>"111001000",
  512=>"111111111",
  513=>"000000000",
  514=>"000001001",
  515=>"000000111",
  516=>"110100110",
  517=>"111111000",
  518=>"000000011",
  519=>"111111111",
  520=>"010011000",
  521=>"111111010",
  522=>"111001001",
  523=>"000100100",
  524=>"011001000",
  525=>"111111101",
  526=>"000000000",
  527=>"101111111",
  528=>"111000000",
  529=>"000000000",
  530=>"111111111",
  531=>"000000001",
  532=>"000001100",
  533=>"110111111",
  534=>"111000000",
  535=>"001001001",
  536=>"001000000",
  537=>"000000000",
  538=>"000001111",
  539=>"111111111",
  540=>"111111111",
  541=>"111111111",
  542=>"111111111",
  543=>"100100100",
  544=>"000000001",
  545=>"110000000",
  546=>"111110111",
  547=>"111000101",
  548=>"000000111",
  549=>"111111111",
  550=>"000000000",
  551=>"111111101",
  552=>"000010111",
  553=>"000000000",
  554=>"000001111",
  555=>"111111111",
  556=>"111111111",
  557=>"000100100",
  558=>"111100000",
  559=>"111100000",
  560=>"011101101",
  561=>"111111111",
  562=>"111001011",
  563=>"111111111",
  564=>"000110110",
  565=>"111111111",
  566=>"000000000",
  567=>"000111100",
  568=>"111111111",
  569=>"111000000",
  570=>"000000000",
  571=>"000000000",
  572=>"000000000",
  573=>"111100100",
  574=>"111111110",
  575=>"000000100",
  576=>"111111000",
  577=>"111111111",
  578=>"000000000",
  579=>"110000011",
  580=>"100000011",
  581=>"110000000",
  582=>"000000000",
  583=>"011111011",
  584=>"000000000",
  585=>"100100100",
  586=>"111111111",
  587=>"111111111",
  588=>"111111111",
  589=>"000000000",
  590=>"010011011",
  591=>"011000001",
  592=>"111100000",
  593=>"111110000",
  594=>"110000011",
  595=>"001010111",
  596=>"000000000",
  597=>"000000000",
  598=>"111111111",
  599=>"000000000",
  600=>"111011011",
  601=>"000000000",
  602=>"111111111",
  603=>"110110110",
  604=>"111111000",
  605=>"001000100",
  606=>"111111001",
  607=>"100000111",
  608=>"010110111",
  609=>"000011011",
  610=>"000001111",
  611=>"000000000",
  612=>"111111111",
  613=>"111110111",
  614=>"111100110",
  615=>"111111111",
  616=>"000000000",
  617=>"111011000",
  618=>"111011111",
  619=>"000111111",
  620=>"111111111",
  621=>"011000000",
  622=>"100000000",
  623=>"111011010",
  624=>"100100110",
  625=>"111000101",
  626=>"111111111",
  627=>"001000000",
  628=>"000100000",
  629=>"000001000",
  630=>"011111111",
  631=>"001000000",
  632=>"000000000",
  633=>"101000111",
  634=>"111011011",
  635=>"000011001",
  636=>"111111111",
  637=>"000000111",
  638=>"111111011",
  639=>"000110111",
  640=>"111111111",
  641=>"000000000",
  642=>"000000000",
  643=>"000111111",
  644=>"111110000",
  645=>"100000101",
  646=>"111100110",
  647=>"000000000",
  648=>"111111111",
  649=>"000000000",
  650=>"001111111",
  651=>"000000111",
  652=>"100110111",
  653=>"000000000",
  654=>"011011111",
  655=>"111111111",
  656=>"000000000",
  657=>"000011010",
  658=>"111001000",
  659=>"111111111",
  660=>"111111000",
  661=>"000000000",
  662=>"111111111",
  663=>"011001111",
  664=>"101110111",
  665=>"111111111",
  666=>"101001001",
  667=>"000111010",
  668=>"000000000",
  669=>"000011111",
  670=>"100011000",
  671=>"000000001",
  672=>"111111011",
  673=>"111000000",
  674=>"111111111",
  675=>"000000000",
  676=>"101111111",
  677=>"000000100",
  678=>"111111000",
  679=>"111111111",
  680=>"110100000",
  681=>"111111111",
  682=>"000010110",
  683=>"111111111",
  684=>"001000000",
  685=>"111111111",
  686=>"000000000",
  687=>"111111111",
  688=>"000000000",
  689=>"000110000",
  690=>"111111111",
  691=>"111011110",
  692=>"000000000",
  693=>"000000000",
  694=>"000111111",
  695=>"000110111",
  696=>"111111111",
  697=>"111111000",
  698=>"000000111",
  699=>"000110111",
  700=>"000000000",
  701=>"110000000",
  702=>"011001011",
  703=>"000000001",
  704=>"111000000",
  705=>"111111111",
  706=>"111001000",
  707=>"111110110",
  708=>"000011111",
  709=>"000000000",
  710=>"111000000",
  711=>"000000000",
  712=>"111110111",
  713=>"111111111",
  714=>"000000100",
  715=>"111010000",
  716=>"111111111",
  717=>"110111111",
  718=>"000000100",
  719=>"000001000",
  720=>"110110000",
  721=>"000000000",
  722=>"000000000",
  723=>"000000000",
  724=>"010000110",
  725=>"100001011",
  726=>"000000000",
  727=>"111000100",
  728=>"111111111",
  729=>"111111111",
  730=>"001101111",
  731=>"111100100",
  732=>"101101111",
  733=>"111111111",
  734=>"000000000",
  735=>"000000000",
  736=>"000000000",
  737=>"000111111",
  738=>"000000000",
  739=>"000000000",
  740=>"000100101",
  741=>"001011111",
  742=>"111111111",
  743=>"111100101",
  744=>"000000000",
  745=>"111100100",
  746=>"111000000",
  747=>"001000000",
  748=>"010000001",
  749=>"111100100",
  750=>"000100101",
  751=>"010000111",
  752=>"000000011",
  753=>"001011001",
  754=>"111011011",
  755=>"000010110",
  756=>"000100111",
  757=>"011101110",
  758=>"111110010",
  759=>"111011111",
  760=>"001000100",
  761=>"111111111",
  762=>"000000100",
  763=>"000000000",
  764=>"101111000",
  765=>"111111100",
  766=>"100000000",
  767=>"010100000",
  768=>"000000000",
  769=>"111111100",
  770=>"110111111",
  771=>"000101011",
  772=>"111000000",
  773=>"111111111",
  774=>"111001001",
  775=>"000001011",
  776=>"111101101",
  777=>"000000000",
  778=>"000000000",
  779=>"111111111",
  780=>"000000000",
  781=>"000000000",
  782=>"111111111",
  783=>"000110011",
  784=>"111000000",
  785=>"000000100",
  786=>"011000000",
  787=>"011000000",
  788=>"011110000",
  789=>"000001000",
  790=>"111011011",
  791=>"011111011",
  792=>"000000001",
  793=>"000000110",
  794=>"000000000",
  795=>"000000000",
  796=>"111111111",
  797=>"001001001",
  798=>"010110010",
  799=>"000000110",
  800=>"111011001",
  801=>"110000000",
  802=>"000100111",
  803=>"111111111",
  804=>"111111111",
  805=>"011111011",
  806=>"111111111",
  807=>"100000101",
  808=>"111111110",
  809=>"111110100",
  810=>"000000000",
  811=>"000111111",
  812=>"110111111",
  813=>"100110110",
  814=>"011011000",
  815=>"001001011",
  816=>"111111111",
  817=>"111001010",
  818=>"111111101",
  819=>"010000000",
  820=>"111111100",
  821=>"111110000",
  822=>"000000000",
  823=>"100110111",
  824=>"111111111",
  825=>"111111001",
  826=>"111111111",
  827=>"010000000",
  828=>"000111000",
  829=>"100000111",
  830=>"111101100",
  831=>"000111001",
  832=>"000000000",
  833=>"111111111",
  834=>"111111111",
  835=>"111111111",
  836=>"111111111",
  837=>"000000110",
  838=>"110111101",
  839=>"111111111",
  840=>"111111111",
  841=>"000000000",
  842=>"111111111",
  843=>"111001111",
  844=>"111111000",
  845=>"000000000",
  846=>"111110011",
  847=>"111111111",
  848=>"111111111",
  849=>"110111111",
  850=>"000000111",
  851=>"011001111",
  852=>"111011000",
  853=>"011011011",
  854=>"000000000",
  855=>"111111110",
  856=>"111111111",
  857=>"111001000",
  858=>"101111000",
  859=>"111000000",
  860=>"111111111",
  861=>"100110100",
  862=>"000000000",
  863=>"001001010",
  864=>"101100100",
  865=>"111111111",
  866=>"111110110",
  867=>"100000000",
  868=>"000000000",
  869=>"111001111",
  870=>"111011011",
  871=>"000100011",
  872=>"110110110",
  873=>"011000111",
  874=>"001000001",
  875=>"111110000",
  876=>"011011110",
  877=>"000010000",
  878=>"111000000",
  879=>"000000111",
  880=>"000000000",
  881=>"111001000",
  882=>"010000100",
  883=>"101111111",
  884=>"001001001",
  885=>"100100100",
  886=>"000000000",
  887=>"111111111",
  888=>"111111110",
  889=>"000000110",
  890=>"111111111",
  891=>"010110111",
  892=>"110001000",
  893=>"101001001",
  894=>"000000000",
  895=>"110000000",
  896=>"111111111",
  897=>"111101000",
  898=>"001001011",
  899=>"000000000",
  900=>"000000000",
  901=>"000000000",
  902=>"000010111",
  903=>"000000000",
  904=>"111001111",
  905=>"000000000",
  906=>"001111111",
  907=>"100000100",
  908=>"111111111",
  909=>"101000000",
  910=>"111000101",
  911=>"000000000",
  912=>"111111000",
  913=>"101000000",
  914=>"000000000",
  915=>"000111010",
  916=>"101000000",
  917=>"000010010",
  918=>"111111111",
  919=>"111111111",
  920=>"000000010",
  921=>"000111001",
  922=>"111111111",
  923=>"000000111",
  924=>"001111111",
  925=>"000000000",
  926=>"011000110",
  927=>"000000000",
  928=>"000011011",
  929=>"111111111",
  930=>"001000011",
  931=>"000000100",
  932=>"000000000",
  933=>"000000000",
  934=>"111011010",
  935=>"000000000",
  936=>"000001011",
  937=>"100100110",
  938=>"111100000",
  939=>"001010000",
  940=>"001000000",
  941=>"011000000",
  942=>"000000000",
  943=>"111111111",
  944=>"111110111",
  945=>"111111111",
  946=>"000000000",
  947=>"010010111",
  948=>"111111000",
  949=>"100100110",
  950=>"111111111",
  951=>"000001111",
  952=>"111000000",
  953=>"000000000",
  954=>"010000000",
  955=>"111111101",
  956=>"111111111",
  957=>"111111111",
  958=>"000000000",
  959=>"001011111",
  960=>"111000100",
  961=>"111111110",
  962=>"011001111",
  963=>"000000000",
  964=>"111000101",
  965=>"001000001",
  966=>"000010000",
  967=>"000000000",
  968=>"111000000",
  969=>"000000111",
  970=>"111111111",
  971=>"111110110",
  972=>"000000000",
  973=>"111111011",
  974=>"000000000",
  975=>"111111101",
  976=>"111111111",
  977=>"111000000",
  978=>"110000000",
  979=>"101111111",
  980=>"011011011",
  981=>"110111111",
  982=>"000100111",
  983=>"011001001",
  984=>"111111111",
  985=>"000000000",
  986=>"000000000",
  987=>"000000100",
  988=>"000001011",
  989=>"000000000",
  990=>"000111011",
  991=>"110100110",
  992=>"111111111",
  993=>"001101000",
  994=>"000110011",
  995=>"000000001",
  996=>"111100100",
  997=>"000000000",
  998=>"000000000",
  999=>"111111111",
  1000=>"111110110",
  1001=>"000000000",
  1002=>"000000000",
  1003=>"111001100",
  1004=>"000000000",
  1005=>"111111011",
  1006=>"000000000",
  1007=>"111110000",
  1008=>"000000100",
  1009=>"011011111",
  1010=>"000001001",
  1011=>"111111010",
  1012=>"111011000",
  1013=>"000000000",
  1014=>"110110111",
  1015=>"000000000",
  1016=>"111111111",
  1017=>"111101111",
  1018=>"110010000",
  1019=>"111111000",
  1020=>"111100111",
  1021=>"011001100",
  1022=>"111111111",
  1023=>"111111110",
  1024=>"010111111",
  1025=>"111111111",
  1026=>"000000000",
  1027=>"101100000",
  1028=>"000000000",
  1029=>"111001101",
  1030=>"000000000",
  1031=>"101000001",
  1032=>"111111111",
  1033=>"000000000",
  1034=>"010111010",
  1035=>"111111101",
  1036=>"110110110",
  1037=>"111111110",
  1038=>"100111111",
  1039=>"000000000",
  1040=>"111111111",
  1041=>"000011111",
  1042=>"111111001",
  1043=>"111111111",
  1044=>"000000000",
  1045=>"110110100",
  1046=>"000000000",
  1047=>"000000000",
  1048=>"000000000",
  1049=>"000100101",
  1050=>"111111111",
  1051=>"110100110",
  1052=>"000000111",
  1053=>"111111110",
  1054=>"111111111",
  1055=>"000000111",
  1056=>"101001111",
  1057=>"110110110",
  1058=>"110110110",
  1059=>"000000000",
  1060=>"000000111",
  1061=>"111000001",
  1062=>"010001101",
  1063=>"000000000",
  1064=>"000000111",
  1065=>"000000000",
  1066=>"011001110",
  1067=>"111111111",
  1068=>"111111000",
  1069=>"000011011",
  1070=>"001001001",
  1071=>"111011011",
  1072=>"111111111",
  1073=>"111011000",
  1074=>"000100000",
  1075=>"000000000",
  1076=>"101001000",
  1077=>"110111110",
  1078=>"111101000",
  1079=>"111001000",
  1080=>"111111000",
  1081=>"011000000",
  1082=>"111111111",
  1083=>"000000000",
  1084=>"000000010",
  1085=>"000000000",
  1086=>"000110110",
  1087=>"111111000",
  1088=>"011001000",
  1089=>"001001111",
  1090=>"001000000",
  1091=>"000000000",
  1092=>"000000000",
  1093=>"000000000",
  1094=>"000000111",
  1095=>"111111111",
  1096=>"111111011",
  1097=>"000000111",
  1098=>"111111100",
  1099=>"101011111",
  1100=>"111101111",
  1101=>"001101101",
  1102=>"000011110",
  1103=>"000000000",
  1104=>"000000000",
  1105=>"111111000",
  1106=>"000000111",
  1107=>"011011100",
  1108=>"000000000",
  1109=>"000001001",
  1110=>"000101110",
  1111=>"011111000",
  1112=>"111111111",
  1113=>"101000000",
  1114=>"000000000",
  1115=>"000000000",
  1116=>"111111111",
  1117=>"000000000",
  1118=>"000000001",
  1119=>"011001100",
  1120=>"111000100",
  1121=>"011111000",
  1122=>"100111111",
  1123=>"000000000",
  1124=>"110110000",
  1125=>"000000000",
  1126=>"000100111",
  1127=>"111111111",
  1128=>"100111111",
  1129=>"010111101",
  1130=>"111010110",
  1131=>"000000000",
  1132=>"100000000",
  1133=>"000000000",
  1134=>"000000000",
  1135=>"001001000",
  1136=>"000000011",
  1137=>"101111000",
  1138=>"111111111",
  1139=>"111111111",
  1140=>"111111111",
  1141=>"010010000",
  1142=>"000000000",
  1143=>"011111001",
  1144=>"011111111",
  1145=>"111101000",
  1146=>"111111010",
  1147=>"000000111",
  1148=>"100100110",
  1149=>"001000000",
  1150=>"000000000",
  1151=>"001011011",
  1152=>"000000000",
  1153=>"111001111",
  1154=>"110111111",
  1155=>"011011000",
  1156=>"111111000",
  1157=>"000000111",
  1158=>"110110111",
  1159=>"000101111",
  1160=>"000110110",
  1161=>"010110000",
  1162=>"100111001",
  1163=>"010111111",
  1164=>"000000000",
  1165=>"000000001",
  1166=>"000000000",
  1167=>"111111111",
  1168=>"000000001",
  1169=>"000000000",
  1170=>"000000001",
  1171=>"000000111",
  1172=>"111111111",
  1173=>"000000000",
  1174=>"000111110",
  1175=>"111111111",
  1176=>"001000000",
  1177=>"000000000",
  1178=>"111111011",
  1179=>"111000000",
  1180=>"111110111",
  1181=>"000001101",
  1182=>"000100111",
  1183=>"111111111",
  1184=>"001000101",
  1185=>"000011110",
  1186=>"001001111",
  1187=>"111111111",
  1188=>"000001001",
  1189=>"001000000",
  1190=>"111001111",
  1191=>"111010000",
  1192=>"000000111",
  1193=>"000000000",
  1194=>"000000000",
  1195=>"110000111",
  1196=>"111110000",
  1197=>"111101111",
  1198=>"100100101",
  1199=>"000100000",
  1200=>"111000000",
  1201=>"000000000",
  1202=>"110110010",
  1203=>"100101111",
  1204=>"100110011",
  1205=>"111111011",
  1206=>"000000000",
  1207=>"111111010",
  1208=>"000000000",
  1209=>"110000000",
  1210=>"101000000",
  1211=>"110100111",
  1212=>"000000000",
  1213=>"001001101",
  1214=>"111111111",
  1215=>"011111001",
  1216=>"100100000",
  1217=>"110000100",
  1218=>"000000000",
  1219=>"111111111",
  1220=>"010111111",
  1221=>"011011000",
  1222=>"000111011",
  1223=>"101101111",
  1224=>"011010010",
  1225=>"000000000",
  1226=>"000000000",
  1227=>"000000000",
  1228=>"111111111",
  1229=>"000110111",
  1230=>"000000000",
  1231=>"000101111",
  1232=>"001001000",
  1233=>"111001000",
  1234=>"000000000",
  1235=>"011111010",
  1236=>"000000000",
  1237=>"110000001",
  1238=>"000100111",
  1239=>"000000101",
  1240=>"001000000",
  1241=>"110110110",
  1242=>"000000111",
  1243=>"000011111",
  1244=>"111111101",
  1245=>"110000000",
  1246=>"000000000",
  1247=>"000000111",
  1248=>"111111011",
  1249=>"000000011",
  1250=>"111111000",
  1251=>"110000011",
  1252=>"111111111",
  1253=>"000000100",
  1254=>"111111111",
  1255=>"111111111",
  1256=>"111111010",
  1257=>"111111111",
  1258=>"001011001",
  1259=>"000010000",
  1260=>"011000000",
  1261=>"101111111",
  1262=>"000000111",
  1263=>"000110111",
  1264=>"000001101",
  1265=>"010000000",
  1266=>"111111111",
  1267=>"101101111",
  1268=>"111111111",
  1269=>"110110101",
  1270=>"000100111",
  1271=>"001111000",
  1272=>"111111110",
  1273=>"000000100",
  1274=>"111101000",
  1275=>"000000100",
  1276=>"000100000",
  1277=>"111111110",
  1278=>"000000000",
  1279=>"111111111",
  1280=>"000000000",
  1281=>"000010001",
  1282=>"000000000",
  1283=>"010111111",
  1284=>"100000000",
  1285=>"100111110",
  1286=>"111101000",
  1287=>"111000100",
  1288=>"011001000",
  1289=>"000000000",
  1290=>"000101111",
  1291=>"000000111",
  1292=>"110100100",
  1293=>"100000000",
  1294=>"000000111",
  1295=>"000111111",
  1296=>"111000101",
  1297=>"011111000",
  1298=>"100000000",
  1299=>"000000001",
  1300=>"010000001",
  1301=>"000000000",
  1302=>"110100100",
  1303=>"011111111",
  1304=>"100001000",
  1305=>"000000100",
  1306=>"111111000",
  1307=>"010110110",
  1308=>"110111110",
  1309=>"000000100",
  1310=>"011001000",
  1311=>"000000111",
  1312=>"000110111",
  1313=>"110001001",
  1314=>"100000000",
  1315=>"111001000",
  1316=>"000001111",
  1317=>"000000000",
  1318=>"010010111",
  1319=>"001111000",
  1320=>"110111110",
  1321=>"111111111",
  1322=>"000000000",
  1323=>"000000111",
  1324=>"000000001",
  1325=>"000000000",
  1326=>"111000010",
  1327=>"000000000",
  1328=>"111111010",
  1329=>"111111111",
  1330=>"111111111",
  1331=>"001000000",
  1332=>"011101111",
  1333=>"111111111",
  1334=>"111111111",
  1335=>"000000000",
  1336=>"000000000",
  1337=>"111111101",
  1338=>"001110111",
  1339=>"111111111",
  1340=>"001000100",
  1341=>"000000111",
  1342=>"000100110",
  1343=>"000000101",
  1344=>"000000000",
  1345=>"000000000",
  1346=>"000000001",
  1347=>"111110110",
  1348=>"001001111",
  1349=>"011000000",
  1350=>"110110000",
  1351=>"000001111",
  1352=>"000000000",
  1353=>"111110010",
  1354=>"001001000",
  1355=>"111100100",
  1356=>"111110000",
  1357=>"111110000",
  1358=>"101101111",
  1359=>"010011111",
  1360=>"011000010",
  1361=>"101100000",
  1362=>"000000000",
  1363=>"111101111",
  1364=>"100000000",
  1365=>"001011011",
  1366=>"000000111",
  1367=>"111111100",
  1368=>"111001001",
  1369=>"000000101",
  1370=>"000001111",
  1371=>"101101111",
  1372=>"110101111",
  1373=>"000000000",
  1374=>"001111111",
  1375=>"110101100",
  1376=>"000111111",
  1377=>"111111110",
  1378=>"101110110",
  1379=>"111100101",
  1380=>"101100000",
  1381=>"000000000",
  1382=>"000000000",
  1383=>"000000011",
  1384=>"110111110",
  1385=>"000001011",
  1386=>"111001000",
  1387=>"100110110",
  1388=>"000011111",
  1389=>"000000111",
  1390=>"111111111",
  1391=>"111100000",
  1392=>"000000001",
  1393=>"001011011",
  1394=>"000010111",
  1395=>"011000000",
  1396=>"111000000",
  1397=>"000000000",
  1398=>"001001111",
  1399=>"110010000",
  1400=>"000000000",
  1401=>"101101000",
  1402=>"000000011",
  1403=>"111111110",
  1404=>"111111011",
  1405=>"001111001",
  1406=>"000000000",
  1407=>"010111110",
  1408=>"100000001",
  1409=>"110100000",
  1410=>"000000000",
  1411=>"000000010",
  1412=>"000010110",
  1413=>"111111111",
  1414=>"111111111",
  1415=>"111111111",
  1416=>"000000111",
  1417=>"001000000",
  1418=>"111111111",
  1419=>"111111111",
  1420=>"111111101",
  1421=>"110110000",
  1422=>"000111111",
  1423=>"000000000",
  1424=>"000000100",
  1425=>"001000111",
  1426=>"001000011",
  1427=>"000110110",
  1428=>"101100111",
  1429=>"000000000",
  1430=>"010011011",
  1431=>"000001001",
  1432=>"111111111",
  1433=>"001000000",
  1434=>"111111111",
  1435=>"111011111",
  1436=>"000000000",
  1437=>"110110000",
  1438=>"111001000",
  1439=>"111111000",
  1440=>"000000000",
  1441=>"111111111",
  1442=>"000000111",
  1443=>"001001101",
  1444=>"000101101",
  1445=>"111111110",
  1446=>"001000111",
  1447=>"000011011",
  1448=>"011011000",
  1449=>"001101111",
  1450=>"000000000",
  1451=>"000000000",
  1452=>"111110100",
  1453=>"111100100",
  1454=>"000000000",
  1455=>"000000000",
  1456=>"010001101",
  1457=>"000000000",
  1458=>"111110111",
  1459=>"100000000",
  1460=>"111101100",
  1461=>"111111000",
  1462=>"111101111",
  1463=>"000000000",
  1464=>"000000111",
  1465=>"011111011",
  1466=>"000000000",
  1467=>"101000000",
  1468=>"100000000",
  1469=>"100000000",
  1470=>"111110100",
  1471=>"111110100",
  1472=>"111111010",
  1473=>"000000000",
  1474=>"000010000",
  1475=>"111111101",
  1476=>"000110100",
  1477=>"100000000",
  1478=>"101101111",
  1479=>"000111111",
  1480=>"000000001",
  1481=>"111100000",
  1482=>"001000000",
  1483=>"000000000",
  1484=>"100001111",
  1485=>"111111111",
  1486=>"111101111",
  1487=>"111110110",
  1488=>"000110111",
  1489=>"000000000",
  1490=>"111101101",
  1491=>"000000011",
  1492=>"000000000",
  1493=>"111111111",
  1494=>"111101001",
  1495=>"011111011",
  1496=>"110000000",
  1497=>"000000000",
  1498=>"000000110",
  1499=>"101100100",
  1500=>"101111101",
  1501=>"001000100",
  1502=>"000100101",
  1503=>"000000000",
  1504=>"111011000",
  1505=>"011111111",
  1506=>"001000110",
  1507=>"111111000",
  1508=>"010110111",
  1509=>"000100000",
  1510=>"111111000",
  1511=>"000000000",
  1512=>"000000000",
  1513=>"110111111",
  1514=>"011111111",
  1515=>"010111111",
  1516=>"111111111",
  1517=>"000000100",
  1518=>"000000111",
  1519=>"000000000",
  1520=>"000000000",
  1521=>"000000000",
  1522=>"111111011",
  1523=>"111111111",
  1524=>"001110110",
  1525=>"111111110",
  1526=>"101111111",
  1527=>"000110111",
  1528=>"011111000",
  1529=>"000000000",
  1530=>"001000000",
  1531=>"100000111",
  1532=>"000001000",
  1533=>"000100111",
  1534=>"111111111",
  1535=>"111111111",
  1536=>"000000000",
  1537=>"111111111",
  1538=>"000001111",
  1539=>"001001100",
  1540=>"100100000",
  1541=>"001001001",
  1542=>"001001001",
  1543=>"101001101",
  1544=>"000000111",
  1545=>"110110000",
  1546=>"111101000",
  1547=>"000010011",
  1548=>"111011110",
  1549=>"000011111",
  1550=>"000000111",
  1551=>"101100110",
  1552=>"000000100",
  1553=>"000000000",
  1554=>"111110110",
  1555=>"100001000",
  1556=>"001000000",
  1557=>"100111100",
  1558=>"011011011",
  1559=>"001001011",
  1560=>"111111001",
  1561=>"111111110",
  1562=>"100101111",
  1563=>"001001000",
  1564=>"000000000",
  1565=>"111110010",
  1566=>"101111101",
  1567=>"111111111",
  1568=>"100001000",
  1569=>"011000000",
  1570=>"111100101",
  1571=>"000000000",
  1572=>"111111111",
  1573=>"111110011",
  1574=>"111001111",
  1575=>"011000110",
  1576=>"011011111",
  1577=>"000000000",
  1578=>"101101111",
  1579=>"110110000",
  1580=>"111000101",
  1581=>"111111111",
  1582=>"011000000",
  1583=>"110111110",
  1584=>"101111000",
  1585=>"000111000",
  1586=>"011010000",
  1587=>"000000000",
  1588=>"010010000",
  1589=>"000000111",
  1590=>"100000000",
  1591=>"111111110",
  1592=>"000000110",
  1593=>"010010010",
  1594=>"000111111",
  1595=>"111000000",
  1596=>"111111111",
  1597=>"111011011",
  1598=>"111100000",
  1599=>"000000101",
  1600=>"000110110",
  1601=>"000001111",
  1602=>"111000000",
  1603=>"011000000",
  1604=>"010111000",
  1605=>"000000000",
  1606=>"111110100",
  1607=>"111110110",
  1608=>"011111011",
  1609=>"111000000",
  1610=>"111111111",
  1611=>"000000000",
  1612=>"111000000",
  1613=>"011111110",
  1614=>"010010111",
  1615=>"100111011",
  1616=>"000000000",
  1617=>"110110000",
  1618=>"011011000",
  1619=>"000001000",
  1620=>"000000000",
  1621=>"110000111",
  1622=>"000000100",
  1623=>"101101111",
  1624=>"110011000",
  1625=>"101101111",
  1626=>"000000111",
  1627=>"100110000",
  1628=>"000000000",
  1629=>"111110010",
  1630=>"111111111",
  1631=>"000111110",
  1632=>"000111111",
  1633=>"000000000",
  1634=>"010010010",
  1635=>"001001111",
  1636=>"111111110",
  1637=>"111111111",
  1638=>"111111000",
  1639=>"011111111",
  1640=>"001000111",
  1641=>"001111111",
  1642=>"101000000",
  1643=>"110110001",
  1644=>"111111100",
  1645=>"000000000",
  1646=>"010110000",
  1647=>"110110000",
  1648=>"011000010",
  1649=>"000000111",
  1650=>"000010000",
  1651=>"010111111",
  1652=>"000000001",
  1653=>"000000000",
  1654=>"111111111",
  1655=>"010010010",
  1656=>"001000000",
  1657=>"001000000",
  1658=>"101101000",
  1659=>"000000000",
  1660=>"110110100",
  1661=>"110110000",
  1662=>"001001000",
  1663=>"111111111",
  1664=>"111111111",
  1665=>"111100100",
  1666=>"000110111",
  1667=>"000100110",
  1668=>"010010110",
  1669=>"000001111",
  1670=>"111110110",
  1671=>"110010000",
  1672=>"111001101",
  1673=>"111001000",
  1674=>"000001101",
  1675=>"100111111",
  1676=>"000010010",
  1677=>"011000000",
  1678=>"000000001",
  1679=>"111110000",
  1680=>"111111111",
  1681=>"000000000",
  1682=>"000010110",
  1683=>"110110000",
  1684=>"111011111",
  1685=>"111111101",
  1686=>"101111111",
  1687=>"111111100",
  1688=>"011011000",
  1689=>"100000000",
  1690=>"001011000",
  1691=>"111000001",
  1692=>"111111011",
  1693=>"000100110",
  1694=>"001000000",
  1695=>"111000011",
  1696=>"000111111",
  1697=>"111111111",
  1698=>"000001101",
  1699=>"011111110",
  1700=>"000000110",
  1701=>"111111111",
  1702=>"110111111",
  1703=>"011111000",
  1704=>"001001101",
  1705=>"000010010",
  1706=>"011000111",
  1707=>"000000100",
  1708=>"111111111",
  1709=>"111111111",
  1710=>"111111111",
  1711=>"011111110",
  1712=>"011111000",
  1713=>"111111111",
  1714=>"110110110",
  1715=>"111111111",
  1716=>"001001111",
  1717=>"000000000",
  1718=>"010000110",
  1719=>"000000001",
  1720=>"111000100",
  1721=>"111111111",
  1722=>"001101101",
  1723=>"111111011",
  1724=>"000000000",
  1725=>"010000001",
  1726=>"100101000",
  1727=>"010111111",
  1728=>"001000100",
  1729=>"111101000",
  1730=>"110000000",
  1731=>"110000000",
  1732=>"111111000",
  1733=>"111111111",
  1734=>"011001000",
  1735=>"010010110",
  1736=>"000011110",
  1737=>"000000100",
  1738=>"000000010",
  1739=>"110000000",
  1740=>"000000100",
  1741=>"000000110",
  1742=>"000000111",
  1743=>"001001101",
  1744=>"000111111",
  1745=>"000010111",
  1746=>"010000000",
  1747=>"111001111",
  1748=>"010111110",
  1749=>"000000000",
  1750=>"000000111",
  1751=>"111111111",
  1752=>"111111000",
  1753=>"111110111",
  1754=>"000000000",
  1755=>"110011111",
  1756=>"001001111",
  1757=>"000110100",
  1758=>"000010000",
  1759=>"000000010",
  1760=>"000000000",
  1761=>"000000000",
  1762=>"000100111",
  1763=>"111111111",
  1764=>"000001011",
  1765=>"001001001",
  1766=>"011110111",
  1767=>"111111100",
  1768=>"000000011",
  1769=>"000000111",
  1770=>"000100000",
  1771=>"100100100",
  1772=>"000000010",
  1773=>"000000010",
  1774=>"010110111",
  1775=>"011110000",
  1776=>"101111111",
  1777=>"111111100",
  1778=>"000001001",
  1779=>"000000000",
  1780=>"000011001",
  1781=>"101110000",
  1782=>"000000010",
  1783=>"111010000",
  1784=>"001011111",
  1785=>"111101000",
  1786=>"001001001",
  1787=>"000000100",
  1788=>"000000000",
  1789=>"111111111",
  1790=>"110110000",
  1791=>"110011001",
  1792=>"111111111",
  1793=>"100100000",
  1794=>"100000111",
  1795=>"010010000",
  1796=>"001001001",
  1797=>"001010100",
  1798=>"000000000",
  1799=>"010000001",
  1800=>"111001000",
  1801=>"111111000",
  1802=>"001000000",
  1803=>"111110111",
  1804=>"000000001",
  1805=>"010000110",
  1806=>"111111111",
  1807=>"111111111",
  1808=>"111111001",
  1809=>"000000000",
  1810=>"000010000",
  1811=>"000000111",
  1812=>"000101101",
  1813=>"000000000",
  1814=>"000110111",
  1815=>"111111111",
  1816=>"001001000",
  1817=>"000000111",
  1818=>"111111111",
  1819=>"011111010",
  1820=>"001001000",
  1821=>"110000000",
  1822=>"000000000",
  1823=>"000000000",
  1824=>"111111111",
  1825=>"111111111",
  1826=>"101111111",
  1827=>"011010100",
  1828=>"111011111",
  1829=>"000010000",
  1830=>"110111001",
  1831=>"111111011",
  1832=>"111111111",
  1833=>"110000000",
  1834=>"000101000",
  1835=>"000000000",
  1836=>"111000000",
  1837=>"100100101",
  1838=>"111111010",
  1839=>"011000100",
  1840=>"000000000",
  1841=>"111111000",
  1842=>"111101111",
  1843=>"001000000",
  1844=>"111101111",
  1845=>"111000000",
  1846=>"011111111",
  1847=>"111000001",
  1848=>"110111011",
  1849=>"101001011",
  1850=>"000111111",
  1851=>"000000100",
  1852=>"000000011",
  1853=>"101001000",
  1854=>"000110010",
  1855=>"111111111",
  1856=>"001001111",
  1857=>"000111111",
  1858=>"111111001",
  1859=>"001101111",
  1860=>"000000111",
  1861=>"000000111",
  1862=>"000000000",
  1863=>"111111111",
  1864=>"000000000",
  1865=>"111111111",
  1866=>"100100000",
  1867=>"000000110",
  1868=>"111111111",
  1869=>"111110111",
  1870=>"000000000",
  1871=>"001011011",
  1872=>"001001111",
  1873=>"000000111",
  1874=>"110110111",
  1875=>"010110110",
  1876=>"100001000",
  1877=>"001001001",
  1878=>"110010110",
  1879=>"110110000",
  1880=>"111111110",
  1881=>"111111111",
  1882=>"111110111",
  1883=>"111001001",
  1884=>"111111111",
  1885=>"000000100",
  1886=>"010110000",
  1887=>"001001001",
  1888=>"111111000",
  1889=>"000000110",
  1890=>"001111111",
  1891=>"110001001",
  1892=>"100100110",
  1893=>"000000000",
  1894=>"000100110",
  1895=>"111111000",
  1896=>"001101111",
  1897=>"000000111",
  1898=>"111100110",
  1899=>"110111111",
  1900=>"000000000",
  1901=>"000000111",
  1902=>"111011111",
  1903=>"000000000",
  1904=>"000000110",
  1905=>"010010000",
  1906=>"111010110",
  1907=>"111100111",
  1908=>"011011000",
  1909=>"000000111",
  1910=>"000010111",
  1911=>"111010001",
  1912=>"001000101",
  1913=>"000000000",
  1914=>"011000000",
  1915=>"000111111",
  1916=>"111111000",
  1917=>"111111110",
  1918=>"000011001",
  1919=>"111111000",
  1920=>"111111001",
  1921=>"111111110",
  1922=>"001000100",
  1923=>"001001101",
  1924=>"000000000",
  1925=>"000100110",
  1926=>"001001000",
  1927=>"111001100",
  1928=>"011010000",
  1929=>"000100000",
  1930=>"100000000",
  1931=>"001101111",
  1932=>"111111111",
  1933=>"111110110",
  1934=>"111110000",
  1935=>"100100100",
  1936=>"000100000",
  1937=>"111110111",
  1938=>"011001010",
  1939=>"000000000",
  1940=>"111101001",
  1941=>"000000010",
  1942=>"011011110",
  1943=>"001001111",
  1944=>"111000010",
  1945=>"001000111",
  1946=>"111111101",
  1947=>"111100100",
  1948=>"111111111",
  1949=>"010010010",
  1950=>"000011111",
  1951=>"111001000",
  1952=>"000000000",
  1953=>"000111111",
  1954=>"000000001",
  1955=>"000111001",
  1956=>"111111001",
  1957=>"001111111",
  1958=>"011111111",
  1959=>"000110111",
  1960=>"011011111",
  1961=>"000011111",
  1962=>"110010111",
  1963=>"001001000",
  1964=>"000100100",
  1965=>"110111111",
  1966=>"000001111",
  1967=>"111011011",
  1968=>"111100111",
  1969=>"111111100",
  1970=>"111111000",
  1971=>"101111111",
  1972=>"110111010",
  1973=>"111111111",
  1974=>"111100000",
  1975=>"101100000",
  1976=>"011001111",
  1977=>"110110111",
  1978=>"111111101",
  1979=>"000110000",
  1980=>"001001101",
  1981=>"111001111",
  1982=>"111111111",
  1983=>"101101111",
  1984=>"110111111",
  1985=>"001000000",
  1986=>"111000001",
  1987=>"011000010",
  1988=>"000001111",
  1989=>"100000001",
  1990=>"111000000",
  1991=>"000000111",
  1992=>"000000001",
  1993=>"111111000",
  1994=>"101111110",
  1995=>"111111000",
  1996=>"111111001",
  1997=>"110000000",
  1998=>"011011110",
  1999=>"111111111",
  2000=>"001011011",
  2001=>"000001001",
  2002=>"011111111",
  2003=>"000000000",
  2004=>"000100101",
  2005=>"011111101",
  2006=>"011000011",
  2007=>"000000000",
  2008=>"101110110",
  2009=>"000000100",
  2010=>"000111111",
  2011=>"000000011",
  2012=>"111110000",
  2013=>"000000101",
  2014=>"000000001",
  2015=>"001000000",
  2016=>"000000111",
  2017=>"111110111",
  2018=>"101101001",
  2019=>"000000000",
  2020=>"011010111",
  2021=>"001000111",
  2022=>"110111111",
  2023=>"000010000",
  2024=>"000000000",
  2025=>"111000000",
  2026=>"000000100",
  2027=>"000000111",
  2028=>"000000000",
  2029=>"000001001",
  2030=>"000000111",
  2031=>"000000000",
  2032=>"111111111",
  2033=>"111110100",
  2034=>"110111010",
  2035=>"000000110",
  2036=>"010010110",
  2037=>"000110101",
  2038=>"111011000",
  2039=>"111111111",
  2040=>"011011111",
  2041=>"101111110",
  2042=>"111111010",
  2043=>"110111111",
  2044=>"110110111",
  2045=>"000110110",
  2046=>"111010000",
  2047=>"111111111",
  2048=>"111010000",
  2049=>"111110000",
  2050=>"000110000",
  2051=>"100101000",
  2052=>"111111111",
  2053=>"110110100",
  2054=>"000000000",
  2055=>"000000000",
  2056=>"000000100",
  2057=>"001111001",
  2058=>"111111000",
  2059=>"011010000",
  2060=>"110110111",
  2061=>"111111001",
  2062=>"111000000",
  2063=>"111111011",
  2064=>"110111110",
  2065=>"111111111",
  2066=>"000000000",
  2067=>"000010010",
  2068=>"000000001",
  2069=>"000000000",
  2070=>"000000011",
  2071=>"111111111",
  2072=>"000000110",
  2073=>"000000000",
  2074=>"111111111",
  2075=>"011000000",
  2076=>"111111111",
  2077=>"111111011",
  2078=>"000000011",
  2079=>"001000000",
  2080=>"000000000",
  2081=>"100110000",
  2082=>"110000011",
  2083=>"111000111",
  2084=>"011000000",
  2085=>"000001001",
  2086=>"000000000",
  2087=>"000000111",
  2088=>"000111111",
  2089=>"000110110",
  2090=>"000000000",
  2091=>"000000001",
  2092=>"000000101",
  2093=>"000111111",
  2094=>"111000000",
  2095=>"010010110",
  2096=>"100000000",
  2097=>"000000110",
  2098=>"011011011",
  2099=>"000000011",
  2100=>"000000000",
  2101=>"001011111",
  2102=>"010000101",
  2103=>"010101101",
  2104=>"111111111",
  2105=>"111111001",
  2106=>"000000000",
  2107=>"111111111",
  2108=>"001000001",
  2109=>"111111110",
  2110=>"111111111",
  2111=>"111111110",
  2112=>"111000101",
  2113=>"011111110",
  2114=>"001000000",
  2115=>"111111000",
  2116=>"100000000",
  2117=>"011111111",
  2118=>"111111000",
  2119=>"000100000",
  2120=>"011001111",
  2121=>"111111111",
  2122=>"000000000",
  2123=>"111000101",
  2124=>"111111111",
  2125=>"001000000",
  2126=>"111111101",
  2127=>"000000000",
  2128=>"010000000",
  2129=>"000000111",
  2130=>"000111000",
  2131=>"000000000",
  2132=>"111100110",
  2133=>"000000000",
  2134=>"111011111",
  2135=>"000000011",
  2136=>"000000001",
  2137=>"111100111",
  2138=>"000010111",
  2139=>"000100110",
  2140=>"000000001",
  2141=>"001011000",
  2142=>"111100000",
  2143=>"000010000",
  2144=>"000000000",
  2145=>"111111111",
  2146=>"111000100",
  2147=>"000000000",
  2148=>"001000000",
  2149=>"000000001",
  2150=>"000000000",
  2151=>"000000000",
  2152=>"111101000",
  2153=>"111010000",
  2154=>"000000000",
  2155=>"000000001",
  2156=>"000000101",
  2157=>"111111011",
  2158=>"110110110",
  2159=>"000111110",
  2160=>"000000000",
  2161=>"000000110",
  2162=>"000110110",
  2163=>"101111111",
  2164=>"000000001",
  2165=>"000011001",
  2166=>"110111111",
  2167=>"000000000",
  2168=>"000000111",
  2169=>"111101111",
  2170=>"000111111",
  2171=>"000000001",
  2172=>"111101101",
  2173=>"110111111",
  2174=>"011111111",
  2175=>"000000000",
  2176=>"111111111",
  2177=>"111111110",
  2178=>"111000111",
  2179=>"111000000",
  2180=>"001001000",
  2181=>"111001111",
  2182=>"000000011",
  2183=>"111111000",
  2184=>"111111000",
  2185=>"000000000",
  2186=>"100000000",
  2187=>"011000011",
  2188=>"000000000",
  2189=>"000000000",
  2190=>"001001111",
  2191=>"001100100",
  2192=>"001011111",
  2193=>"111011111",
  2194=>"110111111",
  2195=>"110110100",
  2196=>"000000000",
  2197=>"000000000",
  2198=>"000000000",
  2199=>"000000000",
  2200=>"111011111",
  2201=>"000000100",
  2202=>"111001111",
  2203=>"000001000",
  2204=>"000100000",
  2205=>"111000000",
  2206=>"011000111",
  2207=>"110110000",
  2208=>"111101000",
  2209=>"011000000",
  2210=>"001000011",
  2211=>"100100000",
  2212=>"110110110",
  2213=>"000000011",
  2214=>"000000000",
  2215=>"000111011",
  2216=>"111001000",
  2217=>"000000101",
  2218=>"111111111",
  2219=>"000000000",
  2220=>"000000000",
  2221=>"000000011",
  2222=>"111001111",
  2223=>"110000000",
  2224=>"000000000",
  2225=>"000111000",
  2226=>"110111011",
  2227=>"000000000",
  2228=>"000001000",
  2229=>"111101000",
  2230=>"000000000",
  2231=>"001000000",
  2232=>"101001111",
  2233=>"111111000",
  2234=>"111111110",
  2235=>"111111001",
  2236=>"001001111",
  2237=>"000000000",
  2238=>"111111111",
  2239=>"111010110",
  2240=>"000000000",
  2241=>"111111111",
  2242=>"111111110",
  2243=>"000111111",
  2244=>"000111111",
  2245=>"000000110",
  2246=>"010111111",
  2247=>"111000000",
  2248=>"000000000",
  2249=>"111111111",
  2250=>"000000110",
  2251=>"011111010",
  2252=>"101110111",
  2253=>"111100101",
  2254=>"000000100",
  2255=>"000000000",
  2256=>"110110011",
  2257=>"000000001",
  2258=>"101000000",
  2259=>"000010111",
  2260=>"000001111",
  2261=>"011001000",
  2262=>"011111111",
  2263=>"111111111",
  2264=>"000000000",
  2265=>"011010000",
  2266=>"000110100",
  2267=>"000000000",
  2268=>"111011111",
  2269=>"111011111",
  2270=>"000000000",
  2271=>"110011001",
  2272=>"110000000",
  2273=>"001000000",
  2274=>"000000000",
  2275=>"111101000",
  2276=>"111110111",
  2277=>"000100101",
  2278=>"000000000",
  2279=>"111111111",
  2280=>"000000000",
  2281=>"000000000",
  2282=>"111111111",
  2283=>"000111001",
  2284=>"000000000",
  2285=>"010010110",
  2286=>"111111111",
  2287=>"000000000",
  2288=>"101111000",
  2289=>"011010000",
  2290=>"111111111",
  2291=>"111010000",
  2292=>"111111111",
  2293=>"000000000",
  2294=>"011000100",
  2295=>"000000000",
  2296=>"000000000",
  2297=>"000000000",
  2298=>"111111111",
  2299=>"111000100",
  2300=>"000001001",
  2301=>"111011011",
  2302=>"110110000",
  2303=>"111100111",
  2304=>"010000000",
  2305=>"111111011",
  2306=>"000000000",
  2307=>"110111111",
  2308=>"111111000",
  2309=>"000000000",
  2310=>"000000111",
  2311=>"000000000",
  2312=>"000000110",
  2313=>"010010010",
  2314=>"111111111",
  2315=>"111000000",
  2316=>"000001111",
  2317=>"110000000",
  2318=>"110111111",
  2319=>"000000000",
  2320=>"000010000",
  2321=>"110110101",
  2322=>"000000111",
  2323=>"110011000",
  2324=>"000010010",
  2325=>"000001000",
  2326=>"001011001",
  2327=>"000000000",
  2328=>"110000010",
  2329=>"111111111",
  2330=>"110110111",
  2331=>"000100000",
  2332=>"011110111",
  2333=>"100111111",
  2334=>"100000000",
  2335=>"000000000",
  2336=>"000000100",
  2337=>"110111111",
  2338=>"010111111",
  2339=>"001001001",
  2340=>"100100000",
  2341=>"010111100",
  2342=>"111001001",
  2343=>"110010101",
  2344=>"000000000",
  2345=>"000000000",
  2346=>"011000000",
  2347=>"111001111",
  2348=>"111111111",
  2349=>"000000001",
  2350=>"000000000",
  2351=>"000001111",
  2352=>"000000110",
  2353=>"111111111",
  2354=>"000000111",
  2355=>"011111110",
  2356=>"000001011",
  2357=>"111111111",
  2358=>"111111111",
  2359=>"111000000",
  2360=>"111100000",
  2361=>"100000111",
  2362=>"001011111",
  2363=>"111111000",
  2364=>"000001011",
  2365=>"100101111",
  2366=>"111111001",
  2367=>"000000111",
  2368=>"000000111",
  2369=>"111100110",
  2370=>"111111110",
  2371=>"011111111",
  2372=>"111111111",
  2373=>"101111000",
  2374=>"000001011",
  2375=>"010011000",
  2376=>"000000011",
  2377=>"000000000",
  2378=>"000000000",
  2379=>"111011011",
  2380=>"010111100",
  2381=>"000100000",
  2382=>"111010000",
  2383=>"111111001",
  2384=>"011011000",
  2385=>"000010000",
  2386=>"000000111",
  2387=>"000000000",
  2388=>"000000000",
  2389=>"111011011",
  2390=>"000000000",
  2391=>"001001000",
  2392=>"001000111",
  2393=>"111011111",
  2394=>"000000000",
  2395=>"111111111",
  2396=>"111111111",
  2397=>"110000000",
  2398=>"111110111",
  2399=>"111111011",
  2400=>"011001111",
  2401=>"100000000",
  2402=>"011010100",
  2403=>"111111111",
  2404=>"000010110",
  2405=>"000000001",
  2406=>"111110100",
  2407=>"111111111",
  2408=>"000000000",
  2409=>"111111100",
  2410=>"111000000",
  2411=>"111011111",
  2412=>"000000000",
  2413=>"111010000",
  2414=>"000000000",
  2415=>"000000110",
  2416=>"000000000",
  2417=>"111111111",
  2418=>"110010000",
  2419=>"011011000",
  2420=>"000110000",
  2421=>"111110000",
  2422=>"000111111",
  2423=>"111000000",
  2424=>"111111110",
  2425=>"000000110",
  2426=>"000000000",
  2427=>"111111010",
  2428=>"111111000",
  2429=>"111111111",
  2430=>"000000111",
  2431=>"000000000",
  2432=>"000001001",
  2433=>"111111111",
  2434=>"111111111",
  2435=>"000000000",
  2436=>"111111111",
  2437=>"000000001",
  2438=>"000100000",
  2439=>"000000001",
  2440=>"111111111",
  2441=>"111111010",
  2442=>"000010011",
  2443=>"000000000",
  2444=>"111111111",
  2445=>"011011010",
  2446=>"000000100",
  2447=>"000011010",
  2448=>"000010011",
  2449=>"111111111",
  2450=>"000000000",
  2451=>"000000100",
  2452=>"111101100",
  2453=>"000000110",
  2454=>"111111111",
  2455=>"111111111",
  2456=>"000100000",
  2457=>"000000111",
  2458=>"000000111",
  2459=>"000001011",
  2460=>"111111110",
  2461=>"010110010",
  2462=>"100110111",
  2463=>"000000000",
  2464=>"000000000",
  2465=>"001001001",
  2466=>"111000100",
  2467=>"111000110",
  2468=>"001001100",
  2469=>"000000100",
  2470=>"000000011",
  2471=>"100000010",
  2472=>"000000000",
  2473=>"000000000",
  2474=>"111111111",
  2475=>"111011000",
  2476=>"000001111",
  2477=>"011001001",
  2478=>"101000001",
  2479=>"000001111",
  2480=>"111101000",
  2481=>"001000000",
  2482=>"111010000",
  2483=>"001001111",
  2484=>"111111000",
  2485=>"000110111",
  2486=>"111110000",
  2487=>"000000000",
  2488=>"111111111",
  2489=>"000000000",
  2490=>"111000000",
  2491=>"111111111",
  2492=>"001111111",
  2493=>"111111111",
  2494=>"101001101",
  2495=>"010011010",
  2496=>"001011010",
  2497=>"000000000",
  2498=>"001111111",
  2499=>"111111111",
  2500=>"111011111",
  2501=>"001001001",
  2502=>"111001000",
  2503=>"111111111",
  2504=>"110111111",
  2505=>"000000000",
  2506=>"010000100",
  2507=>"111000000",
  2508=>"101110111",
  2509=>"000000000",
  2510=>"000001111",
  2511=>"101101111",
  2512=>"000011011",
  2513=>"000001011",
  2514=>"000000000",
  2515=>"111111111",
  2516=>"000000101",
  2517=>"111111111",
  2518=>"111111001",
  2519=>"111110100",
  2520=>"111000000",
  2521=>"111110110",
  2522=>"111111011",
  2523=>"111111111",
  2524=>"000010010",
  2525=>"100000111",
  2526=>"000000000",
  2527=>"111011011",
  2528=>"111111000",
  2529=>"011001000",
  2530=>"000010111",
  2531=>"000000111",
  2532=>"000010000",
  2533=>"100000000",
  2534=>"000000000",
  2535=>"110110000",
  2536=>"011011000",
  2537=>"000000100",
  2538=>"111011011",
  2539=>"000010111",
  2540=>"110001001",
  2541=>"111100111",
  2542=>"100000000",
  2543=>"000000000",
  2544=>"100111000",
  2545=>"100000111",
  2546=>"111111111",
  2547=>"011000000",
  2548=>"000111111",
  2549=>"001111111",
  2550=>"111111011",
  2551=>"100111111",
  2552=>"001111111",
  2553=>"000000000",
  2554=>"010111000",
  2555=>"111011001",
  2556=>"110110111",
  2557=>"100110100",
  2558=>"111111001",
  2559=>"000000000",
  2560=>"100111111",
  2561=>"000000001",
  2562=>"111101000",
  2563=>"111111110",
  2564=>"000000000",
  2565=>"110000000",
  2566=>"111001000",
  2567=>"000000001",
  2568=>"000111100",
  2569=>"000000000",
  2570=>"000000000",
  2571=>"111011000",
  2572=>"000001011",
  2573=>"000000100",
  2574=>"011011111",
  2575=>"111100110",
  2576=>"101101000",
  2577=>"100111110",
  2578=>"001101111",
  2579=>"111111111",
  2580=>"111101000",
  2581=>"111111000",
  2582=>"000000000",
  2583=>"111110001",
  2584=>"000111111",
  2585=>"111000110",
  2586=>"000000100",
  2587=>"011001000",
  2588=>"000000110",
  2589=>"111111001",
  2590=>"011011011",
  2591=>"000000000",
  2592=>"111111000",
  2593=>"111000000",
  2594=>"111111111",
  2595=>"000101101",
  2596=>"000110111",
  2597=>"111100001",
  2598=>"111000000",
  2599=>"000000011",
  2600=>"001000000",
  2601=>"000000000",
  2602=>"100000000",
  2603=>"000000000",
  2604=>"001101111",
  2605=>"000111111",
  2606=>"100111111",
  2607=>"111111111",
  2608=>"111011111",
  2609=>"000000111",
  2610=>"110110000",
  2611=>"000000000",
  2612=>"111010010",
  2613=>"110110110",
  2614=>"000111110",
  2615=>"111111111",
  2616=>"111111111",
  2617=>"111101111",
  2618=>"000000100",
  2619=>"100000000",
  2620=>"000000000",
  2621=>"001001001",
  2622=>"000001111",
  2623=>"001001111",
  2624=>"001000000",
  2625=>"000001111",
  2626=>"000000001",
  2627=>"111111111",
  2628=>"001011000",
  2629=>"111100100",
  2630=>"100111100",
  2631=>"111111100",
  2632=>"110100100",
  2633=>"000001101",
  2634=>"100111111",
  2635=>"011011000",
  2636=>"000000000",
  2637=>"000000000",
  2638=>"111001000",
  2639=>"000111111",
  2640=>"100000000",
  2641=>"111111000",
  2642=>"000000000",
  2643=>"000000100",
  2644=>"000000000",
  2645=>"000000110",
  2646=>"000100000",
  2647=>"000000000",
  2648=>"111111101",
  2649=>"000100100",
  2650=>"111011000",
  2651=>"100000100",
  2652=>"100100111",
  2653=>"110111111",
  2654=>"100011000",
  2655=>"001111111",
  2656=>"000000110",
  2657=>"000000110",
  2658=>"111111111",
  2659=>"000110111",
  2660=>"000110111",
  2661=>"000000000",
  2662=>"101000000",
  2663=>"000000111",
  2664=>"100000000",
  2665=>"000000000",
  2666=>"110010111",
  2667=>"111011000",
  2668=>"100110110",
  2669=>"111111111",
  2670=>"100100000",
  2671=>"111100000",
  2672=>"110110000",
  2673=>"000011111",
  2674=>"110111110",
  2675=>"000000010",
  2676=>"111111011",
  2677=>"111111100",
  2678=>"000000000",
  2679=>"000000000",
  2680=>"100000010",
  2681=>"110111111",
  2682=>"111111101",
  2683=>"110000000",
  2684=>"000100100",
  2685=>"111111100",
  2686=>"111111000",
  2687=>"111111111",
  2688=>"111100000",
  2689=>"100100110",
  2690=>"111111001",
  2691=>"000000001",
  2692=>"111111111",
  2693=>"000000000",
  2694=>"111111111",
  2695=>"111110000",
  2696=>"111011011",
  2697=>"111111111",
  2698=>"111011011",
  2699=>"111001000",
  2700=>"000111111",
  2701=>"000001000",
  2702=>"100000111",
  2703=>"010111111",
  2704=>"111000000",
  2705=>"111010000",
  2706=>"000110111",
  2707=>"001111111",
  2708=>"111111111",
  2709=>"101000001",
  2710=>"111101000",
  2711=>"110000000",
  2712=>"111000000",
  2713=>"111111110",
  2714=>"111100000",
  2715=>"000001000",
  2716=>"100111111",
  2717=>"000010001",
  2718=>"001111111",
  2719=>"111000000",
  2720=>"111111000",
  2721=>"101001000",
  2722=>"000000001",
  2723=>"101001001",
  2724=>"111001001",
  2725=>"111000000",
  2726=>"010110111",
  2727=>"000000000",
  2728=>"000000000",
  2729=>"110000000",
  2730=>"111111111",
  2731=>"001000000",
  2732=>"001001000",
  2733=>"100000111",
  2734=>"111000000",
  2735=>"111111111",
  2736=>"000100100",
  2737=>"001001001",
  2738=>"111111110",
  2739=>"000000010",
  2740=>"001110111",
  2741=>"111110111",
  2742=>"111000000",
  2743=>"111111111",
  2744=>"010010000",
  2745=>"000000000",
  2746=>"110010110",
  2747=>"000000000",
  2748=>"111010000",
  2749=>"111111011",
  2750=>"100111000",
  2751=>"111111000",
  2752=>"000000111",
  2753=>"111011111",
  2754=>"110111001",
  2755=>"000000011",
  2756=>"000110110",
  2757=>"111111111",
  2758=>"111111001",
  2759=>"000000000",
  2760=>"000000000",
  2761=>"000000011",
  2762=>"000000000",
  2763=>"000000000",
  2764=>"111111011",
  2765=>"100001010",
  2766=>"011111001",
  2767=>"111100000",
  2768=>"000000000",
  2769=>"000000100",
  2770=>"101111111",
  2771=>"000000111",
  2772=>"111111010",
  2773=>"111111110",
  2774=>"000101111",
  2775=>"111110111",
  2776=>"101000001",
  2777=>"111011000",
  2778=>"000001000",
  2779=>"000110111",
  2780=>"110001001",
  2781=>"101111111",
  2782=>"111111111",
  2783=>"110110111",
  2784=>"000010000",
  2785=>"000000101",
  2786=>"000111111",
  2787=>"111111111",
  2788=>"000000000",
  2789=>"111000000",
  2790=>"100000100",
  2791=>"001001101",
  2792=>"000101111",
  2793=>"000110110",
  2794=>"000100100",
  2795=>"100001111",
  2796=>"111111111",
  2797=>"111100100",
  2798=>"111111100",
  2799=>"000000000",
  2800=>"000000000",
  2801=>"111111111",
  2802=>"000001111",
  2803=>"000000011",
  2804=>"000001111",
  2805=>"000110111",
  2806=>"000111011",
  2807=>"000000000",
  2808=>"111011000",
  2809=>"111111001",
  2810=>"000000000",
  2811=>"000000000",
  2812=>"100100000",
  2813=>"001001001",
  2814=>"111001000",
  2815=>"000111111",
  2816=>"100000000",
  2817=>"110111000",
  2818=>"000000000",
  2819=>"111101011",
  2820=>"111111111",
  2821=>"000000100",
  2822=>"000001111",
  2823=>"000111111",
  2824=>"000000000",
  2825=>"000000000",
  2826=>"000000000",
  2827=>"111000000",
  2828=>"111000010",
  2829=>"111001000",
  2830=>"110110100",
  2831=>"110111000",
  2832=>"000000001",
  2833=>"000000000",
  2834=>"000000000",
  2835=>"100111111",
  2836=>"000000000",
  2837=>"000000100",
  2838=>"000111111",
  2839=>"000000001",
  2840=>"111011010",
  2841=>"011011000",
  2842=>"000100110",
  2843=>"111111100",
  2844=>"001011011",
  2845=>"111111111",
  2846=>"011111110",
  2847=>"111001001",
  2848=>"100001000",
  2849=>"011000000",
  2850=>"000110111",
  2851=>"000000110",
  2852=>"111111111",
  2853=>"111111111",
  2854=>"111111111",
  2855=>"111011000",
  2856=>"111111000",
  2857=>"000111111",
  2858=>"000111111",
  2859=>"110111101",
  2860=>"100000000",
  2861=>"001011000",
  2862=>"111110111",
  2863=>"000000000",
  2864=>"000000000",
  2865=>"000000000",
  2866=>"000000000",
  2867=>"011000000",
  2868=>"100000000",
  2869=>"000110111",
  2870=>"000110111",
  2871=>"111111001",
  2872=>"100001001",
  2873=>"111111111",
  2874=>"101001111",
  2875=>"000000001",
  2876=>"111111001",
  2877=>"000000000",
  2878=>"000000000",
  2879=>"110010010",
  2880=>"010100111",
  2881=>"000000000",
  2882=>"001001100",
  2883=>"000000101",
  2884=>"000100111",
  2885=>"111111111",
  2886=>"100100100",
  2887=>"101111111",
  2888=>"110110000",
  2889=>"111111111",
  2890=>"001000000",
  2891=>"011011111",
  2892=>"111101101",
  2893=>"001011011",
  2894=>"000001111",
  2895=>"101111111",
  2896=>"111111110",
  2897=>"000001000",
  2898=>"010000111",
  2899=>"100100111",
  2900=>"001000000",
  2901=>"001001001",
  2902=>"110110000",
  2903=>"000000100",
  2904=>"101001111",
  2905=>"001000111",
  2906=>"000000000",
  2907=>"110000000",
  2908=>"111000111",
  2909=>"010111111",
  2910=>"111111001",
  2911=>"000110110",
  2912=>"111111001",
  2913=>"000000000",
  2914=>"100100010",
  2915=>"100111111",
  2916=>"100111111",
  2917=>"111111111",
  2918=>"110000110",
  2919=>"000111111",
  2920=>"111110111",
  2921=>"111111111",
  2922=>"000000000",
  2923=>"100000000",
  2924=>"001011001",
  2925=>"111111110",
  2926=>"000000000",
  2927=>"110111000",
  2928=>"111111010",
  2929=>"111111111",
  2930=>"111111000",
  2931=>"111111101",
  2932=>"000100111",
  2933=>"000000001",
  2934=>"000000111",
  2935=>"000010000",
  2936=>"111101001",
  2937=>"111111010",
  2938=>"000000000",
  2939=>"111111111",
  2940=>"111000000",
  2941=>"111110000",
  2942=>"000001000",
  2943=>"111111111",
  2944=>"010100000",
  2945=>"111000000",
  2946=>"011001000",
  2947=>"111111000",
  2948=>"101111111",
  2949=>"000000000",
  2950=>"111001000",
  2951=>"000001000",
  2952=>"000000000",
  2953=>"000000001",
  2954=>"000101111",
  2955=>"001001111",
  2956=>"000000111",
  2957=>"111011001",
  2958=>"110111000",
  2959=>"111111011",
  2960=>"111111111",
  2961=>"000000000",
  2962=>"000000000",
  2963=>"111111110",
  2964=>"000000100",
  2965=>"001001000",
  2966=>"000111110",
  2967=>"001000000",
  2968=>"000000100",
  2969=>"111111010",
  2970=>"111111111",
  2971=>"110111111",
  2972=>"111100001",
  2973=>"111111111",
  2974=>"011000000",
  2975=>"000100000",
  2976=>"000000000",
  2977=>"110110001",
  2978=>"011111110",
  2979=>"001001000",
  2980=>"000110111",
  2981=>"000000000",
  2982=>"000001011",
  2983=>"111111111",
  2984=>"000000111",
  2985=>"010111110",
  2986=>"001111111",
  2987=>"101111110",
  2988=>"000111111",
  2989=>"000000000",
  2990=>"111011011",
  2991=>"111111111",
  2992=>"000111010",
  2993=>"100110110",
  2994=>"001011010",
  2995=>"110000110",
  2996=>"111111111",
  2997=>"111111111",
  2998=>"000000000",
  2999=>"111011001",
  3000=>"001011000",
  3001=>"111111111",
  3002=>"111000000",
  3003=>"111111001",
  3004=>"101001101",
  3005=>"000000000",
  3006=>"100000000",
  3007=>"000000000",
  3008=>"111111111",
  3009=>"111011111",
  3010=>"000000000",
  3011=>"000110000",
  3012=>"000011111",
  3013=>"000000110",
  3014=>"000000000",
  3015=>"100111111",
  3016=>"100111101",
  3017=>"000000000",
  3018=>"110011010",
  3019=>"110100100",
  3020=>"000000000",
  3021=>"000111111",
  3022=>"000110111",
  3023=>"111111000",
  3024=>"001001000",
  3025=>"000000000",
  3026=>"000011111",
  3027=>"111111101",
  3028=>"000111111",
  3029=>"000001000",
  3030=>"000000000",
  3031=>"000111111",
  3032=>"100000000",
  3033=>"111000100",
  3034=>"000100111",
  3035=>"111000111",
  3036=>"111111101",
  3037=>"111111111",
  3038=>"111100000",
  3039=>"000001011",
  3040=>"110111111",
  3041=>"001000000",
  3042=>"000000011",
  3043=>"100111111",
  3044=>"110100000",
  3045=>"001111111",
  3046=>"000000111",
  3047=>"111111010",
  3048=>"000011110",
  3049=>"110100000",
  3050=>"001101111",
  3051=>"000000000",
  3052=>"100000000",
  3053=>"111010011",
  3054=>"100100000",
  3055=>"000111111",
  3056=>"001001001",
  3057=>"111111000",
  3058=>"111111001",
  3059=>"111101000",
  3060=>"001100000",
  3061=>"101111000",
  3062=>"111100000",
  3063=>"101101111",
  3064=>"111101100",
  3065=>"001101111",
  3066=>"000111111",
  3067=>"111111000",
  3068=>"110000110",
  3069=>"111111001",
  3070=>"000000000",
  3071=>"101001001",
  3072=>"010010110",
  3073=>"001101111",
  3074=>"111000001",
  3075=>"101101111",
  3076=>"001001000",
  3077=>"111111111",
  3078=>"011000000",
  3079=>"111111111",
  3080=>"000000111",
  3081=>"011011011",
  3082=>"100000000",
  3083=>"111100000",
  3084=>"000100110",
  3085=>"000100000",
  3086=>"111111000",
  3087=>"000000111",
  3088=>"111000000",
  3089=>"001011111",
  3090=>"000000111",
  3091=>"110111111",
  3092=>"111111101",
  3093=>"000000111",
  3094=>"000000111",
  3095=>"001100000",
  3096=>"100100000",
  3097=>"000111111",
  3098=>"001000101",
  3099=>"011010000",
  3100=>"111110000",
  3101=>"111100100",
  3102=>"000000000",
  3103=>"111111111",
  3104=>"001001000",
  3105=>"000000000",
  3106=>"100100100",
  3107=>"101000000",
  3108=>"011001001",
  3109=>"111111111",
  3110=>"000000001",
  3111=>"111111000",
  3112=>"000000001",
  3113=>"111000000",
  3114=>"111111111",
  3115=>"111110000",
  3116=>"101001011",
  3117=>"100111111",
  3118=>"110110111",
  3119=>"001001001",
  3120=>"111111000",
  3121=>"000000001",
  3122=>"001001000",
  3123=>"011111111",
  3124=>"000111111",
  3125=>"000000110",
  3126=>"100100110",
  3127=>"000000000",
  3128=>"110111000",
  3129=>"000000110",
  3130=>"000000000",
  3131=>"000000000",
  3132=>"101101001",
  3133=>"100000001",
  3134=>"000010111",
  3135=>"111000011",
  3136=>"000001001",
  3137=>"110111101",
  3138=>"111000110",
  3139=>"111111000",
  3140=>"000001111",
  3141=>"001000000",
  3142=>"000000000",
  3143=>"111000111",
  3144=>"001001001",
  3145=>"111011011",
  3146=>"111111111",
  3147=>"111111111",
  3148=>"111111111",
  3149=>"111111000",
  3150=>"001011011",
  3151=>"000000000",
  3152=>"011000000",
  3153=>"000001001",
  3154=>"111000000",
  3155=>"011110000",
  3156=>"000111000",
  3157=>"011111000",
  3158=>"111000101",
  3159=>"000000000",
  3160=>"111100000",
  3161=>"111000000",
  3162=>"101001101",
  3163=>"111111000",
  3164=>"000000110",
  3165=>"111111111",
  3166=>"000000111",
  3167=>"011000000",
  3168=>"000000000",
  3169=>"000000000",
  3170=>"000000111",
  3171=>"000000000",
  3172=>"000000000",
  3173=>"011000000",
  3174=>"000000111",
  3175=>"010010000",
  3176=>"000101111",
  3177=>"110000000",
  3178=>"111010111",
  3179=>"001001111",
  3180=>"001000111",
  3181=>"000000000",
  3182=>"111001000",
  3183=>"111111000",
  3184=>"111111111",
  3185=>"000111111",
  3186=>"010111111",
  3187=>"000000111",
  3188=>"111001001",
  3189=>"000100110",
  3190=>"100000000",
  3191=>"000000111",
  3192=>"001101111",
  3193=>"000000111",
  3194=>"010111111",
  3195=>"111111110",
  3196=>"000110110",
  3197=>"011000000",
  3198=>"000111111",
  3199=>"111111000",
  3200=>"001111111",
  3201=>"001001001",
  3202=>"111111011",
  3203=>"111101101",
  3204=>"111001011",
  3205=>"111000000",
  3206=>"111000000",
  3207=>"000111111",
  3208=>"000000000",
  3209=>"000000000",
  3210=>"110110110",
  3211=>"111111111",
  3212=>"110010100",
  3213=>"010111001",
  3214=>"101101111",
  3215=>"100110111",
  3216=>"000000111",
  3217=>"111111111",
  3218=>"011000011",
  3219=>"010010010",
  3220=>"000000100",
  3221=>"000111111",
  3222=>"000001001",
  3223=>"101001001",
  3224=>"001000111",
  3225=>"101000110",
  3226=>"001101100",
  3227=>"111100110",
  3228=>"111111101",
  3229=>"101000111",
  3230=>"111001001",
  3231=>"000000011",
  3232=>"001111011",
  3233=>"000000100",
  3234=>"111000100",
  3235=>"101001111",
  3236=>"000010111",
  3237=>"000000111",
  3238=>"000011000",
  3239=>"100111001",
  3240=>"111111000",
  3241=>"000001111",
  3242=>"111000000",
  3243=>"000000001",
  3244=>"110011011",
  3245=>"111111000",
  3246=>"111111111",
  3247=>"111111000",
  3248=>"111000001",
  3249=>"000100111",
  3250=>"110111110",
  3251=>"000000100",
  3252=>"000000000",
  3253=>"111111011",
  3254=>"000000000",
  3255=>"000000111",
  3256=>"100000110",
  3257=>"111111111",
  3258=>"000000111",
  3259=>"111111110",
  3260=>"000000001",
  3261=>"111111011",
  3262=>"100100111",
  3263=>"111111111",
  3264=>"111111110",
  3265=>"001000000",
  3266=>"111100101",
  3267=>"000100100",
  3268=>"111111000",
  3269=>"000000000",
  3270=>"000110000",
  3271=>"111111000",
  3272=>"111110000",
  3273=>"111111111",
  3274=>"000000001",
  3275=>"000110111",
  3276=>"101101111",
  3277=>"000000100",
  3278=>"001001011",
  3279=>"001000111",
  3280=>"111111111",
  3281=>"111000000",
  3282=>"000010000",
  3283=>"101000000",
  3284=>"001001111",
  3285=>"100000000",
  3286=>"000000000",
  3287=>"001001111",
  3288=>"000000110",
  3289=>"111010000",
  3290=>"111111000",
  3291=>"001111101",
  3292=>"111111000",
  3293=>"111111111",
  3294=>"111111010",
  3295=>"000000000",
  3296=>"111111111",
  3297=>"110011000",
  3298=>"000000110",
  3299=>"111111111",
  3300=>"001001000",
  3301=>"111111000",
  3302=>"011111011",
  3303=>"111111111",
  3304=>"000000100",
  3305=>"000110110",
  3306=>"111111100",
  3307=>"101101111",
  3308=>"000111111",
  3309=>"001001001",
  3310=>"000000000",
  3311=>"001000111",
  3312=>"111011100",
  3313=>"000000001",
  3314=>"001101111",
  3315=>"000001000",
  3316=>"100110111",
  3317=>"110100000",
  3318=>"110100001",
  3319=>"101100111",
  3320=>"000000101",
  3321=>"111111000",
  3322=>"111111111",
  3323=>"000000011",
  3324=>"000000110",
  3325=>"111111110",
  3326=>"011000000",
  3327=>"111111000",
  3328=>"001000000",
  3329=>"000001101",
  3330=>"111011011",
  3331=>"100000000",
  3332=>"111101111",
  3333=>"100111111",
  3334=>"001001111",
  3335=>"100000111",
  3336=>"000000111",
  3337=>"000000000",
  3338=>"110110000",
  3339=>"000000110",
  3340=>"100100111",
  3341=>"111111100",
  3342=>"011111000",
  3343=>"000000000",
  3344=>"111111000",
  3345=>"000110111",
  3346=>"000000000",
  3347=>"000100100",
  3348=>"000011111",
  3349=>"000000111",
  3350=>"000111111",
  3351=>"000111000",
  3352=>"000111111",
  3353=>"111101111",
  3354=>"000111100",
  3355=>"111111001",
  3356=>"100110111",
  3357=>"000000001",
  3358=>"111111011",
  3359=>"000000111",
  3360=>"110010000",
  3361=>"111111000",
  3362=>"111111111",
  3363=>"111110111",
  3364=>"100000000",
  3365=>"111001101",
  3366=>"110111000",
  3367=>"011000000",
  3368=>"000000101",
  3369=>"100101111",
  3370=>"000000010",
  3371=>"111110101",
  3372=>"111111000",
  3373=>"111001001",
  3374=>"000000000",
  3375=>"111011000",
  3376=>"111111111",
  3377=>"111111000",
  3378=>"101100110",
  3379=>"000000111",
  3380=>"100000000",
  3381=>"000111000",
  3382=>"000000000",
  3383=>"001001001",
  3384=>"001000000",
  3385=>"101001111",
  3386=>"111001000",
  3387=>"001101111",
  3388=>"001001111",
  3389=>"111111000",
  3390=>"000000101",
  3391=>"000001111",
  3392=>"000000000",
  3393=>"100111111",
  3394=>"111000001",
  3395=>"111111001",
  3396=>"111111000",
  3397=>"111111101",
  3398=>"001001111",
  3399=>"000000101",
  3400=>"000000010",
  3401=>"011000000",
  3402=>"111111111",
  3403=>"000111111",
  3404=>"010010010",
  3405=>"100000111",
  3406=>"000000001",
  3407=>"000000100",
  3408=>"111111000",
  3409=>"000000111",
  3410=>"001100101",
  3411=>"101111111",
  3412=>"100000001",
  3413=>"011011001",
  3414=>"111101111",
  3415=>"001000111",
  3416=>"111111111",
  3417=>"000000000",
  3418=>"000000000",
  3419=>"111111111",
  3420=>"101000000",
  3421=>"100000000",
  3422=>"001111111",
  3423=>"011111100",
  3424=>"101000000",
  3425=>"000000000",
  3426=>"000100011",
  3427=>"111000000",
  3428=>"000100111",
  3429=>"000000111",
  3430=>"000000100",
  3431=>"100100100",
  3432=>"000010111",
  3433=>"111111111",
  3434=>"000000111",
  3435=>"111010100",
  3436=>"001111000",
  3437=>"000000000",
  3438=>"000000000",
  3439=>"000000000",
  3440=>"000000000",
  3441=>"111001001",
  3442=>"000001001",
  3443=>"000000111",
  3444=>"011010001",
  3445=>"000000101",
  3446=>"111111111",
  3447=>"000111000",
  3448=>"111111000",
  3449=>"010010010",
  3450=>"000000111",
  3451=>"011000000",
  3452=>"010000010",
  3453=>"111111000",
  3454=>"000000000",
  3455=>"000000111",
  3456=>"110110110",
  3457=>"000000000",
  3458=>"000000000",
  3459=>"111111111",
  3460=>"100000000",
  3461=>"011111000",
  3462=>"111111111",
  3463=>"111111110",
  3464=>"111111000",
  3465=>"011111110",
  3466=>"000000001",
  3467=>"111111000",
  3468=>"000101111",
  3469=>"100110011",
  3470=>"111111110",
  3471=>"000000010",
  3472=>"000001000",
  3473=>"111111000",
  3474=>"110110111",
  3475=>"000000110",
  3476=>"110110000",
  3477=>"000000011",
  3478=>"111111111",
  3479=>"111111000",
  3480=>"000111000",
  3481=>"011100000",
  3482=>"000000011",
  3483=>"011111111",
  3484=>"111001001",
  3485=>"111001000",
  3486=>"000111111",
  3487=>"000000000",
  3488=>"000011111",
  3489=>"001000001",
  3490=>"000000001",
  3491=>"000000101",
  3492=>"101000000",
  3493=>"110000000",
  3494=>"000000000",
  3495=>"111101101",
  3496=>"011111001",
  3497=>"000000011",
  3498=>"011011111",
  3499=>"000100111",
  3500=>"000000000",
  3501=>"000100111",
  3502=>"000000110",
  3503=>"000000000",
  3504=>"111000000",
  3505=>"000000001",
  3506=>"111111000",
  3507=>"111011111",
  3508=>"001001111",
  3509=>"111110100",
  3510=>"000100111",
  3511=>"110111111",
  3512=>"111001000",
  3513=>"111111111",
  3514=>"000000000",
  3515=>"001000001",
  3516=>"000101011",
  3517=>"100000000",
  3518=>"000000101",
  3519=>"100100100",
  3520=>"000101111",
  3521=>"000000000",
  3522=>"001000000",
  3523=>"110000000",
  3524=>"111111111",
  3525=>"011011111",
  3526=>"111101000",
  3527=>"111111000",
  3528=>"011000000",
  3529=>"000100110",
  3530=>"000000000",
  3531=>"111111000",
  3532=>"000000000",
  3533=>"111111000",
  3534=>"101000001",
  3535=>"011110101",
  3536=>"111111011",
  3537=>"000000111",
  3538=>"111001101",
  3539=>"001111111",
  3540=>"100101000",
  3541=>"111010111",
  3542=>"000000011",
  3543=>"000000001",
  3544=>"111001111",
  3545=>"011001000",
  3546=>"111111111",
  3547=>"111000000",
  3548=>"000000000",
  3549=>"111101000",
  3550=>"101101000",
  3551=>"101111101",
  3552=>"111111000",
  3553=>"111111100",
  3554=>"111111111",
  3555=>"000100111",
  3556=>"001000010",
  3557=>"100101111",
  3558=>"101000111",
  3559=>"000000111",
  3560=>"111110010",
  3561=>"111111010",
  3562=>"000000111",
  3563=>"110111001",
  3564=>"111111110",
  3565=>"011111111",
  3566=>"000100100",
  3567=>"010011000",
  3568=>"111110111",
  3569=>"011101000",
  3570=>"111001000",
  3571=>"111111111",
  3572=>"111000011",
  3573=>"000000001",
  3574=>"100000000",
  3575=>"011010000",
  3576=>"001111000",
  3577=>"000001101",
  3578=>"111111101",
  3579=>"111101001",
  3580=>"110110111",
  3581=>"110111111",
  3582=>"001000000",
  3583=>"000000111",
  3584=>"000000000",
  3585=>"000000110",
  3586=>"000000000",
  3587=>"111111111",
  3588=>"000000000",
  3589=>"000010110",
  3590=>"111111111",
  3591=>"010000000",
  3592=>"111111110",
  3593=>"000000000",
  3594=>"111111111",
  3595=>"110010110",
  3596=>"000000000",
  3597=>"000000000",
  3598=>"000110000",
  3599=>"110110111",
  3600=>"000000000",
  3601=>"111111111",
  3602=>"010000000",
  3603=>"000000000",
  3604=>"111111111",
  3605=>"000000010",
  3606=>"110111111",
  3607=>"111111101",
  3608=>"111011111",
  3609=>"000000000",
  3610=>"000000000",
  3611=>"110001111",
  3612=>"111111111",
  3613=>"000000110",
  3614=>"111111110",
  3615=>"000000000",
  3616=>"110111111",
  3617=>"111111111",
  3618=>"111111111",
  3619=>"011111001",
  3620=>"001001001",
  3621=>"110111111",
  3622=>"110110110",
  3623=>"110111111",
  3624=>"111111111",
  3625=>"011000000",
  3626=>"011000000",
  3627=>"111111111",
  3628=>"000110111",
  3629=>"000010000",
  3630=>"101111000",
  3631=>"011000000",
  3632=>"011011111",
  3633=>"100000100",
  3634=>"111100110",
  3635=>"111111111",
  3636=>"001011001",
  3637=>"000000000",
  3638=>"110100000",
  3639=>"010110010",
  3640=>"000000110",
  3641=>"011000000",
  3642=>"000000100",
  3643=>"011000000",
  3644=>"110000000",
  3645=>"110110100",
  3646=>"010011011",
  3647=>"000111111",
  3648=>"000001001",
  3649=>"100101111",
  3650=>"000000000",
  3651=>"001000110",
  3652=>"110110110",
  3653=>"000000000",
  3654=>"000001000",
  3655=>"000000000",
  3656=>"100100000",
  3657=>"000000000",
  3658=>"001111010",
  3659=>"000000000",
  3660=>"011001000",
  3661=>"000000000",
  3662=>"110000000",
  3663=>"000010000",
  3664=>"000000000",
  3665=>"011111111",
  3666=>"011111111",
  3667=>"111101101",
  3668=>"000110110",
  3669=>"111111111",
  3670=>"111100000",
  3671=>"000100110",
  3672=>"011111001",
  3673=>"000000001",
  3674=>"000000001",
  3675=>"100100100",
  3676=>"000000000",
  3677=>"000001111",
  3678=>"110111100",
  3679=>"000000000",
  3680=>"111000001",
  3681=>"101000000",
  3682=>"000000111",
  3683=>"110000011",
  3684=>"000100000",
  3685=>"111001001",
  3686=>"000000000",
  3687=>"100111111",
  3688=>"100100100",
  3689=>"000000000",
  3690=>"010000110",
  3691=>"111111111",
  3692=>"000000001",
  3693=>"111011010",
  3694=>"000000111",
  3695=>"111111111",
  3696=>"001100111",
  3697=>"001000100",
  3698=>"101100101",
  3699=>"111111110",
  3700=>"000000000",
  3701=>"100111111",
  3702=>"111111111",
  3703=>"000010000",
  3704=>"111111110",
  3705=>"111111000",
  3706=>"000000001",
  3707=>"111111111",
  3708=>"000000000",
  3709=>"100100000",
  3710=>"000000000",
  3711=>"000100101",
  3712=>"000001011",
  3713=>"111111111",
  3714=>"001011000",
  3715=>"111111111",
  3716=>"000000000",
  3717=>"000000000",
  3718=>"011111111",
  3719=>"000000110",
  3720=>"010010000",
  3721=>"001000000",
  3722=>"001000000",
  3723=>"110000000",
  3724=>"111111111",
  3725=>"110000000",
  3726=>"111111111",
  3727=>"111011000",
  3728=>"000000000",
  3729=>"000100100",
  3730=>"111001010",
  3731=>"111111111",
  3732=>"011111110",
  3733=>"000110111",
  3734=>"100000000",
  3735=>"011111111",
  3736=>"000000100",
  3737=>"001001011",
  3738=>"110111111",
  3739=>"111111111",
  3740=>"111000110",
  3741=>"111000000",
  3742=>"000000000",
  3743=>"110110110",
  3744=>"000000110",
  3745=>"011111100",
  3746=>"111111111",
  3747=>"000000011",
  3748=>"100000000",
  3749=>"111101111",
  3750=>"111111100",
  3751=>"000000000",
  3752=>"000100111",
  3753=>"000000100",
  3754=>"111011000",
  3755=>"000001011",
  3756=>"111111111",
  3757=>"011011000",
  3758=>"111111010",
  3759=>"111111000",
  3760=>"000000000",
  3761=>"011110100",
  3762=>"110110111",
  3763=>"111011010",
  3764=>"000101000",
  3765=>"111111111",
  3766=>"110110111",
  3767=>"111111110",
  3768=>"000000010",
  3769=>"111111111",
  3770=>"110010000",
  3771=>"110100100",
  3772=>"100000000",
  3773=>"010111111",
  3774=>"111010000",
  3775=>"111110111",
  3776=>"111111111",
  3777=>"111111111",
  3778=>"000000110",
  3779=>"111111111",
  3780=>"111111111",
  3781=>"011001000",
  3782=>"111001000",
  3783=>"011000000",
  3784=>"100000000",
  3785=>"111111111",
  3786=>"010000100",
  3787=>"000100110",
  3788=>"011010111",
  3789=>"001000100",
  3790=>"010100100",
  3791=>"000000000",
  3792=>"000000000",
  3793=>"110110111",
  3794=>"110000100",
  3795=>"000000000",
  3796=>"010110110",
  3797=>"011111111",
  3798=>"110000000",
  3799=>"101101111",
  3800=>"001101111",
  3801=>"000001001",
  3802=>"000001111",
  3803=>"011000000",
  3804=>"000000000",
  3805=>"110110011",
  3806=>"111111111",
  3807=>"110100100",
  3808=>"000000000",
  3809=>"111111111",
  3810=>"011000111",
  3811=>"111111010",
  3812=>"110110000",
  3813=>"000000010",
  3814=>"000000000",
  3815=>"000000000",
  3816=>"000000000",
  3817=>"000110000",
  3818=>"000000011",
  3819=>"111111111",
  3820=>"000000000",
  3821=>"111111111",
  3822=>"111111000",
  3823=>"000000000",
  3824=>"111000000",
  3825=>"110110111",
  3826=>"111000000",
  3827=>"000000000",
  3828=>"000000000",
  3829=>"001000000",
  3830=>"000110110",
  3831=>"000000100",
  3832=>"011110111",
  3833=>"110000000",
  3834=>"000110110",
  3835=>"000000010",
  3836=>"110000100",
  3837=>"000000000",
  3838=>"111111111",
  3839=>"100000000",
  3840=>"000111110",
  3841=>"111101111",
  3842=>"111101100",
  3843=>"111111111",
  3844=>"111001011",
  3845=>"000000110",
  3846=>"111111111",
  3847=>"010110100",
  3848=>"000000000",
  3849=>"000000100",
  3850=>"111111111",
  3851=>"000000000",
  3852=>"111111111",
  3853=>"000110110",
  3854=>"011110111",
  3855=>"000000000",
  3856=>"000010011",
  3857=>"111111011",
  3858=>"110111111",
  3859=>"111110000",
  3860=>"111111010",
  3861=>"000000001",
  3862=>"100100100",
  3863=>"000000000",
  3864=>"011000000",
  3865=>"111000000",
  3866=>"000110110",
  3867=>"000010110",
  3868=>"111111111",
  3869=>"100000011",
  3870=>"000000000",
  3871=>"111111111",
  3872=>"000011001",
  3873=>"011110111",
  3874=>"000000011",
  3875=>"011111111",
  3876=>"111111111",
  3877=>"001000111",
  3878=>"001001111",
  3879=>"111111111",
  3880=>"011011010",
  3881=>"111111110",
  3882=>"111111111",
  3883=>"000000000",
  3884=>"000110110",
  3885=>"000000000",
  3886=>"110000111",
  3887=>"001001111",
  3888=>"110110110",
  3889=>"110000000",
  3890=>"111111111",
  3891=>"111111011",
  3892=>"000000001",
  3893=>"000000000",
  3894=>"111110111",
  3895=>"111111111",
  3896=>"000000000",
  3897=>"001101111",
  3898=>"110110110",
  3899=>"111111110",
  3900=>"110110110",
  3901=>"000100110",
  3902=>"110111110",
  3903=>"111111100",
  3904=>"011010010",
  3905=>"000100001",
  3906=>"110110100",
  3907=>"111001101",
  3908=>"000000000",
  3909=>"111111111",
  3910=>"111111111",
  3911=>"000000000",
  3912=>"111111111",
  3913=>"111000100",
  3914=>"010010000",
  3915=>"111100000",
  3916=>"010010010",
  3917=>"000000110",
  3918=>"111111111",
  3919=>"111111111",
  3920=>"000000000",
  3921=>"000001101",
  3922=>"010000000",
  3923=>"111111101",
  3924=>"000000000",
  3925=>"100100100",
  3926=>"111111111",
  3927=>"100111010",
  3928=>"000000000",
  3929=>"000000100",
  3930=>"010010010",
  3931=>"000000000",
  3932=>"111111101",
  3933=>"111011000",
  3934=>"011111111",
  3935=>"000000000",
  3936=>"110110100",
  3937=>"111111110",
  3938=>"000100100",
  3939=>"000000000",
  3940=>"001011000",
  3941=>"111111111",
  3942=>"111111111",
  3943=>"111010000",
  3944=>"100010000",
  3945=>"111111111",
  3946=>"110010000",
  3947=>"110000000",
  3948=>"000000000",
  3949=>"110111000",
  3950=>"111101000",
  3951=>"101111111",
  3952=>"111111111",
  3953=>"100000000",
  3954=>"111111111",
  3955=>"011011010",
  3956=>"110100100",
  3957=>"111111111",
  3958=>"111111111",
  3959=>"111111101",
  3960=>"011111000",
  3961=>"101101111",
  3962=>"000000101",
  3963=>"111111111",
  3964=>"000000000",
  3965=>"111001111",
  3966=>"100001111",
  3967=>"111111111",
  3968=>"001001111",
  3969=>"111101111",
  3970=>"000000100",
  3971=>"000000101",
  3972=>"111111111",
  3973=>"000000001",
  3974=>"000000000",
  3975=>"111111111",
  3976=>"000000000",
  3977=>"011001001",
  3978=>"000000000",
  3979=>"111101001",
  3980=>"011010000",
  3981=>"111011011",
  3982=>"001011111",
  3983=>"111111000",
  3984=>"111010000",
  3985=>"111110110",
  3986=>"000000000",
  3987=>"111111111",
  3988=>"111111111",
  3989=>"111111111",
  3990=>"111100000",
  3991=>"100000000",
  3992=>"000000000",
  3993=>"110110110",
  3994=>"000000000",
  3995=>"011011111",
  3996=>"001000001",
  3997=>"111111111",
  3998=>"110010110",
  3999=>"110010000",
  4000=>"111000000",
  4001=>"110100000",
  4002=>"000000110",
  4003=>"000100110",
  4004=>"111100100",
  4005=>"001001101",
  4006=>"000000111",
  4007=>"111110000",
  4008=>"100100000",
  4009=>"000100000",
  4010=>"000000000",
  4011=>"011011000",
  4012=>"000111111",
  4013=>"110000000",
  4014=>"111011000",
  4015=>"000000000",
  4016=>"000000000",
  4017=>"001010110",
  4018=>"111111111",
  4019=>"111111111",
  4020=>"111111111",
  4021=>"001001101",
  4022=>"111000010",
  4023=>"000100111",
  4024=>"010111111",
  4025=>"111111111",
  4026=>"000100000",
  4027=>"010000010",
  4028=>"000000000",
  4029=>"111111111",
  4030=>"000000000",
  4031=>"100100100",
  4032=>"111111101",
  4033=>"000010010",
  4034=>"111111111",
  4035=>"000000000",
  4036=>"111100111",
  4037=>"111100000",
  4038=>"000000000",
  4039=>"000001101",
  4040=>"000000000",
  4041=>"000000111",
  4042=>"000000000",
  4043=>"110011111",
  4044=>"111000000",
  4045=>"111111111",
  4046=>"000000000",
  4047=>"110011001",
  4048=>"000000000",
  4049=>"011111111",
  4050=>"000000000",
  4051=>"111000000",
  4052=>"100100000",
  4053=>"000000000",
  4054=>"110110000",
  4055=>"001000000",
  4056=>"000000110",
  4057=>"010110110",
  4058=>"111111111",
  4059=>"111110100",
  4060=>"111111111",
  4061=>"011000000",
  4062=>"000000111",
  4063=>"000001011",
  4064=>"010000000",
  4065=>"000000110",
  4066=>"101001000",
  4067=>"001000000",
  4068=>"000000000",
  4069=>"000000000",
  4070=>"000000000",
  4071=>"101101111",
  4072=>"000100110",
  4073=>"111000010",
  4074=>"101111111",
  4075=>"111111111",
  4076=>"111000001",
  4077=>"110000110",
  4078=>"011100110",
  4079=>"011111111",
  4080=>"110110100",
  4081=>"011000001",
  4082=>"111100101",
  4083=>"111000001",
  4084=>"000110101",
  4085=>"000000000",
  4086=>"000011011",
  4087=>"111011000",
  4088=>"111000111",
  4089=>"111110110",
  4090=>"111000000",
  4091=>"000000000",
  4092=>"000000000",
  4093=>"110100111",
  4094=>"011111111",
  4095=>"000000000",
  4096=>"111111000",
  4097=>"110000000",
  4098=>"100100000",
  4099=>"101000000",
  4100=>"110110000",
  4101=>"000101100",
  4102=>"000000000",
  4103=>"111011000",
  4104=>"100111111",
  4105=>"000000000",
  4106=>"010000111",
  4107=>"100000000",
  4108=>"110110110",
  4109=>"000001111",
  4110=>"000010010",
  4111=>"111111111",
  4112=>"000000000",
  4113=>"111111111",
  4114=>"000010000",
  4115=>"111110000",
  4116=>"000000000",
  4117=>"000000000",
  4118=>"111111111",
  4119=>"010110100",
  4120=>"000000000",
  4121=>"111111101",
  4122=>"000000111",
  4123=>"111001111",
  4124=>"111111111",
  4125=>"011111111",
  4126=>"011001100",
  4127=>"000100100",
  4128=>"011111111",
  4129=>"000000000",
  4130=>"110111111",
  4131=>"111111000",
  4132=>"000000101",
  4133=>"001001101",
  4134=>"000000111",
  4135=>"000001111",
  4136=>"000000001",
  4137=>"111111111",
  4138=>"011110000",
  4139=>"111111111",
  4140=>"000000000",
  4141=>"111111000",
  4142=>"101101111",
  4143=>"000100111",
  4144=>"111001001",
  4145=>"000011111",
  4146=>"000000000",
  4147=>"000111111",
  4148=>"000000000",
  4149=>"111110110",
  4150=>"000010000",
  4151=>"001101101",
  4152=>"011111111",
  4153=>"110111100",
  4154=>"110111111",
  4155=>"000111111",
  4156=>"000000000",
  4157=>"011010000",
  4158=>"010001111",
  4159=>"000000000",
  4160=>"000010010",
  4161=>"001001000",
  4162=>"011110111",
  4163=>"001001111",
  4164=>"110110110",
  4165=>"000100110",
  4166=>"110100000",
  4167=>"000000000",
  4168=>"111111111",
  4169=>"000100111",
  4170=>"000000000",
  4171=>"111111111",
  4172=>"000001111",
  4173=>"000000000",
  4174=>"000000111",
  4175=>"000000000",
  4176=>"111000000",
  4177=>"000000100",
  4178=>"000000110",
  4179=>"110110110",
  4180=>"000111111",
  4181=>"000111111",
  4182=>"011011111",
  4183=>"000100100",
  4184=>"101000001",
  4185=>"000100111",
  4186=>"111100111",
  4187=>"000000000",
  4188=>"110001001",
  4189=>"000101111",
  4190=>"000100000",
  4191=>"111010011",
  4192=>"101111111",
  4193=>"000000000",
  4194=>"000000000",
  4195=>"111101000",
  4196=>"110110000",
  4197=>"101100000",
  4198=>"111100101",
  4199=>"101000000",
  4200=>"100110010",
  4201=>"111100110",
  4202=>"111111111",
  4203=>"000000000",
  4204=>"111111111",
  4205=>"000000000",
  4206=>"100101101",
  4207=>"111111111",
  4208=>"000110000",
  4209=>"000000000",
  4210=>"011011011",
  4211=>"000111110",
  4212=>"010010000",
  4213=>"000000000",
  4214=>"010111111",
  4215=>"111111111",
  4216=>"100000000",
  4217=>"011111011",
  4218=>"100000000",
  4219=>"000010000",
  4220=>"101001001",
  4221=>"000000000",
  4222=>"100110010",
  4223=>"000000000",
  4224=>"000000100",
  4225=>"111000000",
  4226=>"000000111",
  4227=>"000001001",
  4228=>"000001001",
  4229=>"000000000",
  4230=>"000001001",
  4231=>"111000000",
  4232=>"110111110",
  4233=>"111110000",
  4234=>"111111111",
  4235=>"010110010",
  4236=>"001111101",
  4237=>"000000000",
  4238=>"000100111",
  4239=>"000000000",
  4240=>"001101111",
  4241=>"000000000",
  4242=>"110111111",
  4243=>"100100110",
  4244=>"000111111",
  4245=>"011111000",
  4246=>"000000000",
  4247=>"000000000",
  4248=>"111101100",
  4249=>"011000111",
  4250=>"000110011",
  4251=>"100000001",
  4252=>"111111001",
  4253=>"001000000",
  4254=>"110000110",
  4255=>"001000000",
  4256=>"111111000",
  4257=>"110000011",
  4258=>"111111000",
  4259=>"000000001",
  4260=>"111100110",
  4261=>"111111111",
  4262=>"111101101",
  4263=>"001011001",
  4264=>"111111111",
  4265=>"111111111",
  4266=>"000010000",
  4267=>"111111111",
  4268=>"111011011",
  4269=>"110110000",
  4270=>"111111111",
  4271=>"011111111",
  4272=>"001000000",
  4273=>"111111111",
  4274=>"111011010",
  4275=>"111000000",
  4276=>"100100001",
  4277=>"000000001",
  4278=>"000010111",
  4279=>"111111111",
  4280=>"111111111",
  4281=>"111111010",
  4282=>"111000000",
  4283=>"111100111",
  4284=>"000000100",
  4285=>"111100111",
  4286=>"000111111",
  4287=>"111111011",
  4288=>"110110110",
  4289=>"000000000",
  4290=>"001010000",
  4291=>"100000000",
  4292=>"111001000",
  4293=>"101000000",
  4294=>"111111111",
  4295=>"111100000",
  4296=>"000000111",
  4297=>"000000011",
  4298=>"000000101",
  4299=>"001111111",
  4300=>"111111111",
  4301=>"011000001",
  4302=>"000111111",
  4303=>"000100010",
  4304=>"000000000",
  4305=>"000000000",
  4306=>"000000000",
  4307=>"110000000",
  4308=>"000000000",
  4309=>"111111111",
  4310=>"100000000",
  4311=>"000010111",
  4312=>"000000111",
  4313=>"111111110",
  4314=>"000000111",
  4315=>"111111111",
  4316=>"010111111",
  4317=>"000011111",
  4318=>"111110000",
  4319=>"111111111",
  4320=>"111000000",
  4321=>"001011000",
  4322=>"111101100",
  4323=>"000000000",
  4324=>"000111111",
  4325=>"000000000",
  4326=>"000000000",
  4327=>"011000000",
  4328=>"000000000",
  4329=>"101001000",
  4330=>"111111111",
  4331=>"000000101",
  4332=>"000000000",
  4333=>"111111111",
  4334=>"111111111",
  4335=>"000000000",
  4336=>"111111111",
  4337=>"111111111",
  4338=>"000000000",
  4339=>"000000110",
  4340=>"111111111",
  4341=>"011100100",
  4342=>"110110100",
  4343=>"000000000",
  4344=>"111111111",
  4345=>"100000000",
  4346=>"111011111",
  4347=>"000001001",
  4348=>"110111110",
  4349=>"000000110",
  4350=>"000000000",
  4351=>"000000000",
  4352=>"111111100",
  4353=>"001001001",
  4354=>"111000001",
  4355=>"111111111",
  4356=>"000000000",
  4357=>"001000011",
  4358=>"001111111",
  4359=>"000001111",
  4360=>"100000000",
  4361=>"111100100",
  4362=>"111100101",
  4363=>"111111111",
  4364=>"100000000",
  4365=>"000110000",
  4366=>"000000001",
  4367=>"000000000",
  4368=>"110110101",
  4369=>"111111011",
  4370=>"000000000",
  4371=>"000000101",
  4372=>"000110111",
  4373=>"000000000",
  4374=>"000000000",
  4375=>"111111111",
  4376=>"111111111",
  4377=>"111000000",
  4378=>"000111001",
  4379=>"000000000",
  4380=>"110110100",
  4381=>"111100000",
  4382=>"000000000",
  4383=>"111000000",
  4384=>"001111000",
  4385=>"000000000",
  4386=>"011000110",
  4387=>"010001000",
  4388=>"111111111",
  4389=>"000111111",
  4390=>"011111011",
  4391=>"111100100",
  4392=>"000010111",
  4393=>"000000000",
  4394=>"000011000",
  4395=>"000001011",
  4396=>"000001001",
  4397=>"100100000",
  4398=>"000000000",
  4399=>"000101011",
  4400=>"100001101",
  4401=>"110010001",
  4402=>"111111111",
  4403=>"110110110",
  4404=>"000000110",
  4405=>"101111111",
  4406=>"111111111",
  4407=>"001000001",
  4408=>"000001010",
  4409=>"111000000",
  4410=>"111111111",
  4411=>"101110000",
  4412=>"110110000",
  4413=>"001001011",
  4414=>"000000001",
  4415=>"111000000",
  4416=>"100100000",
  4417=>"001111111",
  4418=>"000000001",
  4419=>"000011111",
  4420=>"000101101",
  4421=>"111111111",
  4422=>"000000000",
  4423=>"000000000",
  4424=>"111101111",
  4425=>"000000001",
  4426=>"111011011",
  4427=>"100100000",
  4428=>"111101111",
  4429=>"000000111",
  4430=>"111000001",
  4431=>"000110110",
  4432=>"000000000",
  4433=>"000000000",
  4434=>"000000000",
  4435=>"111111111",
  4436=>"111111010",
  4437=>"111011011",
  4438=>"000001111",
  4439=>"111110100",
  4440=>"000010011",
  4441=>"000000000",
  4442=>"000110110",
  4443=>"000000000",
  4444=>"000000000",
  4445=>"000000000",
  4446=>"000000011",
  4447=>"001001000",
  4448=>"111111111",
  4449=>"111111011",
  4450=>"011011001",
  4451=>"001001001",
  4452=>"110010000",
  4453=>"000100000",
  4454=>"110000000",
  4455=>"000000101",
  4456=>"011011000",
  4457=>"001001000",
  4458=>"100000000",
  4459=>"100000000",
  4460=>"111111111",
  4461=>"111100111",
  4462=>"110111111",
  4463=>"111101111",
  4464=>"000000000",
  4465=>"111001011",
  4466=>"001111010",
  4467=>"111001101",
  4468=>"000000100",
  4469=>"000110111",
  4470=>"100000111",
  4471=>"111111001",
  4472=>"000000000",
  4473=>"111111101",
  4474=>"000001111",
  4475=>"000000000",
  4476=>"101101111",
  4477=>"000000101",
  4478=>"000000000",
  4479=>"111110110",
  4480=>"011111111",
  4481=>"000000000",
  4482=>"000001001",
  4483=>"000000000",
  4484=>"000001111",
  4485=>"001111100",
  4486=>"110110001",
  4487=>"111111111",
  4488=>"000000000",
  4489=>"001000111",
  4490=>"001111011",
  4491=>"111111111",
  4492=>"000000000",
  4493=>"111010111",
  4494=>"111111111",
  4495=>"111110100",
  4496=>"000000000",
  4497=>"000000000",
  4498=>"011111111",
  4499=>"111111001",
  4500=>"111111111",
  4501=>"001101111",
  4502=>"110000000",
  4503=>"010000000",
  4504=>"000100100",
  4505=>"001000000",
  4506=>"111011101",
  4507=>"101000001",
  4508=>"100000000",
  4509=>"000000010",
  4510=>"001111111",
  4511=>"011111111",
  4512=>"000000000",
  4513=>"000001111",
  4514=>"111101111",
  4515=>"001000100",
  4516=>"111111111",
  4517=>"000000000",
  4518=>"000000100",
  4519=>"011110101",
  4520=>"111111111",
  4521=>"000111111",
  4522=>"111111111",
  4523=>"111000000",
  4524=>"011011111",
  4525=>"000000000",
  4526=>"001000111",
  4527=>"111111111",
  4528=>"000000000",
  4529=>"000000000",
  4530=>"000000000",
  4531=>"000000000",
  4532=>"110110000",
  4533=>"011000111",
  4534=>"010011011",
  4535=>"000000000",
  4536=>"000000000",
  4537=>"111110111",
  4538=>"111111001",
  4539=>"000000000",
  4540=>"111111111",
  4541=>"111111111",
  4542=>"111111100",
  4543=>"000001001",
  4544=>"000001000",
  4545=>"000000000",
  4546=>"000000000",
  4547=>"001101111",
  4548=>"110111111",
  4549=>"110000000",
  4550=>"000000000",
  4551=>"000000000",
  4552=>"111000100",
  4553=>"000000000",
  4554=>"000000100",
  4555=>"100111111",
  4556=>"000001001",
  4557=>"000000111",
  4558=>"000000000",
  4559=>"000000111",
  4560=>"111101001",
  4561=>"101111111",
  4562=>"101001000",
  4563=>"101111111",
  4564=>"000011001",
  4565=>"000110111",
  4566=>"001101001",
  4567=>"011011011",
  4568=>"111011111",
  4569=>"100110010",
  4570=>"000000000",
  4571=>"111111000",
  4572=>"101000100",
  4573=>"100000001",
  4574=>"111011011",
  4575=>"100111111",
  4576=>"111111001",
  4577=>"001001000",
  4578=>"011000000",
  4579=>"111111000",
  4580=>"000000000",
  4581=>"111111111",
  4582=>"000010111",
  4583=>"101000000",
  4584=>"000000000",
  4585=>"000000001",
  4586=>"111111000",
  4587=>"000000000",
  4588=>"111111111",
  4589=>"011010000",
  4590=>"000000000",
  4591=>"000000110",
  4592=>"100100001",
  4593=>"111111011",
  4594=>"010010000",
  4595=>"000000000",
  4596=>"011000001",
  4597=>"001000101",
  4598=>"111111111",
  4599=>"000010100",
  4600=>"000000000",
  4601=>"000000000",
  4602=>"000000000",
  4603=>"000100111",
  4604=>"000000000",
  4605=>"111000000",
  4606=>"000010010",
  4607=>"000000111",
  4608=>"111001101",
  4609=>"100000000",
  4610=>"100101111",
  4611=>"000000000",
  4612=>"011111011",
  4613=>"001100111",
  4614=>"010011010",
  4615=>"111111111",
  4616=>"011000000",
  4617=>"000000000",
  4618=>"000000111",
  4619=>"001001011",
  4620=>"100110110",
  4621=>"001100111",
  4622=>"111111111",
  4623=>"011001000",
  4624=>"111111101",
  4625=>"000000100",
  4626=>"011000000",
  4627=>"000000111",
  4628=>"110000011",
  4629=>"111000000",
  4630=>"110111111",
  4631=>"011011011",
  4632=>"000000000",
  4633=>"000000000",
  4634=>"000000000",
  4635=>"000001111",
  4636=>"111111001",
  4637=>"000100111",
  4638=>"111001001",
  4639=>"001000000",
  4640=>"110111100",
  4641=>"010110110",
  4642=>"100000000",
  4643=>"111111111",
  4644=>"000000001",
  4645=>"000000011",
  4646=>"000100101",
  4647=>"001000000",
  4648=>"001011101",
  4649=>"100100111",
  4650=>"010001111",
  4651=>"000000001",
  4652=>"101101101",
  4653=>"000100111",
  4654=>"000010110",
  4655=>"001000111",
  4656=>"111111111",
  4657=>"000001000",
  4658=>"001000000",
  4659=>"000000000",
  4660=>"011111000",
  4661=>"011011110",
  4662=>"000000011",
  4663=>"001000000",
  4664=>"000000000",
  4665=>"000000000",
  4666=>"111011010",
  4667=>"000000000",
  4668=>"111000000",
  4669=>"111001000",
  4670=>"111111111",
  4671=>"000000000",
  4672=>"111111110",
  4673=>"111010000",
  4674=>"011111111",
  4675=>"100000000",
  4676=>"111001000",
  4677=>"000000001",
  4678=>"010011111",
  4679=>"111100000",
  4680=>"011111111",
  4681=>"011111111",
  4682=>"100000000",
  4683=>"000001100",
  4684=>"011001000",
  4685=>"111011000",
  4686=>"011000000",
  4687=>"010111100",
  4688=>"111111100",
  4689=>"111010111",
  4690=>"011010010",
  4691=>"000000000",
  4692=>"000000000",
  4693=>"000000010",
  4694=>"000000000",
  4695=>"000111111",
  4696=>"000000101",
  4697=>"000000000",
  4698=>"000000000",
  4699=>"010011111",
  4700=>"100000111",
  4701=>"000111001",
  4702=>"111111111",
  4703=>"100100100",
  4704=>"111000000",
  4705=>"000000000",
  4706=>"101111111",
  4707=>"000000001",
  4708=>"001111110",
  4709=>"101101100",
  4710=>"000100111",
  4711=>"001111111",
  4712=>"000000000",
  4713=>"111000000",
  4714=>"000110111",
  4715=>"110110100",
  4716=>"111111111",
  4717=>"000000000",
  4718=>"000000111",
  4719=>"000000000",
  4720=>"000100000",
  4721=>"111111111",
  4722=>"000000110",
  4723=>"111111000",
  4724=>"100000000",
  4725=>"111111110",
  4726=>"000000000",
  4727=>"001011010",
  4728=>"101101111",
  4729=>"101001001",
  4730=>"110000000",
  4731=>"001001111",
  4732=>"100000100",
  4733=>"111101101",
  4734=>"010111110",
  4735=>"000000100",
  4736=>"111001001",
  4737=>"111111111",
  4738=>"111110000",
  4739=>"001000000",
  4740=>"110100100",
  4741=>"111111111",
  4742=>"101001000",
  4743=>"111111111",
  4744=>"000000000",
  4745=>"000000000",
  4746=>"111111111",
  4747=>"111110010",
  4748=>"000100111",
  4749=>"001000000",
  4750=>"000000001",
  4751=>"111111000",
  4752=>"111000111",
  4753=>"000000000",
  4754=>"111111000",
  4755=>"111111001",
  4756=>"111111110",
  4757=>"011011001",
  4758=>"000111111",
  4759=>"000111111",
  4760=>"111011111",
  4761=>"101111111",
  4762=>"111111101",
  4763=>"001001111",
  4764=>"000000000",
  4765=>"011011000",
  4766=>"001001000",
  4767=>"000000000",
  4768=>"111111111",
  4769=>"000000000",
  4770=>"000000111",
  4771=>"111111111",
  4772=>"110110110",
  4773=>"110111111",
  4774=>"111000100",
  4775=>"011100100",
  4776=>"111111111",
  4777=>"111001101",
  4778=>"010111111",
  4779=>"000010010",
  4780=>"000100100",
  4781=>"111111111",
  4782=>"111000000",
  4783=>"001000000",
  4784=>"000000011",
  4785=>"001001101",
  4786=>"111111111",
  4787=>"000000000",
  4788=>"000000000",
  4789=>"011000000",
  4790=>"111111000",
  4791=>"010011111",
  4792=>"111111111",
  4793=>"011111111",
  4794=>"000000000",
  4795=>"001001001",
  4796=>"000001111",
  4797=>"000000000",
  4798=>"000000110",
  4799=>"000000000",
  4800=>"000000001",
  4801=>"101001000",
  4802=>"111111111",
  4803=>"101111000",
  4804=>"111111111",
  4805=>"000000000",
  4806=>"111110010",
  4807=>"000000000",
  4808=>"000111110",
  4809=>"001000000",
  4810=>"110110000",
  4811=>"100000000",
  4812=>"000000000",
  4813=>"001101100",
  4814=>"011111000",
  4815=>"100100000",
  4816=>"000000111",
  4817=>"110000111",
  4818=>"111000000",
  4819=>"000000000",
  4820=>"000110111",
  4821=>"111100111",
  4822=>"100000000",
  4823=>"000000001",
  4824=>"000110111",
  4825=>"000000001",
  4826=>"000100111",
  4827=>"011000111",
  4828=>"000000000",
  4829=>"111000000",
  4830=>"111111111",
  4831=>"011101110",
  4832=>"111111111",
  4833=>"000110111",
  4834=>"100100100",
  4835=>"001000000",
  4836=>"011011001",
  4837=>"010110111",
  4838=>"000000000",
  4839=>"000000000",
  4840=>"111111111",
  4841=>"111111111",
  4842=>"111111111",
  4843=>"000000111",
  4844=>"111001000",
  4845=>"101101101",
  4846=>"111110101",
  4847=>"000011011",
  4848=>"011000000",
  4849=>"000100000",
  4850=>"000000000",
  4851=>"110111111",
  4852=>"111111111",
  4853=>"101101101",
  4854=>"101111100",
  4855=>"111111111",
  4856=>"010111111",
  4857=>"100111101",
  4858=>"111100000",
  4859=>"111111111",
  4860=>"110111111",
  4861=>"111111001",
  4862=>"111110110",
  4863=>"000011001",
  4864=>"000000000",
  4865=>"111100100",
  4866=>"111010000",
  4867=>"111111111",
  4868=>"000100111",
  4869=>"100000011",
  4870=>"101111111",
  4871=>"111111001",
  4872=>"110010011",
  4873=>"000000000",
  4874=>"000110111",
  4875=>"111100100",
  4876=>"111111000",
  4877=>"111111111",
  4878=>"011101111",
  4879=>"000000000",
  4880=>"110111111",
  4881=>"000000000",
  4882=>"111111001",
  4883=>"000000000",
  4884=>"111000000",
  4885=>"000000111",
  4886=>"000000000",
  4887=>"000001011",
  4888=>"001000111",
  4889=>"000100101",
  4890=>"000000000",
  4891=>"000000000",
  4892=>"000100110",
  4893=>"001000111",
  4894=>"000000010",
  4895=>"100100111",
  4896=>"000000000",
  4897=>"000100111",
  4898=>"010111111",
  4899=>"101101000",
  4900=>"000000000",
  4901=>"111110110",
  4902=>"010100100",
  4903=>"000000100",
  4904=>"101111111",
  4905=>"111111111",
  4906=>"011000110",
  4907=>"111101101",
  4908=>"000000000",
  4909=>"000000100",
  4910=>"001000100",
  4911=>"000000101",
  4912=>"001000000",
  4913=>"111111011",
  4914=>"000101111",
  4915=>"111110000",
  4916=>"110000110",
  4917=>"111001000",
  4918=>"111111111",
  4919=>"000000000",
  4920=>"101000000",
  4921=>"001000001",
  4922=>"101000000",
  4923=>"111000000",
  4924=>"000000100",
  4925=>"100000100",
  4926=>"111111111",
  4927=>"000000111",
  4928=>"101100111",
  4929=>"111111000",
  4930=>"001000001",
  4931=>"000111111",
  4932=>"110111100",
  4933=>"000000100",
  4934=>"100100100",
  4935=>"000000001",
  4936=>"000000000",
  4937=>"111111111",
  4938=>"000000000",
  4939=>"110100100",
  4940=>"111111111",
  4941=>"111111110",
  4942=>"010001011",
  4943=>"001000000",
  4944=>"111111111",
  4945=>"000000011",
  4946=>"100100000",
  4947=>"110110110",
  4948=>"001001111",
  4949=>"011011011",
  4950=>"000000000",
  4951=>"111011011",
  4952=>"001111111",
  4953=>"000000000",
  4954=>"111111111",
  4955=>"000011001",
  4956=>"110000000",
  4957=>"111111111",
  4958=>"000000011",
  4959=>"100111000",
  4960=>"000000100",
  4961=>"000111111",
  4962=>"110100111",
  4963=>"111111101",
  4964=>"000000000",
  4965=>"001000000",
  4966=>"110000100",
  4967=>"011111111",
  4968=>"101101101",
  4969=>"100100000",
  4970=>"100100000",
  4971=>"111111100",
  4972=>"000100000",
  4973=>"110000000",
  4974=>"011000000",
  4975=>"111111111",
  4976=>"111111111",
  4977=>"000000000",
  4978=>"110110000",
  4979=>"111001000",
  4980=>"111111110",
  4981=>"111111111",
  4982=>"111001000",
  4983=>"111111110",
  4984=>"101110110",
  4985=>"111001111",
  4986=>"100000111",
  4987=>"111111111",
  4988=>"000000001",
  4989=>"001101011",
  4990=>"101000111",
  4991=>"000101111",
  4992=>"000000000",
  4993=>"111110000",
  4994=>"000000111",
  4995=>"000000000",
  4996=>"001000000",
  4997=>"000010011",
  4998=>"000000111",
  4999=>"111111001",
  5000=>"000000111",
  5001=>"100000000",
  5002=>"111111110",
  5003=>"111110000",
  5004=>"000000101",
  5005=>"000001000",
  5006=>"011011000",
  5007=>"001001011",
  5008=>"000000100",
  5009=>"100111111",
  5010=>"111111111",
  5011=>"000000000",
  5012=>"000110000",
  5013=>"011000010",
  5014=>"000000000",
  5015=>"000000010",
  5016=>"111000000",
  5017=>"100100111",
  5018=>"000111011",
  5019=>"000000110",
  5020=>"000111111",
  5021=>"111111111",
  5022=>"110111111",
  5023=>"000000101",
  5024=>"000000000",
  5025=>"111000000",
  5026=>"100101111",
  5027=>"000100111",
  5028=>"000001101",
  5029=>"111111111",
  5030=>"001000101",
  5031=>"111111111",
  5032=>"000000110",
  5033=>"101111111",
  5034=>"111110110",
  5035=>"111000000",
  5036=>"110111111",
  5037=>"111110110",
  5038=>"100100000",
  5039=>"000001011",
  5040=>"100100111",
  5041=>"000000001",
  5042=>"010110111",
  5043=>"000000101",
  5044=>"101101001",
  5045=>"011011111",
  5046=>"101000100",
  5047=>"000000000",
  5048=>"000000000",
  5049=>"000000000",
  5050=>"111111111",
  5051=>"000000000",
  5052=>"000000000",
  5053=>"000000000",
  5054=>"001110111",
  5055=>"100101100",
  5056=>"011011000",
  5057=>"000000111",
  5058=>"000001111",
  5059=>"000000000",
  5060=>"101100000",
  5061=>"011111101",
  5062=>"000000100",
  5063=>"000000111",
  5064=>"111001101",
  5065=>"011001001",
  5066=>"000000100",
  5067=>"000100000",
  5068=>"010000000",
  5069=>"000000000",
  5070=>"101111111",
  5071=>"111111111",
  5072=>"111000001",
  5073=>"111001101",
  5074=>"110000000",
  5075=>"111111101",
  5076=>"111111111",
  5077=>"000000000",
  5078=>"011011011",
  5079=>"001001001",
  5080=>"100000111",
  5081=>"000000000",
  5082=>"001001011",
  5083=>"000000000",
  5084=>"011111111",
  5085=>"000001011",
  5086=>"000000001",
  5087=>"000001001",
  5088=>"000000000",
  5089=>"000110110",
  5090=>"001000000",
  5091=>"011000000",
  5092=>"000000011",
  5093=>"000000000",
  5094=>"110000000",
  5095=>"111111000",
  5096=>"000000000",
  5097=>"000001000",
  5098=>"100110110",
  5099=>"010111111",
  5100=>"111000101",
  5101=>"111100000",
  5102=>"010010111",
  5103=>"111111111",
  5104=>"000000000",
  5105=>"000000000",
  5106=>"101100111",
  5107=>"100111111",
  5108=>"000000010",
  5109=>"000110111",
  5110=>"111111111",
  5111=>"011011011",
  5112=>"000000011",
  5113=>"101000000",
  5114=>"110111101",
  5115=>"111111111",
  5116=>"111110000",
  5117=>"101111111",
  5118=>"111111111",
  5119=>"111111111",
  5120=>"100110110",
  5121=>"111110111",
  5122=>"111111111",
  5123=>"111111111",
  5124=>"000000000",
  5125=>"000101100",
  5126=>"001000001",
  5127=>"111000111",
  5128=>"000000011",
  5129=>"100110110",
  5130=>"001000000",
  5131=>"111111111",
  5132=>"000000000",
  5133=>"111111111",
  5134=>"111000000",
  5135=>"000000111",
  5136=>"111010000",
  5137=>"000000111",
  5138=>"000001001",
  5139=>"101111111",
  5140=>"100010000",
  5141=>"111111000",
  5142=>"111111111",
  5143=>"110111111",
  5144=>"000000010",
  5145=>"001011011",
  5146=>"111000110",
  5147=>"001000100",
  5148=>"111111110",
  5149=>"000101111",
  5150=>"010111110",
  5151=>"111111001",
  5152=>"000001101",
  5153=>"110111110",
  5154=>"000000000",
  5155=>"011011111",
  5156=>"000010011",
  5157=>"111111111",
  5158=>"001000101",
  5159=>"001011111",
  5160=>"111111111",
  5161=>"110000000",
  5162=>"100100000",
  5163=>"011111100",
  5164=>"001001001",
  5165=>"111111000",
  5166=>"111100111",
  5167=>"111111111",
  5168=>"000000000",
  5169=>"010001001",
  5170=>"011111011",
  5171=>"011110111",
  5172=>"101111011",
  5173=>"000000000",
  5174=>"000000001",
  5175=>"111111000",
  5176=>"111111111",
  5177=>"001111111",
  5178=>"000000000",
  5179=>"111000000",
  5180=>"111101010",
  5181=>"111111111",
  5182=>"011011001",
  5183=>"000000000",
  5184=>"000000000",
  5185=>"000001000",
  5186=>"111011000",
  5187=>"000000000",
  5188=>"010110111",
  5189=>"011011000",
  5190=>"000000111",
  5191=>"000000000",
  5192=>"111011110",
  5193=>"000000000",
  5194=>"111001001",
  5195=>"110111111",
  5196=>"000001010",
  5197=>"001000001",
  5198=>"000000000",
  5199=>"110000000",
  5200=>"000000000",
  5201=>"101000000",
  5202=>"000100000",
  5203=>"111110010",
  5204=>"000101100",
  5205=>"000000011",
  5206=>"010010001",
  5207=>"001000000",
  5208=>"111101111",
  5209=>"000000000",
  5210=>"000001000",
  5211=>"000000000",
  5212=>"111011111",
  5213=>"000111111",
  5214=>"000000111",
  5215=>"111111111",
  5216=>"001100110",
  5217=>"000000001",
  5218=>"000000111",
  5219=>"111001000",
  5220=>"111111000",
  5221=>"111111001",
  5222=>"111111000",
  5223=>"000110101",
  5224=>"111111000",
  5225=>"111111111",
  5226=>"000000011",
  5227=>"000000111",
  5228=>"111111110",
  5229=>"111110110",
  5230=>"111110000",
  5231=>"001111111",
  5232=>"010100100",
  5233=>"100000001",
  5234=>"111111001",
  5235=>"111110000",
  5236=>"000000000",
  5237=>"111111011",
  5238=>"000000011",
  5239=>"000000000",
  5240=>"111111111",
  5241=>"011111111",
  5242=>"000000000",
  5243=>"000110110",
  5244=>"100100000",
  5245=>"000000000",
  5246=>"111111000",
  5247=>"000000000",
  5248=>"001000011",
  5249=>"111111111",
  5250=>"110000000",
  5251=>"000000001",
  5252=>"000000000",
  5253=>"110110000",
  5254=>"001101111",
  5255=>"010111001",
  5256=>"111111100",
  5257=>"100000000",
  5258=>"000000000",
  5259=>"000000000",
  5260=>"000000000",
  5261=>"000000000",
  5262=>"000011111",
  5263=>"111001001",
  5264=>"001011001",
  5265=>"000000110",
  5266=>"000000000",
  5267=>"011001000",
  5268=>"111111111",
  5269=>"000100100",
  5270=>"111111111",
  5271=>"000001001",
  5272=>"000000000",
  5273=>"011111111",
  5274=>"111011010",
  5275=>"011011011",
  5276=>"101000000",
  5277=>"111011000",
  5278=>"000111110",
  5279=>"100000000",
  5280=>"000000000",
  5281=>"110110110",
  5282=>"000000001",
  5283=>"111000001",
  5284=>"001000100",
  5285=>"011000000",
  5286=>"000111111",
  5287=>"100110011",
  5288=>"111011010",
  5289=>"011101111",
  5290=>"100111111",
  5291=>"111111000",
  5292=>"111010110",
  5293=>"000000000",
  5294=>"100111111",
  5295=>"111111111",
  5296=>"011110000",
  5297=>"100111001",
  5298=>"111111111",
  5299=>"000001111",
  5300=>"000100111",
  5301=>"111111000",
  5302=>"010000101",
  5303=>"111011111",
  5304=>"111011111",
  5305=>"000000011",
  5306=>"101000000",
  5307=>"000000000",
  5308=>"000101101",
  5309=>"101101000",
  5310=>"010000000",
  5311=>"011000000",
  5312=>"000000000",
  5313=>"000000111",
  5314=>"001000000",
  5315=>"000111111",
  5316=>"100111110",
  5317=>"110111111",
  5318=>"001000000",
  5319=>"110000001",
  5320=>"111110010",
  5321=>"110000111",
  5322=>"000000000",
  5323=>"110000011",
  5324=>"000001011",
  5325=>"110110110",
  5326=>"011111111",
  5327=>"111010000",
  5328=>"000100111",
  5329=>"000000010",
  5330=>"011000001",
  5331=>"000000000",
  5332=>"011001000",
  5333=>"111111110",
  5334=>"000000111",
  5335=>"110100110",
  5336=>"110110110",
  5337=>"011000000",
  5338=>"100000000",
  5339=>"011111111",
  5340=>"101111111",
  5341=>"100000000",
  5342=>"000000000",
  5343=>"100000000",
  5344=>"000101111",
  5345=>"000000111",
  5346=>"000000100",
  5347=>"000000000",
  5348=>"001000000",
  5349=>"000000001",
  5350=>"000100111",
  5351=>"111000000",
  5352=>"100110000",
  5353=>"000000000",
  5354=>"110111111",
  5355=>"010010010",
  5356=>"111001000",
  5357=>"000000101",
  5358=>"000000100",
  5359=>"110111111",
  5360=>"111111001",
  5361=>"000000000",
  5362=>"111111001",
  5363=>"110111111",
  5364=>"111011000",
  5365=>"000011111",
  5366=>"000110111",
  5367=>"110111000",
  5368=>"000000000",
  5369=>"111000000",
  5370=>"000000001",
  5371=>"000001111",
  5372=>"000001111",
  5373=>"110100100",
  5374=>"000000000",
  5375=>"111110111",
  5376=>"000000000",
  5377=>"010011001",
  5378=>"000000000",
  5379=>"110000000",
  5380=>"111000000",
  5381=>"000000000",
  5382=>"000111111",
  5383=>"000001001",
  5384=>"000110111",
  5385=>"000000000",
  5386=>"000000000",
  5387=>"111111111",
  5388=>"111100111",
  5389=>"000000111",
  5390=>"111111000",
  5391=>"000000111",
  5392=>"000010000",
  5393=>"000000001",
  5394=>"100100111",
  5395=>"111111001",
  5396=>"000000000",
  5397=>"011000000",
  5398=>"100000011",
  5399=>"101111111",
  5400=>"111111001",
  5401=>"001011111",
  5402=>"111111100",
  5403=>"000001111",
  5404=>"010111011",
  5405=>"000000000",
  5406=>"001000000",
  5407=>"111111101",
  5408=>"010000011",
  5409=>"000000000",
  5410=>"111010000",
  5411=>"111111000",
  5412=>"110111111",
  5413=>"101111000",
  5414=>"000000011",
  5415=>"100110111",
  5416=>"010110111",
  5417=>"001000000",
  5418=>"110000000",
  5419=>"111111100",
  5420=>"111110100",
  5421=>"100110000",
  5422=>"111000000",
  5423=>"111111111",
  5424=>"001000000",
  5425=>"110111111",
  5426=>"000001111",
  5427=>"100110110",
  5428=>"111000101",
  5429=>"101011111",
  5430=>"111000000",
  5431=>"000111000",
  5432=>"011111110",
  5433=>"111000111",
  5434=>"111111001",
  5435=>"111011101",
  5436=>"011000000",
  5437=>"000110111",
  5438=>"010111111",
  5439=>"111011000",
  5440=>"111111111",
  5441=>"101111000",
  5442=>"000111111",
  5443=>"000000111",
  5444=>"000001111",
  5445=>"111111111",
  5446=>"011011000",
  5447=>"000000001",
  5448=>"000000000",
  5449=>"000110111",
  5450=>"000000000",
  5451=>"010011111",
  5452=>"111110000",
  5453=>"000000000",
  5454=>"111001111",
  5455=>"100100110",
  5456=>"001001000",
  5457=>"000000000",
  5458=>"100100001",
  5459=>"000000000",
  5460=>"111111000",
  5461=>"011011011",
  5462=>"000000001",
  5463=>"000001111",
  5464=>"100100000",
  5465=>"111111010",
  5466=>"111111111",
  5467=>"000000000",
  5468=>"110111111",
  5469=>"111111000",
  5470=>"111111111",
  5471=>"111011111",
  5472=>"111110110",
  5473=>"000000000",
  5474=>"110111111",
  5475=>"000000000",
  5476=>"111111000",
  5477=>"000000000",
  5478=>"100111111",
  5479=>"111001111",
  5480=>"100100000",
  5481=>"111111000",
  5482=>"000100111",
  5483=>"111111111",
  5484=>"010000000",
  5485=>"010000110",
  5486=>"100000101",
  5487=>"000110000",
  5488=>"111000000",
  5489=>"011111111",
  5490=>"010010110",
  5491=>"000000001",
  5492=>"000000000",
  5493=>"111000100",
  5494=>"111011000",
  5495=>"111111000",
  5496=>"000000111",
  5497=>"000000000",
  5498=>"111000000",
  5499=>"000000110",
  5500=>"011110111",
  5501=>"111110000",
  5502=>"001011001",
  5503=>"000000011",
  5504=>"000000011",
  5505=>"110110111",
  5506=>"000011111",
  5507=>"000000000",
  5508=>"000000000",
  5509=>"000100110",
  5510=>"000000000",
  5511=>"111111111",
  5512=>"000000000",
  5513=>"111110111",
  5514=>"110111001",
  5515=>"000000000",
  5516=>"111001111",
  5517=>"000111111",
  5518=>"000000000",
  5519=>"000000001",
  5520=>"000011110",
  5521=>"111111001",
  5522=>"000100100",
  5523=>"000000000",
  5524=>"000111111",
  5525=>"000000000",
  5526=>"111111010",
  5527=>"000000011",
  5528=>"111111000",
  5529=>"000000000",
  5530=>"000110111",
  5531=>"000000100",
  5532=>"000000000",
  5533=>"011011000",
  5534=>"100101101",
  5535=>"001001000",
  5536=>"000000000",
  5537=>"010100100",
  5538=>"111111111",
  5539=>"011111111",
  5540=>"000000001",
  5541=>"101111000",
  5542=>"111111111",
  5543=>"000000000",
  5544=>"011001001",
  5545=>"110000000",
  5546=>"000000000",
  5547=>"110111111",
  5548=>"011111111",
  5549=>"000101111",
  5550=>"000000100",
  5551=>"000000111",
  5552=>"000010111",
  5553=>"000000000",
  5554=>"000000000",
  5555=>"010111010",
  5556=>"110000111",
  5557=>"001000101",
  5558=>"111001111",
  5559=>"000000111",
  5560=>"000000000",
  5561=>"111111111",
  5562=>"111111110",
  5563=>"010011010",
  5564=>"110110111",
  5565=>"000000000",
  5566=>"001000000",
  5567=>"010011011",
  5568=>"111011111",
  5569=>"111111111",
  5570=>"001000001",
  5571=>"011001111",
  5572=>"000000011",
  5573=>"101111011",
  5574=>"110000000",
  5575=>"000000001",
  5576=>"000000000",
  5577=>"000000000",
  5578=>"110000000",
  5579=>"100101100",
  5580=>"000000111",
  5581=>"111111000",
  5582=>"011111111",
  5583=>"000110111",
  5584=>"000111111",
  5585=>"100101001",
  5586=>"111111111",
  5587=>"111111111",
  5588=>"111111010",
  5589=>"000000000",
  5590=>"101000000",
  5591=>"000000000",
  5592=>"011011001",
  5593=>"111000000",
  5594=>"111111111",
  5595=>"111001000",
  5596=>"000100110",
  5597=>"110000000",
  5598=>"111111000",
  5599=>"110100000",
  5600=>"110111111",
  5601=>"000111111",
  5602=>"101111111",
  5603=>"111111111",
  5604=>"111010000",
  5605=>"111111000",
  5606=>"000000000",
  5607=>"100000100",
  5608=>"000000000",
  5609=>"110110110",
  5610=>"100100111",
  5611=>"011111111",
  5612=>"111111111",
  5613=>"000000111",
  5614=>"111000100",
  5615=>"111111111",
  5616=>"000000001",
  5617=>"000000111",
  5618=>"000111111",
  5619=>"000000000",
  5620=>"111111111",
  5621=>"001000000",
  5622=>"000110110",
  5623=>"111111110",
  5624=>"100111111",
  5625=>"000000000",
  5626=>"000000000",
  5627=>"000000001",
  5628=>"100111111",
  5629=>"001000001",
  5630=>"000000000",
  5631=>"111111111",
  5632=>"001000100",
  5633=>"001001001",
  5634=>"000101101",
  5635=>"000000000",
  5636=>"000000000",
  5637=>"000110110",
  5638=>"000000000",
  5639=>"111111111",
  5640=>"001000000",
  5641=>"001001011",
  5642=>"011010010",
  5643=>"101000001",
  5644=>"110110100",
  5645=>"000000000",
  5646=>"001111111",
  5647=>"000000001",
  5648=>"011011010",
  5649=>"010011001",
  5650=>"000000111",
  5651=>"000000000",
  5652=>"100101001",
  5653=>"000111111",
  5654=>"000001001",
  5655=>"110110000",
  5656=>"000000000",
  5657=>"010000010",
  5658=>"010000000",
  5659=>"000000100",
  5660=>"111011001",
  5661=>"001000001",
  5662=>"110111011",
  5663=>"001111101",
  5664=>"110110110",
  5665=>"100000100",
  5666=>"000001111",
  5667=>"101000000",
  5668=>"110111111",
  5669=>"100101011",
  5670=>"000001011",
  5671=>"111001000",
  5672=>"000110110",
  5673=>"100100101",
  5674=>"011011001",
  5675=>"100101111",
  5676=>"111111111",
  5677=>"111111100",
  5678=>"001000111",
  5679=>"110000011",
  5680=>"111101001",
  5681=>"110110110",
  5682=>"100000001",
  5683=>"010110110",
  5684=>"110110110",
  5685=>"000010011",
  5686=>"111010011",
  5687=>"101001011",
  5688=>"001101100",
  5689=>"011011111",
  5690=>"000011111",
  5691=>"000000000",
  5692=>"001001001",
  5693=>"010011011",
  5694=>"110110110",
  5695=>"111011100",
  5696=>"100001101",
  5697=>"110100100",
  5698=>"000101101",
  5699=>"001000001",
  5700=>"111011011",
  5701=>"000000001",
  5702=>"000111110",
  5703=>"000000000",
  5704=>"110000000",
  5705=>"000001111",
  5706=>"111111111",
  5707=>"111101101",
  5708=>"000101111",
  5709=>"111111100",
  5710=>"110110011",
  5711=>"001000011",
  5712=>"000011010",
  5713=>"111111111",
  5714=>"111111000",
  5715=>"110110110",
  5716=>"111110100",
  5717=>"111101000",
  5718=>"000000101",
  5719=>"110000000",
  5720=>"110110111",
  5721=>"001001101",
  5722=>"001000000",
  5723=>"011011101",
  5724=>"000000010",
  5725=>"000000111",
  5726=>"000000110",
  5727=>"110110100",
  5728=>"100100110",
  5729=>"000000000",
  5730=>"001000010",
  5731=>"011111111",
  5732=>"111111000",
  5733=>"100000000",
  5734=>"000000110",
  5735=>"010111111",
  5736=>"000000000",
  5737=>"111011011",
  5738=>"001001101",
  5739=>"000000111",
  5740=>"000011111",
  5741=>"110111111",
  5742=>"001001001",
  5743=>"000000001",
  5744=>"111000000",
  5745=>"000001111",
  5746=>"010010010",
  5747=>"000001011",
  5748=>"110111010",
  5749=>"000111111",
  5750=>"111111101",
  5751=>"000000000",
  5752=>"000001101",
  5753=>"000001011",
  5754=>"111000100",
  5755=>"000000000",
  5756=>"111111010",
  5757=>"100001101",
  5758=>"000000000",
  5759=>"001111111",
  5760=>"101101000",
  5761=>"100000001",
  5762=>"101100111",
  5763=>"110110110",
  5764=>"010010011",
  5765=>"101100101",
  5766=>"001111101",
  5767=>"001000011",
  5768=>"000000110",
  5769=>"101001011",
  5770=>"111111011",
  5771=>"000000011",
  5772=>"000000000",
  5773=>"101101111",
  5774=>"000000000",
  5775=>"000000000",
  5776=>"111011011",
  5777=>"110110110",
  5778=>"111001011",
  5779=>"001001001",
  5780=>"011101111",
  5781=>"111101000",
  5782=>"101001000",
  5783=>"111111101",
  5784=>"000000110",
  5785=>"001011001",
  5786=>"111001101",
  5787=>"111011000",
  5788=>"111101100",
  5789=>"001001001",
  5790=>"101111101",
  5791=>"100000001",
  5792=>"000001011",
  5793=>"000100010",
  5794=>"011010010",
  5795=>"111111000",
  5796=>"001000000",
  5797=>"001011111",
  5798=>"110000000",
  5799=>"110110111",
  5800=>"000000101",
  5801=>"001000101",
  5802=>"101101101",
  5803=>"010110000",
  5804=>"000000000",
  5805=>"011111111",
  5806=>"111111111",
  5807=>"000000000",
  5808=>"000101111",
  5809=>"000010111",
  5810=>"110010010",
  5811=>"111010000",
  5812=>"110011010",
  5813=>"111111111",
  5814=>"010011011",
  5815=>"111111101",
  5816=>"101101001",
  5817=>"010111111",
  5818=>"001001001",
  5819=>"111001100",
  5820=>"101101001",
  5821=>"110111111",
  5822=>"110111111",
  5823=>"000001000",
  5824=>"010010000",
  5825=>"000000100",
  5826=>"110111000",
  5827=>"111110111",
  5828=>"111111110",
  5829=>"000001101",
  5830=>"001000000",
  5831=>"110110100",
  5832=>"000001111",
  5833=>"001001001",
  5834=>"000000000",
  5835=>"110000000",
  5836=>"000000000",
  5837=>"000000001",
  5838=>"001000001",
  5839=>"000000000",
  5840=>"111111110",
  5841=>"000000010",
  5842=>"110000000",
  5843=>"000000000",
  5844=>"000000000",
  5845=>"111110100",
  5846=>"000000001",
  5847=>"000010011",
  5848=>"010010011",
  5849=>"110110000",
  5850=>"100111111",
  5851=>"000000101",
  5852=>"001101101",
  5853=>"000000000",
  5854=>"010000000",
  5855=>"101001101",
  5856=>"011000110",
  5857=>"010000000",
  5858=>"101111111",
  5859=>"101101101",
  5860=>"100101100",
  5861=>"000000110",
  5862=>"000000010",
  5863=>"000000100",
  5864=>"100000000",
  5865=>"111100111",
  5866=>"101001000",
  5867=>"100111111",
  5868=>"111001001",
  5869=>"101101001",
  5870=>"111011010",
  5871=>"001101101",
  5872=>"100101111",
  5873=>"000000001",
  5874=>"101101111",
  5875=>"101001101",
  5876=>"001001101",
  5877=>"001011011",
  5878=>"110111011",
  5879=>"000110110",
  5880=>"111001111",
  5881=>"111001001",
  5882=>"100110110",
  5883=>"111010010",
  5884=>"111101000",
  5885=>"111011001",
  5886=>"001101100",
  5887=>"000000101",
  5888=>"111000000",
  5889=>"001101001",
  5890=>"110110000",
  5891=>"000000001",
  5892=>"001111111",
  5893=>"011001011",
  5894=>"111111111",
  5895=>"111101111",
  5896=>"111111011",
  5897=>"111111111",
  5898=>"111111001",
  5899=>"000001000",
  5900=>"110110110",
  5901=>"110101101",
  5902=>"000101100",
  5903=>"000110010",
  5904=>"000100111",
  5905=>"111001000",
  5906=>"000000000",
  5907=>"001001010",
  5908=>"000001000",
  5909=>"000000011",
  5910=>"011010110",
  5911=>"011111111",
  5912=>"110110110",
  5913=>"001001000",
  5914=>"001000110",
  5915=>"000000111",
  5916=>"010000110",
  5917=>"000000000",
  5918=>"110111111",
  5919=>"000000000",
  5920=>"000000000",
  5921=>"010110011",
  5922=>"011011010",
  5923=>"000000110",
  5924=>"001001001",
  5925=>"011010110",
  5926=>"110111111",
  5927=>"000000000",
  5928=>"011111011",
  5929=>"100000111",
  5930=>"110110010",
  5931=>"111011000",
  5932=>"101111111",
  5933=>"000110001",
  5934=>"000110000",
  5935=>"000000111",
  5936=>"100110111",
  5937=>"000000011",
  5938=>"110100101",
  5939=>"111111111",
  5940=>"111111110",
  5941=>"110010011",
  5942=>"100101101",
  5943=>"110110111",
  5944=>"010110100",
  5945=>"101001101",
  5946=>"000000000",
  5947=>"011111011",
  5948=>"101101111",
  5949=>"000010000",
  5950=>"111111101",
  5951=>"111101100",
  5952=>"011011000",
  5953=>"111101001",
  5954=>"110111110",
  5955=>"110010000",
  5956=>"100100110",
  5957=>"000000100",
  5958=>"111110111",
  5959=>"111011111",
  5960=>"000011011",
  5961=>"101111101",
  5962=>"101111111",
  5963=>"110110110",
  5964=>"001001001",
  5965=>"001000011",
  5966=>"000000000",
  5967=>"110110100",
  5968=>"110110110",
  5969=>"001100111",
  5970=>"010000111",
  5971=>"111100101",
  5972=>"000010110",
  5973=>"011011011",
  5974=>"101000101",
  5975=>"100010010",
  5976=>"100000000",
  5977=>"100100000",
  5978=>"111100010",
  5979=>"000111111",
  5980=>"001000000",
  5981=>"111001000",
  5982=>"110110110",
  5983=>"110000110",
  5984=>"111101001",
  5985=>"111111111",
  5986=>"010010110",
  5987=>"100100100",
  5988=>"110111111",
  5989=>"111000000",
  5990=>"010100000",
  5991=>"010010010",
  5992=>"111110111",
  5993=>"111110110",
  5994=>"000000000",
  5995=>"001001001",
  5996=>"110110110",
  5997=>"001101111",
  5998=>"001111111",
  5999=>"011000000",
  6000=>"100111111",
  6001=>"111001011",
  6002=>"111110110",
  6003=>"000000000",
  6004=>"111111101",
  6005=>"111111111",
  6006=>"111111111",
  6007=>"000000110",
  6008=>"111111101",
  6009=>"001111001",
  6010=>"110110010",
  6011=>"001001001",
  6012=>"001000100",
  6013=>"111111110",
  6014=>"000000000",
  6015=>"111000000",
  6016=>"110010010",
  6017=>"110110010",
  6018=>"011010000",
  6019=>"000000000",
  6020=>"101101101",
  6021=>"000100101",
  6022=>"000000001",
  6023=>"101110111",
  6024=>"000101000",
  6025=>"110100100",
  6026=>"011111010",
  6027=>"000101101",
  6028=>"001011000",
  6029=>"011011011",
  6030=>"111011010",
  6031=>"010010000",
  6032=>"110111111",
  6033=>"111011111",
  6034=>"111110110",
  6035=>"001001001",
  6036=>"111101111",
  6037=>"100111101",
  6038=>"110110100",
  6039=>"111110110",
  6040=>"101101111",
  6041=>"011011111",
  6042=>"101001111",
  6043=>"000000001",
  6044=>"000000000",
  6045=>"111011011",
  6046=>"111001001",
  6047=>"000111000",
  6048=>"010111111",
  6049=>"000001011",
  6050=>"110000101",
  6051=>"100101111",
  6052=>"111100001",
  6053=>"111101110",
  6054=>"000010010",
  6055=>"111111110",
  6056=>"111011111",
  6057=>"000001111",
  6058=>"001000100",
  6059=>"100100001",
  6060=>"101101101",
  6061=>"001101101",
  6062=>"001001111",
  6063=>"100101101",
  6064=>"001101111",
  6065=>"111000000",
  6066=>"110110011",
  6067=>"010000000",
  6068=>"110011001",
  6069=>"100000000",
  6070=>"001001111",
  6071=>"110110110",
  6072=>"001011011",
  6073=>"110110111",
  6074=>"111110110",
  6075=>"100101000",
  6076=>"001001101",
  6077=>"010000000",
  6078=>"111110110",
  6079=>"011010010",
  6080=>"000000000",
  6081=>"001001101",
  6082=>"000000010",
  6083=>"001000001",
  6084=>"111111111",
  6085=>"110100111",
  6086=>"110110110",
  6087=>"111101101",
  6088=>"100000000",
  6089=>"010011111",
  6090=>"000000110",
  6091=>"111111001",
  6092=>"100010000",
  6093=>"110110010",
  6094=>"111010010",
  6095=>"101111111",
  6096=>"111110110",
  6097=>"100000000",
  6098=>"111111111",
  6099=>"000000000",
  6100=>"111110111",
  6101=>"000000000",
  6102=>"100010011",
  6103=>"011011011",
  6104=>"111111111",
  6105=>"110111101",
  6106=>"101001000",
  6107=>"101101001",
  6108=>"111100000",
  6109=>"110000000",
  6110=>"100100000",
  6111=>"011111111",
  6112=>"000001001",
  6113=>"000000000",
  6114=>"101101001",
  6115=>"010010001",
  6116=>"110000111",
  6117=>"001000000",
  6118=>"011010010",
  6119=>"000001001",
  6120=>"000000000",
  6121=>"111111011",
  6122=>"000110111",
  6123=>"001001101",
  6124=>"100011001",
  6125=>"110110110",
  6126=>"010000000",
  6127=>"101001101",
  6128=>"101101111",
  6129=>"111000011",
  6130=>"101101011",
  6131=>"110110110",
  6132=>"100101011",
  6133=>"001101001",
  6134=>"110111101",
  6135=>"011011110",
  6136=>"110000000",
  6137=>"110000110",
  6138=>"111111111",
  6139=>"110110010",
  6140=>"001111011",
  6141=>"111110001",
  6142=>"000000111",
  6143=>"111111111",
  6144=>"110000000",
  6145=>"110111010",
  6146=>"000000000",
  6147=>"000000000",
  6148=>"111110100",
  6149=>"001001000",
  6150=>"001101111",
  6151=>"111111111",
  6152=>"011111001",
  6153=>"111111111",
  6154=>"110110111",
  6155=>"111011111",
  6156=>"000000100",
  6157=>"100000000",
  6158=>"010001000",
  6159=>"111111111",
  6160=>"111111111",
  6161=>"111111101",
  6162=>"111111111",
  6163=>"111111111",
  6164=>"111111101",
  6165=>"100110110",
  6166=>"111011011",
  6167=>"110110110",
  6168=>"101101111",
  6169=>"101111111",
  6170=>"110100100",
  6171=>"000000001",
  6172=>"111111111",
  6173=>"000111111",
  6174=>"111111111",
  6175=>"100000111",
  6176=>"111111111",
  6177=>"111101000",
  6178=>"000000000",
  6179=>"110000000",
  6180=>"000000001",
  6181=>"001010111",
  6182=>"110100001",
  6183=>"000100111",
  6184=>"111111111",
  6185=>"000000000",
  6186=>"111111111",
  6187=>"111111111",
  6188=>"000000001",
  6189=>"000000000",
  6190=>"110010110",
  6191=>"000000001",
  6192=>"100110111",
  6193=>"111011011",
  6194=>"011111111",
  6195=>"111110000",
  6196=>"100110100",
  6197=>"000100111",
  6198=>"000000000",
  6199=>"111000111",
  6200=>"101001001",
  6201=>"101001011",
  6202=>"000011111",
  6203=>"011111000",
  6204=>"001000000",
  6205=>"100000000",
  6206=>"111011111",
  6207=>"111111111",
  6208=>"011011011",
  6209=>"000011001",
  6210=>"001111111",
  6211=>"100000000",
  6212=>"000000000",
  6213=>"011111111",
  6214=>"000110000",
  6215=>"100100101",
  6216=>"000000000",
  6217=>"100110111",
  6218=>"111111111",
  6219=>"111101000",
  6220=>"111111111",
  6221=>"101000000",
  6222=>"100000100",
  6223=>"000000000",
  6224=>"111111111",
  6225=>"001011000",
  6226=>"111100100",
  6227=>"001111101",
  6228=>"001001001",
  6229=>"111111011",
  6230=>"111001001",
  6231=>"110111111",
  6232=>"111111001",
  6233=>"000000000",
  6234=>"100000000",
  6235=>"111011111",
  6236=>"011111111",
  6237=>"111111000",
  6238=>"111111111",
  6239=>"001001000",
  6240=>"000000000",
  6241=>"110110111",
  6242=>"111110110",
  6243=>"110111111",
  6244=>"111011110",
  6245=>"001000100",
  6246=>"111111111",
  6247=>"001000000",
  6248=>"111111011",
  6249=>"111111111",
  6250=>"111111111",
  6251=>"111111110",
  6252=>"100100100",
  6253=>"100000000",
  6254=>"111111111",
  6255=>"111011000",
  6256=>"100000000",
  6257=>"000000000",
  6258=>"111111111",
  6259=>"000000000",
  6260=>"000101100",
  6261=>"011111111",
  6262=>"000000000",
  6263=>"001101111",
  6264=>"111111011",
  6265=>"111111111",
  6266=>"001000000",
  6267=>"101001011",
  6268=>"000000000",
  6269=>"000111111",
  6270=>"011111111",
  6271=>"000000000",
  6272=>"111111111",
  6273=>"100000111",
  6274=>"110010010",
  6275=>"110001111",
  6276=>"111011011",
  6277=>"000000000",
  6278=>"000000000",
  6279=>"101000010",
  6280=>"000000100",
  6281=>"000100100",
  6282=>"111111111",
  6283=>"100111111",
  6284=>"011111011",
  6285=>"100000000",
  6286=>"100101111",
  6287=>"110111011",
  6288=>"011011111",
  6289=>"001110110",
  6290=>"111111000",
  6291=>"000000100",
  6292=>"000001000",
  6293=>"000000010",
  6294=>"111011100",
  6295=>"000000100",
  6296=>"001001001",
  6297=>"000001000",
  6298=>"110110011",
  6299=>"001011000",
  6300=>"111110111",
  6301=>"111001010",
  6302=>"111111000",
  6303=>"111111111",
  6304=>"110000000",
  6305=>"100001000",
  6306=>"011011010",
  6307=>"000000000",
  6308=>"010111101",
  6309=>"100000011",
  6310=>"111110010",
  6311=>"110100100",
  6312=>"000110111",
  6313=>"111111111",
  6314=>"001001000",
  6315=>"000000111",
  6316=>"101000000",
  6317=>"100000000",
  6318=>"110111011",
  6319=>"000000000",
  6320=>"111111111",
  6321=>"110100111",
  6322=>"111110110",
  6323=>"000000000",
  6324=>"001011000",
  6325=>"111111011",
  6326=>"111111111",
  6327=>"111011011",
  6328=>"100100101",
  6329=>"000000001",
  6330=>"111011111",
  6331=>"000000000",
  6332=>"111110110",
  6333=>"001000111",
  6334=>"010110000",
  6335=>"111001001",
  6336=>"111110110",
  6337=>"100000000",
  6338=>"111110011",
  6339=>"000000000",
  6340=>"000000100",
  6341=>"110110110",
  6342=>"001001111",
  6343=>"111111111",
  6344=>"000000110",
  6345=>"100110100",
  6346=>"011010000",
  6347=>"111111111",
  6348=>"100000000",
  6349=>"100110110",
  6350=>"111111011",
  6351=>"000000000",
  6352=>"000111111",
  6353=>"011011000",
  6354=>"111011011",
  6355=>"111101111",
  6356=>"001001001",
  6357=>"100000111",
  6358=>"111010000",
  6359=>"011001000",
  6360=>"001001000",
  6361=>"111111111",
  6362=>"111111111",
  6363=>"000000000",
  6364=>"100100000",
  6365=>"100100000",
  6366=>"000000000",
  6367=>"111111111",
  6368=>"000000000",
  6369=>"000111010",
  6370=>"111110110",
  6371=>"100000000",
  6372=>"001000000",
  6373=>"000110000",
  6374=>"001001011",
  6375=>"111111111",
  6376=>"111111111",
  6377=>"100001111",
  6378=>"000000001",
  6379=>"111111111",
  6380=>"111111111",
  6381=>"100000110",
  6382=>"001000101",
  6383=>"011111011",
  6384=>"111001001",
  6385=>"101000100",
  6386=>"001000111",
  6387=>"111100001",
  6388=>"000000000",
  6389=>"000000000",
  6390=>"000000000",
  6391=>"000000000",
  6392=>"000000000",
  6393=>"100000000",
  6394=>"000000000",
  6395=>"000100100",
  6396=>"101111111",
  6397=>"011000000",
  6398=>"111000000",
  6399=>"000100000",
  6400=>"100100000",
  6401=>"111001111",
  6402=>"100100100",
  6403=>"111001000",
  6404=>"110000111",
  6405=>"000011000",
  6406=>"000000000",
  6407=>"101111111",
  6408=>"100100111",
  6409=>"000001111",
  6410=>"111111111",
  6411=>"000001001",
  6412=>"100000000",
  6413=>"111111111",
  6414=>"101101011",
  6415=>"000100111",
  6416=>"101010111",
  6417=>"100000000",
  6418=>"011111100",
  6419=>"111111111",
  6420=>"001011001",
  6421=>"000000000",
  6422=>"100101111",
  6423=>"101101101",
  6424=>"110001111",
  6425=>"111111011",
  6426=>"110000100",
  6427=>"000000011",
  6428=>"111111110",
  6429=>"110000000",
  6430=>"001111011",
  6431=>"110000000",
  6432=>"000000000",
  6433=>"111100000",
  6434=>"001111111",
  6435=>"000000000",
  6436=>"001111100",
  6437=>"000001100",
  6438=>"100000001",
  6439=>"000111111",
  6440=>"000111111",
  6441=>"000000000",
  6442=>"100100101",
  6443=>"111111111",
  6444=>"000001111",
  6445=>"100100110",
  6446=>"111010000",
  6447=>"000000000",
  6448=>"011011001",
  6449=>"111111111",
  6450=>"000000000",
  6451=>"111110010",
  6452=>"110000000",
  6453=>"000110100",
  6454=>"111100110",
  6455=>"111110110",
  6456=>"010010010",
  6457=>"111111110",
  6458=>"000000011",
  6459=>"110000101",
  6460=>"111111111",
  6461=>"100000000",
  6462=>"001011011",
  6463=>"101110011",
  6464=>"111000000",
  6465=>"000001001",
  6466=>"100000000",
  6467=>"000110100",
  6468=>"001111000",
  6469=>"111111111",
  6470=>"100111111",
  6471=>"100100100",
  6472=>"111010010",
  6473=>"011000000",
  6474=>"111100000",
  6475=>"000010010",
  6476=>"001001000",
  6477=>"001011001",
  6478=>"100100111",
  6479=>"000100100",
  6480=>"000000000",
  6481=>"111001100",
  6482=>"001111111",
  6483=>"111111111",
  6484=>"110111111",
  6485=>"000010011",
  6486=>"000000111",
  6487=>"000000000",
  6488=>"111100111",
  6489=>"000000000",
  6490=>"100111111",
  6491=>"010010010",
  6492=>"101111011",
  6493=>"000000000",
  6494=>"011011000",
  6495=>"000000000",
  6496=>"011001000",
  6497=>"111101100",
  6498=>"000000001",
  6499=>"000000100",
  6500=>"000000000",
  6501=>"001000000",
  6502=>"110100010",
  6503=>"101001000",
  6504=>"111101101",
  6505=>"001000110",
  6506=>"111111110",
  6507=>"000000000",
  6508=>"000011011",
  6509=>"010000100",
  6510=>"011111111",
  6511=>"111111111",
  6512=>"111111111",
  6513=>"011000011",
  6514=>"000111111",
  6515=>"110111001",
  6516=>"011111111",
  6517=>"001001000",
  6518=>"111000000",
  6519=>"111111101",
  6520=>"000000000",
  6521=>"110110000",
  6522=>"110110111",
  6523=>"000000000",
  6524=>"011011111",
  6525=>"100111111",
  6526=>"100000000",
  6527=>"001000000",
  6528=>"000100110",
  6529=>"111000000",
  6530=>"100011011",
  6531=>"001111111",
  6532=>"000000000",
  6533=>"000000000",
  6534=>"111111111",
  6535=>"000111111",
  6536=>"000000111",
  6537=>"111111111",
  6538=>"001000000",
  6539=>"100111111",
  6540=>"111111111",
  6541=>"100110100",
  6542=>"100100111",
  6543=>"110111011",
  6544=>"111111111",
  6545=>"001000000",
  6546=>"111111111",
  6547=>"000000000",
  6548=>"000000000",
  6549=>"011111000",
  6550=>"011011001",
  6551=>"000000001",
  6552=>"000000000",
  6553=>"011001000",
  6554=>"111101111",
  6555=>"000001001",
  6556=>"101101111",
  6557=>"111111000",
  6558=>"110100000",
  6559=>"111111110",
  6560=>"011011111",
  6561=>"000000001",
  6562=>"100000000",
  6563=>"001011001",
  6564=>"111111111",
  6565=>"111111111",
  6566=>"000000000",
  6567=>"000000000",
  6568=>"000111110",
  6569=>"000000110",
  6570=>"111111001",
  6571=>"100100100",
  6572=>"000010000",
  6573=>"111111111",
  6574=>"011111110",
  6575=>"111111111",
  6576=>"000000000",
  6577=>"111111111",
  6578=>"111111111",
  6579=>"100100000",
  6580=>"000000000",
  6581=>"000100111",
  6582=>"011000000",
  6583=>"000000000",
  6584=>"001000000",
  6585=>"000000000",
  6586=>"100110000",
  6587=>"000100100",
  6588=>"000000000",
  6589=>"000000100",
  6590=>"101100100",
  6591=>"100000011",
  6592=>"100110000",
  6593=>"000000000",
  6594=>"111111011",
  6595=>"000000010",
  6596=>"110001001",
  6597=>"110111001",
  6598=>"111000010",
  6599=>"111110100",
  6600=>"100100100",
  6601=>"111111111",
  6602=>"111001000",
  6603=>"000000000",
  6604=>"011010000",
  6605=>"000000000",
  6606=>"010010000",
  6607=>"000000000",
  6608=>"000101111",
  6609=>"110110010",
  6610=>"011000000",
  6611=>"000000010",
  6612=>"000010000",
  6613=>"011011111",
  6614=>"000000100",
  6615=>"000000000",
  6616=>"001111000",
  6617=>"010001000",
  6618=>"111010000",
  6619=>"111100100",
  6620=>"111101000",
  6621=>"111100000",
  6622=>"111001000",
  6623=>"101001110",
  6624=>"001111110",
  6625=>"000100100",
  6626=>"000000000",
  6627=>"000000000",
  6628=>"100010110",
  6629=>"011111111",
  6630=>"110010010",
  6631=>"001001000",
  6632=>"111111111",
  6633=>"011000000",
  6634=>"000000000",
  6635=>"111001000",
  6636=>"011011010",
  6637=>"000000000",
  6638=>"111110111",
  6639=>"110111111",
  6640=>"011000001",
  6641=>"000011011",
  6642=>"000000000",
  6643=>"111010000",
  6644=>"111100110",
  6645=>"000000001",
  6646=>"100000001",
  6647=>"011110110",
  6648=>"000000000",
  6649=>"000100000",
  6650=>"011001011",
  6651=>"110110111",
  6652=>"000000000",
  6653=>"000000001",
  6654=>"011011011",
  6655=>"001000001",
  6656=>"111100101",
  6657=>"111111011",
  6658=>"000000000",
  6659=>"111111111",
  6660=>"111111111",
  6661=>"111110111",
  6662=>"000000000",
  6663=>"000000000",
  6664=>"111011000",
  6665=>"100000101",
  6666=>"000000000",
  6667=>"000000001",
  6668=>"100100100",
  6669=>"111001001",
  6670=>"110110110",
  6671=>"111111111",
  6672=>"000001000",
  6673=>"011011111",
  6674=>"000000000",
  6675=>"000100111",
  6676=>"000000000",
  6677=>"001001011",
  6678=>"011001000",
  6679=>"011011111",
  6680=>"111111111",
  6681=>"100000100",
  6682=>"000010001",
  6683=>"000001001",
  6684=>"011000000",
  6685=>"101100111",
  6686=>"000000001",
  6687=>"111110111",
  6688=>"000000000",
  6689=>"000000000",
  6690=>"111111100",
  6691=>"010000010",
  6692=>"111101101",
  6693=>"000000001",
  6694=>"111111111",
  6695=>"111111011",
  6696=>"001000000",
  6697=>"000011001",
  6698=>"111100101",
  6699=>"001001101",
  6700=>"111111111",
  6701=>"111110000",
  6702=>"000000000",
  6703=>"100110111",
  6704=>"101111111",
  6705=>"000010000",
  6706=>"000000100",
  6707=>"111111111",
  6708=>"001101111",
  6709=>"111111110",
  6710=>"111111011",
  6711=>"000001000",
  6712=>"000000000",
  6713=>"000001110",
  6714=>"000000100",
  6715=>"000000011",
  6716=>"111111111",
  6717=>"111110111",
  6718=>"111111011",
  6719=>"111111111",
  6720=>"000000000",
  6721=>"001000101",
  6722=>"000110110",
  6723=>"010110111",
  6724=>"111110111",
  6725=>"111111111",
  6726=>"110011000",
  6727=>"111111111",
  6728=>"011011001",
  6729=>"111111111",
  6730=>"111111111",
  6731=>"111111110",
  6732=>"011110000",
  6733=>"111001000",
  6734=>"010011000",
  6735=>"000000000",
  6736=>"000001000",
  6737=>"001000111",
  6738=>"000100000",
  6739=>"001100101",
  6740=>"000000001",
  6741=>"111010011",
  6742=>"001011110",
  6743=>"111111111",
  6744=>"000000000",
  6745=>"111111111",
  6746=>"100100110",
  6747=>"111000000",
  6748=>"010000000",
  6749=>"111111111",
  6750=>"001001101",
  6751=>"111000000",
  6752=>"000000000",
  6753=>"101000000",
  6754=>"011111111",
  6755=>"000000111",
  6756=>"101111111",
  6757=>"111000000",
  6758=>"000000000",
  6759=>"000000000",
  6760=>"100001111",
  6761=>"000000000",
  6762=>"001000000",
  6763=>"000111110",
  6764=>"111001001",
  6765=>"111111111",
  6766=>"111111111",
  6767=>"100100000",
  6768=>"000100111",
  6769=>"000000000",
  6770=>"111111111",
  6771=>"000110111",
  6772=>"011000000",
  6773=>"000000000",
  6774=>"000000000",
  6775=>"101100111",
  6776=>"111001111",
  6777=>"111111100",
  6778=>"000000000",
  6779=>"110000000",
  6780=>"100100100",
  6781=>"111111111",
  6782=>"000000000",
  6783=>"000000001",
  6784=>"000000000",
  6785=>"110111111",
  6786=>"100001001",
  6787=>"011011111",
  6788=>"001011011",
  6789=>"111111111",
  6790=>"111110000",
  6791=>"011010000",
  6792=>"000000000",
  6793=>"111101111",
  6794=>"000000000",
  6795=>"111111111",
  6796=>"111111011",
  6797=>"000000000",
  6798=>"111111110",
  6799=>"110110111",
  6800=>"000000000",
  6801=>"011011001",
  6802=>"000000000",
  6803=>"111111110",
  6804=>"101001001",
  6805=>"010000000",
  6806=>"011001000",
  6807=>"101000100",
  6808=>"101101000",
  6809=>"001011000",
  6810=>"101111111",
  6811=>"001000111",
  6812=>"000000111",
  6813=>"010000001",
  6814=>"000000000",
  6815=>"111111111",
  6816=>"000011011",
  6817=>"011111011",
  6818=>"110000110",
  6819=>"111001000",
  6820=>"111110100",
  6821=>"011000000",
  6822=>"100100000",
  6823=>"011011011",
  6824=>"111011111",
  6825=>"000000000",
  6826=>"111100111",
  6827=>"000000010",
  6828=>"001111100",
  6829=>"100000001",
  6830=>"111111100",
  6831=>"000111011",
  6832=>"111111111",
  6833=>"111011011",
  6834=>"101100100",
  6835=>"000111001",
  6836=>"100111001",
  6837=>"111111000",
  6838=>"000000110",
  6839=>"000100111",
  6840=>"011011101",
  6841=>"000000111",
  6842=>"111111110",
  6843=>"000000110",
  6844=>"111111111",
  6845=>"000000000",
  6846=>"001111111",
  6847=>"111111111",
  6848=>"111100100",
  6849=>"000000000",
  6850=>"111000000",
  6851=>"000000000",
  6852=>"111111111",
  6853=>"101111111",
  6854=>"000100100",
  6855=>"111111111",
  6856=>"000001111",
  6857=>"001010110",
  6858=>"111111011",
  6859=>"000000000",
  6860=>"111111111",
  6861=>"000000000",
  6862=>"000100111",
  6863=>"000001111",
  6864=>"111111011",
  6865=>"111111111",
  6866=>"111011000",
  6867=>"000000000",
  6868=>"111001000",
  6869=>"000111111",
  6870=>"000000110",
  6871=>"000000100",
  6872=>"111111111",
  6873=>"101100000",
  6874=>"111111111",
  6875=>"110000000",
  6876=>"001000000",
  6877=>"111111100",
  6878=>"111111111",
  6879=>"000111000",
  6880=>"100100110",
  6881=>"101011000",
  6882=>"000000000",
  6883=>"000000000",
  6884=>"100100001",
  6885=>"111100000",
  6886=>"111111100",
  6887=>"001111010",
  6888=>"100000000",
  6889=>"000000000",
  6890=>"000100011",
  6891=>"000000000",
  6892=>"111111111",
  6893=>"110100000",
  6894=>"100100111",
  6895=>"000000000",
  6896=>"000000001",
  6897=>"111010100",
  6898=>"111111111",
  6899=>"000000000",
  6900=>"000110111",
  6901=>"111000000",
  6902=>"001000101",
  6903=>"111111111",
  6904=>"000000000",
  6905=>"111111000",
  6906=>"011000001",
  6907=>"000001000",
  6908=>"001011001",
  6909=>"000000110",
  6910=>"000000100",
  6911=>"000000000",
  6912=>"000100100",
  6913=>"110010001",
  6914=>"111100111",
  6915=>"000000000",
  6916=>"111111001",
  6917=>"011011011",
  6918=>"001010000",
  6919=>"011111111",
  6920=>"000000000",
  6921=>"000001111",
  6922=>"001000000",
  6923=>"000000000",
  6924=>"000000000",
  6925=>"111011111",
  6926=>"000000000",
  6927=>"000000000",
  6928=>"011000000",
  6929=>"000000000",
  6930=>"100000000",
  6931=>"111111111",
  6932=>"100111110",
  6933=>"010110111",
  6934=>"000110111",
  6935=>"111111110",
  6936=>"101111111",
  6937=>"111111111",
  6938=>"111011111",
  6939=>"000100110",
  6940=>"110110111",
  6941=>"001000111",
  6942=>"111111011",
  6943=>"000000000",
  6944=>"100100100",
  6945=>"000011010",
  6946=>"100100100",
  6947=>"111111111",
  6948=>"000000000",
  6949=>"100111111",
  6950=>"000100100",
  6951=>"011111111",
  6952=>"000000011",
  6953=>"011111000",
  6954=>"001000000",
  6955=>"000000000",
  6956=>"111111111",
  6957=>"111111011",
  6958=>"111111111",
  6959=>"111111111",
  6960=>"000000010",
  6961=>"111111111",
  6962=>"000111111",
  6963=>"000111111",
  6964=>"111111111",
  6965=>"111011001",
  6966=>"111011011",
  6967=>"111001001",
  6968=>"000000000",
  6969=>"000000000",
  6970=>"100110111",
  6971=>"000000000",
  6972=>"111111111",
  6973=>"001001001",
  6974=>"000111111",
  6975=>"111111111",
  6976=>"111111111",
  6977=>"111111111",
  6978=>"111111111",
  6979=>"111111111",
  6980=>"111111111",
  6981=>"110000000",
  6982=>"010011000",
  6983=>"000000000",
  6984=>"000000000",
  6985=>"111111000",
  6986=>"111111111",
  6987=>"111110110",
  6988=>"000000000",
  6989=>"000000001",
  6990=>"000000000",
  6991=>"111111100",
  6992=>"111110100",
  6993=>"000000000",
  6994=>"111111111",
  6995=>"011111110",
  6996=>"000011111",
  6997=>"011000011",
  6998=>"001001000",
  6999=>"111000001",
  7000=>"111111111",
  7001=>"111111111",
  7002=>"111111111",
  7003=>"000010111",
  7004=>"111111111",
  7005=>"000000000",
  7006=>"001111111",
  7007=>"111111111",
  7008=>"111110111",
  7009=>"011001001",
  7010=>"000000000",
  7011=>"000000000",
  7012=>"100101101",
  7013=>"000000000",
  7014=>"000000000",
  7015=>"110011011",
  7016=>"110010001",
  7017=>"111110111",
  7018=>"111111111",
  7019=>"111111101",
  7020=>"100100110",
  7021=>"111111111",
  7022=>"000000000",
  7023=>"011000000",
  7024=>"000000000",
  7025=>"100000000",
  7026=>"111011111",
  7027=>"111111111",
  7028=>"000100100",
  7029=>"111111001",
  7030=>"001111111",
  7031=>"110111111",
  7032=>"101000000",
  7033=>"000000000",
  7034=>"000000010",
  7035=>"010000000",
  7036=>"101001000",
  7037=>"010110110",
  7038=>"111000101",
  7039=>"111111111",
  7040=>"101000001",
  7041=>"100001000",
  7042=>"111111111",
  7043=>"011100000",
  7044=>"110111111",
  7045=>"111101000",
  7046=>"000000000",
  7047=>"101111110",
  7048=>"000001101",
  7049=>"111111111",
  7050=>"100100110",
  7051=>"000000000",
  7052=>"111111111",
  7053=>"111011111",
  7054=>"101000101",
  7055=>"111101111",
  7056=>"000000000",
  7057=>"111111101",
  7058=>"111111111",
  7059=>"111111111",
  7060=>"010001011",
  7061=>"000000000",
  7062=>"000000000",
  7063=>"000000000",
  7064=>"000001000",
  7065=>"000100100",
  7066=>"000100000",
  7067=>"000000001",
  7068=>"111111111",
  7069=>"111111000",
  7070=>"000100100",
  7071=>"110110000",
  7072=>"110000100",
  7073=>"001000000",
  7074=>"101000000",
  7075=>"010011111",
  7076=>"111110010",
  7077=>"000000000",
  7078=>"001000000",
  7079=>"000000000",
  7080=>"110111111",
  7081=>"110000000",
  7082=>"000000000",
  7083=>"011011011",
  7084=>"000010000",
  7085=>"111001001",
  7086=>"010111111",
  7087=>"111000000",
  7088=>"111001111",
  7089=>"111111110",
  7090=>"110111111",
  7091=>"111111111",
  7092=>"111001000",
  7093=>"110110000",
  7094=>"000000000",
  7095=>"000000001",
  7096=>"000111111",
  7097=>"000000000",
  7098=>"000001000",
  7099=>"000000011",
  7100=>"110110100",
  7101=>"000000000",
  7102=>"111111111",
  7103=>"110110000",
  7104=>"110110110",
  7105=>"101000000",
  7106=>"000000000",
  7107=>"111111111",
  7108=>"111110110",
  7109=>"000000111",
  7110=>"111111111",
  7111=>"100101111",
  7112=>"111110110",
  7113=>"000000000",
  7114=>"111111111",
  7115=>"111111101",
  7116=>"000001111",
  7117=>"111001000",
  7118=>"111111111",
  7119=>"000000110",
  7120=>"000000001",
  7121=>"111111100",
  7122=>"001111000",
  7123=>"111111000",
  7124=>"111111101",
  7125=>"011011111",
  7126=>"000000000",
  7127=>"000110110",
  7128=>"000000011",
  7129=>"000000000",
  7130=>"000001000",
  7131=>"110110010",
  7132=>"000011011",
  7133=>"001000000",
  7134=>"111011111",
  7135=>"011011111",
  7136=>"000000000",
  7137=>"001000000",
  7138=>"001011000",
  7139=>"000000000",
  7140=>"110000111",
  7141=>"101101000",
  7142=>"111011111",
  7143=>"111111111",
  7144=>"111111111",
  7145=>"111111111",
  7146=>"000010010",
  7147=>"001111111",
  7148=>"111111000",
  7149=>"011000000",
  7150=>"000000000",
  7151=>"001000000",
  7152=>"010000000",
  7153=>"111111111",
  7154=>"111111111",
  7155=>"000000101",
  7156=>"001100111",
  7157=>"110100110",
  7158=>"111111111",
  7159=>"110011001",
  7160=>"001111111",
  7161=>"111111111",
  7162=>"000010110",
  7163=>"111111000",
  7164=>"111111111",
  7165=>"111111101",
  7166=>"111000001",
  7167=>"111111000",
  7168=>"000000000",
  7169=>"110111111",
  7170=>"111111111",
  7171=>"000000001",
  7172=>"100100110",
  7173=>"000000000",
  7174=>"110111111",
  7175=>"000000000",
  7176=>"000000000",
  7177=>"001111111",
  7178=>"100000000",
  7179=>"111111111",
  7180=>"001001111",
  7181=>"000000001",
  7182=>"111111111",
  7183=>"000000000",
  7184=>"000001001",
  7185=>"100101111",
  7186=>"000000000",
  7187=>"111111111",
  7188=>"111111011",
  7189=>"001101111",
  7190=>"000000001",
  7191=>"100100100",
  7192=>"111111111",
  7193=>"111111111",
  7194=>"000101111",
  7195=>"100101100",
  7196=>"000110100",
  7197=>"001101111",
  7198=>"000100111",
  7199=>"000011001",
  7200=>"111100000",
  7201=>"000000000",
  7202=>"110110100",
  7203=>"000000001",
  7204=>"001111111",
  7205=>"000000000",
  7206=>"111101111",
  7207=>"011001011",
  7208=>"111111111",
  7209=>"000110010",
  7210=>"111110100",
  7211=>"100100100",
  7212=>"000000000",
  7213=>"100011000",
  7214=>"010010011",
  7215=>"111111111",
  7216=>"101110111",
  7217=>"111111111",
  7218=>"100000000",
  7219=>"000000000",
  7220=>"000000000",
  7221=>"111110000",
  7222=>"111001011",
  7223=>"101100000",
  7224=>"000011001",
  7225=>"110110000",
  7226=>"000000001",
  7227=>"111111110",
  7228=>"000111111",
  7229=>"110000000",
  7230=>"000001001",
  7231=>"000000000",
  7232=>"000111111",
  7233=>"101001001",
  7234=>"011010000",
  7235=>"110111111",
  7236=>"000000000",
  7237=>"111111111",
  7238=>"000000100",
  7239=>"111111011",
  7240=>"011001110",
  7241=>"000100111",
  7242=>"000000000",
  7243=>"010010010",
  7244=>"000000001",
  7245=>"010010011",
  7246=>"111111000",
  7247=>"110110000",
  7248=>"111111111",
  7249=>"000011010",
  7250=>"000111111",
  7251=>"010000000",
  7252=>"111011000",
  7253=>"111001000",
  7254=>"000010110",
  7255=>"110110100",
  7256=>"111111111",
  7257=>"000000011",
  7258=>"000000011",
  7259=>"111111111",
  7260=>"000000000",
  7261=>"000011011",
  7262=>"011111111",
  7263=>"111111111",
  7264=>"111111111",
  7265=>"000000000",
  7266=>"001001101",
  7267=>"101111110",
  7268=>"011111000",
  7269=>"000111111",
  7270=>"111111111",
  7271=>"010111000",
  7272=>"111111111",
  7273=>"111000100",
  7274=>"111111011",
  7275=>"111000000",
  7276=>"110100111",
  7277=>"111111111",
  7278=>"011111111",
  7279=>"000000101",
  7280=>"111000000",
  7281=>"011000000",
  7282=>"100100100",
  7283=>"000000100",
  7284=>"100000000",
  7285=>"111100110",
  7286=>"010011000",
  7287=>"000000000",
  7288=>"111000001",
  7289=>"111101100",
  7290=>"000000000",
  7291=>"011010000",
  7292=>"010110110",
  7293=>"000000000",
  7294=>"000000000",
  7295=>"111111111",
  7296=>"000111111",
  7297=>"000000110",
  7298=>"000000000",
  7299=>"110100000",
  7300=>"000000000",
  7301=>"111111111",
  7302=>"000111111",
  7303=>"011110100",
  7304=>"111111111",
  7305=>"000000000",
  7306=>"110110100",
  7307=>"000111110",
  7308=>"011111111",
  7309=>"011000000",
  7310=>"111111111",
  7311=>"111111111",
  7312=>"000000110",
  7313=>"100100100",
  7314=>"011011000",
  7315=>"000000000",
  7316=>"000000000",
  7317=>"000100000",
  7318=>"000000000",
  7319=>"111111111",
  7320=>"000000000",
  7321=>"111111111",
  7322=>"000000110",
  7323=>"000000000",
  7324=>"111000000",
  7325=>"110111000",
  7326=>"101000011",
  7327=>"110110000",
  7328=>"111001000",
  7329=>"000010000",
  7330=>"110111111",
  7331=>"110111001",
  7332=>"000000000",
  7333=>"011000000",
  7334=>"000000101",
  7335=>"010110000",
  7336=>"011011011",
  7337=>"111111111",
  7338=>"100100100",
  7339=>"010011111",
  7340=>"000000000",
  7341=>"111111111",
  7342=>"000000001",
  7343=>"010001000",
  7344=>"000100111",
  7345=>"111111111",
  7346=>"110110110",
  7347=>"010110111",
  7348=>"110011111",
  7349=>"111110000",
  7350=>"001001001",
  7351=>"000000101",
  7352=>"110111111",
  7353=>"111110111",
  7354=>"000000000",
  7355=>"000000000",
  7356=>"000000000",
  7357=>"100111111",
  7358=>"001001000",
  7359=>"111111111",
  7360=>"111110100",
  7361=>"111111001",
  7362=>"000000001",
  7363=>"111000001",
  7364=>"110111111",
  7365=>"111011011",
  7366=>"111000000",
  7367=>"111111111",
  7368=>"001001011",
  7369=>"111111111",
  7370=>"001000000",
  7371=>"011101111",
  7372=>"011000110",
  7373=>"110110000",
  7374=>"111111111",
  7375=>"000000000",
  7376=>"011111111",
  7377=>"000000001",
  7378=>"000000111",
  7379=>"111110111",
  7380=>"011000000",
  7381=>"111111111",
  7382=>"000000000",
  7383=>"111111111",
  7384=>"000000001",
  7385=>"000100100",
  7386=>"011111111",
  7387=>"010000000",
  7388=>"000000001",
  7389=>"111111111",
  7390=>"111111111",
  7391=>"111100000",
  7392=>"000000111",
  7393=>"000000000",
  7394=>"011111111",
  7395=>"011011011",
  7396=>"111111011",
  7397=>"111111111",
  7398=>"110011001",
  7399=>"001101100",
  7400=>"000000111",
  7401=>"000000000",
  7402=>"111111001",
  7403=>"000000000",
  7404=>"000000000",
  7405=>"000000000",
  7406=>"111111100",
  7407=>"000000000",
  7408=>"100000001",
  7409=>"111111111",
  7410=>"101001111",
  7411=>"001001001",
  7412=>"110111111",
  7413=>"000111111",
  7414=>"111110110",
  7415=>"000000110",
  7416=>"000000111",
  7417=>"111111111",
  7418=>"011011011",
  7419=>"111111100",
  7420=>"001011111",
  7421=>"001000001",
  7422=>"000000000",
  7423=>"111011011",
  7424=>"111111111",
  7425=>"001011011",
  7426=>"000000000",
  7427=>"111111111",
  7428=>"000101111",
  7429=>"111111111",
  7430=>"111111111",
  7431=>"010110000",
  7432=>"000000000",
  7433=>"111111111",
  7434=>"100110111",
  7435=>"111111111",
  7436=>"100111111",
  7437=>"110111111",
  7438=>"111011111",
  7439=>"111111111",
  7440=>"111111000",
  7441=>"000000000",
  7442=>"111111111",
  7443=>"110110111",
  7444=>"111111111",
  7445=>"000000000",
  7446=>"100100000",
  7447=>"111111111",
  7448=>"110010110",
  7449=>"000010010",
  7450=>"000110000",
  7451=>"110110110",
  7452=>"100101011",
  7453=>"000000000",
  7454=>"111111000",
  7455=>"010111111",
  7456=>"001000000",
  7457=>"111111111",
  7458=>"000000000",
  7459=>"111111111",
  7460=>"000000000",
  7461=>"000000101",
  7462=>"000000000",
  7463=>"111001000",
  7464=>"100100111",
  7465=>"111111001",
  7466=>"111111000",
  7467=>"000000000",
  7468=>"111111111",
  7469=>"010000001",
  7470=>"110000111",
  7471=>"111111111",
  7472=>"011001000",
  7473=>"000000000",
  7474=>"110100100",
  7475=>"000000000",
  7476=>"000000011",
  7477=>"000000000",
  7478=>"000100100",
  7479=>"000000001",
  7480=>"001000000",
  7481=>"111111010",
  7482=>"000010000",
  7483=>"001011000",
  7484=>"000010000",
  7485=>"001100111",
  7486=>"100100110",
  7487=>"000000000",
  7488=>"111111110",
  7489=>"011111110",
  7490=>"111111001",
  7491=>"000000110",
  7492=>"000000111",
  7493=>"000110000",
  7494=>"111111111",
  7495=>"000000110",
  7496=>"000000000",
  7497=>"000011111",
  7498=>"111000001",
  7499=>"010110100",
  7500=>"111000000",
  7501=>"000000000",
  7502=>"011000001",
  7503=>"000000000",
  7504=>"111011000",
  7505=>"110000000",
  7506=>"000000000",
  7507=>"000000000",
  7508=>"011010111",
  7509=>"110110000",
  7510=>"000100000",
  7511=>"100100110",
  7512=>"111111111",
  7513=>"011000111",
  7514=>"111111111",
  7515=>"001000111",
  7516=>"001001000",
  7517=>"000000000",
  7518=>"111111111",
  7519=>"100000000",
  7520=>"111111111",
  7521=>"000000000",
  7522=>"001000111",
  7523=>"000000000",
  7524=>"000110000",
  7525=>"000000111",
  7526=>"000111111",
  7527=>"110111111",
  7528=>"001101111",
  7529=>"000000000",
  7530=>"000000000",
  7531=>"000000000",
  7532=>"111111111",
  7533=>"000000111",
  7534=>"111111100",
  7535=>"000110110",
  7536=>"111111111",
  7537=>"110110100",
  7538=>"011000101",
  7539=>"011000000",
  7540=>"110111011",
  7541=>"111001000",
  7542=>"000011011",
  7543=>"110111010",
  7544=>"111111111",
  7545=>"000000001",
  7546=>"100100100",
  7547=>"111111111",
  7548=>"000000001",
  7549=>"111111111",
  7550=>"000000001",
  7551=>"110111111",
  7552=>"111111111",
  7553=>"001000000",
  7554=>"000001000",
  7555=>"111000000",
  7556=>"011000000",
  7557=>"001001011",
  7558=>"000000000",
  7559=>"110110111",
  7560=>"000000001",
  7561=>"000000000",
  7562=>"111111111",
  7563=>"111111111",
  7564=>"010110111",
  7565=>"001001000",
  7566=>"001011111",
  7567=>"111111111",
  7568=>"000000000",
  7569=>"000000111",
  7570=>"011011000",
  7571=>"000000000",
  7572=>"000011111",
  7573=>"111111011",
  7574=>"000000000",
  7575=>"011000100",
  7576=>"111111111",
  7577=>"100100000",
  7578=>"000111111",
  7579=>"111111111",
  7580=>"000000001",
  7581=>"010000100",
  7582=>"000000000",
  7583=>"111111111",
  7584=>"001001001",
  7585=>"100110110",
  7586=>"011011101",
  7587=>"011000000",
  7588=>"111111100",
  7589=>"110111111",
  7590=>"100000101",
  7591=>"000000000",
  7592=>"000000000",
  7593=>"110110100",
  7594=>"000000011",
  7595=>"111010000",
  7596=>"111111111",
  7597=>"000000111",
  7598=>"111110111",
  7599=>"111111111",
  7600=>"000000000",
  7601=>"000010110",
  7602=>"110000001",
  7603=>"111111110",
  7604=>"000000000",
  7605=>"000000111",
  7606=>"000000000",
  7607=>"111111001",
  7608=>"010000000",
  7609=>"000000000",
  7610=>"000000000",
  7611=>"000000111",
  7612=>"111111111",
  7613=>"111011111",
  7614=>"111111110",
  7615=>"001011011",
  7616=>"000000000",
  7617=>"010010000",
  7618=>"110011111",
  7619=>"111111111",
  7620=>"111110111",
  7621=>"111111111",
  7622=>"011000000",
  7623=>"000000000",
  7624=>"000000000",
  7625=>"100110000",
  7626=>"011011001",
  7627=>"000000000",
  7628=>"011011111",
  7629=>"010110111",
  7630=>"000000100",
  7631=>"111111111",
  7632=>"000000000",
  7633=>"111111011",
  7634=>"000000000",
  7635=>"000000000",
  7636=>"001001001",
  7637=>"000000000",
  7638=>"111111000",
  7639=>"111000000",
  7640=>"010100101",
  7641=>"110010000",
  7642=>"000000000",
  7643=>"001001101",
  7644=>"100000100",
  7645=>"111011011",
  7646=>"111111111",
  7647=>"100000000",
  7648=>"000000000",
  7649=>"111111111",
  7650=>"000000000",
  7651=>"111100000",
  7652=>"110100000",
  7653=>"011011000",
  7654=>"000000000",
  7655=>"011111001",
  7656=>"010000000",
  7657=>"000101111",
  7658=>"000000000",
  7659=>"000000100",
  7660=>"110100000",
  7661=>"111111011",
  7662=>"001001111",
  7663=>"111111111",
  7664=>"000000000",
  7665=>"000000000",
  7666=>"000000100",
  7667=>"000000000",
  7668=>"111100000",
  7669=>"111001001",
  7670=>"111111111",
  7671=>"111111001",
  7672=>"001011011",
  7673=>"010100000",
  7674=>"111111111",
  7675=>"011011000",
  7676=>"000000000",
  7677=>"000100000",
  7678=>"101111001",
  7679=>"111110110",
  7680=>"011111111",
  7681=>"000001111",
  7682=>"000000000",
  7683=>"110100111",
  7684=>"000000001",
  7685=>"110111110",
  7686=>"000000000",
  7687=>"111111111",
  7688=>"000000111",
  7689=>"000000111",
  7690=>"111110111",
  7691=>"000000110",
  7692=>"000100110",
  7693=>"111111000",
  7694=>"100110111",
  7695=>"000000000",
  7696=>"110100111",
  7697=>"000000010",
  7698=>"100111000",
  7699=>"000000111",
  7700=>"110000000",
  7701=>"111000000",
  7702=>"000000110",
  7703=>"001001101",
  7704=>"000000111",
  7705=>"001000000",
  7706=>"011010010",
  7707=>"000011111",
  7708=>"010011000",
  7709=>"000000000",
  7710=>"111111000",
  7711=>"000110111",
  7712=>"000000011",
  7713=>"110000000",
  7714=>"000000110",
  7715=>"110100111",
  7716=>"110111111",
  7717=>"000011000",
  7718=>"110110111",
  7719=>"111111111",
  7720=>"000000000",
  7721=>"001000111",
  7722=>"011111011",
  7723=>"000110111",
  7724=>"000000111",
  7725=>"111111000",
  7726=>"101111111",
  7727=>"001111111",
  7728=>"011111111",
  7729=>"000000011",
  7730=>"000001000",
  7731=>"100100000",
  7732=>"000111111",
  7733=>"000001000",
  7734=>"000000001",
  7735=>"000000000",
  7736=>"111111000",
  7737=>"011000111",
  7738=>"000001111",
  7739=>"111111011",
  7740=>"000000010",
  7741=>"101100110",
  7742=>"000110111",
  7743=>"101000110",
  7744=>"011111000",
  7745=>"000111000",
  7746=>"111111111",
  7747=>"111111110",
  7748=>"111000111",
  7749=>"001000110",
  7750=>"111000000",
  7751=>"111000011",
  7752=>"011011011",
  7753=>"000000001",
  7754=>"111111010",
  7755=>"000010000",
  7756=>"000000000",
  7757=>"000000001",
  7758=>"000010011",
  7759=>"111111000",
  7760=>"111000000",
  7761=>"110111010",
  7762=>"000000100",
  7763=>"011111000",
  7764=>"000000000",
  7765=>"111111010",
  7766=>"000000011",
  7767=>"111111101",
  7768=>"000000000",
  7769=>"111000000",
  7770=>"111111110",
  7771=>"010001011",
  7772=>"111111010",
  7773=>"111111111",
  7774=>"001001111",
  7775=>"111111000",
  7776=>"000111111",
  7777=>"111010010",
  7778=>"111111111",
  7779=>"000001111",
  7780=>"011001000",
  7781=>"011111111",
  7782=>"111111000",
  7783=>"010011000",
  7784=>"111001000",
  7785=>"111111111",
  7786=>"001000000",
  7787=>"011111111",
  7788=>"001111111",
  7789=>"111100001",
  7790=>"100000111",
  7791=>"000111111",
  7792=>"111011000",
  7793=>"111001001",
  7794=>"100110110",
  7795=>"111111111",
  7796=>"001000000",
  7797=>"000000000",
  7798=>"111001000",
  7799=>"000000000",
  7800=>"000000111",
  7801=>"011000000",
  7802=>"000101101",
  7803=>"011000000",
  7804=>"000111111",
  7805=>"111110000",
  7806=>"111111111",
  7807=>"000000111",
  7808=>"000000000",
  7809=>"000000111",
  7810=>"010000110",
  7811=>"110110111",
  7812=>"000010111",
  7813=>"001000000",
  7814=>"111111000",
  7815=>"000000111",
  7816=>"111111111",
  7817=>"001001100",
  7818=>"000111111",
  7819=>"111111111",
  7820=>"000000000",
  7821=>"111011000",
  7822=>"000000000",
  7823=>"000000000",
  7824=>"000000011",
  7825=>"101110111",
  7826=>"111111011",
  7827=>"000000000",
  7828=>"111111111",
  7829=>"000111111",
  7830=>"111000000",
  7831=>"111000000",
  7832=>"000000000",
  7833=>"111111111",
  7834=>"111101001",
  7835=>"000000000",
  7836=>"011000000",
  7837=>"000000000",
  7838=>"010011001",
  7839=>"111000000",
  7840=>"000000111",
  7841=>"111100011",
  7842=>"000000000",
  7843=>"111111000",
  7844=>"000011111",
  7845=>"111010000",
  7846=>"111111110",
  7847=>"001111000",
  7848=>"011111111",
  7849=>"000001111",
  7850=>"111001111",
  7851=>"111111111",
  7852=>"111000000",
  7853=>"100111100",
  7854=>"000000111",
  7855=>"100110111",
  7856=>"000111001",
  7857=>"000000001",
  7858=>"000111000",
  7859=>"000000111",
  7860=>"011000000",
  7861=>"000000111",
  7862=>"111111111",
  7863=>"111111111",
  7864=>"011000000",
  7865=>"100000000",
  7866=>"101000001",
  7867=>"001000000",
  7868=>"111000000",
  7869=>"001000000",
  7870=>"000000100",
  7871=>"000101111",
  7872=>"000000000",
  7873=>"110010010",
  7874=>"100100100",
  7875=>"111111111",
  7876=>"000000011",
  7877=>"000101111",
  7878=>"001011000",
  7879=>"011111111",
  7880=>"000111111",
  7881=>"000010111",
  7882=>"000000111",
  7883=>"000100111",
  7884=>"111111011",
  7885=>"000000110",
  7886=>"000000001",
  7887=>"000001000",
  7888=>"000000111",
  7889=>"000000111",
  7890=>"000011011",
  7891=>"000000000",
  7892=>"100000000",
  7893=>"000000111",
  7894=>"110000101",
  7895=>"010011111",
  7896=>"111111000",
  7897=>"110001111",
  7898=>"000000000",
  7899=>"000000000",
  7900=>"111111000",
  7901=>"001000000",
  7902=>"011000000",
  7903=>"011011010",
  7904=>"110000000",
  7905=>"000000011",
  7906=>"111111111",
  7907=>"001000000",
  7908=>"000000000",
  7909=>"011110100",
  7910=>"111111000",
  7911=>"000000000",
  7912=>"000000111",
  7913=>"000000000",
  7914=>"111111111",
  7915=>"001111111",
  7916=>"000111111",
  7917=>"001000111",
  7918=>"000110011",
  7919=>"101001000",
  7920=>"110100110",
  7921=>"000000000",
  7922=>"001001001",
  7923=>"111111011",
  7924=>"111111100",
  7925=>"011111111",
  7926=>"011111101",
  7927=>"111011001",
  7928=>"000000000",
  7929=>"000001001",
  7930=>"111111011",
  7931=>"000000000",
  7932=>"000101000",
  7933=>"110110111",
  7934=>"111000000",
  7935=>"000000000",
  7936=>"000001111",
  7937=>"000000011",
  7938=>"111111011",
  7939=>"011011001",
  7940=>"110000000",
  7941=>"000001010",
  7942=>"001000000",
  7943=>"000111010",
  7944=>"000111110",
  7945=>"000011000",
  7946=>"101000000",
  7947=>"000000000",
  7948=>"011111101",
  7949=>"110100010",
  7950=>"010000000",
  7951=>"111111001",
  7952=>"001111101",
  7953=>"100110010",
  7954=>"111001000",
  7955=>"000000010",
  7956=>"111110000",
  7957=>"111110000",
  7958=>"000100100",
  7959=>"111101000",
  7960=>"111111110",
  7961=>"111001101",
  7962=>"000000111",
  7963=>"010111110",
  7964=>"000000111",
  7965=>"000001100",
  7966=>"110000000",
  7967=>"111111111",
  7968=>"111000000",
  7969=>"000111111",
  7970=>"110000000",
  7971=>"011010011",
  7972=>"000000111",
  7973=>"111111000",
  7974=>"111111111",
  7975=>"111000000",
  7976=>"000000000",
  7977=>"000000000",
  7978=>"111000000",
  7979=>"111111011",
  7980=>"111111111",
  7981=>"100000000",
  7982=>"000000111",
  7983=>"000000100",
  7984=>"011111111",
  7985=>"111111111",
  7986=>"000111000",
  7987=>"111000111",
  7988=>"110100000",
  7989=>"000110011",
  7990=>"111111000",
  7991=>"000000111",
  7992=>"110100000",
  7993=>"111000000",
  7994=>"000000111",
  7995=>"111001000",
  7996=>"111111111",
  7997=>"111110000",
  7998=>"000011111",
  7999=>"000000000",
  8000=>"011001000",
  8001=>"101100100",
  8002=>"001000111",
  8003=>"111000001",
  8004=>"001001000",
  8005=>"111000111",
  8006=>"000000000",
  8007=>"010000000",
  8008=>"111111000",
  8009=>"010010111",
  8010=>"110000111",
  8011=>"011000000",
  8012=>"111010000",
  8013=>"001000000",
  8014=>"111111110",
  8015=>"000001011",
  8016=>"000000001",
  8017=>"111011000",
  8018=>"000111110",
  8019=>"000000001",
  8020=>"010101110",
  8021=>"011111111",
  8022=>"011110100",
  8023=>"111111011",
  8024=>"111111111",
  8025=>"111011111",
  8026=>"111111111",
  8027=>"100000000",
  8028=>"111000111",
  8029=>"111000111",
  8030=>"111110100",
  8031=>"110111111",
  8032=>"000000000",
  8033=>"000100110",
  8034=>"111101001",
  8035=>"110100101",
  8036=>"000001000",
  8037=>"000000100",
  8038=>"000000100",
  8039=>"000111110",
  8040=>"011000000",
  8041=>"000000111",
  8042=>"000000111",
  8043=>"000111001",
  8044=>"000111001",
  8045=>"000000000",
  8046=>"010010000",
  8047=>"111111111",
  8048=>"000011110",
  8049=>"000110010",
  8050=>"011001111",
  8051=>"000000011",
  8052=>"010110000",
  8053=>"111110100",
  8054=>"010010011",
  8055=>"011111111",
  8056=>"000000000",
  8057=>"000111011",
  8058=>"000000000",
  8059=>"000000000",
  8060=>"000000000",
  8061=>"101111111",
  8062=>"000101111",
  8063=>"111000000",
  8064=>"001001000",
  8065=>"111111111",
  8066=>"110111111",
  8067=>"000000111",
  8068=>"000000011",
  8069=>"000100101",
  8070=>"000010110",
  8071=>"110110111",
  8072=>"011000010",
  8073=>"100111101",
  8074=>"111111011",
  8075=>"111011111",
  8076=>"111111011",
  8077=>"011111000",
  8078=>"111111111",
  8079=>"111111110",
  8080=>"000111111",
  8081=>"111111111",
  8082=>"111010000",
  8083=>"010000000",
  8084=>"000000010",
  8085=>"000000000",
  8086=>"000000000",
  8087=>"001111001",
  8088=>"111110000",
  8089=>"010000000",
  8090=>"000000111",
  8091=>"000000110",
  8092=>"101111111",
  8093=>"000011000",
  8094=>"000100100",
  8095=>"000001011",
  8096=>"000111111",
  8097=>"000000011",
  8098=>"101000000",
  8099=>"111111111",
  8100=>"001000110",
  8101=>"110111000",
  8102=>"010010000",
  8103=>"011010111",
  8104=>"100101111",
  8105=>"111111000",
  8106=>"000000101",
  8107=>"101100100",
  8108=>"000111100",
  8109=>"001111111",
  8110=>"010111111",
  8111=>"000000000",
  8112=>"111111111",
  8113=>"000000001",
  8114=>"001111100",
  8115=>"000000000",
  8116=>"000010010",
  8117=>"111100000",
  8118=>"111100000",
  8119=>"111001001",
  8120=>"111111111",
  8121=>"111000000",
  8122=>"000111111",
  8123=>"111000000",
  8124=>"111000110",
  8125=>"001000000",
  8126=>"100000000",
  8127=>"000100000",
  8128=>"111111111",
  8129=>"001001001",
  8130=>"000000000",
  8131=>"111000001",
  8132=>"111111111",
  8133=>"010111110",
  8134=>"111111010",
  8135=>"111000000",
  8136=>"000000100",
  8137=>"111111000",
  8138=>"000101011",
  8139=>"111010111",
  8140=>"111000000",
  8141=>"111111000",
  8142=>"000111111",
  8143=>"111000000",
  8144=>"001011111",
  8145=>"100000000",
  8146=>"011010000",
  8147=>"101111111",
  8148=>"110100001",
  8149=>"000000011",
  8150=>"111111101",
  8151=>"100100011",
  8152=>"000000011",
  8153=>"000001011",
  8154=>"000001111",
  8155=>"000000111",
  8156=>"000101110",
  8157=>"101111000",
  8158=>"111000001",
  8159=>"000100000",
  8160=>"000000000",
  8161=>"000100100",
  8162=>"111111000",
  8163=>"000111100",
  8164=>"011111111",
  8165=>"011000000",
  8166=>"111101110",
  8167=>"111111111",
  8168=>"000000000",
  8169=>"001000001",
  8170=>"000011011",
  8171=>"000111110",
  8172=>"000111111",
  8173=>"100111110",
  8174=>"100000000",
  8175=>"111000000",
  8176=>"000111000",
  8177=>"111111111",
  8178=>"000000000",
  8179=>"101101101",
  8180=>"000000110",
  8181=>"000111111",
  8182=>"000000110",
  8183=>"000000111",
  8184=>"000100111",
  8185=>"000001000",
  8186=>"010000111",
  8187=>"111000000",
  8188=>"000111111",
  8189=>"000111111",
  8190=>"000011000",
  8191=>"000000000",
  8192=>"111011001",
  8193=>"000000000",
  8194=>"111111111",
  8195=>"100000000",
  8196=>"111111111",
  8197=>"011011001",
  8198=>"001000000",
  8199=>"100000001",
  8200=>"000011111",
  8201=>"111111101",
  8202=>"000000000",
  8203=>"000000001",
  8204=>"110100110",
  8205=>"100100001",
  8206=>"000000000",
  8207=>"000101111",
  8208=>"011001011",
  8209=>"000000000",
  8210=>"001000100",
  8211=>"000110110",
  8212=>"001111111",
  8213=>"111111111",
  8214=>"000000000",
  8215=>"110110111",
  8216=>"111110100",
  8217=>"011110100",
  8218=>"111111111",
  8219=>"001001001",
  8220=>"000000000",
  8221=>"000000000",
  8222=>"111111101",
  8223=>"000000000",
  8224=>"000010000",
  8225=>"011000000",
  8226=>"011010000",
  8227=>"111111000",
  8228=>"111100111",
  8229=>"000000001",
  8230=>"111110000",
  8231=>"111110111",
  8232=>"010000000",
  8233=>"100000000",
  8234=>"111111111",
  8235=>"000000000",
  8236=>"110111011",
  8237=>"111111001",
  8238=>"111011011",
  8239=>"000000000",
  8240=>"111111100",
  8241=>"000000000",
  8242=>"000000000",
  8243=>"000000000",
  8244=>"111011000",
  8245=>"111001001",
  8246=>"001011001",
  8247=>"010000100",
  8248=>"111100000",
  8249=>"010000111",
  8250=>"000000011",
  8251=>"000011011",
  8252=>"111111111",
  8253=>"100111111",
  8254=>"111001000",
  8255=>"000000111",
  8256=>"011011011",
  8257=>"101101111",
  8258=>"000111111",
  8259=>"111110000",
  8260=>"001001001",
  8261=>"000000000",
  8262=>"000000000",
  8263=>"111111111",
  8264=>"111100101",
  8265=>"000000000",
  8266=>"100100110",
  8267=>"011111101",
  8268=>"000000100",
  8269=>"111001100",
  8270=>"111011111",
  8271=>"111111000",
  8272=>"000000111",
  8273=>"101111110",
  8274=>"111111110",
  8275=>"000000110",
  8276=>"001111011",
  8277=>"000010110",
  8278=>"000100111",
  8279=>"110111110",
  8280=>"111011111",
  8281=>"111101001",
  8282=>"000111110",
  8283=>"100100100",
  8284=>"011000100",
  8285=>"111110110",
  8286=>"011010110",
  8287=>"000001111",
  8288=>"111111111",
  8289=>"110111111",
  8290=>"000000000",
  8291=>"111100000",
  8292=>"111000000",
  8293=>"011111111",
  8294=>"011000111",
  8295=>"000000000",
  8296=>"000010111",
  8297=>"011111111",
  8298=>"000000000",
  8299=>"000000000",
  8300=>"011000110",
  8301=>"111011000",
  8302=>"000000110",
  8303=>"110000000",
  8304=>"011111111",
  8305=>"000111111",
  8306=>"000000000",
  8307=>"111000001",
  8308=>"000000000",
  8309=>"111111011",
  8310=>"001000000",
  8311=>"000011111",
  8312=>"000011011",
  8313=>"111000000",
  8314=>"111111111",
  8315=>"000111000",
  8316=>"111000000",
  8317=>"000000111",
  8318=>"011001010",
  8319=>"000000000",
  8320=>"000000000",
  8321=>"111111111",
  8322=>"000000110",
  8323=>"000011111",
  8324=>"000001011",
  8325=>"000000000",
  8326=>"000111111",
  8327=>"111110111",
  8328=>"110010111",
  8329=>"100111111",
  8330=>"000000000",
  8331=>"000000000",
  8332=>"000000000",
  8333=>"101111100",
  8334=>"100110111",
  8335=>"111111000",
  8336=>"000000000",
  8337=>"000000000",
  8338=>"001111111",
  8339=>"111001000",
  8340=>"000010000",
  8341=>"111111101",
  8342=>"000000000",
  8343=>"111110000",
  8344=>"000011110",
  8345=>"111111111",
  8346=>"000000000",
  8347=>"111111011",
  8348=>"000000100",
  8349=>"011001011",
  8350=>"000000000",
  8351=>"100101101",
  8352=>"011111000",
  8353=>"111011000",
  8354=>"000000001",
  8355=>"111111111",
  8356=>"110110110",
  8357=>"000100111",
  8358=>"000000000",
  8359=>"100100110",
  8360=>"111111000",
  8361=>"111011111",
  8362=>"000000000",
  8363=>"111001111",
  8364=>"111111111",
  8365=>"110101000",
  8366=>"111111111",
  8367=>"010001000",
  8368=>"000011001",
  8369=>"000110111",
  8370=>"110110000",
  8371=>"000000000",
  8372=>"001000000",
  8373=>"000000000",
  8374=>"000000000",
  8375=>"000000000",
  8376=>"000111101",
  8377=>"110100100",
  8378=>"111001000",
  8379=>"000010110",
  8380=>"111011010",
  8381=>"110010111",
  8382=>"000000000",
  8383=>"000011000",
  8384=>"010000000",
  8385=>"111111111",
  8386=>"011111001",
  8387=>"110110000",
  8388=>"111011011",
  8389=>"111111010",
  8390=>"111111110",
  8391=>"000000000",
  8392=>"000000000",
  8393=>"100101101",
  8394=>"001001110",
  8395=>"111111000",
  8396=>"111111111",
  8397=>"100100000",
  8398=>"000010010",
  8399=>"111111101",
  8400=>"001011111",
  8401=>"111111010",
  8402=>"111111111",
  8403=>"111111111",
  8404=>"001101111",
  8405=>"000100000",
  8406=>"111110000",
  8407=>"001000001",
  8408=>"000000000",
  8409=>"100111101",
  8410=>"000000010",
  8411=>"000011110",
  8412=>"111111111",
  8413=>"110100000",
  8414=>"111110000",
  8415=>"000001001",
  8416=>"000000000",
  8417=>"000011001",
  8418=>"111011000",
  8419=>"011011111",
  8420=>"111111111",
  8421=>"000100100",
  8422=>"111111111",
  8423=>"110111000",
  8424=>"111111111",
  8425=>"000000000",
  8426=>"000111111",
  8427=>"111111111",
  8428=>"111111111",
  8429=>"000100111",
  8430=>"111111111",
  8431=>"100111000",
  8432=>"010011110",
  8433=>"000000100",
  8434=>"111010110",
  8435=>"011110100",
  8436=>"001011000",
  8437=>"101111101",
  8438=>"010000000",
  8439=>"000000010",
  8440=>"111111111",
  8441=>"001000000",
  8442=>"110111111",
  8443=>"010010001",
  8444=>"110110110",
  8445=>"000000100",
  8446=>"111111111",
  8447=>"000000000",
  8448=>"000000000",
  8449=>"110100100",
  8450=>"100100000",
  8451=>"111111111",
  8452=>"100110110",
  8453=>"110111011",
  8454=>"000000000",
  8455=>"110111001",
  8456=>"110110001",
  8457=>"000000000",
  8458=>"011011111",
  8459=>"001000101",
  8460=>"111111100",
  8461=>"000000000",
  8462=>"110000000",
  8463=>"000000010",
  8464=>"000000110",
  8465=>"000000000",
  8466=>"111111111",
  8467=>"000000001",
  8468=>"111111101",
  8469=>"111011011",
  8470=>"111111111",
  8471=>"000000000",
  8472=>"111101001",
  8473=>"000111000",
  8474=>"000001001",
  8475=>"000100111",
  8476=>"111111111",
  8477=>"111011111",
  8478=>"000000001",
  8479=>"111001000",
  8480=>"000000000",
  8481=>"000000000",
  8482=>"000000111",
  8483=>"000000000",
  8484=>"100110000",
  8485=>"000000111",
  8486=>"111111111",
  8487=>"000000000",
  8488=>"111111000",
  8489=>"001111111",
  8490=>"110011000",
  8491=>"000000000",
  8492=>"000000000",
  8493=>"110011101",
  8494=>"111100000",
  8495=>"000000000",
  8496=>"000110011",
  8497=>"011011000",
  8498=>"010000000",
  8499=>"100100000",
  8500=>"000000000",
  8501=>"111011000",
  8502=>"111111111",
  8503=>"000111011",
  8504=>"000000000",
  8505=>"000000100",
  8506=>"111000000",
  8507=>"111111111",
  8508=>"111011011",
  8509=>"001001000",
  8510=>"110000000",
  8511=>"000000000",
  8512=>"101000000",
  8513=>"010111111",
  8514=>"001011111",
  8515=>"000000000",
  8516=>"010000111",
  8517=>"010000111",
  8518=>"000000000",
  8519=>"000100100",
  8520=>"000000000",
  8521=>"111111000",
  8522=>"000001011",
  8523=>"000000100",
  8524=>"000000000",
  8525=>"110111001",
  8526=>"011011001",
  8527=>"000000000",
  8528=>"111111111",
  8529=>"000000000",
  8530=>"000010110",
  8531=>"110110000",
  8532=>"111111111",
  8533=>"001001011",
  8534=>"000000000",
  8535=>"100110000",
  8536=>"011000000",
  8537=>"000000000",
  8538=>"000110000",
  8539=>"000000101",
  8540=>"100000000",
  8541=>"000000000",
  8542=>"000011111",
  8543=>"110110000",
  8544=>"111100001",
  8545=>"111111111",
  8546=>"101000100",
  8547=>"111000010",
  8548=>"000100000",
  8549=>"000000000",
  8550=>"111111111",
  8551=>"000000100",
  8552=>"111111100",
  8553=>"000000000",
  8554=>"111111111",
  8555=>"110000001",
  8556=>"100110111",
  8557=>"000000000",
  8558=>"111111010",
  8559=>"111100100",
  8560=>"000000000",
  8561=>"010000000",
  8562=>"111011010",
  8563=>"100110100",
  8564=>"111111111",
  8565=>"111101001",
  8566=>"111111111",
  8567=>"111111111",
  8568=>"111111111",
  8569=>"111111011",
  8570=>"000000000",
  8571=>"001011111",
  8572=>"000000001",
  8573=>"011000000",
  8574=>"000010111",
  8575=>"111110000",
  8576=>"000110111",
  8577=>"011011011",
  8578=>"000000000",
  8579=>"100100000",
  8580=>"111111100",
  8581=>"001001011",
  8582=>"000011111",
  8583=>"111111000",
  8584=>"000000100",
  8585=>"111111111",
  8586=>"000000000",
  8587=>"110110011",
  8588=>"001011111",
  8589=>"110100110",
  8590=>"010000011",
  8591=>"111111000",
  8592=>"000000000",
  8593=>"000000000",
  8594=>"000000000",
  8595=>"100100110",
  8596=>"000011111",
  8597=>"000010000",
  8598=>"011011011",
  8599=>"111111111",
  8600=>"010000000",
  8601=>"010000000",
  8602=>"111111111",
  8603=>"000000000",
  8604=>"010000111",
  8605=>"111111111",
  8606=>"111000011",
  8607=>"000000000",
  8608=>"000000000",
  8609=>"110110110",
  8610=>"000111111",
  8611=>"111111111",
  8612=>"000110111",
  8613=>"000111111",
  8614=>"000000000",
  8615=>"110010000",
  8616=>"000010010",
  8617=>"110111111",
  8618=>"111011111",
  8619=>"111111001",
  8620=>"111111111",
  8621=>"001111011",
  8622=>"100111110",
  8623=>"111111111",
  8624=>"000000000",
  8625=>"111111110",
  8626=>"000000000",
  8627=>"000010010",
  8628=>"011010000",
  8629=>"111111111",
  8630=>"111111111",
  8631=>"000001000",
  8632=>"000111111",
  8633=>"000111111",
  8634=>"111111111",
  8635=>"000000000",
  8636=>"000000000",
  8637=>"100001001",
  8638=>"111011001",
  8639=>"111111111",
  8640=>"111111111",
  8641=>"000000000",
  8642=>"000000000",
  8643=>"000000000",
  8644=>"000000100",
  8645=>"001001011",
  8646=>"111111111",
  8647=>"000000000",
  8648=>"000110111",
  8649=>"001011011",
  8650=>"000000101",
  8651=>"111111111",
  8652=>"110000000",
  8653=>"011011111",
  8654=>"001000001",
  8655=>"000000010",
  8656=>"111111011",
  8657=>"011111111",
  8658=>"111001001",
  8659=>"000000000",
  8660=>"000000000",
  8661=>"011111111",
  8662=>"001111001",
  8663=>"000001111",
  8664=>"001000101",
  8665=>"000000000",
  8666=>"000000000",
  8667=>"111011011",
  8668=>"000000000",
  8669=>"010010000",
  8670=>"000000000",
  8671=>"111111111",
  8672=>"111111111",
  8673=>"110111100",
  8674=>"000000000",
  8675=>"111111111",
  8676=>"111111111",
  8677=>"111111111",
  8678=>"000100000",
  8679=>"000000000",
  8680=>"111000000",
  8681=>"000000000",
  8682=>"101000000",
  8683=>"000000001",
  8684=>"101001001",
  8685=>"001101101",
  8686=>"110111111",
  8687=>"111111100",
  8688=>"111111111",
  8689=>"010010010",
  8690=>"111000111",
  8691=>"101111011",
  8692=>"011111111",
  8693=>"000001001",
  8694=>"111111111",
  8695=>"111110000",
  8696=>"101010000",
  8697=>"000101110",
  8698=>"000000001",
  8699=>"000000000",
  8700=>"000110111",
  8701=>"000000000",
  8702=>"000011011",
  8703=>"000000001",
  8704=>"111111111",
  8705=>"111111110",
  8706=>"000000000",
  8707=>"000000000",
  8708=>"100100001",
  8709=>"000100101",
  8710=>"001111111",
  8711=>"000000000",
  8712=>"000011000",
  8713=>"110111111",
  8714=>"111010000",
  8715=>"000000000",
  8716=>"000000001",
  8717=>"000000000",
  8718=>"000001001",
  8719=>"000101101",
  8720=>"000000000",
  8721=>"000000001",
  8722=>"000011110",
  8723=>"000000000",
  8724=>"111111000",
  8725=>"000000101",
  8726=>"000000000",
  8727=>"001000000",
  8728=>"110110110",
  8729=>"111111110",
  8730=>"000000000",
  8731=>"111111111",
  8732=>"000000000",
  8733=>"111000000",
  8734=>"111111111",
  8735=>"000110111",
  8736=>"111111111",
  8737=>"000000000",
  8738=>"110101001",
  8739=>"111111111",
  8740=>"111111111",
  8741=>"000100111",
  8742=>"000000000",
  8743=>"000111011",
  8744=>"100000000",
  8745=>"000000000",
  8746=>"111111111",
  8747=>"001011000",
  8748=>"100100001",
  8749=>"000100000",
  8750=>"111111110",
  8751=>"000000001",
  8752=>"111111111",
  8753=>"000111111",
  8754=>"001001000",
  8755=>"000000000",
  8756=>"000000000",
  8757=>"111011011",
  8758=>"000000000",
  8759=>"001101111",
  8760=>"001001000",
  8761=>"000111111",
  8762=>"111111111",
  8763=>"110010000",
  8764=>"001001111",
  8765=>"011110110",
  8766=>"011011011",
  8767=>"111111111",
  8768=>"000000000",
  8769=>"000011111",
  8770=>"101000000",
  8771=>"111111010",
  8772=>"111111111",
  8773=>"111111111",
  8774=>"000000110",
  8775=>"111111110",
  8776=>"111111111",
  8777=>"000000000",
  8778=>"111011001",
  8779=>"010000000",
  8780=>"111111111",
  8781=>"111111111",
  8782=>"110110111",
  8783=>"000001001",
  8784=>"001111111",
  8785=>"111111111",
  8786=>"000000000",
  8787=>"000000000",
  8788=>"000000000",
  8789=>"110110100",
  8790=>"010110111",
  8791=>"111111111",
  8792=>"111111111",
  8793=>"111101100",
  8794=>"000010010",
  8795=>"010111111",
  8796=>"111111111",
  8797=>"100001000",
  8798=>"111111100",
  8799=>"001000000",
  8800=>"100100010",
  8801=>"000000100",
  8802=>"001000000",
  8803=>"111111010",
  8804=>"111111111",
  8805=>"110110010",
  8806=>"000110111",
  8807=>"110111111",
  8808=>"000000000",
  8809=>"000000000",
  8810=>"110110000",
  8811=>"000000000",
  8812=>"000000000",
  8813=>"111111111",
  8814=>"111111111",
  8815=>"111111000",
  8816=>"000000000",
  8817=>"111111111",
  8818=>"110010000",
  8819=>"101100101",
  8820=>"000000000",
  8821=>"000000000",
  8822=>"111111100",
  8823=>"000000000",
  8824=>"111001000",
  8825=>"111111111",
  8826=>"000000000",
  8827=>"000000000",
  8828=>"110110110",
  8829=>"000000000",
  8830=>"111000000",
  8831=>"000000000",
  8832=>"111111111",
  8833=>"111111111",
  8834=>"001000000",
  8835=>"001011011",
  8836=>"000000101",
  8837=>"111111101",
  8838=>"111111111",
  8839=>"110111111",
  8840=>"000000000",
  8841=>"000000100",
  8842=>"111111111",
  8843=>"110110111",
  8844=>"111111111",
  8845=>"110110100",
  8846=>"110110100",
  8847=>"000000000",
  8848=>"111111111",
  8849=>"000100000",
  8850=>"000000011",
  8851=>"111111111",
  8852=>"000000000",
  8853=>"011011011",
  8854=>"111111111",
  8855=>"000000001",
  8856=>"000000000",
  8857=>"100110110",
  8858=>"111111111",
  8859=>"110000001",
  8860=>"001101000",
  8861=>"111110110",
  8862=>"110000100",
  8863=>"111111101",
  8864=>"000010100",
  8865=>"010011001",
  8866=>"000000000",
  8867=>"111111101",
  8868=>"000000000",
  8869=>"000110110",
  8870=>"000000000",
  8871=>"011110110",
  8872=>"000000000",
  8873=>"000000001",
  8874=>"101101100",
  8875=>"000000101",
  8876=>"000000000",
  8877=>"111101101",
  8878=>"000000001",
  8879=>"111110000",
  8880=>"001111000",
  8881=>"001001000",
  8882=>"000001000",
  8883=>"000000101",
  8884=>"010111111",
  8885=>"001011001",
  8886=>"000001000",
  8887=>"011111111",
  8888=>"111111110",
  8889=>"000000000",
  8890=>"000011011",
  8891=>"000000000",
  8892=>"100111111",
  8893=>"000000000",
  8894=>"111111110",
  8895=>"111111111",
  8896=>"001000000",
  8897=>"111111111",
  8898=>"111111111",
  8899=>"111111111",
  8900=>"111111111",
  8901=>"000000000",
  8902=>"011000000",
  8903=>"000111000",
  8904=>"000000000",
  8905=>"000000000",
  8906=>"000000101",
  8907=>"000000000",
  8908=>"000000000",
  8909=>"111111111",
  8910=>"000000000",
  8911=>"000000000",
  8912=>"110000000",
  8913=>"111111111",
  8914=>"111111111",
  8915=>"000000000",
  8916=>"111111111",
  8917=>"110000000",
  8918=>"000000010",
  8919=>"101111111",
  8920=>"111111111",
  8921=>"110110000",
  8922=>"111011111",
  8923=>"000000000",
  8924=>"111111111",
  8925=>"000000000",
  8926=>"000000000",
  8927=>"111111111",
  8928=>"111101110",
  8929=>"000000000",
  8930=>"111010011",
  8931=>"000000000",
  8932=>"111101000",
  8933=>"100111111",
  8934=>"000111111",
  8935=>"011100000",
  8936=>"111111111",
  8937=>"111110100",
  8938=>"101100000",
  8939=>"110110100",
  8940=>"111111111",
  8941=>"001000000",
  8942=>"111111111",
  8943=>"000000111",
  8944=>"111111001",
  8945=>"111111111",
  8946=>"101100111",
  8947=>"000011011",
  8948=>"000000000",
  8949=>"000011001",
  8950=>"001100111",
  8951=>"000000000",
  8952=>"111111011",
  8953=>"111111111",
  8954=>"000000000",
  8955=>"000000000",
  8956=>"000000110",
  8957=>"001001111",
  8958=>"000101111",
  8959=>"010010000",
  8960=>"000000000",
  8961=>"000000000",
  8962=>"000111111",
  8963=>"000011111",
  8964=>"000000000",
  8965=>"111111111",
  8966=>"000000000",
  8967=>"111111111",
  8968=>"010111000",
  8969=>"000000000",
  8970=>"001001000",
  8971=>"111111111",
  8972=>"000001000",
  8973=>"000011111",
  8974=>"000000011",
  8975=>"000000000",
  8976=>"111111111",
  8977=>"000000000",
  8978=>"000000100",
  8979=>"000000000",
  8980=>"111101111",
  8981=>"101111000",
  8982=>"101001101",
  8983=>"111111000",
  8984=>"110110100",
  8985=>"111010010",
  8986=>"111111001",
  8987=>"000010111",
  8988=>"111111111",
  8989=>"001100101",
  8990=>"000001001",
  8991=>"000000000",
  8992=>"011111001",
  8993=>"111111111",
  8994=>"000000000",
  8995=>"000000000",
  8996=>"000000000",
  8997=>"001010000",
  8998=>"011011011",
  8999=>"100100000",
  9000=>"100111111",
  9001=>"000000011",
  9002=>"110111000",
  9003=>"111111111",
  9004=>"011111111",
  9005=>"100000000",
  9006=>"111111111",
  9007=>"000110000",
  9008=>"000000001",
  9009=>"111111111",
  9010=>"111011111",
  9011=>"110110000",
  9012=>"000001010",
  9013=>"110110110",
  9014=>"000100000",
  9015=>"000000000",
  9016=>"001001000",
  9017=>"101000000",
  9018=>"000000000",
  9019=>"011000000",
  9020=>"000101111",
  9021=>"111100100",
  9022=>"011011111",
  9023=>"111111111",
  9024=>"111100100",
  9025=>"000000000",
  9026=>"000000000",
  9027=>"100100101",
  9028=>"111111111",
  9029=>"000000000",
  9030=>"000000000",
  9031=>"000000100",
  9032=>"000000000",
  9033=>"011000000",
  9034=>"111010000",
  9035=>"100110100",
  9036=>"110000000",
  9037=>"111111101",
  9038=>"000000000",
  9039=>"111111111",
  9040=>"110111111",
  9041=>"110110110",
  9042=>"111000000",
  9043=>"100111110",
  9044=>"001000000",
  9045=>"011001011",
  9046=>"000000000",
  9047=>"111101111",
  9048=>"111111111",
  9049=>"111111001",
  9050=>"011111111",
  9051=>"001010000",
  9052=>"000110111",
  9053=>"000000000",
  9054=>"000000000",
  9055=>"000000001",
  9056=>"000000000",
  9057=>"000000111",
  9058=>"011111100",
  9059=>"111111111",
  9060=>"111011011",
  9061=>"000000001",
  9062=>"111000000",
  9063=>"111111110",
  9064=>"010111011",
  9065=>"111110111",
  9066=>"111111111",
  9067=>"000000000",
  9068=>"100000000",
  9069=>"000000001",
  9070=>"100111111",
  9071=>"000000000",
  9072=>"000000100",
  9073=>"000000010",
  9074=>"000111111",
  9075=>"111111111",
  9076=>"001111111",
  9077=>"000000000",
  9078=>"000000000",
  9079=>"000000000",
  9080=>"101001000",
  9081=>"000000000",
  9082=>"111111110",
  9083=>"000001011",
  9084=>"101110111",
  9085=>"000000000",
  9086=>"000001011",
  9087=>"101000101",
  9088=>"001001000",
  9089=>"111111001",
  9090=>"011111111",
  9091=>"000000111",
  9092=>"000000000",
  9093=>"111111111",
  9094=>"111110110",
  9095=>"000000000",
  9096=>"111111101",
  9097=>"001001000",
  9098=>"111111111",
  9099=>"000000000",
  9100=>"101111111",
  9101=>"000000101",
  9102=>"111111111",
  9103=>"000000011",
  9104=>"000000000",
  9105=>"000000111",
  9106=>"000000000",
  9107=>"000011111",
  9108=>"000000000",
  9109=>"000000000",
  9110=>"001000001",
  9111=>"001111000",
  9112=>"101111011",
  9113=>"011111111",
  9114=>"000000000",
  9115=>"000000000",
  9116=>"111111111",
  9117=>"000000000",
  9118=>"001001000",
  9119=>"111000000",
  9120=>"000011000",
  9121=>"011011000",
  9122=>"000000111",
  9123=>"111111111",
  9124=>"001111111",
  9125=>"111111011",
  9126=>"111111111",
  9127=>"010110111",
  9128=>"111111111",
  9129=>"001111111",
  9130=>"000000111",
  9131=>"000000000",
  9132=>"011001111",
  9133=>"000000000",
  9134=>"000010010",
  9135=>"111110000",
  9136=>"111110000",
  9137=>"000111011",
  9138=>"111111100",
  9139=>"001101100",
  9140=>"001001101",
  9141=>"000010000",
  9142=>"000100100",
  9143=>"111111111",
  9144=>"100100111",
  9145=>"000000000",
  9146=>"000100110",
  9147=>"000100111",
  9148=>"000000000",
  9149=>"111011000",
  9150=>"110111111",
  9151=>"001011101",
  9152=>"100000111",
  9153=>"000000000",
  9154=>"000000000",
  9155=>"111111011",
  9156=>"111100000",
  9157=>"000000001",
  9158=>"110111000",
  9159=>"000000000",
  9160=>"000000000",
  9161=>"011011011",
  9162=>"111101111",
  9163=>"111111000",
  9164=>"000000000",
  9165=>"111111111",
  9166=>"010000111",
  9167=>"010011011",
  9168=>"000000000",
  9169=>"111111101",
  9170=>"110111111",
  9171=>"111000000",
  9172=>"111111111",
  9173=>"111101000",
  9174=>"101100000",
  9175=>"011111100",
  9176=>"111101101",
  9177=>"000000100",
  9178=>"000000000",
  9179=>"011000000",
  9180=>"000001111",
  9181=>"111001001",
  9182=>"111111111",
  9183=>"111111111",
  9184=>"100100000",
  9185=>"111111111",
  9186=>"000100110",
  9187=>"111111111",
  9188=>"111100001",
  9189=>"000010110",
  9190=>"111000101",
  9191=>"111111000",
  9192=>"100101101",
  9193=>"000000011",
  9194=>"000000000",
  9195=>"000000000",
  9196=>"000000001",
  9197=>"000000110",
  9198=>"001001001",
  9199=>"111111101",
  9200=>"000000000",
  9201=>"111111111",
  9202=>"011001001",
  9203=>"110111111",
  9204=>"111111111",
  9205=>"111111111",
  9206=>"011111111",
  9207=>"100100110",
  9208=>"000000000",
  9209=>"100101111",
  9210=>"111111111",
  9211=>"111111001",
  9212=>"001001001",
  9213=>"000111111",
  9214=>"000000000",
  9215=>"111110110",
  9216=>"000101110",
  9217=>"000000000",
  9218=>"101000000",
  9219=>"111111111",
  9220=>"110000000",
  9221=>"000000110",
  9222=>"000000000",
  9223=>"111111111",
  9224=>"000000111",
  9225=>"111111000",
  9226=>"000000000",
  9227=>"001011011",
  9228=>"000110110",
  9229=>"111000000",
  9230=>"110111111",
  9231=>"011000000",
  9232=>"000000110",
  9233=>"100111111",
  9234=>"000011011",
  9235=>"000000000",
  9236=>"111011000",
  9237=>"111111101",
  9238=>"111110100",
  9239=>"000000001",
  9240=>"000000111",
  9241=>"001001011",
  9242=>"100000000",
  9243=>"011111111",
  9244=>"000000100",
  9245=>"011100111",
  9246=>"011001010",
  9247=>"111110100",
  9248=>"101000000",
  9249=>"100100001",
  9250=>"110110110",
  9251=>"111111000",
  9252=>"001111111",
  9253=>"000100111",
  9254=>"000000000",
  9255=>"111011100",
  9256=>"000000111",
  9257=>"000000111",
  9258=>"000000000",
  9259=>"110110000",
  9260=>"000000000",
  9261=>"111111000",
  9262=>"000000000",
  9263=>"000010111",
  9264=>"000000000",
  9265=>"000000000",
  9266=>"100111011",
  9267=>"100100100",
  9268=>"000000000",
  9269=>"010000000",
  9270=>"100000111",
  9271=>"111111011",
  9272=>"011111110",
  9273=>"111000100",
  9274=>"000000011",
  9275=>"000111100",
  9276=>"000000111",
  9277=>"111000000",
  9278=>"110111000",
  9279=>"001000000",
  9280=>"001111111",
  9281=>"111111001",
  9282=>"111111111",
  9283=>"111000000",
  9284=>"110111111",
  9285=>"001011111",
  9286=>"111000000",
  9287=>"000000111",
  9288=>"000000011",
  9289=>"000000000",
  9290=>"111111110",
  9291=>"100000111",
  9292=>"011001000",
  9293=>"000111111",
  9294=>"000000000",
  9295=>"000010000",
  9296=>"111000000",
  9297=>"111111100",
  9298=>"000000111",
  9299=>"000000001",
  9300=>"000000000",
  9301=>"000000000",
  9302=>"001000111",
  9303=>"111111111",
  9304=>"000000000",
  9305=>"111011001",
  9306=>"111110000",
  9307=>"000110100",
  9308=>"111111010",
  9309=>"001011111",
  9310=>"001010111",
  9311=>"111111111",
  9312=>"111000000",
  9313=>"111111000",
  9314=>"001110111",
  9315=>"000000000",
  9316=>"000000000",
  9317=>"100000000",
  9318=>"111111111",
  9319=>"000000001",
  9320=>"111111111",
  9321=>"100000110",
  9322=>"111010000",
  9323=>"000000111",
  9324=>"000010010",
  9325=>"111001000",
  9326=>"011000001",
  9327=>"000000001",
  9328=>"100110000",
  9329=>"111000000",
  9330=>"111111100",
  9331=>"111000111",
  9332=>"000000000",
  9333=>"000000000",
  9334=>"111000111",
  9335=>"000000110",
  9336=>"100000001",
  9337=>"000000000",
  9338=>"000000011",
  9339=>"011000000",
  9340=>"011001000",
  9341=>"010111011",
  9342=>"000000111",
  9343=>"000111111",
  9344=>"111000000",
  9345=>"001000001",
  9346=>"010110110",
  9347=>"100000001",
  9348=>"000001111",
  9349=>"100000000",
  9350=>"100000100",
  9351=>"000000011",
  9352=>"001001111",
  9353=>"010000000",
  9354=>"000111111",
  9355=>"000000111",
  9356=>"000001111",
  9357=>"110111111",
  9358=>"001001111",
  9359=>"110110111",
  9360=>"000000000",
  9361=>"111111111",
  9362=>"000111111",
  9363=>"111110101",
  9364=>"011000111",
  9365=>"000111011",
  9366=>"111010000",
  9367=>"111000010",
  9368=>"000111000",
  9369=>"100101111",
  9370=>"000000010",
  9371=>"110000000",
  9372=>"000000000",
  9373=>"110100000",
  9374=>"000000001",
  9375=>"000000000",
  9376=>"111101111",
  9377=>"111000000",
  9378=>"000000000",
  9379=>"111111111",
  9380=>"000011111",
  9381=>"000000110",
  9382=>"000111111",
  9383=>"111100100",
  9384=>"111000000",
  9385=>"000111111",
  9386=>"111000100",
  9387=>"110111111",
  9388=>"000001011",
  9389=>"111111110",
  9390=>"110000001",
  9391=>"101111011",
  9392=>"000000000",
  9393=>"111001100",
  9394=>"111111111",
  9395=>"000000000",
  9396=>"111100100",
  9397=>"111111111",
  9398=>"011111111",
  9399=>"011110011",
  9400=>"111000101",
  9401=>"001111111",
  9402=>"100000000",
  9403=>"111110000",
  9404=>"000000000",
  9405=>"000000000",
  9406=>"011110000",
  9407=>"001000000",
  9408=>"001001011",
  9409=>"010000100",
  9410=>"000100100",
  9411=>"001000101",
  9412=>"001000000",
  9413=>"000111110",
  9414=>"000000000",
  9415=>"100001101",
  9416=>"110110000",
  9417=>"000000000",
  9418=>"001001111",
  9419=>"000010110",
  9420=>"111110100",
  9421=>"111101000",
  9422=>"000110111",
  9423=>"000000100",
  9424=>"000000000",
  9425=>"000000000",
  9426=>"000010111",
  9427=>"000000000",
  9428=>"111101111",
  9429=>"111000000",
  9430=>"011000000",
  9431=>"000000111",
  9432=>"000000000",
  9433=>"000000000",
  9434=>"111100000",
  9435=>"011111110",
  9436=>"111111011",
  9437=>"011001000",
  9438=>"111111000",
  9439=>"000000000",
  9440=>"000000000",
  9441=>"000000111",
  9442=>"101100111",
  9443=>"111000000",
  9444=>"111111001",
  9445=>"111010100",
  9446=>"111010111",
  9447=>"110110111",
  9448=>"000000111",
  9449=>"111001001",
  9450=>"111100000",
  9451=>"000011111",
  9452=>"000000111",
  9453=>"011010000",
  9454=>"000100101",
  9455=>"101000000",
  9456=>"000001000",
  9457=>"011000000",
  9458=>"111111101",
  9459=>"111111111",
  9460=>"111111000",
  9461=>"001111110",
  9462=>"100110100",
  9463=>"111111111",
  9464=>"111011111",
  9465=>"011111111",
  9466=>"111110111",
  9467=>"111111111",
  9468=>"110111111",
  9469=>"011010000",
  9470=>"111111111",
  9471=>"111001000",
  9472=>"000000101",
  9473=>"011111110",
  9474=>"001001000",
  9475=>"111110000",
  9476=>"000000000",
  9477=>"100000000",
  9478=>"111000000",
  9479=>"001000111",
  9480=>"111111000",
  9481=>"111111000",
  9482=>"111000000",
  9483=>"111111001",
  9484=>"001000000",
  9485=>"000001111",
  9486=>"011101111",
  9487=>"111111111",
  9488=>"111100000",
  9489=>"001011111",
  9490=>"001000000",
  9491=>"111110000",
  9492=>"011111000",
  9493=>"010000111",
  9494=>"110110110",
  9495=>"001111111",
  9496=>"111111111",
  9497=>"111110110",
  9498=>"011000010",
  9499=>"000010011",
  9500=>"000100110",
  9501=>"000000001",
  9502=>"010000000",
  9503=>"111111111",
  9504=>"111011001",
  9505=>"111111000",
  9506=>"111111111",
  9507=>"100111111",
  9508=>"000011111",
  9509=>"000110111",
  9510=>"010000010",
  9511=>"100110011",
  9512=>"011000000",
  9513=>"000000000",
  9514=>"100000000",
  9515=>"110100010",
  9516=>"001000000",
  9517=>"000111111",
  9518=>"000000110",
  9519=>"010000100",
  9520=>"111111111",
  9521=>"000000001",
  9522=>"111000111",
  9523=>"111001000",
  9524=>"111110110",
  9525=>"111000110",
  9526=>"111000100",
  9527=>"111000000",
  9528=>"100110000",
  9529=>"101000100",
  9530=>"000000000",
  9531=>"111100000",
  9532=>"010011111",
  9533=>"000000111",
  9534=>"000000010",
  9535=>"111111001",
  9536=>"111000000",
  9537=>"000000011",
  9538=>"111101010",
  9539=>"111000000",
  9540=>"111000000",
  9541=>"000000000",
  9542=>"000111100",
  9543=>"110000000",
  9544=>"001011111",
  9545=>"000000110",
  9546=>"000000110",
  9547=>"100100001",
  9548=>"011010000",
  9549=>"100000000",
  9550=>"011011000",
  9551=>"100110111",
  9552=>"110111111",
  9553=>"111111111",
  9554=>"111111111",
  9555=>"101111111",
  9556=>"000011101",
  9557=>"011000111",
  9558=>"111110110",
  9559=>"111111111",
  9560=>"000001111",
  9561=>"100000000",
  9562=>"111111111",
  9563=>"000111111",
  9564=>"000100100",
  9565=>"001000000",
  9566=>"101000000",
  9567=>"110110111",
  9568=>"111000000",
  9569=>"011111111",
  9570=>"110000111",
  9571=>"000000111",
  9572=>"000000101",
  9573=>"111000000",
  9574=>"111111010",
  9575=>"000000001",
  9576=>"000000000",
  9577=>"100000000",
  9578=>"000000000",
  9579=>"111001000",
  9580=>"011111111",
  9581=>"100000000",
  9582=>"111011011",
  9583=>"000011111",
  9584=>"000011111",
  9585=>"110000010",
  9586=>"111000000",
  9587=>"000111000",
  9588=>"111111111",
  9589=>"111111000",
  9590=>"001110000",
  9591=>"011101111",
  9592=>"111000000",
  9593=>"111111111",
  9594=>"000011011",
  9595=>"111111000",
  9596=>"000001011",
  9597=>"000000000",
  9598=>"111111000",
  9599=>"001000000",
  9600=>"111111001",
  9601=>"111111111",
  9602=>"000010111",
  9603=>"000000000",
  9604=>"001111011",
  9605=>"111100000",
  9606=>"001011001",
  9607=>"000000000",
  9608=>"111000000",
  9609=>"000011000",
  9610=>"000000000",
  9611=>"110111000",
  9612=>"111111111",
  9613=>"000110000",
  9614=>"000000000",
  9615=>"000000000",
  9616=>"111111111",
  9617=>"000000000",
  9618=>"100111111",
  9619=>"001011111",
  9620=>"111111111",
  9621=>"000000000",
  9622=>"000000000",
  9623=>"111011001",
  9624=>"000000111",
  9625=>"110010011",
  9626=>"111100000",
  9627=>"111111000",
  9628=>"000001111",
  9629=>"111111111",
  9630=>"000000000",
  9631=>"000000010",
  9632=>"010011000",
  9633=>"110011001",
  9634=>"000000001",
  9635=>"111100000",
  9636=>"111000110",
  9637=>"000000100",
  9638=>"100000000",
  9639=>"111000011",
  9640=>"000000100",
  9641=>"000111111",
  9642=>"000111110",
  9643=>"111111101",
  9644=>"000000001",
  9645=>"101000000",
  9646=>"011000000",
  9647=>"000011000",
  9648=>"000000001",
  9649=>"011000000",
  9650=>"000000000",
  9651=>"000000001",
  9652=>"111111111",
  9653=>"111111101",
  9654=>"100111111",
  9655=>"000000010",
  9656=>"110000000",
  9657=>"101100111",
  9658=>"011011111",
  9659=>"010000100",
  9660=>"000000000",
  9661=>"111000001",
  9662=>"000000000",
  9663=>"001000000",
  9664=>"111110000",
  9665=>"000000000",
  9666=>"100000010",
  9667=>"111001011",
  9668=>"000100101",
  9669=>"011011000",
  9670=>"000000000",
  9671=>"111000000",
  9672=>"000101111",
  9673=>"111011110",
  9674=>"111001111",
  9675=>"000000100",
  9676=>"000000111",
  9677=>"011001001",
  9678=>"111111011",
  9679=>"100110110",
  9680=>"000000000",
  9681=>"001011010",
  9682=>"100000001",
  9683=>"111011011",
  9684=>"100110111",
  9685=>"011000000",
  9686=>"101000000",
  9687=>"001001000",
  9688=>"111000000",
  9689=>"111000000",
  9690=>"001111111",
  9691=>"111110110",
  9692=>"000000100",
  9693=>"101111001",
  9694=>"001000000",
  9695=>"000000110",
  9696=>"000000000",
  9697=>"000001000",
  9698=>"000001001",
  9699=>"101111111",
  9700=>"111011111",
  9701=>"000000111",
  9702=>"111111011",
  9703=>"001011011",
  9704=>"100100100",
  9705=>"110010000",
  9706=>"110000001",
  9707=>"000011111",
  9708=>"100100110",
  9709=>"111111001",
  9710=>"100110111",
  9711=>"110000000",
  9712=>"000110110",
  9713=>"000011011",
  9714=>"101000001",
  9715=>"110000000",
  9716=>"011111111",
  9717=>"000000000",
  9718=>"111010000",
  9719=>"001001110",
  9720=>"101111111",
  9721=>"000000000",
  9722=>"000110000",
  9723=>"000000111",
  9724=>"000000000",
  9725=>"111111010",
  9726=>"000000111",
  9727=>"011000000",
  9728=>"111000000",
  9729=>"000000000",
  9730=>"000000000",
  9731=>"000001110",
  9732=>"000011000",
  9733=>"111000000",
  9734=>"000101111",
  9735=>"110000000",
  9736=>"111111111",
  9737=>"000010000",
  9738=>"000100111",
  9739=>"011000001",
  9740=>"000100111",
  9741=>"000111010",
  9742=>"100000101",
  9743=>"000000000",
  9744=>"011001111",
  9745=>"000111111",
  9746=>"001111111",
  9747=>"111001001",
  9748=>"100000111",
  9749=>"000000000",
  9750=>"000000000",
  9751=>"101001011",
  9752=>"000000100",
  9753=>"001001111",
  9754=>"111000000",
  9755=>"011111100",
  9756=>"000000000",
  9757=>"110111100",
  9758=>"000001000",
  9759=>"110111000",
  9760=>"000000000",
  9761=>"100100000",
  9762=>"000100001",
  9763=>"000010111",
  9764=>"000000000",
  9765=>"111111001",
  9766=>"110110111",
  9767=>"111101001",
  9768=>"010100000",
  9769=>"000000000",
  9770=>"111111111",
  9771=>"110110111",
  9772=>"111101111",
  9773=>"111111000",
  9774=>"000000111",
  9775=>"111111110",
  9776=>"111100000",
  9777=>"000111111",
  9778=>"011001001",
  9779=>"111111100",
  9780=>"000000101",
  9781=>"000111111",
  9782=>"000000001",
  9783=>"011000000",
  9784=>"000100110",
  9785=>"101100000",
  9786=>"000000010",
  9787=>"001000010",
  9788=>"000000000",
  9789=>"111111110",
  9790=>"000001110",
  9791=>"000000000",
  9792=>"011101110",
  9793=>"000011011",
  9794=>"000000000",
  9795=>"110100000",
  9796=>"000000000",
  9797=>"001001111",
  9798=>"000000000",
  9799=>"111111111",
  9800=>"001000000",
  9801=>"111100011",
  9802=>"111111111",
  9803=>"000000111",
  9804=>"110110000",
  9805=>"000000011",
  9806=>"111000000",
  9807=>"111111111",
  9808=>"000000101",
  9809=>"111111111",
  9810=>"000100100",
  9811=>"000001000",
  9812=>"000111000",
  9813=>"000000000",
  9814=>"110111111",
  9815=>"000111111",
  9816=>"110110000",
  9817=>"101000100",
  9818=>"111111000",
  9819=>"110100000",
  9820=>"001000110",
  9821=>"111111000",
  9822=>"000100101",
  9823=>"000110111",
  9824=>"001111111",
  9825=>"000000000",
  9826=>"000000011",
  9827=>"000000000",
  9828=>"000000110",
  9829=>"000000111",
  9830=>"111111111",
  9831=>"000000000",
  9832=>"000000000",
  9833=>"111000111",
  9834=>"111111000",
  9835=>"001001001",
  9836=>"000001111",
  9837=>"111111111",
  9838=>"000000011",
  9839=>"100100011",
  9840=>"111111111",
  9841=>"000000001",
  9842=>"000000000",
  9843=>"010000100",
  9844=>"101000000",
  9845=>"111000000",
  9846=>"001000000",
  9847=>"000000111",
  9848=>"100000000",
  9849=>"000000000",
  9850=>"010111111",
  9851=>"000000110",
  9852=>"110110100",
  9853=>"110111000",
  9854=>"000000111",
  9855=>"000000101",
  9856=>"000000000",
  9857=>"100100101",
  9858=>"000000000",
  9859=>"111000011",
  9860=>"000010000",
  9861=>"000000110",
  9862=>"111110000",
  9863=>"011110000",
  9864=>"000000000",
  9865=>"111000000",
  9866=>"000001111",
  9867=>"000000111",
  9868=>"000000100",
  9869=>"110110010",
  9870=>"000000101",
  9871=>"000000010",
  9872=>"000000111",
  9873=>"000000000",
  9874=>"000000111",
  9875=>"111111111",
  9876=>"000110000",
  9877=>"000000001",
  9878=>"100000000",
  9879=>"111111000",
  9880=>"000000111",
  9881=>"100000111",
  9882=>"001000000",
  9883=>"111111000",
  9884=>"000000000",
  9885=>"000000000",
  9886=>"111111111",
  9887=>"000000000",
  9888=>"111111000",
  9889=>"000000000",
  9890=>"000000000",
  9891=>"011111001",
  9892=>"000110111",
  9893=>"111111001",
  9894=>"111000000",
  9895=>"100110000",
  9896=>"110100111",
  9897=>"010000000",
  9898=>"111111011",
  9899=>"000000111",
  9900=>"000111111",
  9901=>"000111100",
  9902=>"000000101",
  9903=>"000110100",
  9904=>"110100110",
  9905=>"100100100",
  9906=>"111111111",
  9907=>"000000000",
  9908=>"111110110",
  9909=>"111000110",
  9910=>"110111111",
  9911=>"111111111",
  9912=>"100000000",
  9913=>"100111111",
  9914=>"000011111",
  9915=>"100110111",
  9916=>"000000000",
  9917=>"111011011",
  9918=>"111011111",
  9919=>"011111111",
  9920=>"000011000",
  9921=>"000000000",
  9922=>"000110111",
  9923=>"101101000",
  9924=>"100101010",
  9925=>"110111000",
  9926=>"010011111",
  9927=>"100110000",
  9928=>"111101110",
  9929=>"001000111",
  9930=>"000000000",
  9931=>"000100101",
  9932=>"000000000",
  9933=>"000000000",
  9934=>"000001111",
  9935=>"000000111",
  9936=>"110100000",
  9937=>"111111111",
  9938=>"000111111",
  9939=>"000000101",
  9940=>"001000000",
  9941=>"001111111",
  9942=>"000000111",
  9943=>"101100101",
  9944=>"111111110",
  9945=>"100000001",
  9946=>"000000111",
  9947=>"101000111",
  9948=>"111111011",
  9949=>"111110110",
  9950=>"011011011",
  9951=>"000000001",
  9952=>"000000000",
  9953=>"101000111",
  9954=>"000000000",
  9955=>"100100101",
  9956=>"000111111",
  9957=>"110111001",
  9958=>"000000111",
  9959=>"000100111",
  9960=>"111000111",
  9961=>"111111111",
  9962=>"111000111",
  9963=>"000000101",
  9964=>"000000011",
  9965=>"101101111",
  9966=>"010100011",
  9967=>"000010000",
  9968=>"111111011",
  9969=>"111000101",
  9970=>"111111001",
  9971=>"001101111",
  9972=>"111000000",
  9973=>"000100111",
  9974=>"000000011",
  9975=>"111100000",
  9976=>"111111110",
  9977=>"001001011",
  9978=>"110111100",
  9979=>"110000000",
  9980=>"111000111",
  9981=>"010010010",
  9982=>"000001011",
  9983=>"100000111",
  9984=>"100000000",
  9985=>"101000000",
  9986=>"000000000",
  9987=>"000000001",
  9988=>"100100000",
  9989=>"000110111",
  9990=>"111111000",
  9991=>"111110010",
  9992=>"011000000",
  9993=>"111111111",
  9994=>"110000000",
  9995=>"011111011",
  9996=>"000000110",
  9997=>"000011010",
  9998=>"110111000",
  9999=>"000011000",
  10000=>"000000001",
  10001=>"000000100",
  10002=>"101000000",
  10003=>"010010001",
  10004=>"111111011",
  10005=>"111000000",
  10006=>"111011000",
  10007=>"000000111",
  10008=>"111111100",
  10009=>"000000000",
  10010=>"001100000",
  10011=>"000000000",
  10012=>"111111000",
  10013=>"111101000",
  10014=>"000011111",
  10015=>"000100001",
  10016=>"111111011",
  10017=>"010000000",
  10018=>"001011111",
  10019=>"111111111",
  10020=>"111010000",
  10021=>"111111001",
  10022=>"000000000",
  10023=>"001000011",
  10024=>"000000000",
  10025=>"111111100",
  10026=>"111111000",
  10027=>"101000000",
  10028=>"111111001",
  10029=>"000110110",
  10030=>"111000000",
  10031=>"000000100",
  10032=>"111110000",
  10033=>"111000000",
  10034=>"001111110",
  10035=>"111010111",
  10036=>"000000111",
  10037=>"000001000",
  10038=>"111111111",
  10039=>"111000000",
  10040=>"111111000",
  10041=>"111111100",
  10042=>"000000111",
  10043=>"111111111",
  10044=>"001001100",
  10045=>"000000000",
  10046=>"010111000",
  10047=>"101001111",
  10048=>"101111011",
  10049=>"101101100",
  10050=>"111110110",
  10051=>"110000000",
  10052=>"111111000",
  10053=>"100100111",
  10054=>"000000000",
  10055=>"111100111",
  10056=>"110111111",
  10057=>"000000000",
  10058=>"000000001",
  10059=>"011011000",
  10060=>"000000000",
  10061=>"111001111",
  10062=>"111111001",
  10063=>"000000111",
  10064=>"001001001",
  10065=>"000000111",
  10066=>"111010000",
  10067=>"000000111",
  10068=>"000000000",
  10069=>"001011001",
  10070=>"111111011",
  10071=>"111111111",
  10072=>"111111000",
  10073=>"111011011",
  10074=>"000000001",
  10075=>"000000111",
  10076=>"101000000",
  10077=>"011111111",
  10078=>"100000000",
  10079=>"001001101",
  10080=>"000000000",
  10081=>"000000111",
  10082=>"111110110",
  10083=>"000000001",
  10084=>"111111000",
  10085=>"000000100",
  10086=>"000111111",
  10087=>"000100001",
  10088=>"110110000",
  10089=>"000111011",
  10090=>"010000100",
  10091=>"111111111",
  10092=>"110111110",
  10093=>"000000111",
  10094=>"011011111",
  10095=>"000000111",
  10096=>"011110111",
  10097=>"100111111",
  10098=>"000111111",
  10099=>"011111111",
  10100=>"000111111",
  10101=>"000000001",
  10102=>"000000111",
  10103=>"000111001",
  10104=>"111000001",
  10105=>"011111110",
  10106=>"111100111",
  10107=>"000000000",
  10108=>"111111000",
  10109=>"100000000",
  10110=>"111111111",
  10111=>"001001100",
  10112=>"111101011",
  10113=>"000111111",
  10114=>"000000111",
  10115=>"000000100",
  10116=>"111010011",
  10117=>"000000000",
  10118=>"111111000",
  10119=>"111010101",
  10120=>"100000111",
  10121=>"000111011",
  10122=>"000110111",
  10123=>"111111100",
  10124=>"111111111",
  10125=>"001111111",
  10126=>"000000111",
  10127=>"000000100",
  10128=>"111111000",
  10129=>"111110110",
  10130=>"111010110",
  10131=>"101100111",
  10132=>"000000000",
  10133=>"000011011",
  10134=>"000000000",
  10135=>"100110110",
  10136=>"000000000",
  10137=>"111111111",
  10138=>"010111000",
  10139=>"100111110",
  10140=>"111111001",
  10141=>"000000000",
  10142=>"000000000",
  10143=>"000000010",
  10144=>"000111111",
  10145=>"000100000",
  10146=>"000100101",
  10147=>"111101000",
  10148=>"100110111",
  10149=>"010000000",
  10150=>"000010110",
  10151=>"000000111",
  10152=>"111001000",
  10153=>"101111111",
  10154=>"100100001",
  10155=>"000000000",
  10156=>"000000000",
  10157=>"111111000",
  10158=>"111111111",
  10159=>"111111001",
  10160=>"111101111",
  10161=>"000111111",
  10162=>"000000111",
  10163=>"111101111",
  10164=>"000000000",
  10165=>"000000000",
  10166=>"111000001",
  10167=>"111111111",
  10168=>"000000110",
  10169=>"011111111",
  10170=>"000000100",
  10171=>"101101001",
  10172=>"011000000",
  10173=>"101000101",
  10174=>"111000000",
  10175=>"000100111",
  10176=>"111111000",
  10177=>"111111000",
  10178=>"111111110",
  10179=>"000000011",
  10180=>"111111100",
  10181=>"001000100",
  10182=>"000111111",
  10183=>"100001000",
  10184=>"101000111",
  10185=>"110010000",
  10186=>"101000100",
  10187=>"110100000",
  10188=>"101000000",
  10189=>"110000000",
  10190=>"000000000",
  10191=>"010011000",
  10192=>"000000000",
  10193=>"100100111",
  10194=>"000000000",
  10195=>"000011111",
  10196=>"001000000",
  10197=>"010111111",
  10198=>"100110111",
  10199=>"000111111",
  10200=>"000100100",
  10201=>"110111100",
  10202=>"111110000",
  10203=>"111111100",
  10204=>"001011110",
  10205=>"000100111",
  10206=>"001010000",
  10207=>"000000100",
  10208=>"000001000",
  10209=>"111000000",
  10210=>"111111111",
  10211=>"111000000",
  10212=>"000000001",
  10213=>"111111111",
  10214=>"000000100",
  10215=>"111111000",
  10216=>"011111100",
  10217=>"000000000",
  10218=>"111111000",
  10219=>"111111111",
  10220=>"000000000",
  10221=>"000111111",
  10222=>"000000000",
  10223=>"000011111",
  10224=>"000000111",
  10225=>"000111111",
  10226=>"111111111",
  10227=>"000000000",
  10228=>"111111000",
  10229=>"000000001",
  10230=>"111000000",
  10231=>"000001111",
  10232=>"110100000",
  10233=>"000100000",
  10234=>"011111111",
  10235=>"111100000",
  10236=>"011000000",
  10237=>"111111001",
  10238=>"001101111",
  10239=>"110111111",
  10240=>"000000001",
  10241=>"011000111",
  10242=>"000000101",
  10243=>"111111111",
  10244=>"000101111",
  10245=>"111111111",
  10246=>"111111111",
  10247=>"111111111",
  10248=>"000000000",
  10249=>"000000000",
  10250=>"110100111",
  10251=>"100100100",
  10252=>"001001111",
  10253=>"001001011",
  10254=>"000110110",
  10255=>"000000000",
  10256=>"100111000",
  10257=>"100000000",
  10258=>"100100100",
  10259=>"000111110",
  10260=>"001000000",
  10261=>"001011001",
  10262=>"000000000",
  10263=>"001001000",
  10264=>"111000000",
  10265=>"001001000",
  10266=>"000000110",
  10267=>"000000000",
  10268=>"000000000",
  10269=>"000000000",
  10270=>"110110110",
  10271=>"001000000",
  10272=>"011000000",
  10273=>"000000000",
  10274=>"111010011",
  10275=>"110111111",
  10276=>"011110110",
  10277=>"111101100",
  10278=>"110000000",
  10279=>"111111111",
  10280=>"000011110",
  10281=>"010111111",
  10282=>"001000000",
  10283=>"100000000",
  10284=>"000000000",
  10285=>"111111111",
  10286=>"111001000",
  10287=>"111111000",
  10288=>"011111111",
  10289=>"101100110",
  10290=>"000100110",
  10291=>"100111011",
  10292=>"111111111",
  10293=>"100000001",
  10294=>"100110110",
  10295=>"000000100",
  10296=>"001101001",
  10297=>"111111111",
  10298=>"110111111",
  10299=>"000000001",
  10300=>"111001001",
  10301=>"000000111",
  10302=>"111100100",
  10303=>"001111111",
  10304=>"000000000",
  10305=>"111001001",
  10306=>"011000111",
  10307=>"000110111",
  10308=>"011111111",
  10309=>"001000000",
  10310=>"111111000",
  10311=>"001001001",
  10312=>"111111111",
  10313=>"000000011",
  10314=>"000000001",
  10315=>"111111110",
  10316=>"011000001",
  10317=>"111111100",
  10318=>"000111111",
  10319=>"111111111",
  10320=>"000000000",
  10321=>"000011010",
  10322=>"000000001",
  10323=>"000000100",
  10324=>"100101111",
  10325=>"111111110",
  10326=>"000010111",
  10327=>"111111111",
  10328=>"111000000",
  10329=>"111001111",
  10330=>"110111111",
  10331=>"101111111",
  10332=>"111111111",
  10333=>"000011000",
  10334=>"000001011",
  10335=>"001000000",
  10336=>"000111111",
  10337=>"100111111",
  10338=>"000111111",
  10339=>"100100010",
  10340=>"100100000",
  10341=>"001000110",
  10342=>"011111111",
  10343=>"111111111",
  10344=>"101000000",
  10345=>"000000100",
  10346=>"000000000",
  10347=>"000000000",
  10348=>"000001011",
  10349=>"110111000",
  10350=>"111111010",
  10351=>"111111111",
  10352=>"000000110",
  10353=>"000100010",
  10354=>"000000001",
  10355=>"011111111",
  10356=>"001001000",
  10357=>"000100000",
  10358=>"001001111",
  10359=>"100100000",
  10360=>"011111111",
  10361=>"000000000",
  10362=>"111001001",
  10363=>"111111111",
  10364=>"100000100",
  10365=>"111101100",
  10366=>"000001111",
  10367=>"100000000",
  10368=>"000000000",
  10369=>"000111111",
  10370=>"000001111",
  10371=>"000000000",
  10372=>"000000000",
  10373=>"100100111",
  10374=>"000000000",
  10375=>"000000000",
  10376=>"001111111",
  10377=>"100100000",
  10378=>"111111111",
  10379=>"101000000",
  10380=>"000101000",
  10381=>"111000111",
  10382=>"000010111",
  10383=>"000000100",
  10384=>"000000000",
  10385=>"000000001",
  10386=>"000000000",
  10387=>"111111111",
  10388=>"111110110",
  10389=>"111111111",
  10390=>"111111001",
  10391=>"000000000",
  10392=>"011001001",
  10393=>"000000000",
  10394=>"000000000",
  10395=>"000000000",
  10396=>"011001001",
  10397=>"011110110",
  10398=>"000000000",
  10399=>"101110010",
  10400=>"000001011",
  10401=>"100000010",
  10402=>"000000000",
  10403=>"111000000",
  10404=>"101111111",
  10405=>"000100000",
  10406=>"111111111",
  10407=>"100110000",
  10408=>"111111111",
  10409=>"100000100",
  10410=>"000000000",
  10411=>"111001111",
  10412=>"000000111",
  10413=>"000000000",
  10414=>"001111111",
  10415=>"000010100",
  10416=>"110000000",
  10417=>"110110101",
  10418=>"100101101",
  10419=>"010111111",
  10420=>"000000000",
  10421=>"111101001",
  10422=>"000111111",
  10423=>"000000000",
  10424=>"000000000",
  10425=>"011000000",
  10426=>"100100110",
  10427=>"000000000",
  10428=>"001000000",
  10429=>"000000000",
  10430=>"000000000",
  10431=>"000000000",
  10432=>"000000000",
  10433=>"000100111",
  10434=>"001111111",
  10435=>"111110111",
  10436=>"000000111",
  10437=>"011110111",
  10438=>"000100110",
  10439=>"111111111",
  10440=>"111110100",
  10441=>"111111111",
  10442=>"000000011",
  10443=>"111111111",
  10444=>"101111110",
  10445=>"110111010",
  10446=>"000000000",
  10447=>"111110111",
  10448=>"111111111",
  10449=>"111010000",
  10450=>"110111110",
  10451=>"001001111",
  10452=>"000000011",
  10453=>"000000010",
  10454=>"000000111",
  10455=>"000000110",
  10456=>"000000000",
  10457=>"111111111",
  10458=>"000000001",
  10459=>"111111111",
  10460=>"111111111",
  10461=>"111111011",
  10462=>"001001011",
  10463=>"100110110",
  10464=>"000000100",
  10465=>"000000111",
  10466=>"000000111",
  10467=>"111111111",
  10468=>"000000000",
  10469=>"101101101",
  10470=>"101000001",
  10471=>"111111111",
  10472=>"000000100",
  10473=>"111101101",
  10474=>"000100100",
  10475=>"111111111",
  10476=>"000000000",
  10477=>"000000000",
  10478=>"011000111",
  10479=>"111000001",
  10480=>"110111000",
  10481=>"001001000",
  10482=>"000000000",
  10483=>"100100100",
  10484=>"111101000",
  10485=>"000000000",
  10486=>"000100111",
  10487=>"111111111",
  10488=>"000000000",
  10489=>"000000000",
  10490=>"101100111",
  10491=>"000100100",
  10492=>"110111110",
  10493=>"111111111",
  10494=>"000111001",
  10495=>"101111100",
  10496=>"011000011",
  10497=>"001001111",
  10498=>"111110000",
  10499=>"111111000",
  10500=>"100000000",
  10501=>"000011111",
  10502=>"111111111",
  10503=>"000000100",
  10504=>"001111111",
  10505=>"000000000",
  10506=>"110000000",
  10507=>"011000000",
  10508=>"000000100",
  10509=>"000000000",
  10510=>"111111011",
  10511=>"111111111",
  10512=>"111111000",
  10513=>"110110111",
  10514=>"011011111",
  10515=>"000000000",
  10516=>"111011000",
  10517=>"000010111",
  10518=>"011111111",
  10519=>"011011111",
  10520=>"100100000",
  10521=>"000000000",
  10522=>"011111111",
  10523=>"011111100",
  10524=>"001001000",
  10525=>"111110111",
  10526=>"111111111",
  10527=>"111001111",
  10528=>"111110111",
  10529=>"111111101",
  10530=>"001011011",
  10531=>"000000100",
  10532=>"111111000",
  10533=>"111111011",
  10534=>"101001000",
  10535=>"000000000",
  10536=>"011010010",
  10537=>"000000000",
  10538=>"111111111",
  10539=>"000000111",
  10540=>"000101111",
  10541=>"110111110",
  10542=>"000111111",
  10543=>"100110111",
  10544=>"000000000",
  10545=>"111111111",
  10546=>"000000001",
  10547=>"111000000",
  10548=>"011000000",
  10549=>"001001111",
  10550=>"111111011",
  10551=>"111011010",
  10552=>"000000000",
  10553=>"111101011",
  10554=>"111001001",
  10555=>"100100000",
  10556=>"011011011",
  10557=>"111110111",
  10558=>"111010000",
  10559=>"000110000",
  10560=>"000000110",
  10561=>"000100000",
  10562=>"111111111",
  10563=>"011111111",
  10564=>"010000000",
  10565=>"111110111",
  10566=>"111110110",
  10567=>"101100010",
  10568=>"011000001",
  10569=>"000000000",
  10570=>"000000000",
  10571=>"011001001",
  10572=>"110000000",
  10573=>"000000000",
  10574=>"000000000",
  10575=>"100000100",
  10576=>"101000000",
  10577=>"001111100",
  10578=>"000000011",
  10579=>"000000000",
  10580=>"000000100",
  10581=>"011001011",
  10582=>"000000000",
  10583=>"111111111",
  10584=>"111111111",
  10585=>"000001000",
  10586=>"110100100",
  10587=>"100110111",
  10588=>"011111100",
  10589=>"100111111",
  10590=>"000011010",
  10591=>"000000000",
  10592=>"001100000",
  10593=>"000010010",
  10594=>"011000000",
  10595=>"011001011",
  10596=>"001000000",
  10597=>"000000000",
  10598=>"111111000",
  10599=>"111111011",
  10600=>"000000000",
  10601=>"100000101",
  10602=>"011000100",
  10603=>"111111101",
  10604=>"110111111",
  10605=>"101100010",
  10606=>"011000110",
  10607=>"000000000",
  10608=>"000010011",
  10609=>"000000000",
  10610=>"111011000",
  10611=>"010110000",
  10612=>"000000000",
  10613=>"000000000",
  10614=>"111111111",
  10615=>"111111111",
  10616=>"000000000",
  10617=>"011111111",
  10618=>"001000011",
  10619=>"000010011",
  10620=>"000110111",
  10621=>"000001111",
  10622=>"011000000",
  10623=>"000000000",
  10624=>"110110110",
  10625=>"000010011",
  10626=>"000000000",
  10627=>"111011011",
  10628=>"000000000",
  10629=>"000100100",
  10630=>"100101001",
  10631=>"111111111",
  10632=>"111011111",
  10633=>"000101111",
  10634=>"000000000",
  10635=>"111111111",
  10636=>"001000000",
  10637=>"010111111",
  10638=>"010110000",
  10639=>"111111000",
  10640=>"000100111",
  10641=>"111111001",
  10642=>"000000000",
  10643=>"000110110",
  10644=>"111111111",
  10645=>"000000000",
  10646=>"000001101",
  10647=>"111111111",
  10648=>"000100111",
  10649=>"000000000",
  10650=>"011111111",
  10651=>"111111111",
  10652=>"111111111",
  10653=>"111111111",
  10654=>"000111100",
  10655=>"000000000",
  10656=>"000111001",
  10657=>"000000110",
  10658=>"000000010",
  10659=>"111111001",
  10660=>"001111111",
  10661=>"111111111",
  10662=>"000001000",
  10663=>"000000000",
  10664=>"000000000",
  10665=>"001111111",
  10666=>"001000001",
  10667=>"100111111",
  10668=>"000000000",
  10669=>"111111111",
  10670=>"110110000",
  10671=>"000000101",
  10672=>"000000000",
  10673=>"000000000",
  10674=>"000111011",
  10675=>"011011000",
  10676=>"011011001",
  10677=>"011100000",
  10678=>"000001100",
  10679=>"111111111",
  10680=>"110100110",
  10681=>"111111111",
  10682=>"011000000",
  10683=>"001001001",
  10684=>"001000000",
  10685=>"001100001",
  10686=>"001011001",
  10687=>"111110100",
  10688=>"111111111",
  10689=>"111011111",
  10690=>"111111111",
  10691=>"000000000",
  10692=>"001111111",
  10693=>"110000111",
  10694=>"000100000",
  10695=>"111111111",
  10696=>"100111111",
  10697=>"000000000",
  10698=>"000000111",
  10699=>"000000110",
  10700=>"111110111",
  10701=>"110100101",
  10702=>"110000000",
  10703=>"100111001",
  10704=>"111111111",
  10705=>"011001111",
  10706=>"110111110",
  10707=>"111100111",
  10708=>"110110110",
  10709=>"011000000",
  10710=>"000001011",
  10711=>"111000011",
  10712=>"000000000",
  10713=>"000110000",
  10714=>"101111111",
  10715=>"100111111",
  10716=>"111111001",
  10717=>"000000100",
  10718=>"110000000",
  10719=>"001000000",
  10720=>"110110110",
  10721=>"010010110",
  10722=>"011000100",
  10723=>"111111111",
  10724=>"111111111",
  10725=>"100111111",
  10726=>"001001001",
  10727=>"111111110",
  10728=>"000000000",
  10729=>"111111000",
  10730=>"011111111",
  10731=>"000100100",
  10732=>"000100110",
  10733=>"000000100",
  10734=>"111111111",
  10735=>"000100000",
  10736=>"111100100",
  10737=>"000000111",
  10738=>"111111111",
  10739=>"010111000",
  10740=>"111111111",
  10741=>"101000000",
  10742=>"000000100",
  10743=>"000110010",
  10744=>"100000000",
  10745=>"110110111",
  10746=>"000010001",
  10747=>"000000000",
  10748=>"111111011",
  10749=>"000000010",
  10750=>"000010000",
  10751=>"000000011",
  10752=>"000000111",
  10753=>"111111100",
  10754=>"101100111",
  10755=>"100000000",
  10756=>"111111111",
  10757=>"111100111",
  10758=>"111111111",
  10759=>"000000111",
  10760=>"111111000",
  10761=>"111110110",
  10762=>"111111111",
  10763=>"100100000",
  10764=>"111100100",
  10765=>"000000101",
  10766=>"011111111",
  10767=>"000000000",
  10768=>"111111000",
  10769=>"101000000",
  10770=>"110100100",
  10771=>"000000000",
  10772=>"111111111",
  10773=>"001111111",
  10774=>"000110111",
  10775=>"001011001",
  10776=>"111111011",
  10777=>"000000000",
  10778=>"001000000",
  10779=>"111000110",
  10780=>"111011011",
  10781=>"111001111",
  10782=>"000000000",
  10783=>"111010110",
  10784=>"000000000",
  10785=>"000000000",
  10786=>"100110000",
  10787=>"000001111",
  10788=>"000000000",
  10789=>"111111111",
  10790=>"000000000",
  10791=>"101111111",
  10792=>"011111111",
  10793=>"000000000",
  10794=>"111111111",
  10795=>"111000000",
  10796=>"111111111",
  10797=>"111111000",
  10798=>"111111111",
  10799=>"110010011",
  10800=>"011111000",
  10801=>"000000000",
  10802=>"000000000",
  10803=>"111111011",
  10804=>"000000000",
  10805=>"000000000",
  10806=>"000000000",
  10807=>"000111111",
  10808=>"000000000",
  10809=>"000111100",
  10810=>"111111111",
  10811=>"000000000",
  10812=>"111100111",
  10813=>"000000000",
  10814=>"101110110",
  10815=>"111111111",
  10816=>"000011011",
  10817=>"000000010",
  10818=>"111111111",
  10819=>"111111111",
  10820=>"000000001",
  10821=>"000000000",
  10822=>"111111111",
  10823=>"111011000",
  10824=>"010010011",
  10825=>"000000000",
  10826=>"110111111",
  10827=>"000000000",
  10828=>"100100111",
  10829=>"111101000",
  10830=>"000100111",
  10831=>"111111111",
  10832=>"000100101",
  10833=>"000000000",
  10834=>"111111111",
  10835=>"000000000",
  10836=>"111111111",
  10837=>"000000000",
  10838=>"100100101",
  10839=>"000000100",
  10840=>"011010000",
  10841=>"000000000",
  10842=>"000000100",
  10843=>"110110111",
  10844=>"111110111",
  10845=>"000010011",
  10846=>"000011010",
  10847=>"011011001",
  10848=>"001000000",
  10849=>"111101001",
  10850=>"000000000",
  10851=>"111111111",
  10852=>"000000000",
  10853=>"101000100",
  10854=>"100000011",
  10855=>"111111111",
  10856=>"011100000",
  10857=>"001101111",
  10858=>"011011111",
  10859=>"000001010",
  10860=>"011011111",
  10861=>"000000000",
  10862=>"100110111",
  10863=>"000110110",
  10864=>"000000001",
  10865=>"000001000",
  10866=>"000000000",
  10867=>"000100111",
  10868=>"111111111",
  10869=>"111100000",
  10870=>"111111000",
  10871=>"000000000",
  10872=>"100000000",
  10873=>"000101111",
  10874=>"000000011",
  10875=>"000000000",
  10876=>"100000110",
  10877=>"111111111",
  10878=>"011011000",
  10879=>"001000001",
  10880=>"000000001",
  10881=>"000000000",
  10882=>"110000000",
  10883=>"000000000",
  10884=>"000000000",
  10885=>"010110111",
  10886=>"000001000",
  10887=>"000000000",
  10888=>"000000111",
  10889=>"000100000",
  10890=>"000111010",
  10891=>"111000000",
  10892=>"000011001",
  10893=>"101010000",
  10894=>"110111111",
  10895=>"111111111",
  10896=>"110111111",
  10897=>"101000000",
  10898=>"001000001",
  10899=>"000000000",
  10900=>"111111111",
  10901=>"110111111",
  10902=>"000001111",
  10903=>"000000000",
  10904=>"111000000",
  10905=>"000000000",
  10906=>"111101000",
  10907=>"000000000",
  10908=>"101111111",
  10909=>"111110000",
  10910=>"111111111",
  10911=>"111111111",
  10912=>"000000000",
  10913=>"100000000",
  10914=>"111111111",
  10915=>"000000000",
  10916=>"111111111",
  10917=>"011011111",
  10918=>"101011111",
  10919=>"000000000",
  10920=>"000100110",
  10921=>"111111011",
  10922=>"000000000",
  10923=>"101111001",
  10924=>"000000001",
  10925=>"111110111",
  10926=>"111111110",
  10927=>"000000001",
  10928=>"000000000",
  10929=>"001000000",
  10930=>"000000110",
  10931=>"011111000",
  10932=>"111111001",
  10933=>"111111000",
  10934=>"000111101",
  10935=>"111000101",
  10936=>"110110111",
  10937=>"111111111",
  10938=>"001001011",
  10939=>"111111101",
  10940=>"000000000",
  10941=>"110111111",
  10942=>"000010111",
  10943=>"111111001",
  10944=>"110110111",
  10945=>"111111111",
  10946=>"111111111",
  10947=>"000000000",
  10948=>"000000000",
  10949=>"000000001",
  10950=>"000000010",
  10951=>"000000110",
  10952=>"011111111",
  10953=>"111111111",
  10954=>"001000100",
  10955=>"111111111",
  10956=>"000000000",
  10957=>"000000000",
  10958=>"000101101",
  10959=>"000100111",
  10960=>"111111110",
  10961=>"011001110",
  10962=>"100110100",
  10963=>"001000101",
  10964=>"111111101",
  10965=>"000001011",
  10966=>"000000111",
  10967=>"000000010",
  10968=>"011111111",
  10969=>"111111010",
  10970=>"010111111",
  10971=>"111111111",
  10972=>"000000000",
  10973=>"110110110",
  10974=>"001111010",
  10975=>"110111111",
  10976=>"111111111",
  10977=>"000000100",
  10978=>"111111110",
  10979=>"000011111",
  10980=>"101101100",
  10981=>"111000001",
  10982=>"000000000",
  10983=>"111111000",
  10984=>"111111110",
  10985=>"111100000",
  10986=>"111111011",
  10987=>"000000001",
  10988=>"000000100",
  10989=>"111111011",
  10990=>"000000000",
  10991=>"000100110",
  10992=>"000111111",
  10993=>"110000000",
  10994=>"000000001",
  10995=>"001000000",
  10996=>"111111111",
  10997=>"111111010",
  10998=>"000010111",
  10999=>"111111111",
  11000=>"111111101",
  11001=>"000000000",
  11002=>"000000101",
  11003=>"111111111",
  11004=>"100000101",
  11005=>"111111111",
  11006=>"001001000",
  11007=>"010010011",
  11008=>"011001001",
  11009=>"001001101",
  11010=>"000000000",
  11011=>"111111001",
  11012=>"000000111",
  11013=>"110111111",
  11014=>"111110100",
  11015=>"000000101",
  11016=>"111011011",
  11017=>"000000000",
  11018=>"000000000",
  11019=>"111111111",
  11020=>"000000000",
  11021=>"110000000",
  11022=>"011011011",
  11023=>"111111111",
  11024=>"111101101",
  11025=>"100000100",
  11026=>"111111111",
  11027=>"000000000",
  11028=>"000000111",
  11029=>"111000000",
  11030=>"100111111",
  11031=>"000000000",
  11032=>"101001001",
  11033=>"111011000",
  11034=>"111001101",
  11035=>"000000000",
  11036=>"000000000",
  11037=>"111000000",
  11038=>"000000000",
  11039=>"111011011",
  11040=>"000000100",
  11041=>"000000000",
  11042=>"111111000",
  11043=>"000000100",
  11044=>"011000001",
  11045=>"111111111",
  11046=>"111011111",
  11047=>"101101111",
  11048=>"000000000",
  11049=>"000000000",
  11050=>"111100111",
  11051=>"111111010",
  11052=>"000001001",
  11053=>"111000000",
  11054=>"111111111",
  11055=>"001000000",
  11056=>"000001111",
  11057=>"111111001",
  11058=>"111000000",
  11059=>"000010111",
  11060=>"111111111",
  11061=>"111001000",
  11062=>"110100000",
  11063=>"000011111",
  11064=>"000000000",
  11065=>"111001011",
  11066=>"111111111",
  11067=>"111111111",
  11068=>"111001001",
  11069=>"110111111",
  11070=>"001100110",
  11071=>"011111011",
  11072=>"000000000",
  11073=>"110111111",
  11074=>"111111111",
  11075=>"111111111",
  11076=>"000000110",
  11077=>"111000000",
  11078=>"111111111",
  11079=>"000000000",
  11080=>"000000000",
  11081=>"011111011",
  11082=>"111110111",
  11083=>"000000000",
  11084=>"000000000",
  11085=>"000000000",
  11086=>"000000000",
  11087=>"000010011",
  11088=>"000000100",
  11089=>"111111111",
  11090=>"111111011",
  11091=>"000000111",
  11092=>"011001000",
  11093=>"000000001",
  11094=>"100100110",
  11095=>"110100000",
  11096=>"111111111",
  11097=>"111111100",
  11098=>"111111111",
  11099=>"110100000",
  11100=>"100100010",
  11101=>"000000000",
  11102=>"000101101",
  11103=>"111000000",
  11104=>"111111011",
  11105=>"100000111",
  11106=>"000100000",
  11107=>"101101111",
  11108=>"000000000",
  11109=>"000000100",
  11110=>"101000111",
  11111=>"111011000",
  11112=>"000001011",
  11113=>"000001111",
  11114=>"000010110",
  11115=>"111111100",
  11116=>"000000000",
  11117=>"101111000",
  11118=>"111111111",
  11119=>"111111111",
  11120=>"111000000",
  11121=>"000000000",
  11122=>"100000111",
  11123=>"100111000",
  11124=>"000000100",
  11125=>"011011000",
  11126=>"011011100",
  11127=>"010000100",
  11128=>"000000000",
  11129=>"111101111",
  11130=>"111111111",
  11131=>"111111111",
  11132=>"111111111",
  11133=>"111111111",
  11134=>"000000000",
  11135=>"111111111",
  11136=>"000100111",
  11137=>"010000000",
  11138=>"000111111",
  11139=>"000011111",
  11140=>"110010000",
  11141=>"111111000",
  11142=>"111000000",
  11143=>"000000000",
  11144=>"000001101",
  11145=>"111111011",
  11146=>"000000101",
  11147=>"111000111",
  11148=>"000000000",
  11149=>"100100001",
  11150=>"111111111",
  11151=>"000000001",
  11152=>"000110110",
  11153=>"000001001",
  11154=>"100000100",
  11155=>"000000000",
  11156=>"111111111",
  11157=>"000110010",
  11158=>"111111111",
  11159=>"111111111",
  11160=>"000000111",
  11161=>"110100100",
  11162=>"111000000",
  11163=>"000000000",
  11164=>"000000101",
  11165=>"011000000",
  11166=>"000000000",
  11167=>"111111111",
  11168=>"000010111",
  11169=>"000110111",
  11170=>"000000111",
  11171=>"000011111",
  11172=>"000001111",
  11173=>"111111000",
  11174=>"111111111",
  11175=>"001000000",
  11176=>"110000000",
  11177=>"000000111",
  11178=>"111111110",
  11179=>"101000000",
  11180=>"000111111",
  11181=>"000000000",
  11182=>"001000011",
  11183=>"000011111",
  11184=>"111111111",
  11185=>"111111001",
  11186=>"000000000",
  11187=>"000000000",
  11188=>"000000001",
  11189=>"111111111",
  11190=>"000000111",
  11191=>"000000011",
  11192=>"111111111",
  11193=>"111111111",
  11194=>"111111111",
  11195=>"001001101",
  11196=>"000000000",
  11197=>"000000110",
  11198=>"101111110",
  11199=>"110111111",
  11200=>"110110111",
  11201=>"011000000",
  11202=>"011111111",
  11203=>"000000000",
  11204=>"110100000",
  11205=>"100100111",
  11206=>"110000111",
  11207=>"100000000",
  11208=>"011000000",
  11209=>"011111110",
  11210=>"000000111",
  11211=>"100000000",
  11212=>"111111000",
  11213=>"111000001",
  11214=>"000000110",
  11215=>"000000000",
  11216=>"100100000",
  11217=>"011111111",
  11218=>"111111111",
  11219=>"110110111",
  11220=>"000111111",
  11221=>"010000001",
  11222=>"011011001",
  11223=>"001001001",
  11224=>"111111111",
  11225=>"100100000",
  11226=>"000000110",
  11227=>"000000000",
  11228=>"111111111",
  11229=>"101000110",
  11230=>"111111111",
  11231=>"011111111",
  11232=>"000000000",
  11233=>"001000001",
  11234=>"111111111",
  11235=>"100111111",
  11236=>"110110111",
  11237=>"111111111",
  11238=>"100111111",
  11239=>"001111000",
  11240=>"111111111",
  11241=>"111111000",
  11242=>"011000110",
  11243=>"000000101",
  11244=>"000000000",
  11245=>"111111001",
  11246=>"000000000",
  11247=>"111111011",
  11248=>"111111011",
  11249=>"000000000",
  11250=>"111010011",
  11251=>"000000000",
  11252=>"111111111",
  11253=>"000000000",
  11254=>"111000000",
  11255=>"111100111",
  11256=>"000000000",
  11257=>"001111111",
  11258=>"001000000",
  11259=>"000000011",
  11260=>"110111000",
  11261=>"000000000",
  11262=>"000100111",
  11263=>"011011001",
  11264=>"000000000",
  11265=>"010000000",
  11266=>"111000000",
  11267=>"000000000",
  11268=>"001001111",
  11269=>"001000111",
  11270=>"111111110",
  11271=>"111111001",
  11272=>"000000111",
  11273=>"111111111",
  11274=>"111101100",
  11275=>"000111111",
  11276=>"011011011",
  11277=>"110000011",
  11278=>"011111011",
  11279=>"110111111",
  11280=>"110000000",
  11281=>"111000000",
  11282=>"100000000",
  11283=>"110111111",
  11284=>"000000000",
  11285=>"110100000",
  11286=>"000000000",
  11287=>"011111111",
  11288=>"101000001",
  11289=>"001001011",
  11290=>"111111001",
  11291=>"100101110",
  11292=>"111000000",
  11293=>"100000000",
  11294=>"101001110",
  11295=>"000111111",
  11296=>"100110000",
  11297=>"100110100",
  11298=>"001001001",
  11299=>"001011011",
  11300=>"111111111",
  11301=>"010000001",
  11302=>"000000000",
  11303=>"100111111",
  11304=>"001001000",
  11305=>"011111000",
  11306=>"111111111",
  11307=>"100000001",
  11308=>"000000111",
  11309=>"000100111",
  11310=>"111100111",
  11311=>"100111111",
  11312=>"110111010",
  11313=>"001001000",
  11314=>"011011011",
  11315=>"000000110",
  11316=>"000000000",
  11317=>"100100100",
  11318=>"000000000",
  11319=>"011000000",
  11320=>"000000101",
  11321=>"111111001",
  11322=>"111111111",
  11323=>"111111000",
  11324=>"100000000",
  11325=>"100110100",
  11326=>"111111111",
  11327=>"110000000",
  11328=>"111111111",
  11329=>"001011111",
  11330=>"111000000",
  11331=>"000000011",
  11332=>"001001101",
  11333=>"000000000",
  11334=>"111011000",
  11335=>"111111111",
  11336=>"011100111",
  11337=>"111111111",
  11338=>"000000101",
  11339=>"100111111",
  11340=>"001001111",
  11341=>"111101001",
  11342=>"100111111",
  11343=>"010111110",
  11344=>"101000011",
  11345=>"000000000",
  11346=>"111111000",
  11347=>"001000010",
  11348=>"111101101",
  11349=>"110010110",
  11350=>"101000000",
  11351=>"111000000",
  11352=>"000010010",
  11353=>"010100111",
  11354=>"110110110",
  11355=>"110011011",
  11356=>"001001001",
  11357=>"000000000",
  11358=>"000001111",
  11359=>"111111011",
  11360=>"111011100",
  11361=>"000111000",
  11362=>"001100110",
  11363=>"001111111",
  11364=>"000001101",
  11365=>"011000000",
  11366=>"000000000",
  11367=>"111100100",
  11368=>"010000010",
  11369=>"010111111",
  11370=>"000000100",
  11371=>"110111111",
  11372=>"000000000",
  11373=>"110110010",
  11374=>"111111111",
  11375=>"000000000",
  11376=>"000000111",
  11377=>"001000000",
  11378=>"000000011",
  11379=>"111111011",
  11380=>"111111111",
  11381=>"000000110",
  11382=>"111111110",
  11383=>"000101111",
  11384=>"000100101",
  11385=>"001111111",
  11386=>"111111111",
  11387=>"111111111",
  11388=>"000000110",
  11389=>"000000000",
  11390=>"111111010",
  11391=>"110100000",
  11392=>"001111111",
  11393=>"000000000",
  11394=>"000111111",
  11395=>"000000100",
  11396=>"111111111",
  11397=>"000000010",
  11398=>"000000001",
  11399=>"111111111",
  11400=>"000100110",
  11401=>"111111000",
  11402=>"111111111",
  11403=>"001101101",
  11404=>"111111011",
  11405=>"110111000",
  11406=>"111011000",
  11407=>"100000000",
  11408=>"000000000",
  11409=>"111001111",
  11410=>"111100000",
  11411=>"010111111",
  11412=>"001000011",
  11413=>"000110100",
  11414=>"111111111",
  11415=>"011111111",
  11416=>"111111010",
  11417=>"111111111",
  11418=>"100100101",
  11419=>"011011111",
  11420=>"000100100",
  11421=>"001101111",
  11422=>"111111011",
  11423=>"000000000",
  11424=>"110011011",
  11425=>"011110010",
  11426=>"000000111",
  11427=>"000000001",
  11428=>"001001011",
  11429=>"011010101",
  11430=>"000000000",
  11431=>"101001001",
  11432=>"000011000",
  11433=>"000000111",
  11434=>"000111111",
  11435=>"111111111",
  11436=>"010110111",
  11437=>"110111111",
  11438=>"000011011",
  11439=>"000000111",
  11440=>"111111111",
  11441=>"000101111",
  11442=>"000001000",
  11443=>"011000000",
  11444=>"110110110",
  11445=>"111111100",
  11446=>"000111011",
  11447=>"000000000",
  11448=>"000000100",
  11449=>"011111111",
  11450=>"001100101",
  11451=>"111111111",
  11452=>"111111110",
  11453=>"111110100",
  11454=>"001001111",
  11455=>"000000111",
  11456=>"000000000",
  11457=>"110000000",
  11458=>"111110000",
  11459=>"000000000",
  11460=>"001000000",
  11461=>"010011010",
  11462=>"000000000",
  11463=>"000111001",
  11464=>"111111111",
  11465=>"000000000",
  11466=>"110100111",
  11467=>"110110110",
  11468=>"010011111",
  11469=>"000000110",
  11470=>"000000111",
  11471=>"100011011",
  11472=>"111111111",
  11473=>"000001001",
  11474=>"000000111",
  11475=>"000000101",
  11476=>"111111101",
  11477=>"101000000",
  11478=>"000000000",
  11479=>"000000111",
  11480=>"011111011",
  11481=>"001001000",
  11482=>"001001000",
  11483=>"111111111",
  11484=>"000000000",
  11485=>"111111111",
  11486=>"000000000",
  11487=>"100111101",
  11488=>"111111111",
  11489=>"000000000",
  11490=>"000111111",
  11491=>"000111111",
  11492=>"101101101",
  11493=>"011010001",
  11494=>"111111000",
  11495=>"111111001",
  11496=>"011011101",
  11497=>"000100111",
  11498=>"111111111",
  11499=>"000000000",
  11500=>"000000010",
  11501=>"000011011",
  11502=>"000000000",
  11503=>"111011010",
  11504=>"010111111",
  11505=>"000011011",
  11506=>"011011111",
  11507=>"000110110",
  11508=>"110110111",
  11509=>"011011111",
  11510=>"111011111",
  11511=>"011010011",
  11512=>"000110111",
  11513=>"000000000",
  11514=>"011111000",
  11515=>"001001111",
  11516=>"100101111",
  11517=>"110111111",
  11518=>"000011011",
  11519=>"110100100",
  11520=>"000001111",
  11521=>"000011111",
  11522=>"111111010",
  11523=>"110101111",
  11524=>"111111111",
  11525=>"010010000",
  11526=>"111110110",
  11527=>"000101111",
  11528=>"111010001",
  11529=>"011001001",
  11530=>"110111110",
  11531=>"101000001",
  11532=>"000000010",
  11533=>"110111111",
  11534=>"000000010",
  11535=>"010011001",
  11536=>"001011001",
  11537=>"010010001",
  11538=>"111100111",
  11539=>"000001111",
  11540=>"001001001",
  11541=>"101000000",
  11542=>"100110110",
  11543=>"011001101",
  11544=>"001001000",
  11545=>"111001111",
  11546=>"111111111",
  11547=>"110000100",
  11548=>"110111110",
  11549=>"111000000",
  11550=>"101101101",
  11551=>"111011011",
  11552=>"100110110",
  11553=>"001000100",
  11554=>"000101111",
  11555=>"110100101",
  11556=>"011000000",
  11557=>"101111111",
  11558=>"100000000",
  11559=>"111111111",
  11560=>"111000000",
  11561=>"110111111",
  11562=>"111000000",
  11563=>"111111011",
  11564=>"011011001",
  11565=>"110110110",
  11566=>"000000000",
  11567=>"000010000",
  11568=>"111111000",
  11569=>"111111011",
  11570=>"001000000",
  11571=>"010110100",
  11572=>"000001011",
  11573=>"001000000",
  11574=>"000000011",
  11575=>"000000010",
  11576=>"000000000",
  11577=>"010010010",
  11578=>"100111001",
  11579=>"001001001",
  11580=>"100000000",
  11581=>"000000000",
  11582=>"111000000",
  11583=>"111110100",
  11584=>"111111000",
  11585=>"111111000",
  11586=>"000000001",
  11587=>"000110110",
  11588=>"011111000",
  11589=>"011010000",
  11590=>"000000100",
  11591=>"111111111",
  11592=>"000100110",
  11593=>"011011011",
  11594=>"011111111",
  11595=>"001011010",
  11596=>"110111110",
  11597=>"000000000",
  11598=>"111111010",
  11599=>"000000000",
  11600=>"010110010",
  11601=>"111111111",
  11602=>"111100110",
  11603=>"001101111",
  11604=>"111000000",
  11605=>"111111111",
  11606=>"110111111",
  11607=>"111111111",
  11608=>"000000000",
  11609=>"010000000",
  11610=>"101100111",
  11611=>"111111100",
  11612=>"100000010",
  11613=>"101000001",
  11614=>"011111110",
  11615=>"010000000",
  11616=>"011000111",
  11617=>"111000100",
  11618=>"011000001",
  11619=>"000000001",
  11620=>"011011111",
  11621=>"101000000",
  11622=>"010100000",
  11623=>"100000000",
  11624=>"110111111",
  11625=>"000011011",
  11626=>"011011011",
  11627=>"111011001",
  11628=>"001000000",
  11629=>"000000100",
  11630=>"110100110",
  11631=>"111111111",
  11632=>"000000000",
  11633=>"111111111",
  11634=>"000001111",
  11635=>"111100100",
  11636=>"000000000",
  11637=>"100100100",
  11638=>"110010011",
  11639=>"000000001",
  11640=>"000000000",
  11641=>"111111010",
  11642=>"000000110",
  11643=>"000110111",
  11644=>"011110010",
  11645=>"010001000",
  11646=>"000000011",
  11647=>"001000100",
  11648=>"010000000",
  11649=>"110010111",
  11650=>"100000000",
  11651=>"111111000",
  11652=>"000000111",
  11653=>"000000000",
  11654=>"000110110",
  11655=>"000001011",
  11656=>"000000000",
  11657=>"011011010",
  11658=>"001111111",
  11659=>"000111000",
  11660=>"111101111",
  11661=>"100110111",
  11662=>"111000000",
  11663=>"000001011",
  11664=>"011000000",
  11665=>"110111010",
  11666=>"000101111",
  11667=>"100100000",
  11668=>"000000111",
  11669=>"000111110",
  11670=>"001011111",
  11671=>"011011001",
  11672=>"100101111",
  11673=>"111111111",
  11674=>"000110111",
  11675=>"000110000",
  11676=>"000000000",
  11677=>"111011000",
  11678=>"000000100",
  11679=>"000000000",
  11680=>"000100111",
  11681=>"110001001",
  11682=>"011111111",
  11683=>"000011001",
  11684=>"000011011",
  11685=>"001000000",
  11686=>"000001111",
  11687=>"111101101",
  11688=>"011001001",
  11689=>"010000000",
  11690=>"010011011",
  11691=>"001111100",
  11692=>"000000000",
  11693=>"111111001",
  11694=>"000110111",
  11695=>"100011000",
  11696=>"001111111",
  11697=>"000000000",
  11698=>"000000000",
  11699=>"000010010",
  11700=>"111111111",
  11701=>"011000000",
  11702=>"011000110",
  11703=>"000001001",
  11704=>"000011111",
  11705=>"001111111",
  11706=>"111000000",
  11707=>"111100000",
  11708=>"000000000",
  11709=>"001001011",
  11710=>"111111111",
  11711=>"101001001",
  11712=>"100110111",
  11713=>"001000000",
  11714=>"000000000",
  11715=>"110111010",
  11716=>"000000110",
  11717=>"110110110",
  11718=>"101100100",
  11719=>"111000000",
  11720=>"100001001",
  11721=>"111000000",
  11722=>"011000000",
  11723=>"011010010",
  11724=>"111111000",
  11725=>"110111010",
  11726=>"000000000",
  11727=>"000110111",
  11728=>"101001111",
  11729=>"011111100",
  11730=>"010110100",
  11731=>"000000000",
  11732=>"000111111",
  11733=>"110100001",
  11734=>"111111101",
  11735=>"111101111",
  11736=>"000000000",
  11737=>"111111100",
  11738=>"001000000",
  11739=>"000100111",
  11740=>"011010000",
  11741=>"111111110",
  11742=>"000000000",
  11743=>"100101110",
  11744=>"111111110",
  11745=>"111110000",
  11746=>"000000000",
  11747=>"000000000",
  11748=>"000001000",
  11749=>"000000000",
  11750=>"111111011",
  11751=>"000000000",
  11752=>"111011011",
  11753=>"100110000",
  11754=>"000011011",
  11755=>"000000000",
  11756=>"011001000",
  11757=>"011011001",
  11758=>"000001001",
  11759=>"110111111",
  11760=>"000000111",
  11761=>"000000111",
  11762=>"101110111",
  11763=>"000000000",
  11764=>"000000000",
  11765=>"000000000",
  11766=>"000000111",
  11767=>"111110111",
  11768=>"000010000",
  11769=>"010011010",
  11770=>"111110000",
  11771=>"111111000",
  11772=>"101100000",
  11773=>"100111110",
  11774=>"000100111",
  11775=>"000000111",
  11776=>"000000000",
  11777=>"111000001",
  11778=>"111111111",
  11779=>"100000000",
  11780=>"111111111",
  11781=>"001111111",
  11782=>"011000000",
  11783=>"000000111",
  11784=>"011111010",
  11785=>"000111000",
  11786=>"000000000",
  11787=>"110000000",
  11788=>"110111000",
  11789=>"111111000",
  11790=>"111111011",
  11791=>"000000000",
  11792=>"000000000",
  11793=>"010111110",
  11794=>"000000000",
  11795=>"000111111",
  11796=>"000000010",
  11797=>"111111000",
  11798=>"111001000",
  11799=>"100100100",
  11800=>"111100100",
  11801=>"001000000",
  11802=>"111101100",
  11803=>"011000101",
  11804=>"000000000",
  11805=>"101000000",
  11806=>"000111111",
  11807=>"000000011",
  11808=>"000011100",
  11809=>"111100110",
  11810=>"000010110",
  11811=>"111000111",
  11812=>"010111111",
  11813=>"111111000",
  11814=>"000000100",
  11815=>"000000000",
  11816=>"111111111",
  11817=>"111111000",
  11818=>"111111000",
  11819=>"111000100",
  11820=>"111111111",
  11821=>"000111000",
  11822=>"001000001",
  11823=>"000000001",
  11824=>"000000000",
  11825=>"011111111",
  11826=>"000100110",
  11827=>"100000100",
  11828=>"000000000",
  11829=>"000111111",
  11830=>"000000100",
  11831=>"000000100",
  11832=>"111111111",
  11833=>"000000001",
  11834=>"011001111",
  11835=>"101000000",
  11836=>"000000000",
  11837=>"000000111",
  11838=>"001111100",
  11839=>"111111111",
  11840=>"000000001",
  11841=>"111101001",
  11842=>"111111111",
  11843=>"000000111",
  11844=>"000011001",
  11845=>"000000110",
  11846=>"111010000",
  11847=>"000001011",
  11848=>"000000111",
  11849=>"000000111",
  11850=>"111000001",
  11851=>"001010111",
  11852=>"110111111",
  11853=>"100111111",
  11854=>"101001000",
  11855=>"111111000",
  11856=>"011000000",
  11857=>"100000000",
  11858=>"000010000",
  11859=>"110110110",
  11860=>"000100000",
  11861=>"110110000",
  11862=>"000000111",
  11863=>"000111111",
  11864=>"000111111",
  11865=>"101100111",
  11866=>"101111101",
  11867=>"000000111",
  11868=>"111011000",
  11869=>"000000001",
  11870=>"000110111",
  11871=>"111110000",
  11872=>"111000000",
  11873=>"100110111",
  11874=>"001111001",
  11875=>"011000000",
  11876=>"010000111",
  11877=>"010010010",
  11878=>"100100110",
  11879=>"110110111",
  11880=>"000110010",
  11881=>"111111111",
  11882=>"111110111",
  11883=>"000000001",
  11884=>"111011000",
  11885=>"111000000",
  11886=>"000000000",
  11887=>"000000000",
  11888=>"100111110",
  11889=>"000111111",
  11890=>"001111111",
  11891=>"111111100",
  11892=>"000110100",
  11893=>"000110111",
  11894=>"100111111",
  11895=>"111111000",
  11896=>"000000000",
  11897=>"111111010",
  11898=>"000000101",
  11899=>"111000100",
  11900=>"110100010",
  11901=>"000000000",
  11902=>"101111001",
  11903=>"000101100",
  11904=>"111111111",
  11905=>"001111110",
  11906=>"000000000",
  11907=>"111100000",
  11908=>"111111111",
  11909=>"111000000",
  11910=>"000101111",
  11911=>"111111000",
  11912=>"000000100",
  11913=>"000000000",
  11914=>"111111001",
  11915=>"100000000",
  11916=>"111110000",
  11917=>"001111111",
  11918=>"000110111",
  11919=>"111110000",
  11920=>"000000110",
  11921=>"100000000",
  11922=>"010111000",
  11923=>"000000000",
  11924=>"000000000",
  11925=>"011110111",
  11926=>"000000000",
  11927=>"111111111",
  11928=>"000000001",
  11929=>"011000110",
  11930=>"111010000",
  11931=>"011111000",
  11932=>"000000111",
  11933=>"001000000",
  11934=>"000000111",
  11935=>"111111000",
  11936=>"111111111",
  11937=>"100010000",
  11938=>"111111011",
  11939=>"111111111",
  11940=>"110111111",
  11941=>"111011111",
  11942=>"100111111",
  11943=>"000001111",
  11944=>"000000000",
  11945=>"000000100",
  11946=>"000000000",
  11947=>"000000111",
  11948=>"110110000",
  11949=>"000101111",
  11950=>"000000000",
  11951=>"111001000",
  11952=>"011011000",
  11953=>"000110110",
  11954=>"111111010",
  11955=>"000111111",
  11956=>"100000100",
  11957=>"111111111",
  11958=>"010011100",
  11959=>"111111000",
  11960=>"001001111",
  11961=>"011101111",
  11962=>"000000001",
  11963=>"000011111",
  11964=>"000000111",
  11965=>"111111000",
  11966=>"000000000",
  11967=>"000110111",
  11968=>"000000000",
  11969=>"111100000",
  11970=>"000111111",
  11971=>"111111111",
  11972=>"111000000",
  11973=>"010011000",
  11974=>"111111111",
  11975=>"010111111",
  11976=>"111111111",
  11977=>"000000111",
  11978=>"111110111",
  11979=>"001001111",
  11980=>"000000001",
  11981=>"000000001",
  11982=>"000000001",
  11983=>"000000000",
  11984=>"000000111",
  11985=>"111111111",
  11986=>"000000000",
  11987=>"000010000",
  11988=>"100000010",
  11989=>"100110110",
  11990=>"000000000",
  11991=>"111111000",
  11992=>"111111111",
  11993=>"000000011",
  11994=>"000000000",
  11995=>"110111000",
  11996=>"000000011",
  11997=>"111000000",
  11998=>"010000000",
  11999=>"011111111",
  12000=>"111011000",
  12001=>"111101000",
  12002=>"000000100",
  12003=>"000111111",
  12004=>"111000000",
  12005=>"000001111",
  12006=>"001111111",
  12007=>"000111000",
  12008=>"000000001",
  12009=>"000000110",
  12010=>"111000000",
  12011=>"000111111",
  12012=>"000000010",
  12013=>"111000000",
  12014=>"110110111",
  12015=>"111000000",
  12016=>"111000000",
  12017=>"000000111",
  12018=>"000000111",
  12019=>"110111000",
  12020=>"000000000",
  12021=>"001101000",
  12022=>"000011011",
  12023=>"111111111",
  12024=>"010110111",
  12025=>"000111111",
  12026=>"111111111",
  12027=>"000111111",
  12028=>"111001000",
  12029=>"011011001",
  12030=>"111111011",
  12031=>"001000000",
  12032=>"001000001",
  12033=>"000101101",
  12034=>"000000111",
  12035=>"111111111",
  12036=>"111000000",
  12037=>"001001000",
  12038=>"000000111",
  12039=>"000101111",
  12040=>"001000000",
  12041=>"000111111",
  12042=>"111000111",
  12043=>"111111000",
  12044=>"111100111",
  12045=>"000000000",
  12046=>"111111100",
  12047=>"000000000",
  12048=>"000000111",
  12049=>"111111000",
  12050=>"111000000",
  12051=>"000000000",
  12052=>"111111000",
  12053=>"000000100",
  12054=>"011011000",
  12055=>"000100111",
  12056=>"011010111",
  12057=>"111000000",
  12058=>"110000111",
  12059=>"000000111",
  12060=>"001000000",
  12061=>"000000111",
  12062=>"000111111",
  12063=>"000000000",
  12064=>"000100111",
  12065=>"111111111",
  12066=>"000000000",
  12067=>"111111111",
  12068=>"110000111",
  12069=>"000000000",
  12070=>"111111000",
  12071=>"001111000",
  12072=>"000111111",
  12073=>"000000111",
  12074=>"111111011",
  12075=>"000101000",
  12076=>"000000111",
  12077=>"000011001",
  12078=>"000000000",
  12079=>"000000000",
  12080=>"111111000",
  12081=>"000000000",
  12082=>"000010000",
  12083=>"111000000",
  12084=>"000001111",
  12085=>"000100000",
  12086=>"000000001",
  12087=>"111000000",
  12088=>"001011111",
  12089=>"111000000",
  12090=>"000110111",
  12091=>"000000001",
  12092=>"000000111",
  12093=>"000000111",
  12094=>"100000000",
  12095=>"101000011",
  12096=>"000100111",
  12097=>"000000000",
  12098=>"000000000",
  12099=>"010111010",
  12100=>"111111111",
  12101=>"111000111",
  12102=>"000110111",
  12103=>"000000111",
  12104=>"000000111",
  12105=>"000000011",
  12106=>"011000111",
  12107=>"010110010",
  12108=>"000000000",
  12109=>"111111011",
  12110=>"111000011",
  12111=>"011001011",
  12112=>"000011111",
  12113=>"111011000",
  12114=>"000000111",
  12115=>"111111111",
  12116=>"110111011",
  12117=>"011111111",
  12118=>"000000000",
  12119=>"111010111",
  12120=>"000000000",
  12121=>"111000000",
  12122=>"000111111",
  12123=>"111111111",
  12124=>"111000000",
  12125=>"000110111",
  12126=>"000000000",
  12127=>"100100000",
  12128=>"111000000",
  12129=>"000111111",
  12130=>"000111011",
  12131=>"111000000",
  12132=>"111111111",
  12133=>"000001111",
  12134=>"000111010",
  12135=>"110111111",
  12136=>"000110111",
  12137=>"111000000",
  12138=>"000000000",
  12139=>"111001000",
  12140=>"000000010",
  12141=>"111111111",
  12142=>"111111110",
  12143=>"010111111",
  12144=>"000000111",
  12145=>"000111111",
  12146=>"000000111",
  12147=>"001001000",
  12148=>"000000001",
  12149=>"001111111",
  12150=>"000000000",
  12151=>"100100100",
  12152=>"000000000",
  12153=>"110111111",
  12154=>"001000100",
  12155=>"000111000",
  12156=>"000111111",
  12157=>"111111111",
  12158=>"000011111",
  12159=>"111111000",
  12160=>"110000000",
  12161=>"000111111",
  12162=>"000000011",
  12163=>"111000111",
  12164=>"100000000",
  12165=>"111111110",
  12166=>"000000110",
  12167=>"111000001",
  12168=>"100000000",
  12169=>"000000001",
  12170=>"011111010",
  12171=>"111100111",
  12172=>"111111111",
  12173=>"001001111",
  12174=>"000000000",
  12175=>"000000000",
  12176=>"000001000",
  12177=>"100110111",
  12178=>"001011101",
  12179=>"000000111",
  12180=>"111111111",
  12181=>"010111010",
  12182=>"101101000",
  12183=>"110111111",
  12184=>"111111111",
  12185=>"000000000",
  12186=>"001000111",
  12187=>"111111110",
  12188=>"000000111",
  12189=>"000010000",
  12190=>"000000000",
  12191=>"111101000",
  12192=>"000010111",
  12193=>"100100111",
  12194=>"000000000",
  12195=>"111111001",
  12196=>"111000000",
  12197=>"111110000",
  12198=>"100000000",
  12199=>"100000011",
  12200=>"111001000",
  12201=>"000000111",
  12202=>"111000111",
  12203=>"000000000",
  12204=>"010110000",
  12205=>"000000110",
  12206=>"001000000",
  12207=>"111111101",
  12208=>"000000000",
  12209=>"000000110",
  12210=>"111111000",
  12211=>"000000000",
  12212=>"101000000",
  12213=>"000000111",
  12214=>"111000100",
  12215=>"111111000",
  12216=>"000100111",
  12217=>"100000111",
  12218=>"000111111",
  12219=>"111100100",
  12220=>"111001000",
  12221=>"000000000",
  12222=>"000001001",
  12223=>"100110111",
  12224=>"111111111",
  12225=>"110010000",
  12226=>"000110000",
  12227=>"111111000",
  12228=>"000011111",
  12229=>"111111001",
  12230=>"000001111",
  12231=>"000111111",
  12232=>"000011001",
  12233=>"000111111",
  12234=>"000000000",
  12235=>"000000110",
  12236=>"111111011",
  12237=>"000111111",
  12238=>"000000000",
  12239=>"111111000",
  12240=>"000000000",
  12241=>"000001001",
  12242=>"000110000",
  12243=>"111100111",
  12244=>"011001011",
  12245=>"101100100",
  12246=>"010111111",
  12247=>"000010011",
  12248=>"111011000",
  12249=>"000010110",
  12250=>"000000100",
  12251=>"111000000",
  12252=>"000000000",
  12253=>"001000000",
  12254=>"000000000",
  12255=>"110110111",
  12256=>"111111010",
  12257=>"111111111",
  12258=>"000000000",
  12259=>"000000111",
  12260=>"100000011",
  12261=>"011101111",
  12262=>"111001000",
  12263=>"000111111",
  12264=>"111111000",
  12265=>"111111000",
  12266=>"111000000",
  12267=>"000011111",
  12268=>"000000000",
  12269=>"000110111",
  12270=>"000000001",
  12271=>"000111111",
  12272=>"000111111",
  12273=>"001111111",
  12274=>"111111111",
  12275=>"001000010",
  12276=>"111111111",
  12277=>"000000001",
  12278=>"110111111",
  12279=>"001001000",
  12280=>"000000111",
  12281=>"000000111",
  12282=>"000001000",
  12283=>"000111000",
  12284=>"000000000",
  12285=>"000111111",
  12286=>"111000000",
  12287=>"110000000",
  12288=>"100000000",
  12289=>"000000000",
  12290=>"100000000",
  12291=>"111111111",
  12292=>"111111111",
  12293=>"100000100",
  12294=>"000000000",
  12295=>"001000000",
  12296=>"000000000",
  12297=>"111100000",
  12298=>"111111111",
  12299=>"011111111",
  12300=>"110110110",
  12301=>"000000000",
  12302=>"100100100",
  12303=>"001001000",
  12304=>"111111111",
  12305=>"011111111",
  12306=>"000000000",
  12307=>"111111111",
  12308=>"111100111",
  12309=>"000100000",
  12310=>"111001011",
  12311=>"011011011",
  12312=>"000000101",
  12313=>"101000000",
  12314=>"001001000",
  12315=>"111100100",
  12316=>"100000000",
  12317=>"111111111",
  12318=>"111110111",
  12319=>"001000110",
  12320=>"111000001",
  12321=>"110110110",
  12322=>"000000000",
  12323=>"111111011",
  12324=>"000000000",
  12325=>"000000000",
  12326=>"111111111",
  12327=>"011111111",
  12328=>"100100111",
  12329=>"110110011",
  12330=>"000000111",
  12331=>"000111111",
  12332=>"001101100",
  12333=>"111101000",
  12334=>"110110111",
  12335=>"101100100",
  12336=>"100111111",
  12337=>"011001000",
  12338=>"110110000",
  12339=>"110111111",
  12340=>"000000000",
  12341=>"111001110",
  12342=>"100000111",
  12343=>"001001001",
  12344=>"001001001",
  12345=>"011010000",
  12346=>"111111111",
  12347=>"000000000",
  12348=>"101100100",
  12349=>"111110111",
  12350=>"111111000",
  12351=>"000000000",
  12352=>"011011100",
  12353=>"001000000",
  12354=>"001111111",
  12355=>"110110111",
  12356=>"111111111",
  12357=>"000000001",
  12358=>"111111011",
  12359=>"100100000",
  12360=>"111111111",
  12361=>"110111000",
  12362=>"110110110",
  12363=>"111111111",
  12364=>"111110010",
  12365=>"011111110",
  12366=>"010010111",
  12367=>"100111111",
  12368=>"111000000",
  12369=>"111110000",
  12370=>"001001000",
  12371=>"000000110",
  12372=>"100100110",
  12373=>"000000000",
  12374=>"011011001",
  12375=>"110011011",
  12376=>"011100110",
  12377=>"000000000",
  12378=>"001100000",
  12379=>"011001111",
  12380=>"100100111",
  12381=>"111000001",
  12382=>"001111111",
  12383=>"001001001",
  12384=>"111101100",
  12385=>"000000000",
  12386=>"001101111",
  12387=>"000000000",
  12388=>"011010000",
  12389=>"111011011",
  12390=>"001111111",
  12391=>"011011111",
  12392=>"101111110",
  12393=>"111111111",
  12394=>"111111011",
  12395=>"000010010",
  12396=>"011011011",
  12397=>"111110110",
  12398=>"111101101",
  12399=>"111111111",
  12400=>"000000000",
  12401=>"010000000",
  12402=>"011011011",
  12403=>"111111011",
  12404=>"000000000",
  12405=>"111000000",
  12406=>"111111111",
  12407=>"000000000",
  12408=>"000100100",
  12409=>"010000100",
  12410=>"000000000",
  12411=>"000000000",
  12412=>"100100100",
  12413=>"101001111",
  12414=>"000000000",
  12415=>"101000000",
  12416=>"000000001",
  12417=>"000001011",
  12418=>"000000101",
  12419=>"111101111",
  12420=>"100100100",
  12421=>"000000000",
  12422=>"000000001",
  12423=>"111110100",
  12424=>"000100010",
  12425=>"111011111",
  12426=>"111111000",
  12427=>"000000000",
  12428=>"111111111",
  12429=>"000000000",
  12430=>"100000111",
  12431=>"000000000",
  12432=>"001101111",
  12433=>"100001011",
  12434=>"000000111",
  12435=>"000001101",
  12436=>"000000000",
  12437=>"111111111",
  12438=>"000000000",
  12439=>"000000000",
  12440=>"111111111",
  12441=>"100111111",
  12442=>"000000000",
  12443=>"101101101",
  12444=>"111001001",
  12445=>"000001011",
  12446=>"110000000",
  12447=>"000000100",
  12448=>"011111000",
  12449=>"000111111",
  12450=>"001101101",
  12451=>"000000000",
  12452=>"000001001",
  12453=>"010111111",
  12454=>"000000000",
  12455=>"000000100",
  12456=>"111111111",
  12457=>"000000100",
  12458=>"000000000",
  12459=>"000000000",
  12460=>"001111011",
  12461=>"101100100",
  12462=>"000000000",
  12463=>"001000000",
  12464=>"100110111",
  12465=>"100101101",
  12466=>"110111110",
  12467=>"001110110",
  12468=>"011110111",
  12469=>"000000000",
  12470=>"000111111",
  12471=>"001000000",
  12472=>"000000100",
  12473=>"000101111",
  12474=>"000000000",
  12475=>"100010110",
  12476=>"100000000",
  12477=>"100010000",
  12478=>"100000111",
  12479=>"111011111",
  12480=>"000000000",
  12481=>"111011001",
  12482=>"111111011",
  12483=>"000000010",
  12484=>"011111111",
  12485=>"100010111",
  12486=>"000000000",
  12487=>"101111111",
  12488=>"111111111",
  12489=>"100001011",
  12490=>"001101101",
  12491=>"011011000",
  12492=>"000000000",
  12493=>"111111111",
  12494=>"111111111",
  12495=>"111111111",
  12496=>"111111111",
  12497=>"111100100",
  12498=>"111110110",
  12499=>"110100101",
  12500=>"001101101",
  12501=>"111110000",
  12502=>"000001111",
  12503=>"011001001",
  12504=>"000000000",
  12505=>"111111110",
  12506=>"000000000",
  12507=>"000000000",
  12508=>"000000000",
  12509=>"100100111",
  12510=>"111111111",
  12511=>"000000110",
  12512=>"110100000",
  12513=>"000001001",
  12514=>"111111110",
  12515=>"000000000",
  12516=>"111001111",
  12517=>"000100100",
  12518=>"111111001",
  12519=>"101001000",
  12520=>"100111111",
  12521=>"000000000",
  12522=>"000000000",
  12523=>"000000000",
  12524=>"111000100",
  12525=>"001001001",
  12526=>"110110110",
  12527=>"111110100",
  12528=>"111000000",
  12529=>"000000000",
  12530=>"110010010",
  12531=>"111011000",
  12532=>"000000000",
  12533=>"000110110",
  12534=>"000100000",
  12535=>"110111111",
  12536=>"100000000",
  12537=>"000000110",
  12538=>"000100100",
  12539=>"111111101",
  12540=>"110110111",
  12541=>"110110110",
  12542=>"011111010",
  12543=>"111111101",
  12544=>"100000000",
  12545=>"101101101",
  12546=>"111001100",
  12547=>"000000000",
  12548=>"000000000",
  12549=>"000000110",
  12550=>"011011100",
  12551=>"010011001",
  12552=>"001011011",
  12553=>"000000000",
  12554=>"110111111",
  12555=>"001000110",
  12556=>"100000000",
  12557=>"000001011",
  12558=>"111011000",
  12559=>"001111000",
  12560=>"111110111",
  12561=>"111011111",
  12562=>"000000010",
  12563=>"000000000",
  12564=>"000000101",
  12565=>"111110111",
  12566=>"111111111",
  12567=>"110100100",
  12568=>"111111111",
  12569=>"000000000",
  12570=>"001001111",
  12571=>"000110111",
  12572=>"100100100",
  12573=>"001000011",
  12574=>"111101000",
  12575=>"000000111",
  12576=>"011001011",
  12577=>"000111111",
  12578=>"001011011",
  12579=>"011011101",
  12580=>"101100111",
  12581=>"111011111",
  12582=>"000000000",
  12583=>"111001111",
  12584=>"100011111",
  12585=>"111111111",
  12586=>"011000111",
  12587=>"000000000",
  12588=>"111111111",
  12589=>"111111110",
  12590=>"100100111",
  12591=>"111110100",
  12592=>"111111110",
  12593=>"100001001",
  12594=>"000000000",
  12595=>"111111111",
  12596=>"111111110",
  12597=>"000010000",
  12598=>"000010100",
  12599=>"100000000",
  12600=>"000000000",
  12601=>"000000000",
  12602=>"000100111",
  12603=>"001000000",
  12604=>"000000000",
  12605=>"000100011",
  12606=>"111111011",
  12607=>"111110000",
  12608=>"000000000",
  12609=>"001001001",
  12610=>"001011111",
  12611=>"110000111",
  12612=>"111111100",
  12613=>"111111111",
  12614=>"111100011",
  12615=>"000000000",
  12616=>"100111111",
  12617=>"001000101",
  12618=>"001000001",
  12619=>"100100110",
  12620=>"111100111",
  12621=>"111111111",
  12622=>"110111110",
  12623=>"100111111",
  12624=>"000000000",
  12625=>"000000110",
  12626=>"111000001",
  12627=>"111001001",
  12628=>"100111111",
  12629=>"001011011",
  12630=>"011011010",
  12631=>"001110100",
  12632=>"000000001",
  12633=>"000101111",
  12634=>"111000000",
  12635=>"000000000",
  12636=>"111111111",
  12637=>"111111111",
  12638=>"110000111",
  12639=>"111011001",
  12640=>"001011011",
  12641=>"000000000",
  12642=>"100100100",
  12643=>"000000111",
  12644=>"000000000",
  12645=>"100100000",
  12646=>"111110111",
  12647=>"100100111",
  12648=>"101100101",
  12649=>"100000110",
  12650=>"000000001",
  12651=>"000100010",
  12652=>"000000111",
  12653=>"100100000",
  12654=>"000000000",
  12655=>"111101000",
  12656=>"000000110",
  12657=>"000000000",
  12658=>"101100100",
  12659=>"110111000",
  12660=>"011111011",
  12661=>"111110100",
  12662=>"111111111",
  12663=>"101111111",
  12664=>"011000000",
  12665=>"111111110",
  12666=>"001001111",
  12667=>"000010110",
  12668=>"101001001",
  12669=>"000000101",
  12670=>"000100000",
  12671=>"000000100",
  12672=>"000001111",
  12673=>"000111111",
  12674=>"110110110",
  12675=>"111111011",
  12676=>"001101101",
  12677=>"010010010",
  12678=>"011111111",
  12679=>"000000111",
  12680=>"111111111",
  12681=>"000000000",
  12682=>"110111111",
  12683=>"110111111",
  12684=>"111101111",
  12685=>"100100100",
  12686=>"100000000",
  12687=>"111111111",
  12688=>"001000001",
  12689=>"001000001",
  12690=>"111100101",
  12691=>"100100100",
  12692=>"000100000",
  12693=>"011011011",
  12694=>"001000001",
  12695=>"110111111",
  12696=>"000001001",
  12697=>"011101000",
  12698=>"000000000",
  12699=>"010011111",
  12700=>"001111001",
  12701=>"110111110",
  12702=>"000000011",
  12703=>"000100100",
  12704=>"011111111",
  12705=>"011001001",
  12706=>"000000111",
  12707=>"011011000",
  12708=>"000001001",
  12709=>"000010010",
  12710=>"111110100",
  12711=>"000000000",
  12712=>"000000000",
  12713=>"000001011",
  12714=>"111111111",
  12715=>"000000000",
  12716=>"000000111",
  12717=>"000011011",
  12718=>"001000100",
  12719=>"000000000",
  12720=>"011110000",
  12721=>"000000001",
  12722=>"011000000",
  12723=>"111001000",
  12724=>"101000000",
  12725=>"111000100",
  12726=>"100000100",
  12727=>"110111111",
  12728=>"111111110",
  12729=>"110111111",
  12730=>"111111100",
  12731=>"100100001",
  12732=>"001000000",
  12733=>"111111111",
  12734=>"100000000",
  12735=>"101100100",
  12736=>"011011000",
  12737=>"101100111",
  12738=>"000000000",
  12739=>"101001000",
  12740=>"111011111",
  12741=>"000100111",
  12742=>"100000000",
  12743=>"000000111",
  12744=>"100000000",
  12745=>"110111111",
  12746=>"100000001",
  12747=>"100000110",
  12748=>"000010000",
  12749=>"111111111",
  12750=>"000000000",
  12751=>"011111111",
  12752=>"000000100",
  12753=>"111111111",
  12754=>"111001000",
  12755=>"111011011",
  12756=>"111101100",
  12757=>"111000100",
  12758=>"111111111",
  12759=>"111111000",
  12760=>"100100101",
  12761=>"010110111",
  12762=>"100000111",
  12763=>"001000100",
  12764=>"000111001",
  12765=>"000111011",
  12766=>"111111110",
  12767=>"101111111",
  12768=>"110111111",
  12769=>"111000111",
  12770=>"000000010",
  12771=>"100101111",
  12772=>"000000111",
  12773=>"001000001",
  12774=>"111110010",
  12775=>"011011111",
  12776=>"100100001",
  12777=>"000110111",
  12778=>"111110111",
  12779=>"111111111",
  12780=>"110110111",
  12781=>"000010000",
  12782=>"000000000",
  12783=>"111111111",
  12784=>"000000000",
  12785=>"100101000",
  12786=>"010011111",
  12787=>"100000100",
  12788=>"000000000",
  12789=>"111111011",
  12790=>"110111111",
  12791=>"110111100",
  12792=>"011011011",
  12793=>"000000000",
  12794=>"110111111",
  12795=>"010000000",
  12796=>"000010000",
  12797=>"011111111",
  12798=>"000000000",
  12799=>"111111110",
  12800=>"100001001",
  12801=>"111000000",
  12802=>"000000111",
  12803=>"001001010",
  12804=>"011000000",
  12805=>"000000100",
  12806=>"000000000",
  12807=>"000110111",
  12808=>"111111010",
  12809=>"001000111",
  12810=>"001000100",
  12811=>"111111011",
  12812=>"110111100",
  12813=>"111000000",
  12814=>"001001101",
  12815=>"000000000",
  12816=>"110111110",
  12817=>"000000101",
  12818=>"001001111",
  12819=>"110111111",
  12820=>"101011111",
  12821=>"111111111",
  12822=>"111110010",
  12823=>"110110010",
  12824=>"100100110",
  12825=>"011111111",
  12826=>"001000001",
  12827=>"011011000",
  12828=>"111111101",
  12829=>"000000000",
  12830=>"111100100",
  12831=>"111111000",
  12832=>"010111111",
  12833=>"001001000",
  12834=>"110110110",
  12835=>"111110000",
  12836=>"001000000",
  12837=>"000001010",
  12838=>"000000000",
  12839=>"111111000",
  12840=>"000110000",
  12841=>"000000000",
  12842=>"000000111",
  12843=>"000000111",
  12844=>"110110110",
  12845=>"000100000",
  12846=>"011011000",
  12847=>"100110011",
  12848=>"001101111",
  12849=>"111111001",
  12850=>"101001000",
  12851=>"010000000",
  12852=>"001001000",
  12853=>"011011111",
  12854=>"011011000",
  12855=>"000100111",
  12856=>"100000000",
  12857=>"010110110",
  12858=>"000000000",
  12859=>"001000111",
  12860=>"111111011",
  12861=>"111110110",
  12862=>"100011110",
  12863=>"000000000",
  12864=>"010111111",
  12865=>"110111011",
  12866=>"110110111",
  12867=>"011111010",
  12868=>"000000000",
  12869=>"101101000",
  12870=>"000000000",
  12871=>"111111000",
  12872=>"011111101",
  12873=>"001000111",
  12874=>"000010000",
  12875=>"011001000",
  12876=>"111110010",
  12877=>"000010000",
  12878=>"000000111",
  12879=>"101110111",
  12880=>"110100000",
  12881=>"111110000",
  12882=>"000000111",
  12883=>"100111111",
  12884=>"000000000",
  12885=>"010011001",
  12886=>"111011011",
  12887=>"000000000",
  12888=>"000000010",
  12889=>"101101111",
  12890=>"111000011",
  12891=>"110110110",
  12892=>"101101111",
  12893=>"111111011",
  12894=>"000111111",
  12895=>"110111010",
  12896=>"011000000",
  12897=>"000110111",
  12898=>"111011111",
  12899=>"110000000",
  12900=>"111011000",
  12901=>"000010111",
  12902=>"111110111",
  12903=>"111111111",
  12904=>"011001101",
  12905=>"011111111",
  12906=>"111111111",
  12907=>"011011000",
  12908=>"000000000",
  12909=>"101000100",
  12910=>"111001001",
  12911=>"111000000",
  12912=>"110000001",
  12913=>"111111011",
  12914=>"011000001",
  12915=>"111111111",
  12916=>"111110100",
  12917=>"110000000",
  12918=>"000000000",
  12919=>"011110000",
  12920=>"011000000",
  12921=>"000000000",
  12922=>"111111100",
  12923=>"000001111",
  12924=>"111110110",
  12925=>"011011111",
  12926=>"111000000",
  12927=>"000000000",
  12928=>"110111110",
  12929=>"000000000",
  12930=>"000010111",
  12931=>"000011101",
  12932=>"001001101",
  12933=>"000101111",
  12934=>"110110000",
  12935=>"000000000",
  12936=>"100000111",
  12937=>"101000111",
  12938=>"100100000",
  12939=>"110110111",
  12940=>"010110011",
  12941=>"000010010",
  12942=>"110110111",
  12943=>"110110111",
  12944=>"111100111",
  12945=>"011011000",
  12946=>"111110010",
  12947=>"000000000",
  12948=>"000011000",
  12949=>"000100000",
  12950=>"111001000",
  12951=>"100000100",
  12952=>"000000000",
  12953=>"111111111",
  12954=>"001000000",
  12955=>"011110000",
  12956=>"000000000",
  12957=>"111110000",
  12958=>"000000000",
  12959=>"111011010",
  12960=>"101101111",
  12961=>"100111111",
  12962=>"000000000",
  12963=>"111111111",
  12964=>"000000000",
  12965=>"000000000",
  12966=>"111000000",
  12967=>"110110110",
  12968=>"000000000",
  12969=>"111111111",
  12970=>"001111111",
  12971=>"110111111",
  12972=>"011011010",
  12973=>"111111000",
  12974=>"111110111",
  12975=>"111111111",
  12976=>"000000000",
  12977=>"101011011",
  12978=>"111111011",
  12979=>"101000001",
  12980=>"111111111",
  12981=>"110111111",
  12982=>"011111010",
  12983=>"110111011",
  12984=>"110000000",
  12985=>"000000101",
  12986=>"000000000",
  12987=>"010110111",
  12988=>"001101111",
  12989=>"000000000",
  12990=>"000000000",
  12991=>"111111111",
  12992=>"110100000",
  12993=>"001000000",
  12994=>"000011111",
  12995=>"010110010",
  12996=>"111110111",
  12997=>"000110111",
  12998=>"000111111",
  12999=>"000000001",
  13000=>"111111111",
  13001=>"001000000",
  13002=>"000000001",
  13003=>"001000000",
  13004=>"111000000",
  13005=>"111111111",
  13006=>"111111111",
  13007=>"011111111",
  13008=>"000011111",
  13009=>"111110010",
  13010=>"110110111",
  13011=>"000000111",
  13012=>"111110110",
  13013=>"000000011",
  13014=>"101000000",
  13015=>"111111000",
  13016=>"000000000",
  13017=>"111111111",
  13018=>"100000110",
  13019=>"000000110",
  13020=>"101101111",
  13021=>"000000000",
  13022=>"000000000",
  13023=>"000000111",
  13024=>"000100110",
  13025=>"111111011",
  13026=>"111111100",
  13027=>"000000001",
  13028=>"000000000",
  13029=>"011011011",
  13030=>"111111110",
  13031=>"000000000",
  13032=>"111111111",
  13033=>"000000001",
  13034=>"000000000",
  13035=>"110000110",
  13036=>"111000000",
  13037=>"000000000",
  13038=>"111111111",
  13039=>"000100111",
  13040=>"111111111",
  13041=>"000111111",
  13042=>"001001101",
  13043=>"000000000",
  13044=>"000000000",
  13045=>"101111111",
  13046=>"100000000",
  13047=>"101101011",
  13048=>"110000000",
  13049=>"001100000",
  13050=>"000000000",
  13051=>"001100000",
  13052=>"010011000",
  13053=>"110100111",
  13054=>"011010000",
  13055=>"111111111",
  13056=>"010000000",
  13057=>"111111111",
  13058=>"100101000",
  13059=>"000000011",
  13060=>"111000000",
  13061=>"100000000",
  13062=>"110111100",
  13063=>"110000011",
  13064=>"111001111",
  13065=>"111111111",
  13066=>"110111010",
  13067=>"110000000",
  13068=>"010100000",
  13069=>"101000000",
  13070=>"100111011",
  13071=>"111111110",
  13072=>"000000000",
  13073=>"110010011",
  13074=>"000010111",
  13075=>"111001111",
  13076=>"110010111",
  13077=>"100110111",
  13078=>"001101111",
  13079=>"000010010",
  13080=>"100001011",
  13081=>"000111111",
  13082=>"111111111",
  13083=>"110110110",
  13084=>"111111110",
  13085=>"111110000",
  13086=>"010111110",
  13087=>"000100000",
  13088=>"010011011",
  13089=>"000111111",
  13090=>"000000000",
  13091=>"000000000",
  13092=>"000000011",
  13093=>"000000000",
  13094=>"000110110",
  13095=>"110110111",
  13096=>"110111001",
  13097=>"000000010",
  13098=>"100110011",
  13099=>"111110110",
  13100=>"110111100",
  13101=>"001110110",
  13102=>"000000111",
  13103=>"001000001",
  13104=>"001011011",
  13105=>"001010101",
  13106=>"110111111",
  13107=>"110110111",
  13108=>"111100000",
  13109=>"110100110",
  13110=>"001000001",
  13111=>"000000000",
  13112=>"000000100",
  13113=>"111111111",
  13114=>"111111111",
  13115=>"101001000",
  13116=>"111000000",
  13117=>"000011001",
  13118=>"111011000",
  13119=>"000000111",
  13120=>"100000000",
  13121=>"101000111",
  13122=>"010110011",
  13123=>"111100100",
  13124=>"001000001",
  13125=>"001000000",
  13126=>"100101111",
  13127=>"000000000",
  13128=>"111100101",
  13129=>"010110110",
  13130=>"000110110",
  13131=>"000000000",
  13132=>"110111111",
  13133=>"000000000",
  13134=>"000000111",
  13135=>"101000000",
  13136=>"111111011",
  13137=>"000000000",
  13138=>"101111111",
  13139=>"001010010",
  13140=>"111111110",
  13141=>"001000001",
  13142=>"000000101",
  13143=>"001010000",
  13144=>"100000001",
  13145=>"010110111",
  13146=>"110000000",
  13147=>"100011001",
  13148=>"111111111",
  13149=>"111001011",
  13150=>"100110111",
  13151=>"111110000",
  13152=>"100111001",
  13153=>"111111111",
  13154=>"111111111",
  13155=>"010000000",
  13156=>"000000000",
  13157=>"000000001",
  13158=>"000000000",
  13159=>"000000000",
  13160=>"111110111",
  13161=>"111100000",
  13162=>"011010000",
  13163=>"000000000",
  13164=>"001000000",
  13165=>"000000001",
  13166=>"000111011",
  13167=>"111000111",
  13168=>"101000000",
  13169=>"001001001",
  13170=>"111111111",
  13171=>"011011000",
  13172=>"111000001",
  13173=>"111111111",
  13174=>"011011011",
  13175=>"000000000",
  13176=>"111111111",
  13177=>"000000000",
  13178=>"001000100",
  13179=>"000010001",
  13180=>"000110111",
  13181=>"111111111",
  13182=>"111101111",
  13183=>"111111100",
  13184=>"110110110",
  13185=>"010110111",
  13186=>"111000000",
  13187=>"000000000",
  13188=>"111111110",
  13189=>"001001000",
  13190=>"111111111",
  13191=>"100000000",
  13192=>"111101111",
  13193=>"111011011",
  13194=>"111111000",
  13195=>"000100111",
  13196=>"110110111",
  13197=>"001111100",
  13198=>"100000000",
  13199=>"000000000",
  13200=>"000011011",
  13201=>"111111111",
  13202=>"111101001",
  13203=>"111101000",
  13204=>"110000000",
  13205=>"010010000",
  13206=>"111111111",
  13207=>"001001001",
  13208=>"000000000",
  13209=>"010110110",
  13210=>"111111011",
  13211=>"000000111",
  13212=>"000000000",
  13213=>"110110010",
  13214=>"000000000",
  13215=>"110110111",
  13216=>"000000000",
  13217=>"111100111",
  13218=>"000000001",
  13219=>"000000111",
  13220=>"000100000",
  13221=>"111111111",
  13222=>"000000001",
  13223=>"111011011",
  13224=>"000111100",
  13225=>"110010000",
  13226=>"101001001",
  13227=>"000000000",
  13228=>"000000000",
  13229=>"010110110",
  13230=>"001111010",
  13231=>"101001001",
  13232=>"000000000",
  13233=>"011111111",
  13234=>"000111010",
  13235=>"011011111",
  13236=>"010000000",
  13237=>"000000010",
  13238=>"000001111",
  13239=>"000000000",
  13240=>"000000011",
  13241=>"011111011",
  13242=>"010110111",
  13243=>"110110100",
  13244=>"110111111",
  13245=>"111000000",
  13246=>"100111111",
  13247=>"111100100",
  13248=>"000000000",
  13249=>"111000000",
  13250=>"111110111",
  13251=>"111110010",
  13252=>"110110000",
  13253=>"001011111",
  13254=>"000011001",
  13255=>"010000101",
  13256=>"001000000",
  13257=>"000000111",
  13258=>"111111101",
  13259=>"010000000",
  13260=>"111111011",
  13261=>"111110111",
  13262=>"001111111",
  13263=>"000000111",
  13264=>"110100000",
  13265=>"001001111",
  13266=>"001000000",
  13267=>"000110000",
  13268=>"011111000",
  13269=>"011010000",
  13270=>"000000000",
  13271=>"000000000",
  13272=>"000000000",
  13273=>"000100110",
  13274=>"111111111",
  13275=>"111111111",
  13276=>"000000000",
  13277=>"110110011",
  13278=>"111111011",
  13279=>"111101000",
  13280=>"111101111",
  13281=>"000000000",
  13282=>"101101101",
  13283=>"001000111",
  13284=>"110111000",
  13285=>"001000000",
  13286=>"110100111",
  13287=>"000000000",
  13288=>"000000001",
  13289=>"111111110",
  13290=>"000111111",
  13291=>"011111001",
  13292=>"110111011",
  13293=>"001001001",
  13294=>"000000000",
  13295=>"000001011",
  13296=>"000000000",
  13297=>"011111111",
  13298=>"000000000",
  13299=>"000000000",
  13300=>"110110010",
  13301=>"001101100",
  13302=>"111001000",
  13303=>"001101111",
  13304=>"100110100",
  13305=>"110011011",
  13306=>"000010010",
  13307=>"111111111",
  13308=>"000000000",
  13309=>"010111111",
  13310=>"111000000",
  13311=>"100000101",
  13312=>"000000000",
  13313=>"110000000",
  13314=>"011111111",
  13315=>"000000000",
  13316=>"111111111",
  13317=>"101001111",
  13318=>"000111111",
  13319=>"001001001",
  13320=>"100000110",
  13321=>"111111111",
  13322=>"100100111",
  13323=>"000000000",
  13324=>"000000000",
  13325=>"101001001",
  13326=>"000000000",
  13327=>"111011000",
  13328=>"000000000",
  13329=>"000000001",
  13330=>"001011001",
  13331=>"000000000",
  13332=>"111011001",
  13333=>"000001110",
  13334=>"111100110",
  13335=>"011001001",
  13336=>"000000000",
  13337=>"011011010",
  13338=>"000000001",
  13339=>"111000100",
  13340=>"110100000",
  13341=>"000100000",
  13342=>"111011111",
  13343=>"000001111",
  13344=>"000000011",
  13345=>"110110110",
  13346=>"111111110",
  13347=>"100100000",
  13348=>"000111000",
  13349=>"000000000",
  13350=>"111111111",
  13351=>"111101001",
  13352=>"111111101",
  13353=>"010010100",
  13354=>"000000000",
  13355=>"001000101",
  13356=>"111111001",
  13357=>"111111111",
  13358=>"110000000",
  13359=>"001011100",
  13360=>"111111111",
  13361=>"000110000",
  13362=>"111011011",
  13363=>"010010000",
  13364=>"111111111",
  13365=>"000000000",
  13366=>"111110111",
  13367=>"001101111",
  13368=>"000000000",
  13369=>"100110110",
  13370=>"000101111",
  13371=>"111110000",
  13372=>"101101111",
  13373=>"001001000",
  13374=>"000000000",
  13375=>"111111111",
  13376=>"000111100",
  13377=>"111111111",
  13378=>"001111100",
  13379=>"111111111",
  13380=>"000000000",
  13381=>"110000000",
  13382=>"000000100",
  13383=>"111111111",
  13384=>"010010000",
  13385=>"111111111",
  13386=>"111111111",
  13387=>"111111111",
  13388=>"001111111",
  13389=>"111111111",
  13390=>"001001001",
  13391=>"111111111",
  13392=>"100110111",
  13393=>"111111111",
  13394=>"110111111",
  13395=>"000000000",
  13396=>"000111100",
  13397=>"111111111",
  13398=>"111000100",
  13399=>"000000000",
  13400=>"000100100",
  13401=>"111101101",
  13402=>"111000111",
  13403=>"111111111",
  13404=>"000000000",
  13405=>"000110110",
  13406=>"000001000",
  13407=>"110000000",
  13408=>"000000000",
  13409=>"110100100",
  13410=>"111111000",
  13411=>"111111111",
  13412=>"001001110",
  13413=>"010000010",
  13414=>"110000100",
  13415=>"111111111",
  13416=>"101001000",
  13417=>"010000000",
  13418=>"111111111",
  13419=>"100000000",
  13420=>"000000000",
  13421=>"111111110",
  13422=>"111111011",
  13423=>"100100000",
  13424=>"011011111",
  13425=>"011111111",
  13426=>"000000000",
  13427=>"000000000",
  13428=>"010110100",
  13429=>"111111111",
  13430=>"111000010",
  13431=>"000000101",
  13432=>"111111111",
  13433=>"100110100",
  13434=>"000000000",
  13435=>"011111111",
  13436=>"100110110",
  13437=>"111111111",
  13438=>"000000000",
  13439=>"000000000",
  13440=>"001111101",
  13441=>"000000000",
  13442=>"111000111",
  13443=>"000000000",
  13444=>"111011111",
  13445=>"000000100",
  13446=>"000001101",
  13447=>"111111111",
  13448=>"100000011",
  13449=>"000000000",
  13450=>"000100100",
  13451=>"000000000",
  13452=>"111110000",
  13453=>"000000011",
  13454=>"011000000",
  13455=>"000000100",
  13456=>"011111111",
  13457=>"000001111",
  13458=>"001000000",
  13459=>"100100000",
  13460=>"011010000",
  13461=>"000010000",
  13462=>"111111111",
  13463=>"111111111",
  13464=>"000111111",
  13465=>"111111111",
  13466=>"110110110",
  13467=>"000001111",
  13468=>"011111111",
  13469=>"001000111",
  13470=>"000010000",
  13471=>"111111111",
  13472=>"010010000",
  13473=>"000000000",
  13474=>"000000000",
  13475=>"111100100",
  13476=>"000010010",
  13477=>"111111000",
  13478=>"111111111",
  13479=>"011011011",
  13480=>"000000000",
  13481=>"111111111",
  13482=>"000000000",
  13483=>"111111110",
  13484=>"111101111",
  13485=>"110100000",
  13486=>"000001111",
  13487=>"110111111",
  13488=>"000111101",
  13489=>"110110111",
  13490=>"110111111",
  13491=>"011000000",
  13492=>"111100000",
  13493=>"000001111",
  13494=>"100110111",
  13495=>"001001001",
  13496=>"111101011",
  13497=>"001001101",
  13498=>"000100011",
  13499=>"111111111",
  13500=>"000000000",
  13501=>"111111111",
  13502=>"000000000",
  13503=>"000010000",
  13504=>"001111111",
  13505=>"010111111",
  13506=>"000000001",
  13507=>"111111111",
  13508=>"111101111",
  13509=>"111111111",
  13510=>"111111111",
  13511=>"000110111",
  13512=>"100000111",
  13513=>"111111000",
  13514=>"000000110",
  13515=>"111111111",
  13516=>"000000000",
  13517=>"000000000",
  13518=>"111000000",
  13519=>"011011000",
  13520=>"001001111",
  13521=>"110100101",
  13522=>"000000000",
  13523=>"100001001",
  13524=>"000000000",
  13525=>"000000001",
  13526=>"000000000",
  13527=>"101101111",
  13528=>"111111100",
  13529=>"110111011",
  13530=>"111111111",
  13531=>"001111100",
  13532=>"000000100",
  13533=>"111111111",
  13534=>"001000000",
  13535=>"001000011",
  13536=>"111000000",
  13537=>"010110110",
  13538=>"111111001",
  13539=>"111111011",
  13540=>"000000000",
  13541=>"111111111",
  13542=>"000000010",
  13543=>"000000000",
  13544=>"111001111",
  13545=>"000000000",
  13546=>"000001000",
  13547=>"000000000",
  13548=>"000000000",
  13549=>"001000110",
  13550=>"111111111",
  13551=>"000111111",
  13552=>"111100100",
  13553=>"000100001",
  13554=>"000000000",
  13555=>"000000000",
  13556=>"000111111",
  13557=>"001000011",
  13558=>"001000000",
  13559=>"000000000",
  13560=>"000010011",
  13561=>"000000000",
  13562=>"000000000",
  13563=>"000101000",
  13564=>"111111111",
  13565=>"011011001",
  13566=>"111000100",
  13567=>"000001000",
  13568=>"011001111",
  13569=>"111100100",
  13570=>"000000110",
  13571=>"001001111",
  13572=>"111111111",
  13573=>"011011111",
  13574=>"100100110",
  13575=>"000110111",
  13576=>"000111110",
  13577=>"000000111",
  13578=>"111100111",
  13579=>"111111111",
  13580=>"001001011",
  13581=>"000000011",
  13582=>"111111111",
  13583=>"000000000",
  13584=>"000000000",
  13585=>"001000000",
  13586=>"111011000",
  13587=>"000000000",
  13588=>"000001111",
  13589=>"111111111",
  13590=>"111111100",
  13591=>"000000110",
  13592=>"111011001",
  13593=>"000010110",
  13594=>"011011000",
  13595=>"111111111",
  13596=>"111111111",
  13597=>"100000000",
  13598=>"000100111",
  13599=>"010011111",
  13600=>"001100000",
  13601=>"000000000",
  13602=>"000000000",
  13603=>"000000000",
  13604=>"000000000",
  13605=>"000000000",
  13606=>"000000010",
  13607=>"001101111",
  13608=>"000000000",
  13609=>"000000000",
  13610=>"111111111",
  13611=>"000000000",
  13612=>"111111111",
  13613=>"000000000",
  13614=>"000000001",
  13615=>"000000011",
  13616=>"111111111",
  13617=>"100100110",
  13618=>"001011111",
  13619=>"111000000",
  13620=>"111111111",
  13621=>"000000000",
  13622=>"000110111",
  13623=>"111100111",
  13624=>"111111111",
  13625=>"111011000",
  13626=>"111111010",
  13627=>"001000000",
  13628=>"111111111",
  13629=>"000000000",
  13630=>"110110111",
  13631=>"000000000",
  13632=>"111111100",
  13633=>"010101000",
  13634=>"000111111",
  13635=>"100110110",
  13636=>"100000000",
  13637=>"000100100",
  13638=>"110000000",
  13639=>"000000000",
  13640=>"000000000",
  13641=>"111011111",
  13642=>"110101111",
  13643=>"111111111",
  13644=>"101101111",
  13645=>"000000000",
  13646=>"000000001",
  13647=>"000010000",
  13648=>"110110000",
  13649=>"001001111",
  13650=>"010010010",
  13651=>"110100000",
  13652=>"100111111",
  13653=>"011011011",
  13654=>"111110111",
  13655=>"111000000",
  13656=>"111111111",
  13657=>"000000101",
  13658=>"111000100",
  13659=>"000000000",
  13660=>"011011011",
  13661=>"000000100",
  13662=>"000000011",
  13663=>"111011000",
  13664=>"111111111",
  13665=>"000000000",
  13666=>"001011111",
  13667=>"000000000",
  13668=>"000110000",
  13669=>"000000000",
  13670=>"000000010",
  13671=>"111111111",
  13672=>"111111110",
  13673=>"111010000",
  13674=>"110110110",
  13675=>"111111100",
  13676=>"000000000",
  13677=>"000000001",
  13678=>"100010000",
  13679=>"111111111",
  13680=>"111111110",
  13681=>"000000000",
  13682=>"110110110",
  13683=>"000000000",
  13684=>"000011111",
  13685=>"000100000",
  13686=>"000000001",
  13687=>"000000000",
  13688=>"000000000",
  13689=>"000011001",
  13690=>"111111111",
  13691=>"000111110",
  13692=>"101110111",
  13693=>"111111111",
  13694=>"000000000",
  13695=>"111111111",
  13696=>"000000001",
  13697=>"110100110",
  13698=>"010000000",
  13699=>"111111111",
  13700=>"111111000",
  13701=>"001000011",
  13702=>"111101111",
  13703=>"000000000",
  13704=>"010011111",
  13705=>"111001111",
  13706=>"000100000",
  13707=>"111111000",
  13708=>"111111111",
  13709=>"001100100",
  13710=>"000000000",
  13711=>"000000000",
  13712=>"000011011",
  13713=>"000000000",
  13714=>"001111111",
  13715=>"111111001",
  13716=>"111111111",
  13717=>"000001001",
  13718=>"100000100",
  13719=>"000000000",
  13720=>"111000000",
  13721=>"110110110",
  13722=>"000000000",
  13723=>"000000000",
  13724=>"011111000",
  13725=>"111111111",
  13726=>"000001001",
  13727=>"110110110",
  13728=>"111111111",
  13729=>"001000100",
  13730=>"000110100",
  13731=>"001001011",
  13732=>"111111101",
  13733=>"111111111",
  13734=>"011001111",
  13735=>"111101000",
  13736=>"000000000",
  13737=>"010000100",
  13738=>"000000111",
  13739=>"000010000",
  13740=>"111111111",
  13741=>"111100000",
  13742=>"000000111",
  13743=>"100100001",
  13744=>"000000000",
  13745=>"100110000",
  13746=>"111111000",
  13747=>"011000000",
  13748=>"000000110",
  13749=>"111011000",
  13750=>"100000000",
  13751=>"110100000",
  13752=>"111111111",
  13753=>"000000110",
  13754=>"000000000",
  13755=>"000100100",
  13756=>"111111010",
  13757=>"100110110",
  13758=>"001001000",
  13759=>"101111111",
  13760=>"000000000",
  13761=>"000111111",
  13762=>"000000000",
  13763=>"000000100",
  13764=>"011111001",
  13765=>"111011011",
  13766=>"011111101",
  13767=>"111110110",
  13768=>"000000100",
  13769=>"000000000",
  13770=>"000000111",
  13771=>"111111111",
  13772=>"100000000",
  13773=>"000000000",
  13774=>"001100011",
  13775=>"111110110",
  13776=>"111001011",
  13777=>"100111011",
  13778=>"111000000",
  13779=>"100010000",
  13780=>"011010001",
  13781=>"000000000",
  13782=>"000001110",
  13783=>"000000000",
  13784=>"000100111",
  13785=>"011111111",
  13786=>"000000000",
  13787=>"000000000",
  13788=>"000110100",
  13789=>"111110111",
  13790=>"000000001",
  13791=>"000100111",
  13792=>"001000000",
  13793=>"110110110",
  13794=>"000000001",
  13795=>"000000000",
  13796=>"111111111",
  13797=>"000000000",
  13798=>"011011000",
  13799=>"101000000",
  13800=>"111101111",
  13801=>"111111111",
  13802=>"101000110",
  13803=>"000000000",
  13804=>"100100111",
  13805=>"001000000",
  13806=>"111001000",
  13807=>"000100100",
  13808=>"000000000",
  13809=>"000100100",
  13810=>"000000000",
  13811=>"000000000",
  13812=>"111111100",
  13813=>"011111111",
  13814=>"110110000",
  13815=>"110110110",
  13816=>"001000110",
  13817=>"100110111",
  13818=>"111100000",
  13819=>"000000000",
  13820=>"100000100",
  13821=>"001001110",
  13822=>"000010110",
  13823=>"000100100",
  13824=>"001111111",
  13825=>"011111111",
  13826=>"111011111",
  13827=>"000000000",
  13828=>"011000000",
  13829=>"111110100",
  13830=>"001111111",
  13831=>"110111111",
  13832=>"000110000",
  13833=>"011111111",
  13834=>"011101000",
  13835=>"111011111",
  13836=>"000000000",
  13837=>"001000000",
  13838=>"000000000",
  13839=>"111111111",
  13840=>"111111000",
  13841=>"110101000",
  13842=>"011111111",
  13843=>"111111110",
  13844=>"001011000",
  13845=>"101001111",
  13846=>"110110111",
  13847=>"011111111",
  13848=>"111111011",
  13849=>"111001100",
  13850=>"000000000",
  13851=>"111110100",
  13852=>"001000000",
  13853=>"000110111",
  13854=>"100100101",
  13855=>"110000000",
  13856=>"111000000",
  13857=>"001110110",
  13858=>"110100110",
  13859=>"000111111",
  13860=>"000000000",
  13861=>"011000000",
  13862=>"000000000",
  13863=>"111001000",
  13864=>"000000000",
  13865=>"101000000",
  13866=>"111101111",
  13867=>"000000000",
  13868=>"111001001",
  13869=>"111111010",
  13870=>"000101101",
  13871=>"011001001",
  13872=>"001000001",
  13873=>"000111111",
  13874=>"011001000",
  13875=>"011011000",
  13876=>"111000000",
  13877=>"000111110",
  13878=>"010001000",
  13879=>"011000000",
  13880=>"000000000",
  13881=>"000000000",
  13882=>"000000000",
  13883=>"111111000",
  13884=>"010000000",
  13885=>"111111111",
  13886=>"110110111",
  13887=>"111001001",
  13888=>"000000000",
  13889=>"011000000",
  13890=>"000000000",
  13891=>"100000101",
  13892=>"110110110",
  13893=>"100110111",
  13894=>"001111000",
  13895=>"000000000",
  13896=>"000001000",
  13897=>"100101000",
  13898=>"000001111",
  13899=>"111011000",
  13900=>"001001000",
  13901=>"000000000",
  13902=>"010111111",
  13903=>"111000000",
  13904=>"111111100",
  13905=>"000010111",
  13906=>"011000110",
  13907=>"000110111",
  13908=>"000000000",
  13909=>"000000000",
  13910=>"011000101",
  13911=>"111111001",
  13912=>"111111111",
  13913=>"111001101",
  13914=>"010110111",
  13915=>"001000000",
  13916=>"001001111",
  13917=>"000000000",
  13918=>"000111111",
  13919=>"111000000",
  13920=>"111101000",
  13921=>"000000000",
  13922=>"111111110",
  13923=>"000000011",
  13924=>"001000000",
  13925=>"111100000",
  13926=>"000111111",
  13927=>"111100101",
  13928=>"111111000",
  13929=>"111001000",
  13930=>"000000000",
  13931=>"100110000",
  13932=>"011110111",
  13933=>"111000101",
  13934=>"111000000",
  13935=>"000000000",
  13936=>"000111111",
  13937=>"111111001",
  13938=>"000011000",
  13939=>"110111111",
  13940=>"000000000",
  13941=>"111111010",
  13942=>"001001000",
  13943=>"001001001",
  13944=>"111111111",
  13945=>"110111000",
  13946=>"111111111",
  13947=>"001000100",
  13948=>"000111110",
  13949=>"111111011",
  13950=>"111111000",
  13951=>"000000000",
  13952=>"000111111",
  13953=>"110000000",
  13954=>"100000000",
  13955=>"000001001",
  13956=>"000001101",
  13957=>"111000000",
  13958=>"110100111",
  13959=>"000000000",
  13960=>"000000111",
  13961=>"111111111",
  13962=>"110111001",
  13963=>"111111111",
  13964=>"011111111",
  13965=>"110010000",
  13966=>"011000000",
  13967=>"000111110",
  13968=>"110111111",
  13969=>"111111000",
  13970=>"111111111",
  13971=>"111110000",
  13972=>"000000000",
  13973=>"101111111",
  13974=>"011000000",
  13975=>"000000111",
  13976=>"001111111",
  13977=>"110111101",
  13978=>"000000000",
  13979=>"111011000",
  13980=>"111111011",
  13981=>"111000000",
  13982=>"000000000",
  13983=>"000000111",
  13984=>"111000000",
  13985=>"111111001",
  13986=>"000001111",
  13987=>"110111111",
  13988=>"110000110",
  13989=>"000000000",
  13990=>"000011111",
  13991=>"100110011",
  13992=>"000000000",
  13993=>"001111111",
  13994=>"000111111",
  13995=>"111111101",
  13996=>"110111001",
  13997=>"111101000",
  13998=>"101101000",
  13999=>"000000000",
  14000=>"000000000",
  14001=>"001000000",
  14002=>"110111111",
  14003=>"111111001",
  14004=>"110000001",
  14005=>"111001000",
  14006=>"000000010",
  14007=>"000000011",
  14008=>"000000110",
  14009=>"100101100",
  14010=>"111000000",
  14011=>"010000001",
  14012=>"000110000",
  14013=>"111111000",
  14014=>"101110111",
  14015=>"111100000",
  14016=>"001101000",
  14017=>"111111100",
  14018=>"111111100",
  14019=>"000000011",
  14020=>"111000000",
  14021=>"011011111",
  14022=>"111101101",
  14023=>"111000001",
  14024=>"111000000",
  14025=>"111101101",
  14026=>"101001001",
  14027=>"010011000",
  14028=>"011111111",
  14029=>"011000000",
  14030=>"000101101",
  14031=>"111111000",
  14032=>"000000000",
  14033=>"110100000",
  14034=>"000111111",
  14035=>"000000111",
  14036=>"000110111",
  14037=>"000010011",
  14038=>"000110111",
  14039=>"001000101",
  14040=>"000111111",
  14041=>"000100100",
  14042=>"000000000",
  14043=>"000110111",
  14044=>"111111011",
  14045=>"000000111",
  14046=>"111000000",
  14047=>"000001111",
  14048=>"111000000",
  14049=>"111000000",
  14050=>"110110110",
  14051=>"111011000",
  14052=>"111000000",
  14053=>"100000001",
  14054=>"110010010",
  14055=>"111100100",
  14056=>"111011001",
  14057=>"111001111",
  14058=>"100111111",
  14059=>"101111111",
  14060=>"000000011",
  14061=>"000000111",
  14062=>"000000000",
  14063=>"000111111",
  14064=>"111111001",
  14065=>"000000010",
  14066=>"110111111",
  14067=>"000000000",
  14068=>"011010111",
  14069=>"101111000",
  14070=>"000100110",
  14071=>"101000000",
  14072=>"111011000",
  14073=>"000000100",
  14074=>"010011000",
  14075=>"100000000",
  14076=>"100000000",
  14077=>"110000000",
  14078=>"000000001",
  14079=>"000000000",
  14080=>"000000000",
  14081=>"110100000",
  14082=>"111111111",
  14083=>"010000011",
  14084=>"000001000",
  14085=>"000110111",
  14086=>"000010000",
  14087=>"000110111",
  14088=>"001111001",
  14089=>"000000000",
  14090=>"111111111",
  14091=>"000111101",
  14092=>"111101101",
  14093=>"000110111",
  14094=>"101101100",
  14095=>"100110000",
  14096=>"111111100",
  14097=>"000000000",
  14098=>"000000101",
  14099=>"111111111",
  14100=>"110111010",
  14101=>"101111111",
  14102=>"001000000",
  14103=>"111111011",
  14104=>"001001000",
  14105=>"111000000",
  14106=>"111111100",
  14107=>"000000000",
  14108=>"110000000",
  14109=>"000011111",
  14110=>"000000011",
  14111=>"001101001",
  14112=>"000000110",
  14113=>"111111111",
  14114=>"101100000",
  14115=>"000110111",
  14116=>"000000000",
  14117=>"111000011",
  14118=>"000000011",
  14119=>"111111111",
  14120=>"001000001",
  14121=>"111100000",
  14122=>"111000000",
  14123=>"111000000",
  14124=>"000000000",
  14125=>"111111111",
  14126=>"111111111",
  14127=>"111110011",
  14128=>"011111111",
  14129=>"111111011",
  14130=>"110111111",
  14131=>"011111111",
  14132=>"111111111",
  14133=>"000000111",
  14134=>"101101111",
  14135=>"101000100",
  14136=>"000000000",
  14137=>"000100100",
  14138=>"001100001",
  14139=>"111110110",
  14140=>"000011010",
  14141=>"000000000",
  14142=>"111111101",
  14143=>"111111111",
  14144=>"000000000",
  14145=>"000100101",
  14146=>"000000000",
  14147=>"000000101",
  14148=>"000010111",
  14149=>"000000000",
  14150=>"101111100",
  14151=>"111111011",
  14152=>"111000000",
  14153=>"111001001",
  14154=>"111111000",
  14155=>"111000000",
  14156=>"101001000",
  14157=>"010111011",
  14158=>"011000000",
  14159=>"001011011",
  14160=>"110000010",
  14161=>"000000010",
  14162=>"111111100",
  14163=>"111111111",
  14164=>"001000000",
  14165=>"101010001",
  14166=>"000110000",
  14167=>"111001000",
  14168=>"011111110",
  14169=>"011000111",
  14170=>"000000011",
  14171=>"011110000",
  14172=>"111001001",
  14173=>"111101000",
  14174=>"111111101",
  14175=>"010011001",
  14176=>"000111111",
  14177=>"000000110",
  14178=>"001000000",
  14179=>"010111111",
  14180=>"000100110",
  14181=>"111001000",
  14182=>"010111111",
  14183=>"111111001",
  14184=>"111101000",
  14185=>"000000010",
  14186=>"111111100",
  14187=>"000001001",
  14188=>"110101001",
  14189=>"000000111",
  14190=>"000100111",
  14191=>"010010110",
  14192=>"111000000",
  14193=>"110110010",
  14194=>"111000000",
  14195=>"000011011",
  14196=>"111111111",
  14197=>"111111111",
  14198=>"000000000",
  14199=>"000000001",
  14200=>"000000010",
  14201=>"101100000",
  14202=>"111101000",
  14203=>"110110000",
  14204=>"000000000",
  14205=>"100101111",
  14206=>"000100000",
  14207=>"000000111",
  14208=>"111001101",
  14209=>"011000000",
  14210=>"001011111",
  14211=>"111001000",
  14212=>"111011111",
  14213=>"110100000",
  14214=>"111101000",
  14215=>"100110111",
  14216=>"101111111",
  14217=>"000110100",
  14218=>"111001101",
  14219=>"111100110",
  14220=>"111111111",
  14221=>"000100110",
  14222=>"001000000",
  14223=>"000000000",
  14224=>"111111111",
  14225=>"000110110",
  14226=>"001111111",
  14227=>"001110110",
  14228=>"111111111",
  14229=>"110110000",
  14230=>"111111111",
  14231=>"011011010",
  14232=>"011000100",
  14233=>"111101000",
  14234=>"111111100",
  14235=>"111111111",
  14236=>"000010011",
  14237=>"111001000",
  14238=>"100110110",
  14239=>"000111000",
  14240=>"111100000",
  14241=>"111111111",
  14242=>"111101000",
  14243=>"000010111",
  14244=>"000101000",
  14245=>"111111110",
  14246=>"000000111",
  14247=>"111111000",
  14248=>"110000100",
  14249=>"000110111",
  14250=>"000000000",
  14251=>"000000000",
  14252=>"001111111",
  14253=>"000000000",
  14254=>"111000111",
  14255=>"000001001",
  14256=>"000000011",
  14257=>"111111111",
  14258=>"000100000",
  14259=>"111010111",
  14260=>"111111111",
  14261=>"111111100",
  14262=>"000000000",
  14263=>"111000000",
  14264=>"000000000",
  14265=>"011001001",
  14266=>"100101111",
  14267=>"000000111",
  14268=>"000000000",
  14269=>"011001000",
  14270=>"111100000",
  14271=>"111000000",
  14272=>"000000000",
  14273=>"111111111",
  14274=>"110111111",
  14275=>"000000010",
  14276=>"110111000",
  14277=>"001001001",
  14278=>"111000000",
  14279=>"110000000",
  14280=>"000000000",
  14281=>"110110110",
  14282=>"000000000",
  14283=>"000000111",
  14284=>"000111111",
  14285=>"000110111",
  14286=>"000001101",
  14287=>"000110111",
  14288=>"111000000",
  14289=>"111111111",
  14290=>"111111110",
  14291=>"110100101",
  14292=>"001011111",
  14293=>"000111111",
  14294=>"111101000",
  14295=>"000000000",
  14296=>"000000000",
  14297=>"000010111",
  14298=>"111111110",
  14299=>"110111000",
  14300=>"000000000",
  14301=>"111110110",
  14302=>"000000000",
  14303=>"111100001",
  14304=>"001000000",
  14305=>"111111111",
  14306=>"110111111",
  14307=>"111111100",
  14308=>"110000000",
  14309=>"000010000",
  14310=>"100100000",
  14311=>"000010111",
  14312=>"000001000",
  14313=>"001000000",
  14314=>"111111000",
  14315=>"000101111",
  14316=>"011001111",
  14317=>"110100001",
  14318=>"000101001",
  14319=>"111111011",
  14320=>"111111111",
  14321=>"111111111",
  14322=>"000001100",
  14323=>"111111011",
  14324=>"000011000",
  14325=>"000111111",
  14326=>"000000000",
  14327=>"110101001",
  14328=>"000001111",
  14329=>"000001001",
  14330=>"000000110",
  14331=>"111110110",
  14332=>"100000000",
  14333=>"101001000",
  14334=>"011001001",
  14335=>"000001111",
  14336=>"011101001",
  14337=>"000000000",
  14338=>"101001001",
  14339=>"111110100",
  14340=>"000000100",
  14341=>"111001111",
  14342=>"000000000",
  14343=>"000000000",
  14344=>"111100010",
  14345=>"111110100",
  14346=>"000000001",
  14347=>"011000011",
  14348=>"000000000",
  14349=>"011111101",
  14350=>"000110111",
  14351=>"111111111",
  14352=>"111111101",
  14353=>"011110100",
  14354=>"100000001",
  14355=>"111001000",
  14356=>"111111111",
  14357=>"111111010",
  14358=>"000000000",
  14359=>"011001000",
  14360=>"111111001",
  14361=>"110100000",
  14362=>"111000000",
  14363=>"111100100",
  14364=>"111111011",
  14365=>"000000000",
  14366=>"100100100",
  14367=>"000111111",
  14368=>"111111111",
  14369=>"011010000",
  14370=>"111110100",
  14371=>"000010111",
  14372=>"111111111",
  14373=>"001000000",
  14374=>"111111111",
  14375=>"001011000",
  14376=>"111101000",
  14377=>"000000000",
  14378=>"000000000",
  14379=>"000111111",
  14380=>"111111111",
  14381=>"111100000",
  14382=>"111111111",
  14383=>"000000001",
  14384=>"011011111",
  14385=>"000000000",
  14386=>"111111001",
  14387=>"010110100",
  14388=>"110100001",
  14389=>"000000000",
  14390=>"111111111",
  14391=>"101101001",
  14392=>"000001000",
  14393=>"111101111",
  14394=>"000000000",
  14395=>"111000000",
  14396=>"101111111",
  14397=>"000000000",
  14398=>"000000000",
  14399=>"001000000",
  14400=>"001111111",
  14401=>"111110010",
  14402=>"000000000",
  14403=>"111111110",
  14404=>"101001011",
  14405=>"000000000",
  14406=>"111011111",
  14407=>"111111111",
  14408=>"000010000",
  14409=>"000000100",
  14410=>"000000101",
  14411=>"111111111",
  14412=>"000000001",
  14413=>"000000111",
  14414=>"011000000",
  14415=>"111111111",
  14416=>"111011000",
  14417=>"100000000",
  14418=>"111000000",
  14419=>"000111111",
  14420=>"000000000",
  14421=>"000000000",
  14422=>"000001000",
  14423=>"000000000",
  14424=>"111111000",
  14425=>"111101001",
  14426=>"111111111",
  14427=>"111111111",
  14428=>"000000000",
  14429=>"111111111",
  14430=>"111111111",
  14431=>"000111000",
  14432=>"000000000",
  14433=>"110010111",
  14434=>"111111111",
  14435=>"011001010",
  14436=>"110000000",
  14437=>"111111111",
  14438=>"111111111",
  14439=>"000000000",
  14440=>"001111111",
  14441=>"111111111",
  14442=>"111111000",
  14443=>"000000011",
  14444=>"000000000",
  14445=>"001001111",
  14446=>"111111111",
  14447=>"100100100",
  14448=>"000000111",
  14449=>"111111111",
  14450=>"111100101",
  14451=>"101101001",
  14452=>"111111111",
  14453=>"111111101",
  14454=>"000000000",
  14455=>"000000000",
  14456=>"011001001",
  14457=>"000000001",
  14458=>"000000000",
  14459=>"111111111",
  14460=>"100100100",
  14461=>"000000000",
  14462=>"000001001",
  14463=>"111111111",
  14464=>"111111011",
  14465=>"011001100",
  14466=>"111110100",
  14467=>"000100100",
  14468=>"000000000",
  14469=>"111101111",
  14470=>"000000000",
  14471=>"000000000",
  14472=>"111111111",
  14473=>"111000000",
  14474=>"000000000",
  14475=>"011010000",
  14476=>"100000000",
  14477=>"010000000",
  14478=>"000000100",
  14479=>"010010000",
  14480=>"111111111",
  14481=>"111111111",
  14482=>"111001111",
  14483=>"111110010",
  14484=>"001101111",
  14485=>"110010000",
  14486=>"001011111",
  14487=>"111111111",
  14488=>"111111111",
  14489=>"000000000",
  14490=>"001001100",
  14491=>"111100111",
  14492=>"111000111",
  14493=>"111001001",
  14494=>"100111101",
  14495=>"111111111",
  14496=>"001000000",
  14497=>"111010110",
  14498=>"111111111",
  14499=>"111111111",
  14500=>"000000000",
  14501=>"011001001",
  14502=>"111111111",
  14503=>"110110100",
  14504=>"111101100",
  14505=>"111111000",
  14506=>"000010010",
  14507=>"110000000",
  14508=>"111011000",
  14509=>"100100100",
  14510=>"000000000",
  14511=>"111111111",
  14512=>"111111111",
  14513=>"100100000",
  14514=>"111111111",
  14515=>"000000000",
  14516=>"111011011",
  14517=>"110000111",
  14518=>"000000100",
  14519=>"110110000",
  14520=>"001001001",
  14521=>"001000000",
  14522=>"000000100",
  14523=>"001000000",
  14524=>"111111111",
  14525=>"011000000",
  14526=>"000010000",
  14527=>"101000001",
  14528=>"000000000",
  14529=>"001001011",
  14530=>"111111111",
  14531=>"000000000",
  14532=>"111111111",
  14533=>"111111111",
  14534=>"111111111",
  14535=>"000001001",
  14536=>"111000000",
  14537=>"000000100",
  14538=>"000110111",
  14539=>"100110111",
  14540=>"111111111",
  14541=>"111111111",
  14542=>"111000000",
  14543=>"000000000",
  14544=>"111100101",
  14545=>"000000100",
  14546=>"000000000",
  14547=>"101100111",
  14548=>"110111000",
  14549=>"111111111",
  14550=>"110111011",
  14551=>"101101101",
  14552=>"000000000",
  14553=>"001001101",
  14554=>"000000000",
  14555=>"111111111",
  14556=>"111101100",
  14557=>"111111111",
  14558=>"111111111",
  14559=>"110111111",
  14560=>"000000000",
  14561=>"110110111",
  14562=>"111000111",
  14563=>"011011110",
  14564=>"110000000",
  14565=>"111101111",
  14566=>"111110111",
  14567=>"001001011",
  14568=>"000000111",
  14569=>"000000000",
  14570=>"100000100",
  14571=>"101111111",
  14572=>"111111111",
  14573=>"000110111",
  14574=>"000010111",
  14575=>"000000000",
  14576=>"001111111",
  14577=>"111111101",
  14578=>"111111111",
  14579=>"000000101",
  14580=>"000010000",
  14581=>"100100100",
  14582=>"011000000",
  14583=>"000000111",
  14584=>"111111000",
  14585=>"000000000",
  14586=>"000000000",
  14587=>"000111111",
  14588=>"011111011",
  14589=>"001100100",
  14590=>"011000100",
  14591=>"000000000",
  14592=>"000000000",
  14593=>"101000000",
  14594=>"011111111",
  14595=>"100000000",
  14596=>"111111111",
  14597=>"000000000",
  14598=>"110111111",
  14599=>"001111111",
  14600=>"000111000",
  14601=>"000000011",
  14602=>"111101101",
  14603=>"000111001",
  14604=>"111001101",
  14605=>"000000011",
  14606=>"111111111",
  14607=>"101100010",
  14608=>"110010111",
  14609=>"000100100",
  14610=>"111001001",
  14611=>"111011101",
  14612=>"000000000",
  14613=>"111000100",
  14614=>"101101000",
  14615=>"001011111",
  14616=>"111111011",
  14617=>"111111011",
  14618=>"111000101",
  14619=>"111100111",
  14620=>"111111111",
  14621=>"000000010",
  14622=>"010011000",
  14623=>"000000100",
  14624=>"000001001",
  14625=>"011000111",
  14626=>"000111111",
  14627=>"000111111",
  14628=>"110000000",
  14629=>"111111111",
  14630=>"000111011",
  14631=>"000111111",
  14632=>"011000000",
  14633=>"000000000",
  14634=>"111111111",
  14635=>"000111111",
  14636=>"001111111",
  14637=>"000000001",
  14638=>"100000000",
  14639=>"000000000",
  14640=>"011011111",
  14641=>"111111001",
  14642=>"111000000",
  14643=>"111011011",
  14644=>"000000000",
  14645=>"000001001",
  14646=>"111001101",
  14647=>"000000000",
  14648=>"111111000",
  14649=>"111111111",
  14650=>"000101111",
  14651=>"000000110",
  14652=>"110100000",
  14653=>"111000001",
  14654=>"000010111",
  14655=>"011011110",
  14656=>"111111011",
  14657=>"000000001",
  14658=>"000000000",
  14659=>"111111001",
  14660=>"111111111",
  14661=>"000001100",
  14662=>"000000000",
  14663=>"111111000",
  14664=>"111111111",
  14665=>"010010000",
  14666=>"101100000",
  14667=>"111011111",
  14668=>"000000000",
  14669=>"100110010",
  14670=>"011100000",
  14671=>"111011011",
  14672=>"000000000",
  14673=>"111111111",
  14674=>"110111111",
  14675=>"111010110",
  14676=>"111101111",
  14677=>"011011011",
  14678=>"000000011",
  14679=>"000000000",
  14680=>"110000011",
  14681=>"111111111",
  14682=>"111111000",
  14683=>"000000000",
  14684=>"001001111",
  14685=>"111111111",
  14686=>"001100110",
  14687=>"001011111",
  14688=>"111111111",
  14689=>"000000111",
  14690=>"101001011",
  14691=>"000000000",
  14692=>"111111111",
  14693=>"111111111",
  14694=>"001011011",
  14695=>"001011001",
  14696=>"110100100",
  14697=>"000001111",
  14698=>"001011111",
  14699=>"100000101",
  14700=>"000000011",
  14701=>"000011011",
  14702=>"000110111",
  14703=>"000000100",
  14704=>"000000001",
  14705=>"000000000",
  14706=>"111100100",
  14707=>"011000000",
  14708=>"111111111",
  14709=>"010000100",
  14710=>"111000111",
  14711=>"000101111",
  14712=>"111100000",
  14713=>"000000000",
  14714=>"111111111",
  14715=>"110110100",
  14716=>"111111000",
  14717=>"001001111",
  14718=>"111101111",
  14719=>"000000000",
  14720=>"000000010",
  14721=>"110100001",
  14722=>"000100100",
  14723=>"001011111",
  14724=>"000000000",
  14725=>"111111111",
  14726=>"111110000",
  14727=>"000000000",
  14728=>"001000000",
  14729=>"000000001",
  14730=>"111001111",
  14731=>"100000111",
  14732=>"111111111",
  14733=>"111110111",
  14734=>"000000000",
  14735=>"000000000",
  14736=>"111000000",
  14737=>"111100100",
  14738=>"000000101",
  14739=>"010011000",
  14740=>"001000100",
  14741=>"000000000",
  14742=>"111100101",
  14743=>"000000000",
  14744=>"111000111",
  14745=>"111111111",
  14746=>"000011011",
  14747=>"000000000",
  14748=>"111111111",
  14749=>"111110111",
  14750=>"000000000",
  14751=>"000011111",
  14752=>"011000000",
  14753=>"100100100",
  14754=>"000000000",
  14755=>"011001001",
  14756=>"001101000",
  14757=>"001000000",
  14758=>"000000000",
  14759=>"111010011",
  14760=>"000000000",
  14761=>"001001111",
  14762=>"110110110",
  14763=>"000110110",
  14764=>"000000000",
  14765=>"000111111",
  14766=>"011111111",
  14767=>"000000001",
  14768=>"111111111",
  14769=>"111001000",
  14770=>"111111001",
  14771=>"000000000",
  14772=>"000000000",
  14773=>"000101111",
  14774=>"001011000",
  14775=>"000111011",
  14776=>"111000111",
  14777=>"111111111",
  14778=>"111111100",
  14779=>"111111000",
  14780=>"111111111",
  14781=>"111111000",
  14782=>"000000100",
  14783=>"101101101",
  14784=>"110010000",
  14785=>"101001000",
  14786=>"000000000",
  14787=>"001001100",
  14788=>"001011001",
  14789=>"111000101",
  14790=>"111001000",
  14791=>"000000000",
  14792=>"000010100",
  14793=>"000000111",
  14794=>"101101101",
  14795=>"000000000",
  14796=>"111111000",
  14797=>"000000000",
  14798=>"111101101",
  14799=>"111110100",
  14800=>"111001001",
  14801=>"011001111",
  14802=>"000000000",
  14803=>"000000000",
  14804=>"001000011",
  14805=>"111000001",
  14806=>"111111111",
  14807=>"000000011",
  14808=>"111111101",
  14809=>"111111110",
  14810=>"000000000",
  14811=>"000000001",
  14812=>"000001001",
  14813=>"000000000",
  14814=>"111111111",
  14815=>"010110110",
  14816=>"000000000",
  14817=>"111101101",
  14818=>"000000000",
  14819=>"111101001",
  14820=>"000000000",
  14821=>"111011001",
  14822=>"000001001",
  14823=>"000000000",
  14824=>"111001000",
  14825=>"000000100",
  14826=>"110111111",
  14827=>"100111100",
  14828=>"111111011",
  14829=>"011011101",
  14830=>"101000011",
  14831=>"001101111",
  14832=>"101001000",
  14833=>"110011111",
  14834=>"000000000",
  14835=>"111101101",
  14836=>"000000000",
  14837=>"111111001",
  14838=>"111111110",
  14839=>"001000111",
  14840=>"001111111",
  14841=>"111001001",
  14842=>"000001001",
  14843=>"001001101",
  14844=>"000000000",
  14845=>"000000110",
  14846=>"000000100",
  14847=>"000000000",
  14848=>"101111111",
  14849=>"000110000",
  14850=>"111111111",
  14851=>"110010000",
  14852=>"101111000",
  14853=>"011010000",
  14854=>"110111111",
  14855=>"111101111",
  14856=>"101000000",
  14857=>"000000111",
  14858=>"000100110",
  14859=>"111111111",
  14860=>"110111111",
  14861=>"000000000",
  14862=>"001111111",
  14863=>"110111100",
  14864=>"111011001",
  14865=>"110110111",
  14866=>"111100101",
  14867=>"000000000",
  14868=>"100000000",
  14869=>"111011101",
  14870=>"000000000",
  14871=>"111000000",
  14872=>"000100011",
  14873=>"000000000",
  14874=>"001000001",
  14875=>"100111100",
  14876=>"001111111",
  14877=>"110010000",
  14878=>"011011011",
  14879=>"110100000",
  14880=>"000001111",
  14881=>"110111000",
  14882=>"000001111",
  14883=>"000000111",
  14884=>"111111011",
  14885=>"110111111",
  14886=>"001111011",
  14887=>"000000100",
  14888=>"111000000",
  14889=>"111111111",
  14890=>"001000000",
  14891=>"111111111",
  14892=>"000110111",
  14893=>"000000001",
  14894=>"000000110",
  14895=>"111111101",
  14896=>"000111110",
  14897=>"000001000",
  14898=>"111111000",
  14899=>"111111110",
  14900=>"000011011",
  14901=>"110110110",
  14902=>"000000100",
  14903=>"110111011",
  14904=>"001000111",
  14905=>"111110000",
  14906=>"111111100",
  14907=>"001111111",
  14908=>"101000000",
  14909=>"111111000",
  14910=>"000000111",
  14911=>"000000000",
  14912=>"010010000",
  14913=>"000001001",
  14914=>"000000110",
  14915=>"111111000",
  14916=>"001111111",
  14917=>"001100100",
  14918=>"000110011",
  14919=>"000000000",
  14920=>"100111101",
  14921=>"000001111",
  14922=>"111111000",
  14923=>"011111111",
  14924=>"000010011",
  14925=>"111100000",
  14926=>"110110000",
  14927=>"001001100",
  14928=>"100100000",
  14929=>"110010000",
  14930=>"000000000",
  14931=>"101101100",
  14932=>"110100000",
  14933=>"100100100",
  14934=>"100101001",
  14935=>"000000001",
  14936=>"011001000",
  14937=>"111001111",
  14938=>"111111001",
  14939=>"100000111",
  14940=>"101010111",
  14941=>"011000000",
  14942=>"111001000",
  14943=>"110110110",
  14944=>"111111111",
  14945=>"001000000",
  14946=>"001111111",
  14947=>"001111111",
  14948=>"111110100",
  14949=>"100110110",
  14950=>"000000000",
  14951=>"000000001",
  14952=>"001011000",
  14953=>"111000010",
  14954=>"000000000",
  14955=>"011001000",
  14956=>"001001101",
  14957=>"000000000",
  14958=>"000000001",
  14959=>"100111001",
  14960=>"000000000",
  14961=>"000000011",
  14962=>"001111111",
  14963=>"000110110",
  14964=>"000000011",
  14965=>"100000010",
  14966=>"000001111",
  14967=>"011000110",
  14968=>"011000000",
  14969=>"000000000",
  14970=>"111101000",
  14971=>"000000000",
  14972=>"110000000",
  14973=>"110110011",
  14974=>"001000000",
  14975=>"111011000",
  14976=>"000000111",
  14977=>"000000001",
  14978=>"001011011",
  14979=>"111111000",
  14980=>"001001100",
  14981=>"000000000",
  14982=>"011001111",
  14983=>"111111101",
  14984=>"110111110",
  14985=>"000100000",
  14986=>"111111110",
  14987=>"000101111",
  14988=>"000001111",
  14989=>"000000111",
  14990=>"100000011",
  14991=>"000000000",
  14992=>"000000111",
  14993=>"000000000",
  14994=>"111110000",
  14995=>"011000000",
  14996=>"110000111",
  14997=>"000110111",
  14998=>"111111111",
  14999=>"111011001",
  15000=>"000000001",
  15001=>"111111010",
  15002=>"110100110",
  15003=>"000001000",
  15004=>"110100000",
  15005=>"110110010",
  15006=>"111111111",
  15007=>"010110110",
  15008=>"000110111",
  15009=>"001111011",
  15010=>"110110110",
  15011=>"111111010",
  15012=>"111111011",
  15013=>"110101101",
  15014=>"000100000",
  15015=>"001011011",
  15016=>"111111101",
  15017=>"000000100",
  15018=>"010000000",
  15019=>"000011001",
  15020=>"000100100",
  15021=>"100100011",
  15022=>"000000001",
  15023=>"011111011",
  15024=>"111111111",
  15025=>"111100001",
  15026=>"001111000",
  15027=>"000101111",
  15028=>"111010000",
  15029=>"000000000",
  15030=>"110110111",
  15031=>"111111010",
  15032=>"000001011",
  15033=>"111111111",
  15034=>"111011001",
  15035=>"111110000",
  15036=>"101001100",
  15037=>"000000111",
  15038=>"111100110",
  15039=>"111111111",
  15040=>"111101000",
  15041=>"000001001",
  15042=>"000000101",
  15043=>"111011111",
  15044=>"000101111",
  15045=>"001001001",
  15046=>"001000011",
  15047=>"100111000",
  15048=>"010011011",
  15049=>"111111110",
  15050=>"110010000",
  15051=>"000000000",
  15052=>"011111000",
  15053=>"001101100",
  15054=>"100010000",
  15055=>"000000110",
  15056=>"000100000",
  15057=>"000010001",
  15058=>"111111110",
  15059=>"111111110",
  15060=>"011001000",
  15061=>"111110011",
  15062=>"000000001",
  15063=>"111111011",
  15064=>"100110011",
  15065=>"110111111",
  15066=>"110111111",
  15067=>"111111111",
  15068=>"001000000",
  15069=>"100000100",
  15070=>"001000000",
  15071=>"000000000",
  15072=>"101001111",
  15073=>"000000001",
  15074=>"111100100",
  15075=>"000110100",
  15076=>"000011011",
  15077=>"011000000",
  15078=>"110110111",
  15079=>"000000111",
  15080=>"111111000",
  15081=>"001111111",
  15082=>"111111011",
  15083=>"111111111",
  15084=>"111100101",
  15085=>"110111111",
  15086=>"111000000",
  15087=>"111111111",
  15088=>"000000000",
  15089=>"111101101",
  15090=>"111100111",
  15091=>"110110110",
  15092=>"110000011",
  15093=>"101100100",
  15094=>"111111011",
  15095=>"011001000",
  15096=>"000111111",
  15097=>"111111000",
  15098=>"100100000",
  15099=>"001000100",
  15100=>"110110111",
  15101=>"001000000",
  15102=>"000000011",
  15103=>"010111110",
  15104=>"000000001",
  15105=>"000000100",
  15106=>"001000000",
  15107=>"111110000",
  15108=>"110110110",
  15109=>"000110111",
  15110=>"001000000",
  15111=>"111111001",
  15112=>"000001000",
  15113=>"001000001",
  15114=>"111100101",
  15115=>"111001011",
  15116=>"100100111",
  15117=>"000000100",
  15118=>"011111000",
  15119=>"111001100",
  15120=>"100000011",
  15121=>"000000100",
  15122=>"000000000",
  15123=>"001111111",
  15124=>"000001011",
  15125=>"111111111",
  15126=>"000110111",
  15127=>"100100111",
  15128=>"111110110",
  15129=>"111111100",
  15130=>"110111000",
  15131=>"000000111",
  15132=>"101101101",
  15133=>"000001000",
  15134=>"000000000",
  15135=>"000010111",
  15136=>"100111000",
  15137=>"000000000",
  15138=>"000000000",
  15139=>"000000110",
  15140=>"000010010",
  15141=>"110111111",
  15142=>"011011000",
  15143=>"110111000",
  15144=>"001111111",
  15145=>"011011111",
  15146=>"111111111",
  15147=>"001000000",
  15148=>"000000000",
  15149=>"001001001",
  15150=>"111100000",
  15151=>"000000001",
  15152=>"110110000",
  15153=>"100110110",
  15154=>"000000001",
  15155=>"000000111",
  15156=>"000000000",
  15157=>"011110110",
  15158=>"111111000",
  15159=>"011001001",
  15160=>"110010000",
  15161=>"100000001",
  15162=>"110000000",
  15163=>"011001000",
  15164=>"000000100",
  15165=>"110111110",
  15166=>"111001000",
  15167=>"110110100",
  15168=>"111000000",
  15169=>"100111000",
  15170=>"111111000",
  15171=>"000000001",
  15172=>"001100000",
  15173=>"100000000",
  15174=>"100110110",
  15175=>"001111011",
  15176=>"000000000",
  15177=>"111111100",
  15178=>"000110110",
  15179=>"011011001",
  15180=>"011110000",
  15181=>"001011000",
  15182=>"000000001",
  15183=>"000111111",
  15184=>"111000000",
  15185=>"110100111",
  15186=>"111110011",
  15187=>"001000000",
  15188=>"111101100",
  15189=>"011011011",
  15190=>"000000001",
  15191=>"100110111",
  15192=>"111111010",
  15193=>"000010011",
  15194=>"000111100",
  15195=>"111010000",
  15196=>"110000001",
  15197=>"001001001",
  15198=>"110100000",
  15199=>"000000110",
  15200=>"001011000",
  15201=>"000111000",
  15202=>"001001000",
  15203=>"000000001",
  15204=>"100100110",
  15205=>"010010000",
  15206=>"000000111",
  15207=>"110100110",
  15208=>"001001001",
  15209=>"100100000",
  15210=>"001101111",
  15211=>"110000000",
  15212=>"100111110",
  15213=>"010111111",
  15214=>"000111000",
  15215=>"001111100",
  15216=>"001001000",
  15217=>"000000000",
  15218=>"000111111",
  15219=>"111111111",
  15220=>"110000010",
  15221=>"010010111",
  15222=>"000000000",
  15223=>"111111000",
  15224=>"111111001",
  15225=>"101000000",
  15226=>"100110000",
  15227=>"000010100",
  15228=>"110110110",
  15229=>"011111111",
  15230=>"000000001",
  15231=>"000000111",
  15232=>"000111011",
  15233=>"010010011",
  15234=>"100110111",
  15235=>"100111000",
  15236=>"111111110",
  15237=>"111011011",
  15238=>"000000011",
  15239=>"000000111",
  15240=>"000000111",
  15241=>"111111000",
  15242=>"110110000",
  15243=>"000000000",
  15244=>"101111111",
  15245=>"100111011",
  15246=>"110011111",
  15247=>"000000111",
  15248=>"000000000",
  15249=>"101111111",
  15250=>"110110110",
  15251=>"000000111",
  15252=>"111111111",
  15253=>"000000010",
  15254=>"111111010",
  15255=>"111111000",
  15256=>"001001000",
  15257=>"000000000",
  15258=>"111111010",
  15259=>"111111110",
  15260=>"000000000",
  15261=>"110111110",
  15262=>"110011111",
  15263=>"111111111",
  15264=>"000000000",
  15265=>"011011001",
  15266=>"111111001",
  15267=>"111111001",
  15268=>"000000001",
  15269=>"111111100",
  15270=>"011111000",
  15271=>"101100000",
  15272=>"001001001",
  15273=>"111111100",
  15274=>"000000011",
  15275=>"110000100",
  15276=>"111111111",
  15277=>"001000100",
  15278=>"000110111",
  15279=>"000000110",
  15280=>"111110101",
  15281=>"101101111",
  15282=>"110111110",
  15283=>"110111110",
  15284=>"000000000",
  15285=>"000000000",
  15286=>"100000111",
  15287=>"000100000",
  15288=>"111111110",
  15289=>"100111111",
  15290=>"100110111",
  15291=>"110111011",
  15292=>"001011011",
  15293=>"000000111",
  15294=>"001011110",
  15295=>"000101111",
  15296=>"100100111",
  15297=>"000000000",
  15298=>"000000000",
  15299=>"111111111",
  15300=>"011011111",
  15301=>"100110111",
  15302=>"000000010",
  15303=>"000001110",
  15304=>"111011000",
  15305=>"000111111",
  15306=>"111110010",
  15307=>"000110110",
  15308=>"110000100",
  15309=>"011111001",
  15310=>"111111000",
  15311=>"110110000",
  15312=>"111000000",
  15313=>"111000000",
  15314=>"000110111",
  15315=>"111011111",
  15316=>"101101001",
  15317=>"000010110",
  15318=>"110100111",
  15319=>"111111111",
  15320=>"000000000",
  15321=>"000000010",
  15322=>"111010000",
  15323=>"111011000",
  15324=>"111111111",
  15325=>"111111011",
  15326=>"100111101",
  15327=>"001011111",
  15328=>"001001111",
  15329=>"110110000",
  15330=>"111111111",
  15331=>"110110111",
  15332=>"111111111",
  15333=>"111111110",
  15334=>"110111111",
  15335=>"111000000",
  15336=>"010010111",
  15337=>"110100000",
  15338=>"000000000",
  15339=>"111111000",
  15340=>"111101101",
  15341=>"011011010",
  15342=>"001001000",
  15343=>"001001111",
  15344=>"111111111",
  15345=>"000000000",
  15346=>"000000100",
  15347=>"001000000",
  15348=>"111001000",
  15349=>"100100111",
  15350=>"110110110",
  15351=>"000000000",
  15352=>"111000000",
  15353=>"110110000",
  15354=>"110111110",
  15355=>"111111101",
  15356=>"111111000",
  15357=>"000001001",
  15358=>"000100100",
  15359=>"011000100",
  15360=>"000000000",
  15361=>"111111001",
  15362=>"101001111",
  15363=>"000000100",
  15364=>"111111101",
  15365=>"000011111",
  15366=>"000000000",
  15367=>"111111111",
  15368=>"000000000",
  15369=>"110000000",
  15370=>"000000000",
  15371=>"000011000",
  15372=>"000111000",
  15373=>"000000000",
  15374=>"100000000",
  15375=>"110110111",
  15376=>"111001000",
  15377=>"010000111",
  15378=>"000000000",
  15379=>"111111011",
  15380=>"000011000",
  15381=>"111111111",
  15382=>"111111101",
  15383=>"000000000",
  15384=>"111110111",
  15385=>"111000000",
  15386=>"000001110",
  15387=>"111111111",
  15388=>"000000000",
  15389=>"111111001",
  15390=>"111000000",
  15391=>"111111001",
  15392=>"001001111",
  15393=>"111111100",
  15394=>"000000000",
  15395=>"111011011",
  15396=>"000000100",
  15397=>"000010000",
  15398=>"001101111",
  15399=>"111001000",
  15400=>"000000000",
  15401=>"001001111",
  15402=>"000000000",
  15403=>"111111111",
  15404=>"000000000",
  15405=>"000000001",
  15406=>"111111111",
  15407=>"011111010",
  15408=>"001011001",
  15409=>"000000000",
  15410=>"100100100",
  15411=>"111111111",
  15412=>"000000000",
  15413=>"100101111",
  15414=>"000000000",
  15415=>"000000000",
  15416=>"101101111",
  15417=>"111101001",
  15418=>"000000000",
  15419=>"000000000",
  15420=>"111001000",
  15421=>"000000000",
  15422=>"110110000",
  15423=>"111111111",
  15424=>"111101011",
  15425=>"111111110",
  15426=>"111000000",
  15427=>"000000000",
  15428=>"111111010",
  15429=>"111111111",
  15430=>"000000001",
  15431=>"111111111",
  15432=>"000000011",
  15433=>"111111110",
  15434=>"000000000",
  15435=>"000000000",
  15436=>"110111111",
  15437=>"000100110",
  15438=>"000000000",
  15439=>"001111111",
  15440=>"011111000",
  15441=>"010000000",
  15442=>"001101100",
  15443=>"101001111",
  15444=>"000000000",
  15445=>"000000000",
  15446=>"111111111",
  15447=>"111111111",
  15448=>"011011011",
  15449=>"000000000",
  15450=>"111111111",
  15451=>"111011111",
  15452=>"000000000",
  15453=>"011111111",
  15454=>"111111011",
  15455=>"100001011",
  15456=>"011111111",
  15457=>"000000000",
  15458=>"111100001",
  15459=>"000000000",
  15460=>"000000000",
  15461=>"111111111",
  15462=>"110110111",
  15463=>"000000000",
  15464=>"000000011",
  15465=>"111111011",
  15466=>"001000000",
  15467=>"000010001",
  15468=>"001000000",
  15469=>"111111111",
  15470=>"111000111",
  15471=>"110110110",
  15472=>"111111111",
  15473=>"111111111",
  15474=>"000000000",
  15475=>"100000011",
  15476=>"000000000",
  15477=>"111111110",
  15478=>"000000000",
  15479=>"111001111",
  15480=>"111101000",
  15481=>"101101111",
  15482=>"001000000",
  15483=>"001000000",
  15484=>"100000000",
  15485=>"000000000",
  15486=>"010111000",
  15487=>"111111111",
  15488=>"111111111",
  15489=>"111111000",
  15490=>"000011011",
  15491=>"100000000",
  15492=>"000000000",
  15493=>"111101001",
  15494=>"000101100",
  15495=>"000000000",
  15496=>"000000000",
  15497=>"111110110",
  15498=>"011001000",
  15499=>"000000000",
  15500=>"111111111",
  15501=>"110111111",
  15502=>"111111000",
  15503=>"000000000",
  15504=>"000010000",
  15505=>"111111111",
  15506=>"000110100",
  15507=>"100000000",
  15508=>"111000000",
  15509=>"110111101",
  15510=>"000000000",
  15511=>"000000000",
  15512=>"001000000",
  15513=>"111111111",
  15514=>"111111111",
  15515=>"111011011",
  15516=>"000110110",
  15517=>"100001001",
  15518=>"100110100",
  15519=>"000000000",
  15520=>"010111011",
  15521=>"111111111",
  15522=>"111111111",
  15523=>"111111111",
  15524=>"000100100",
  15525=>"110110110",
  15526=>"111001000",
  15527=>"000010111",
  15528=>"001000100",
  15529=>"000000000",
  15530=>"111000111",
  15531=>"000000000",
  15532=>"001000000",
  15533=>"100000111",
  15534=>"111111111",
  15535=>"000010000",
  15536=>"111111111",
  15537=>"111101011",
  15538=>"110111111",
  15539=>"111111100",
  15540=>"111111111",
  15541=>"000001001",
  15542=>"111111111",
  15543=>"000000000",
  15544=>"111111111",
  15545=>"000000010",
  15546=>"001111111",
  15547=>"001111100",
  15548=>"111111111",
  15549=>"100100000",
  15550=>"000000111",
  15551=>"110110111",
  15552=>"000100100",
  15553=>"111111111",
  15554=>"000000000",
  15555=>"000000001",
  15556=>"001010110",
  15557=>"100001000",
  15558=>"101111111",
  15559=>"000000100",
  15560=>"001001101",
  15561=>"101000000",
  15562=>"000100000",
  15563=>"011011011",
  15564=>"100100000",
  15565=>"000000100",
  15566=>"110000000",
  15567=>"111111011",
  15568=>"111110111",
  15569=>"000000000",
  15570=>"000000000",
  15571=>"000000000",
  15572=>"000000000",
  15573=>"000110000",
  15574=>"101000111",
  15575=>"000000001",
  15576=>"100111111",
  15577=>"111000000",
  15578=>"000111010",
  15579=>"000000000",
  15580=>"000000000",
  15581=>"100100100",
  15582=>"010000000",
  15583=>"000000010",
  15584=>"011111111",
  15585=>"011011111",
  15586=>"000111011",
  15587=>"000000000",
  15588=>"000000000",
  15589=>"100100100",
  15590=>"000000000",
  15591=>"111111111",
  15592=>"111111011",
  15593=>"101111111",
  15594=>"101001101",
  15595=>"000000000",
  15596=>"111111111",
  15597=>"001000000",
  15598=>"000000000",
  15599=>"000001000",
  15600=>"111100000",
  15601=>"000000000",
  15602=>"111111111",
  15603=>"000000001",
  15604=>"000000000",
  15605=>"111111111",
  15606=>"111100000",
  15607=>"111111111",
  15608=>"100000000",
  15609=>"000100100",
  15610=>"100100001",
  15611=>"000000100",
  15612=>"110100101",
  15613=>"000000000",
  15614=>"111111111",
  15615=>"000000000",
  15616=>"000000000",
  15617=>"101100100",
  15618=>"111111111",
  15619=>"001000000",
  15620=>"110110000",
  15621=>"111111111",
  15622=>"111111001",
  15623=>"111111111",
  15624=>"001001000",
  15625=>"011011001",
  15626=>"000000000",
  15627=>"110110100",
  15628=>"100000100",
  15629=>"000000100",
  15630=>"000000000",
  15631=>"000000000",
  15632=>"000001111",
  15633=>"000000000",
  15634=>"100100110",
  15635=>"100111001",
  15636=>"000000000",
  15637=>"111000111",
  15638=>"000000100",
  15639=>"000000000",
  15640=>"111111111",
  15641=>"110110111",
  15642=>"000100111",
  15643=>"000100110",
  15644=>"111111100",
  15645=>"000000111",
  15646=>"000010000",
  15647=>"000010000",
  15648=>"000000000",
  15649=>"000000001",
  15650=>"111111110",
  15651=>"100100110",
  15652=>"111001001",
  15653=>"000000011",
  15654=>"000000000",
  15655=>"000100000",
  15656=>"000100100",
  15657=>"111111010",
  15658=>"000110111",
  15659=>"000000000",
  15660=>"111111111",
  15661=>"111100100",
  15662=>"001011111",
  15663=>"100000001",
  15664=>"111111000",
  15665=>"111111111",
  15666=>"000000111",
  15667=>"111011010",
  15668=>"000000111",
  15669=>"000000100",
  15670=>"100100000",
  15671=>"111111111",
  15672=>"000000000",
  15673=>"000000000",
  15674=>"000000000",
  15675=>"111000000",
  15676=>"000000000",
  15677=>"000000000",
  15678=>"000001000",
  15679=>"101111000",
  15680=>"111111000",
  15681=>"000000000",
  15682=>"000001000",
  15683=>"000000000",
  15684=>"111000111",
  15685=>"000000000",
  15686=>"000000000",
  15687=>"110110010",
  15688=>"110100100",
  15689=>"000000000",
  15690=>"111111010",
  15691=>"000001111",
  15692=>"000000000",
  15693=>"111100111",
  15694=>"000000000",
  15695=>"110111001",
  15696=>"000101101",
  15697=>"111111111",
  15698=>"000000111",
  15699=>"111111111",
  15700=>"000000110",
  15701=>"000000000",
  15702=>"110000110",
  15703=>"110110000",
  15704=>"101111111",
  15705=>"111111011",
  15706=>"111000000",
  15707=>"000000000",
  15708=>"000001000",
  15709=>"000000000",
  15710=>"111111010",
  15711=>"111011111",
  15712=>"111111000",
  15713=>"011111111",
  15714=>"100000000",
  15715=>"000000000",
  15716=>"110100110",
  15717=>"101111110",
  15718=>"000000000",
  15719=>"101001001",
  15720=>"111111111",
  15721=>"001000000",
  15722=>"111100110",
  15723=>"111101001",
  15724=>"111101001",
  15725=>"111111111",
  15726=>"010111111",
  15727=>"111111011",
  15728=>"111111111",
  15729=>"000000000",
  15730=>"110000000",
  15731=>"111001100",
  15732=>"111111111",
  15733=>"000000000",
  15734=>"000000000",
  15735=>"011011011",
  15736=>"000000011",
  15737=>"111111000",
  15738=>"101111111",
  15739=>"000001101",
  15740=>"110010110",
  15741=>"111111111",
  15742=>"000001001",
  15743=>"000000000",
  15744=>"111111111",
  15745=>"111111111",
  15746=>"111111111",
  15747=>"000010000",
  15748=>"111111110",
  15749=>"011001111",
  15750=>"010000100",
  15751=>"111111111",
  15752=>"000000000",
  15753=>"101001001",
  15754=>"000011011",
  15755=>"011001011",
  15756=>"100000000",
  15757=>"111111111",
  15758=>"110111011",
  15759=>"001001011",
  15760=>"000000000",
  15761=>"111111111",
  15762=>"100000000",
  15763=>"000000000",
  15764=>"000000000",
  15765=>"000010010",
  15766=>"111001000",
  15767=>"000000000",
  15768=>"111001000",
  15769=>"111111111",
  15770=>"111111101",
  15771=>"011011000",
  15772=>"000000000",
  15773=>"001111111",
  15774=>"111111001",
  15775=>"011111110",
  15776=>"000010110",
  15777=>"111110111",
  15778=>"111111001",
  15779=>"000000000",
  15780=>"000000000",
  15781=>"111111010",
  15782=>"111111000",
  15783=>"000000000",
  15784=>"000000000",
  15785=>"111111011",
  15786=>"000000000",
  15787=>"100000000",
  15788=>"000000001",
  15789=>"000000000",
  15790=>"000111111",
  15791=>"111111111",
  15792=>"111001011",
  15793=>"000000100",
  15794=>"011011000",
  15795=>"111111111",
  15796=>"000110100",
  15797=>"000001000",
  15798=>"111110101",
  15799=>"101111111",
  15800=>"000000000",
  15801=>"101101100",
  15802=>"100100111",
  15803=>"000111101",
  15804=>"111111111",
  15805=>"100100001",
  15806=>"000000000",
  15807=>"101100101",
  15808=>"000000000",
  15809=>"101000000",
  15810=>"111111111",
  15811=>"000000000",
  15812=>"111111011",
  15813=>"100001000",
  15814=>"111111010",
  15815=>"010110100",
  15816=>"000000000",
  15817=>"000011111",
  15818=>"111010000",
  15819=>"000000000",
  15820=>"110000000",
  15821=>"101011111",
  15822=>"111101111",
  15823=>"111111111",
  15824=>"111001001",
  15825=>"000000000",
  15826=>"111111101",
  15827=>"000000000",
  15828=>"101000000",
  15829=>"000000000",
  15830=>"111001011",
  15831=>"011011111",
  15832=>"111101111",
  15833=>"000010000",
  15834=>"001000001",
  15835=>"111111111",
  15836=>"111111111",
  15837=>"011000000",
  15838=>"111100010",
  15839=>"001111111",
  15840=>"111001000",
  15841=>"111111111",
  15842=>"111111000",
  15843=>"010000000",
  15844=>"111111011",
  15845=>"010000000",
  15846=>"100110111",
  15847=>"010110110",
  15848=>"101111111",
  15849=>"010111111",
  15850=>"111001111",
  15851=>"111100100",
  15852=>"001001000",
  15853=>"000000000",
  15854=>"011001001",
  15855=>"111011001",
  15856=>"110110011",
  15857=>"100111111",
  15858=>"111111111",
  15859=>"111010110",
  15860=>"111111111",
  15861=>"001000100",
  15862=>"100000000",
  15863=>"101111010",
  15864=>"000000000",
  15865=>"100110100",
  15866=>"000000000",
  15867=>"000100100",
  15868=>"101111111",
  15869=>"001001100",
  15870=>"111111111",
  15871=>"111111111",
  15872=>"111011111",
  15873=>"111011100",
  15874=>"000000000",
  15875=>"001111111",
  15876=>"111000010",
  15877=>"100000101",
  15878=>"000000000",
  15879=>"001011111",
  15880=>"000000001",
  15881=>"111111000",
  15882=>"000000111",
  15883=>"111110000",
  15884=>"001111000",
  15885=>"000000000",
  15886=>"000000101",
  15887=>"000011111",
  15888=>"100111110",
  15889=>"000000001",
  15890=>"001100100",
  15891=>"100110110",
  15892=>"000000000",
  15893=>"000000000",
  15894=>"111110110",
  15895=>"001000000",
  15896=>"011010000",
  15897=>"000000110",
  15898=>"001110000",
  15899=>"000000000",
  15900=>"111111000",
  15901=>"111100000",
  15902=>"111001000",
  15903=>"111111000",
  15904=>"000000011",
  15905=>"111110110",
  15906=>"011111110",
  15907=>"000000000",
  15908=>"111111111",
  15909=>"000100111",
  15910=>"001000000",
  15911=>"111000000",
  15912=>"001010111",
  15913=>"000000000",
  15914=>"011111000",
  15915=>"111111111",
  15916=>"101000010",
  15917=>"000111111",
  15918=>"000000000",
  15919=>"000000000",
  15920=>"111111111",
  15921=>"000000011",
  15922=>"110110000",
  15923=>"100111001",
  15924=>"100111111",
  15925=>"101001001",
  15926=>"111111111",
  15927=>"111111010",
  15928=>"110111011",
  15929=>"111110000",
  15930=>"000011000",
  15931=>"111111111",
  15932=>"111111111",
  15933=>"111100000",
  15934=>"000110111",
  15935=>"101111110",
  15936=>"000000100",
  15937=>"111111001",
  15938=>"000000011",
  15939=>"111000000",
  15940=>"111111110",
  15941=>"001011110",
  15942=>"000000001",
  15943=>"111111000",
  15944=>"100000001",
  15945=>"001101111",
  15946=>"111111000",
  15947=>"111000001",
  15948=>"111111101",
  15949=>"100100111",
  15950=>"111000000",
  15951=>"000001110",
  15952=>"011000000",
  15953=>"000100000",
  15954=>"000001001",
  15955=>"000111111",
  15956=>"000101111",
  15957=>"000000000",
  15958=>"011111000",
  15959=>"000011011",
  15960=>"111111111",
  15961=>"001101111",
  15962=>"110000111",
  15963=>"110000000",
  15964=>"111111000",
  15965=>"111111100",
  15966=>"011011111",
  15967=>"100100100",
  15968=>"011000001",
  15969=>"000000000",
  15970=>"111111111",
  15971=>"000000000",
  15972=>"000110110",
  15973=>"111111111",
  15974=>"001111111",
  15975=>"000001111",
  15976=>"111001000",
  15977=>"111100000",
  15978=>"111010000",
  15979=>"000111111",
  15980=>"001011011",
  15981=>"001000111",
  15982=>"001001000",
  15983=>"010000000",
  15984=>"111111000",
  15985=>"111001111",
  15986=>"100111111",
  15987=>"001001011",
  15988=>"001101001",
  15989=>"000000110",
  15990=>"111000000",
  15991=>"000000000",
  15992=>"100000111",
  15993=>"101101100",
  15994=>"100110000",
  15995=>"111100100",
  15996=>"111111011",
  15997=>"111111110",
  15998=>"111111111",
  15999=>"000000000",
  16000=>"000000000",
  16001=>"000111111",
  16002=>"000000000",
  16003=>"000000001",
  16004=>"111000100",
  16005=>"100111111",
  16006=>"111011111",
  16007=>"000111011",
  16008=>"111111111",
  16009=>"100110000",
  16010=>"000000000",
  16011=>"000111111",
  16012=>"000000111",
  16013=>"000000001",
  16014=>"000100000",
  16015=>"111111111",
  16016=>"000000000",
  16017=>"000101111",
  16018=>"000111110",
  16019=>"000000000",
  16020=>"000111111",
  16021=>"101111101",
  16022=>"100000111",
  16023=>"111111111",
  16024=>"000000001",
  16025=>"000100111",
  16026=>"100000000",
  16027=>"111100000",
  16028=>"110110000",
  16029=>"111000000",
  16030=>"111000111",
  16031=>"111011001",
  16032=>"111011111",
  16033=>"001011111",
  16034=>"001001001",
  16035=>"111000000",
  16036=>"000001000",
  16037=>"011000001",
  16038=>"001111011",
  16039=>"011110111",
  16040=>"111111111",
  16041=>"000001111",
  16042=>"101000011",
  16043=>"111111000",
  16044=>"111111000",
  16045=>"110110100",
  16046=>"000000111",
  16047=>"000101000",
  16048=>"111100001",
  16049=>"000100100",
  16050=>"010111011",
  16051=>"111100000",
  16052=>"100110110",
  16053=>"111000000",
  16054=>"111001000",
  16055=>"110000011",
  16056=>"011011111",
  16057=>"000000111",
  16058=>"111100000",
  16059=>"011000001",
  16060=>"111111111",
  16061=>"010011111",
  16062=>"111111001",
  16063=>"000100101",
  16064=>"111111111",
  16065=>"111010000",
  16066=>"000111101",
  16067=>"000011111",
  16068=>"011000000",
  16069=>"000001111",
  16070=>"000000111",
  16071=>"111111111",
  16072=>"100000000",
  16073=>"110001111",
  16074=>"011000011",
  16075=>"100100100",
  16076=>"111000111",
  16077=>"111111111",
  16078=>"000000100",
  16079=>"000000001",
  16080=>"111011001",
  16081=>"011011111",
  16082=>"001101100",
  16083=>"101000000",
  16084=>"001001011",
  16085=>"101011001",
  16086=>"100100000",
  16087=>"000011011",
  16088=>"001101111",
  16089=>"110000000",
  16090=>"000000000",
  16091=>"111000000",
  16092=>"110110111",
  16093=>"000010000",
  16094=>"000101100",
  16095=>"110111111",
  16096=>"101100111",
  16097=>"100000111",
  16098=>"000000111",
  16099=>"111000000",
  16100=>"000100111",
  16101=>"011011110",
  16102=>"000110110",
  16103=>"000111111",
  16104=>"111000000",
  16105=>"001000000",
  16106=>"011011000",
  16107=>"111000011",
  16108=>"110000000",
  16109=>"111111110",
  16110=>"111010000",
  16111=>"111011001",
  16112=>"011000000",
  16113=>"000000000",
  16114=>"111111000",
  16115=>"111111100",
  16116=>"000000111",
  16117=>"000001001",
  16118=>"110110100",
  16119=>"000001111",
  16120=>"111111111",
  16121=>"000000001",
  16122=>"101000000",
  16123=>"001111111",
  16124=>"000001011",
  16125=>"001101110",
  16126=>"111111011",
  16127=>"111111110",
  16128=>"000000011",
  16129=>"011111111",
  16130=>"011111011",
  16131=>"000000000",
  16132=>"111001001",
  16133=>"011111000",
  16134=>"011100110",
  16135=>"100110100",
  16136=>"111111100",
  16137=>"100100000",
  16138=>"111000000",
  16139=>"101111111",
  16140=>"011001001",
  16141=>"000111111",
  16142=>"000101111",
  16143=>"111111011",
  16144=>"111010111",
  16145=>"111111110",
  16146=>"011001011",
  16147=>"110110100",
  16148=>"000000111",
  16149=>"111000011",
  16150=>"100110100",
  16151=>"000000000",
  16152=>"100110100",
  16153=>"000000111",
  16154=>"000111111",
  16155=>"111111111",
  16156=>"000111110",
  16157=>"111100111",
  16158=>"111011111",
  16159=>"000001111",
  16160=>"110000000",
  16161=>"111111101",
  16162=>"111111110",
  16163=>"000110111",
  16164=>"111011111",
  16165=>"111100100",
  16166=>"000111111",
  16167=>"111100000",
  16168=>"001001111",
  16169=>"111000000",
  16170=>"001001000",
  16171=>"111111100",
  16172=>"000000000",
  16173=>"000001000",
  16174=>"000000000",
  16175=>"000000111",
  16176=>"011011111",
  16177=>"001111111",
  16178=>"001111111",
  16179=>"000000111",
  16180=>"111111011",
  16181=>"111100100",
  16182=>"111101001",
  16183=>"111011010",
  16184=>"000111000",
  16185=>"111101111",
  16186=>"100100111",
  16187=>"111011000",
  16188=>"011000000",
  16189=>"111001000",
  16190=>"010000000",
  16191=>"000000000",
  16192=>"100000000",
  16193=>"111100000",
  16194=>"001000000",
  16195=>"000100111",
  16196=>"000111111",
  16197=>"010111111",
  16198=>"010000110",
  16199=>"111110111",
  16200=>"111111111",
  16201=>"111011000",
  16202=>"011011111",
  16203=>"111111111",
  16204=>"111111010",
  16205=>"000111111",
  16206=>"011011111",
  16207=>"011111111",
  16208=>"011001100",
  16209=>"110100100",
  16210=>"000101111",
  16211=>"111000000",
  16212=>"111111111",
  16213=>"001110000",
  16214=>"000000000",
  16215=>"101000111",
  16216=>"011000000",
  16217=>"101001111",
  16218=>"000000111",
  16219=>"100101111",
  16220=>"111000001",
  16221=>"000000000",
  16222=>"011001100",
  16223=>"100101111",
  16224=>"000100111",
  16225=>"000111111",
  16226=>"111111000",
  16227=>"100000111",
  16228=>"000100110",
  16229=>"111100000",
  16230=>"011000000",
  16231=>"001000000",
  16232=>"111110110",
  16233=>"000000000",
  16234=>"111111011",
  16235=>"100100000",
  16236=>"001001111",
  16237=>"100100111",
  16238=>"111001001",
  16239=>"111000000",
  16240=>"011011111",
  16241=>"100000000",
  16242=>"111111011",
  16243=>"000011011",
  16244=>"111111001",
  16245=>"111111111",
  16246=>"000001011",
  16247=>"000000000",
  16248=>"111111010",
  16249=>"000000111",
  16250=>"000000000",
  16251=>"111000000",
  16252=>"000111111",
  16253=>"000000111",
  16254=>"111111111",
  16255=>"111111011",
  16256=>"100000100",
  16257=>"000000000",
  16258=>"100000001",
  16259=>"011000000",
  16260=>"111111011",
  16261=>"000000000",
  16262=>"000000000",
  16263=>"110000000",
  16264=>"000000000",
  16265=>"000101111",
  16266=>"000000101",
  16267=>"001000000",
  16268=>"111111111",
  16269=>"000000100",
  16270=>"000000000",
  16271=>"000110111",
  16272=>"110111000",
  16273=>"111111111",
  16274=>"100111001",
  16275=>"000000100",
  16276=>"001111111",
  16277=>"000011011",
  16278=>"000000010",
  16279=>"100000000",
  16280=>"000000111",
  16281=>"000000000",
  16282=>"111000000",
  16283=>"111111000",
  16284=>"000000000",
  16285=>"000101001",
  16286=>"000110111",
  16287=>"000101111",
  16288=>"000000111",
  16289=>"000000001",
  16290=>"111111001",
  16291=>"111100001",
  16292=>"000000100",
  16293=>"001101111",
  16294=>"111011000",
  16295=>"000011111",
  16296=>"000000000",
  16297=>"000111111",
  16298=>"000000010",
  16299=>"101100111",
  16300=>"111111111",
  16301=>"011000100",
  16302=>"000000000",
  16303=>"111000011",
  16304=>"111110000",
  16305=>"100000000",
  16306=>"110010110",
  16307=>"011111111",
  16308=>"001000100",
  16309=>"000000000",
  16310=>"111111111",
  16311=>"000010011",
  16312=>"111000000",
  16313=>"111010000",
  16314=>"000000111",
  16315=>"000000000",
  16316=>"111001001",
  16317=>"111000001",
  16318=>"101101000",
  16319=>"110100001",
  16320=>"111111000",
  16321=>"000111000",
  16322=>"000000000",
  16323=>"111010000",
  16324=>"111111111",
  16325=>"111111000",
  16326=>"111000000",
  16327=>"100111111",
  16328=>"000000111",
  16329=>"000000000",
  16330=>"111000001",
  16331=>"110110000",
  16332=>"000000001",
  16333=>"001111111",
  16334=>"111011011",
  16335=>"111000000",
  16336=>"000000000",
  16337=>"111000110",
  16338=>"000000011",
  16339=>"111111111",
  16340=>"111110100",
  16341=>"000000000",
  16342=>"111111000",
  16343=>"100110000",
  16344=>"111111111",
  16345=>"000000000",
  16346=>"000111111",
  16347=>"011011010",
  16348=>"100110000",
  16349=>"111111111",
  16350=>"011001000",
  16351=>"111001001",
  16352=>"000000000",
  16353=>"011011111",
  16354=>"000111011",
  16355=>"111110111",
  16356=>"000111111",
  16357=>"110000000",
  16358=>"111011000",
  16359=>"001100101",
  16360=>"000000000",
  16361=>"111111111",
  16362=>"011010111",
  16363=>"000000111",
  16364=>"111111111",
  16365=>"001100100",
  16366=>"000111111",
  16367=>"111111111",
  16368=>"100100000",
  16369=>"111100100",
  16370=>"011000111",
  16371=>"110111111",
  16372=>"101100000",
  16373=>"000111111",
  16374=>"000001111",
  16375=>"110000010",
  16376=>"100111111",
  16377=>"001001111",
  16378=>"111001001",
  16379=>"111111111",
  16380=>"001001001",
  16381=>"011111111",
  16382=>"110000000",
  16383=>"000000100",
  16384=>"000000101",
  16385=>"111000000",
  16386=>"111000000",
  16387=>"000110110",
  16388=>"000000000",
  16389=>"001000001",
  16390=>"101001011",
  16391=>"000000101",
  16392=>"111000100",
  16393=>"000111111",
  16394=>"000000000",
  16395=>"101100000",
  16396=>"011111110",
  16397=>"111001000",
  16398=>"111111111",
  16399=>"111111111",
  16400=>"101001111",
  16401=>"000001111",
  16402=>"111100011",
  16403=>"101111111",
  16404=>"111111000",
  16405=>"110100100",
  16406=>"000000000",
  16407=>"110000000",
  16408=>"000001011",
  16409=>"000111111",
  16410=>"111110101",
  16411=>"100000000",
  16412=>"000100111",
  16413=>"101111111",
  16414=>"100111111",
  16415=>"111111101",
  16416=>"111111111",
  16417=>"111111110",
  16418=>"111111111",
  16419=>"111111110",
  16420=>"111101000",
  16421=>"111111111",
  16422=>"000000000",
  16423=>"101111100",
  16424=>"000000000",
  16425=>"111111011",
  16426=>"000000000",
  16427=>"111111000",
  16428=>"110111000",
  16429=>"000110000",
  16430=>"001101000",
  16431=>"100111111",
  16432=>"110111001",
  16433=>"000111111",
  16434=>"000100110",
  16435=>"111111111",
  16436=>"000100100",
  16437=>"011110110",
  16438=>"000000010",
  16439=>"000000010",
  16440=>"111111000",
  16441=>"110111100",
  16442=>"011111000",
  16443=>"010111111",
  16444=>"000000000",
  16445=>"000111011",
  16446=>"000000111",
  16447=>"011000001",
  16448=>"111111000",
  16449=>"110111100",
  16450=>"111111111",
  16451=>"011111000",
  16452=>"111111111",
  16453=>"111101111",
  16454=>"111111111",
  16455=>"111111111",
  16456=>"000000000",
  16457=>"001011111",
  16458=>"101100000",
  16459=>"001011111",
  16460=>"001001000",
  16461=>"111011011",
  16462=>"101111011",
  16463=>"001010110",
  16464=>"111000000",
  16465=>"001000000",
  16466=>"111111111",
  16467=>"100110000",
  16468=>"000001001",
  16469=>"110100100",
  16470=>"000110000",
  16471=>"001000000",
  16472=>"000100100",
  16473=>"100100100",
  16474=>"101000100",
  16475=>"111011110",
  16476=>"001000011",
  16477=>"110000100",
  16478=>"011111000",
  16479=>"000001001",
  16480=>"000000000",
  16481=>"111011001",
  16482=>"000000011",
  16483=>"111111111",
  16484=>"110100011",
  16485=>"101111111",
  16486=>"010011000",
  16487=>"111110000",
  16488=>"000000000",
  16489=>"100111111",
  16490=>"111000000",
  16491=>"000111111",
  16492=>"000000000",
  16493=>"111111111",
  16494=>"001000101",
  16495=>"101000111",
  16496=>"111111111",
  16497=>"111100110",
  16498=>"011111011",
  16499=>"111111111",
  16500=>"100000111",
  16501=>"111111000",
  16502=>"111111001",
  16503=>"000111001",
  16504=>"111011000",
  16505=>"111111000",
  16506=>"110100110",
  16507=>"111100100",
  16508=>"110111000",
  16509=>"001000111",
  16510=>"101110110",
  16511=>"000000000",
  16512=>"000000000",
  16513=>"101111111",
  16514=>"111001000",
  16515=>"111111011",
  16516=>"111111110",
  16517=>"000100111",
  16518=>"001000010",
  16519=>"111111111",
  16520=>"101011111",
  16521=>"101000000",
  16522=>"111111011",
  16523=>"000000111",
  16524=>"000000111",
  16525=>"000100000",
  16526=>"111111111",
  16527=>"111111100",
  16528=>"111111111",
  16529=>"000001111",
  16530=>"101100100",
  16531=>"111000000",
  16532=>"000000000",
  16533=>"001001000",
  16534=>"000000100",
  16535=>"111100100",
  16536=>"001000001",
  16537=>"111110000",
  16538=>"001000000",
  16539=>"111001100",
  16540=>"111100111",
  16541=>"001000001",
  16542=>"000000111",
  16543=>"111001001",
  16544=>"111011111",
  16545=>"000000000",
  16546=>"000111111",
  16547=>"100000000",
  16548=>"000011111",
  16549=>"011011011",
  16550=>"011000111",
  16551=>"011111011",
  16552=>"000000000",
  16553=>"111001000",
  16554=>"000000000",
  16555=>"000111111",
  16556=>"111110111",
  16557=>"010010000",
  16558=>"111000000",
  16559=>"111111101",
  16560=>"000000000",
  16561=>"111011011",
  16562=>"010111010",
  16563=>"000101111",
  16564=>"111000000",
  16565=>"000000001",
  16566=>"000111111",
  16567=>"111000000",
  16568=>"000100100",
  16569=>"011000111",
  16570=>"000000000",
  16571=>"001000000",
  16572=>"110111000",
  16573=>"001000100",
  16574=>"111111111",
  16575=>"101101111",
  16576=>"000000001",
  16577=>"111111110",
  16578=>"000000111",
  16579=>"111011001",
  16580=>"000000000",
  16581=>"111111000",
  16582=>"000010000",
  16583=>"000101111",
  16584=>"000000100",
  16585=>"111011001",
  16586=>"000000000",
  16587=>"111111011",
  16588=>"000000011",
  16589=>"001011100",
  16590=>"000010000",
  16591=>"001011100",
  16592=>"001000000",
  16593=>"111111111",
  16594=>"000101111",
  16595=>"100000011",
  16596=>"000110111",
  16597=>"111111110",
  16598=>"001001000",
  16599=>"000000000",
  16600=>"011011111",
  16601=>"011111000",
  16602=>"010011000",
  16603=>"111111111",
  16604=>"111001000",
  16605=>"000000000",
  16606=>"111111001",
  16607=>"000000111",
  16608=>"000000111",
  16609=>"111000000",
  16610=>"100110111",
  16611=>"111000111",
  16612=>"100111111",
  16613=>"111110111",
  16614=>"111111100",
  16615=>"100000000",
  16616=>"000000111",
  16617=>"001000101",
  16618=>"111011010",
  16619=>"111001001",
  16620=>"111111111",
  16621=>"100000000",
  16622=>"000111000",
  16623=>"111101100",
  16624=>"001000000",
  16625=>"001011111",
  16626=>"111111101",
  16627=>"101111110",
  16628=>"000000000",
  16629=>"000111111",
  16630=>"000001111",
  16631=>"000111111",
  16632=>"111111000",
  16633=>"000000000",
  16634=>"110110000",
  16635=>"001101000",
  16636=>"001000110",
  16637=>"000000111",
  16638=>"111000000",
  16639=>"111111110",
  16640=>"000011111",
  16641=>"010010011",
  16642=>"110111111",
  16643=>"111110111",
  16644=>"111111001",
  16645=>"000000000",
  16646=>"100100100",
  16647=>"001000000",
  16648=>"000100101",
  16649=>"000000011",
  16650=>"000000000",
  16651=>"111111000",
  16652=>"000010010",
  16653=>"111111111",
  16654=>"000111111",
  16655=>"100111101",
  16656=>"000000001",
  16657=>"001111111",
  16658=>"000000000",
  16659=>"111011111",
  16660=>"111000000",
  16661=>"011100100",
  16662=>"010111111",
  16663=>"111101000",
  16664=>"000001011",
  16665=>"000111111",
  16666=>"111011000",
  16667=>"001000110",
  16668=>"001001111",
  16669=>"111001111",
  16670=>"000000111",
  16671=>"111111111",
  16672=>"000100100",
  16673=>"000000101",
  16674=>"110111111",
  16675=>"000000000",
  16676=>"000000110",
  16677=>"111111011",
  16678=>"001011000",
  16679=>"100000001",
  16680=>"000110111",
  16681=>"111111111",
  16682=>"111000100",
  16683=>"110110111",
  16684=>"111111011",
  16685=>"000001011",
  16686=>"111111001",
  16687=>"110000000",
  16688=>"011001000",
  16689=>"001000000",
  16690=>"001111011",
  16691=>"000100111",
  16692=>"111111011",
  16693=>"000100100",
  16694=>"111010011",
  16695=>"000011001",
  16696=>"111011000",
  16697=>"111000000",
  16698=>"000111111",
  16699=>"000001001",
  16700=>"010000000",
  16701=>"010000000",
  16702=>"000111111",
  16703=>"111000000",
  16704=>"111110100",
  16705=>"111111000",
  16706=>"111111111",
  16707=>"000000000",
  16708=>"011111111",
  16709=>"100111011",
  16710=>"001001111",
  16711=>"100111111",
  16712=>"101111111",
  16713=>"111111011",
  16714=>"000000000",
  16715=>"011011000",
  16716=>"111100111",
  16717=>"111110100",
  16718=>"101111111",
  16719=>"000000100",
  16720=>"111110100",
  16721=>"000101111",
  16722=>"101101100",
  16723=>"011111010",
  16724=>"000000000",
  16725=>"000010011",
  16726=>"000000000",
  16727=>"001001000",
  16728=>"000001000",
  16729=>"111111111",
  16730=>"111111100",
  16731=>"100100001",
  16732=>"100101101",
  16733=>"000111111",
  16734=>"100001001",
  16735=>"111001111",
  16736=>"000000000",
  16737=>"111000000",
  16738=>"001101111",
  16739=>"000000000",
  16740=>"011111110",
  16741=>"001000000",
  16742=>"111000100",
  16743=>"111001000",
  16744=>"001111100",
  16745=>"100001000",
  16746=>"111110000",
  16747=>"010011001",
  16748=>"111111000",
  16749=>"000100100",
  16750=>"111111111",
  16751=>"011111111",
  16752=>"111111011",
  16753=>"000010000",
  16754=>"000000100",
  16755=>"000111111",
  16756=>"000000000",
  16757=>"111111000",
  16758=>"000110110",
  16759=>"111000111",
  16760=>"000000000",
  16761=>"111111110",
  16762=>"000000111",
  16763=>"100100100",
  16764=>"000101111",
  16765=>"111110000",
  16766=>"001101111",
  16767=>"111111110",
  16768=>"111011011",
  16769=>"110111111",
  16770=>"110000111",
  16771=>"000000101",
  16772=>"111100000",
  16773=>"000000001",
  16774=>"111111100",
  16775=>"011001111",
  16776=>"011011010",
  16777=>"011011000",
  16778=>"000000100",
  16779=>"000000000",
  16780=>"000000000",
  16781=>"000110010",
  16782=>"111111000",
  16783=>"111110000",
  16784=>"011001000",
  16785=>"011000000",
  16786=>"000000000",
  16787=>"111000000",
  16788=>"011111101",
  16789=>"000000000",
  16790=>"000000000",
  16791=>"001110110",
  16792=>"000111111",
  16793=>"000000000",
  16794=>"000000001",
  16795=>"100000110",
  16796=>"000110111",
  16797=>"111001000",
  16798=>"100000000",
  16799=>"100111111",
  16800=>"111111011",
  16801=>"000100100",
  16802=>"000000100",
  16803=>"101000000",
  16804=>"111111011",
  16805=>"000101000",
  16806=>"111000000",
  16807=>"000000011",
  16808=>"111001011",
  16809=>"000000000",
  16810=>"000000111",
  16811=>"000000111",
  16812=>"011000000",
  16813=>"111111111",
  16814=>"000111100",
  16815=>"001000000",
  16816=>"100000110",
  16817=>"000000000",
  16818=>"000000001",
  16819=>"111000000",
  16820=>"001101111",
  16821=>"111111000",
  16822=>"111111001",
  16823=>"111111111",
  16824=>"111000111",
  16825=>"001110111",
  16826=>"000000000",
  16827=>"100100101",
  16828=>"000100101",
  16829=>"011001011",
  16830=>"000000000",
  16831=>"111110000",
  16832=>"111011011",
  16833=>"000000000",
  16834=>"001001000",
  16835=>"000000000",
  16836=>"100111000",
  16837=>"100110110",
  16838=>"111010000",
  16839=>"000011001",
  16840=>"000000001",
  16841=>"111000111",
  16842=>"000000000",
  16843=>"011000000",
  16844=>"000110111",
  16845=>"110000000",
  16846=>"000000000",
  16847=>"111111111",
  16848=>"111000111",
  16849=>"110111011",
  16850=>"000001111",
  16851=>"000000011",
  16852=>"000110010",
  16853=>"000001000",
  16854=>"000000000",
  16855=>"000110011",
  16856=>"000001111",
  16857=>"100000111",
  16858=>"000111111",
  16859=>"000000000",
  16860=>"111011000",
  16861=>"101000000",
  16862=>"110100000",
  16863=>"001011011",
  16864=>"111011000",
  16865=>"001001101",
  16866=>"100111111",
  16867=>"000000010",
  16868=>"111110110",
  16869=>"000110100",
  16870=>"111111011",
  16871=>"000101101",
  16872=>"010011000",
  16873=>"111111111",
  16874=>"000011111",
  16875=>"011000000",
  16876=>"111111000",
  16877=>"000111100",
  16878=>"111111000",
  16879=>"000000000",
  16880=>"000101111",
  16881=>"011001011",
  16882=>"001000001",
  16883=>"111111111",
  16884=>"000110000",
  16885=>"111011011",
  16886=>"000000000",
  16887=>"000011011",
  16888=>"111111111",
  16889=>"110000000",
  16890=>"001001111",
  16891=>"100000001",
  16892=>"000100111",
  16893=>"111110100",
  16894=>"111011000",
  16895=>"000111111",
  16896=>"001001000",
  16897=>"000000111",
  16898=>"111111111",
  16899=>"000000111",
  16900=>"011000000",
  16901=>"100000000",
  16902=>"001000000",
  16903=>"111111111",
  16904=>"000000001",
  16905=>"000000110",
  16906=>"111111111",
  16907=>"011111111",
  16908=>"111100111",
  16909=>"011111111",
  16910=>"011010110",
  16911=>"000000000",
  16912=>"000000000",
  16913=>"111011111",
  16914=>"001000000",
  16915=>"000000000",
  16916=>"110111111",
  16917=>"000000000",
  16918=>"000001001",
  16919=>"000000000",
  16920=>"111111110",
  16921=>"100001001",
  16922=>"111001100",
  16923=>"001001001",
  16924=>"011000000",
  16925=>"101111001",
  16926=>"111110100",
  16927=>"111111111",
  16928=>"000000000",
  16929=>"001000010",
  16930=>"001001111",
  16931=>"110100000",
  16932=>"111100000",
  16933=>"000000000",
  16934=>"111111111",
  16935=>"100000000",
  16936=>"111011011",
  16937=>"000000000",
  16938=>"100101101",
  16939=>"111110111",
  16940=>"111111110",
  16941=>"110000000",
  16942=>"000000110",
  16943=>"110001001",
  16944=>"111000000",
  16945=>"110000000",
  16946=>"111111111",
  16947=>"000000111",
  16948=>"100110100",
  16949=>"000000100",
  16950=>"000000000",
  16951=>"000000100",
  16952=>"111111111",
  16953=>"100000000",
  16954=>"000011011",
  16955=>"111111000",
  16956=>"110100000",
  16957=>"111000000",
  16958=>"111111111",
  16959=>"111111111",
  16960=>"001000000",
  16961=>"010110000",
  16962=>"111111111",
  16963=>"000000111",
  16964=>"000000000",
  16965=>"000000000",
  16966=>"000000111",
  16967=>"111111111",
  16968=>"000000000",
  16969=>"000110110",
  16970=>"110000111",
  16971=>"101000111",
  16972=>"111111111",
  16973=>"110110111",
  16974=>"000000000",
  16975=>"010110000",
  16976=>"000110110",
  16977=>"001000110",
  16978=>"000000000",
  16979=>"100100100",
  16980=>"000011111",
  16981=>"111000000",
  16982=>"001000000",
  16983=>"110111111",
  16984=>"111100000",
  16985=>"000000101",
  16986=>"110000110",
  16987=>"001001000",
  16988=>"000000000",
  16989=>"111011000",
  16990=>"000000000",
  16991=>"111111011",
  16992=>"000000000",
  16993=>"111111000",
  16994=>"100010010",
  16995=>"111111111",
  16996=>"000000000",
  16997=>"101111111",
  16998=>"111111111",
  16999=>"111111111",
  17000=>"000100111",
  17001=>"000111111",
  17002=>"010010010",
  17003=>"111110000",
  17004=>"010011000",
  17005=>"000010111",
  17006=>"000000010",
  17007=>"000000000",
  17008=>"000000010",
  17009=>"000000111",
  17010=>"101100110",
  17011=>"111111000",
  17012=>"000000000",
  17013=>"111111000",
  17014=>"000000111",
  17015=>"011111011",
  17016=>"111111111",
  17017=>"000000000",
  17018=>"111111011",
  17019=>"111111111",
  17020=>"100100000",
  17021=>"000000000",
  17022=>"111111111",
  17023=>"011111010",
  17024=>"110111111",
  17025=>"111111010",
  17026=>"010110111",
  17027=>"000000000",
  17028=>"000001111",
  17029=>"111110110",
  17030=>"000000000",
  17031=>"111111111",
  17032=>"100000000",
  17033=>"111111011",
  17034=>"000000000",
  17035=>"000000000",
  17036=>"000000000",
  17037=>"011111110",
  17038=>"111111110",
  17039=>"010110010",
  17040=>"001000000",
  17041=>"000010000",
  17042=>"111111111",
  17043=>"011101111",
  17044=>"000000000",
  17045=>"000111111",
  17046=>"001000001",
  17047=>"000000110",
  17048=>"011111111",
  17049=>"000001001",
  17050=>"111110011",
  17051=>"000000000",
  17052=>"000000000",
  17053=>"100000000",
  17054=>"000000000",
  17055=>"111111111",
  17056=>"010000000",
  17057=>"111111111",
  17058=>"111001001",
  17059=>"110100111",
  17060=>"111001011",
  17061=>"111000111",
  17062=>"111111110",
  17063=>"011111110",
  17064=>"001000000",
  17065=>"101111111",
  17066=>"000001001",
  17067=>"110001000",
  17068=>"011000001",
  17069=>"000011110",
  17070=>"100001001",
  17071=>"000110111",
  17072=>"000010000",
  17073=>"000100110",
  17074=>"100000110",
  17075=>"111100100",
  17076=>"111000000",
  17077=>"111011010",
  17078=>"111111000",
  17079=>"001000000",
  17080=>"111111111",
  17081=>"111111111",
  17082=>"111111011",
  17083=>"100000110",
  17084=>"111111111",
  17085=>"101111111",
  17086=>"111000101",
  17087=>"000000000",
  17088=>"111111111",
  17089=>"111011111",
  17090=>"000000000",
  17091=>"000000000",
  17092=>"111111010",
  17093=>"000000000",
  17094=>"101011111",
  17095=>"000000000",
  17096=>"000110110",
  17097=>"000001111",
  17098=>"111110110",
  17099=>"000010000",
  17100=>"000001111",
  17101=>"001101100",
  17102=>"000010110",
  17103=>"000000000",
  17104=>"111111111",
  17105=>"000000000",
  17106=>"011001001",
  17107=>"000000000",
  17108=>"001000000",
  17109=>"111111111",
  17110=>"111111000",
  17111=>"000001000",
  17112=>"000000010",
  17113=>"111111111",
  17114=>"000000000",
  17115=>"011000011",
  17116=>"111111111",
  17117=>"111111111",
  17118=>"111111011",
  17119=>"111011011",
  17120=>"000000000",
  17121=>"000001000",
  17122=>"000000111",
  17123=>"001000000",
  17124=>"111100111",
  17125=>"000100100",
  17126=>"111111111",
  17127=>"111111111",
  17128=>"111111111",
  17129=>"000000000",
  17130=>"000000111",
  17131=>"111111111",
  17132=>"000111111",
  17133=>"110110111",
  17134=>"111111111",
  17135=>"000000000",
  17136=>"000111100",
  17137=>"111111111",
  17138=>"111111000",
  17139=>"100110100",
  17140=>"000000000",
  17141=>"001101100",
  17142=>"001101001",
  17143=>"000000000",
  17144=>"111101101",
  17145=>"000000000",
  17146=>"111011011",
  17147=>"000000000",
  17148=>"100110110",
  17149=>"000100111",
  17150=>"111000000",
  17151=>"111111001",
  17152=>"000000000",
  17153=>"001011011",
  17154=>"000000111",
  17155=>"001000000",
  17156=>"111111111",
  17157=>"001000010",
  17158=>"100000000",
  17159=>"000000000",
  17160=>"000000000",
  17161=>"000000100",
  17162=>"000100110",
  17163=>"001011011",
  17164=>"111111111",
  17165=>"000000000",
  17166=>"001000000",
  17167=>"110111101",
  17168=>"011111111",
  17169=>"110100111",
  17170=>"110000000",
  17171=>"111101111",
  17172=>"011011000",
  17173=>"001111111",
  17174=>"001001000",
  17175=>"111011111",
  17176=>"010000000",
  17177=>"000000000",
  17178=>"111111111",
  17179=>"011111111",
  17180=>"001001001",
  17181=>"111001000",
  17182=>"001011111",
  17183=>"110111011",
  17184=>"110110000",
  17185=>"111111111",
  17186=>"111111011",
  17187=>"000000000",
  17188=>"111111111",
  17189=>"000111111",
  17190=>"000010111",
  17191=>"101000110",
  17192=>"111111111",
  17193=>"000000000",
  17194=>"100100110",
  17195=>"000110110",
  17196=>"000101111",
  17197=>"000000000",
  17198=>"111000100",
  17199=>"000000000",
  17200=>"100001001",
  17201=>"010110111",
  17202=>"110111111",
  17203=>"010000000",
  17204=>"000000000",
  17205=>"000000000",
  17206=>"010111110",
  17207=>"000100100",
  17208=>"000000000",
  17209=>"000000000",
  17210=>"111111111",
  17211=>"111110111",
  17212=>"111111111",
  17213=>"111111111",
  17214=>"111111111",
  17215=>"111111111",
  17216=>"001000000",
  17217=>"111111111",
  17218=>"000000111",
  17219=>"000000000",
  17220=>"000000000",
  17221=>"000000000",
  17222=>"001000001",
  17223=>"111111110",
  17224=>"111101111",
  17225=>"000000111",
  17226=>"000000110",
  17227=>"010111111",
  17228=>"100100100",
  17229=>"000000000",
  17230=>"001111101",
  17231=>"111100100",
  17232=>"111111101",
  17233=>"111111111",
  17234=>"110110111",
  17235=>"111111111",
  17236=>"111000000",
  17237=>"001001011",
  17238=>"000000000",
  17239=>"110100111",
  17240=>"001000000",
  17241=>"000000101",
  17242=>"000000001",
  17243=>"011000000",
  17244=>"000000000",
  17245=>"111111111",
  17246=>"000001110",
  17247=>"000000000",
  17248=>"011111111",
  17249=>"000000001",
  17250=>"001001111",
  17251=>"000000000",
  17252=>"110110110",
  17253=>"000001011",
  17254=>"111111111",
  17255=>"000010010",
  17256=>"111101000",
  17257=>"000000000",
  17258=>"111111111",
  17259=>"000000000",
  17260=>"000000000",
  17261=>"100100000",
  17262=>"000011111",
  17263=>"111110100",
  17264=>"000000000",
  17265=>"101001001",
  17266=>"000000111",
  17267=>"111111111",
  17268=>"000000000",
  17269=>"001001011",
  17270=>"111111111",
  17271=>"000000000",
  17272=>"111111111",
  17273=>"000100000",
  17274=>"000000000",
  17275=>"000000000",
  17276=>"111111111",
  17277=>"000000000",
  17278=>"010011011",
  17279=>"000000000",
  17280=>"111110100",
  17281=>"000010010",
  17282=>"000000000",
  17283=>"001000000",
  17284=>"111111111",
  17285=>"000000001",
  17286=>"000000000",
  17287=>"000000010",
  17288=>"010111111",
  17289=>"000000000",
  17290=>"111001000",
  17291=>"111111111",
  17292=>"111111111",
  17293=>"000000100",
  17294=>"111000011",
  17295=>"000000000",
  17296=>"000000100",
  17297=>"000000000",
  17298=>"000011111",
  17299=>"011011011",
  17300=>"000000000",
  17301=>"010111000",
  17302=>"111011111",
  17303=>"011010100",
  17304=>"101000000",
  17305=>"001001001",
  17306=>"000011111",
  17307=>"111111111",
  17308=>"100111111",
  17309=>"100000100",
  17310=>"001000000",
  17311=>"011001001",
  17312=>"111001000",
  17313=>"000000111",
  17314=>"000000000",
  17315=>"111111111",
  17316=>"011111111",
  17317=>"011010000",
  17318=>"111111111",
  17319=>"111011001",
  17320=>"111100000",
  17321=>"000111111",
  17322=>"000000000",
  17323=>"001000000",
  17324=>"000000000",
  17325=>"100000000",
  17326=>"111101001",
  17327=>"010111111",
  17328=>"010000110",
  17329=>"000111100",
  17330=>"110111111",
  17331=>"000000000",
  17332=>"110111111",
  17333=>"111111111",
  17334=>"000000001",
  17335=>"000100000",
  17336=>"000000111",
  17337=>"110100000",
  17338=>"000000000",
  17339=>"000000000",
  17340=>"000000001",
  17341=>"000000111",
  17342=>"111111111",
  17343=>"001000010",
  17344=>"111111111",
  17345=>"111111111",
  17346=>"111111111",
  17347=>"111100000",
  17348=>"000000001",
  17349=>"111111000",
  17350=>"011011000",
  17351=>"111001001",
  17352=>"100000000",
  17353=>"011000000",
  17354=>"000000111",
  17355=>"110000000",
  17356=>"100000000",
  17357=>"111111111",
  17358=>"000000001",
  17359=>"111111111",
  17360=>"000000000",
  17361=>"001001000",
  17362=>"000000100",
  17363=>"001000000",
  17364=>"000000000",
  17365=>"011000101",
  17366=>"010000011",
  17367=>"011011011",
  17368=>"000000000",
  17369=>"000010010",
  17370=>"100110111",
  17371=>"111010000",
  17372=>"100100110",
  17373=>"111011000",
  17374=>"111111111",
  17375=>"111111110",
  17376=>"111110110",
  17377=>"000000000",
  17378=>"000000000",
  17379=>"000000100",
  17380=>"101101111",
  17381=>"111111101",
  17382=>"001111000",
  17383=>"100000111",
  17384=>"000000000",
  17385=>"111111111",
  17386=>"000000000",
  17387=>"111111111",
  17388=>"111111111",
  17389=>"000100100",
  17390=>"000010010",
  17391=>"000000000",
  17392=>"111100000",
  17393=>"000000110",
  17394=>"111111001",
  17395=>"001110110",
  17396=>"000000000",
  17397=>"000100000",
  17398=>"111111111",
  17399=>"000010111",
  17400=>"111111000",
  17401=>"100101001",
  17402=>"111111111",
  17403=>"000000000",
  17404=>"000000000",
  17405=>"000000001",
  17406=>"000000000",
  17407=>"001000000",
  17408=>"111111111",
  17409=>"111010000",
  17410=>"000000000",
  17411=>"000001100",
  17412=>"000000000",
  17413=>"111111111",
  17414=>"001001000",
  17415=>"100000111",
  17416=>"111011011",
  17417=>"111011001",
  17418=>"000011001",
  17419=>"111001100",
  17420=>"000100100",
  17421=>"111001100",
  17422=>"100101111",
  17423=>"010000000",
  17424=>"000111011",
  17425=>"000111111",
  17426=>"000000000",
  17427=>"000000000",
  17428=>"111011000",
  17429=>"000000000",
  17430=>"011111111",
  17431=>"010000011",
  17432=>"110000000",
  17433=>"111100000",
  17434=>"110011110",
  17435=>"011011111",
  17436=>"111101111",
  17437=>"111100000",
  17438=>"000000011",
  17439=>"000000000",
  17440=>"111111111",
  17441=>"110010111",
  17442=>"110111111",
  17443=>"111100111",
  17444=>"000011010",
  17445=>"001001000",
  17446=>"000000000",
  17447=>"011011001",
  17448=>"100000001",
  17449=>"000010111",
  17450=>"111111111",
  17451=>"000010111",
  17452=>"000000000",
  17453=>"000111111",
  17454=>"001011000",
  17455=>"111111111",
  17456=>"110110100",
  17457=>"000000000",
  17458=>"000000010",
  17459=>"000000000",
  17460=>"110111111",
  17461=>"111111010",
  17462=>"000101111",
  17463=>"000000000",
  17464=>"000001111",
  17465=>"101111111",
  17466=>"000000000",
  17467=>"000000111",
  17468=>"111100111",
  17469=>"000000101",
  17470=>"000111111",
  17471=>"111000000",
  17472=>"011111111",
  17473=>"000100011",
  17474=>"011111000",
  17475=>"000000111",
  17476=>"001001000",
  17477=>"111111111",
  17478=>"010000100",
  17479=>"000000000",
  17480=>"111111111",
  17481=>"111111111",
  17482=>"111111101",
  17483=>"111000110",
  17484=>"110101101",
  17485=>"000000000",
  17486=>"000000000",
  17487=>"000111111",
  17488=>"000111111",
  17489=>"111100101",
  17490=>"011011000",
  17491=>"011011000",
  17492=>"011000000",
  17493=>"010000000",
  17494=>"111000000",
  17495=>"111111111",
  17496=>"000000000",
  17497=>"111111111",
  17498=>"000000000",
  17499=>"011111011",
  17500=>"100101111",
  17501=>"000010111",
  17502=>"100000110",
  17503=>"000001001",
  17504=>"111111000",
  17505=>"110000000",
  17506=>"110111111",
  17507=>"111111011",
  17508=>"001011111",
  17509=>"011011000",
  17510=>"000000111",
  17511=>"000000110",
  17512=>"100100111",
  17513=>"000010111",
  17514=>"111111110",
  17515=>"000000100",
  17516=>"111111111",
  17517=>"000000000",
  17518=>"111100111",
  17519=>"000011111",
  17520=>"000000000",
  17521=>"000101111",
  17522=>"011111001",
  17523=>"100000000",
  17524=>"000000000",
  17525=>"000000000",
  17526=>"011001000",
  17527=>"000111111",
  17528=>"110111111",
  17529=>"101111000",
  17530=>"000000000",
  17531=>"111100111",
  17532=>"111111101",
  17533=>"001111111",
  17534=>"001001000",
  17535=>"000000000",
  17536=>"000000000",
  17537=>"000000000",
  17538=>"111111111",
  17539=>"000001001",
  17540=>"111111111",
  17541=>"000000000",
  17542=>"000000111",
  17543=>"110000111",
  17544=>"111000000",
  17545=>"111101111",
  17546=>"000000000",
  17547=>"111011011",
  17548=>"010111111",
  17549=>"100111111",
  17550=>"111111111",
  17551=>"111111111",
  17552=>"111111011",
  17553=>"111000000",
  17554=>"111000000",
  17555=>"000000000",
  17556=>"000110100",
  17557=>"010111110",
  17558=>"111111111",
  17559=>"111110000",
  17560=>"111111000",
  17561=>"111111011",
  17562=>"111111011",
  17563=>"000000000",
  17564=>"000000001",
  17565=>"000000000",
  17566=>"111111111",
  17567=>"000000000",
  17568=>"111111000",
  17569=>"111100100",
  17570=>"010000000",
  17571=>"000001000",
  17572=>"000000000",
  17573=>"111111000",
  17574=>"010000000",
  17575=>"111110110",
  17576=>"111100000",
  17577=>"100000000",
  17578=>"000000000",
  17579=>"111101111",
  17580=>"001001001",
  17581=>"111111100",
  17582=>"001100110",
  17583=>"000011011",
  17584=>"000000000",
  17585=>"000000000",
  17586=>"111111111",
  17587=>"111111101",
  17588=>"111100101",
  17589=>"111111111",
  17590=>"011111111",
  17591=>"111111011",
  17592=>"000000000",
  17593=>"111110111",
  17594=>"000000001",
  17595=>"000000100",
  17596=>"000000111",
  17597=>"111010000",
  17598=>"111111111",
  17599=>"011111110",
  17600=>"011111111",
  17601=>"001011011",
  17602=>"000000000",
  17603=>"000000000",
  17604=>"111111000",
  17605=>"111111111",
  17606=>"010000111",
  17607=>"000111111",
  17608=>"000000000",
  17609=>"111111100",
  17610=>"001000101",
  17611=>"000000100",
  17612=>"000000100",
  17613=>"000000000",
  17614=>"000000111",
  17615=>"000000000",
  17616=>"000000000",
  17617=>"010001111",
  17618=>"011111111",
  17619=>"000000000",
  17620=>"000000000",
  17621=>"000001000",
  17622=>"100000000",
  17623=>"000100111",
  17624=>"000001111",
  17625=>"110010000",
  17626=>"000000101",
  17627=>"001001000",
  17628=>"111001111",
  17629=>"111111101",
  17630=>"000000000",
  17631=>"110000000",
  17632=>"001001001",
  17633=>"001010111",
  17634=>"000111111",
  17635=>"111000000",
  17636=>"111000000",
  17637=>"000000000",
  17638=>"111111110",
  17639=>"111000000",
  17640=>"111111111",
  17641=>"000001111",
  17642=>"111011111",
  17643=>"110000111",
  17644=>"000111111",
  17645=>"001111110",
  17646=>"111111111",
  17647=>"111111101",
  17648=>"000000000",
  17649=>"111111111",
  17650=>"001000000",
  17651=>"001001111",
  17652=>"000000011",
  17653=>"110110000",
  17654=>"001000001",
  17655=>"000000111",
  17656=>"111111010",
  17657=>"000000000",
  17658=>"001000000",
  17659=>"001111111",
  17660=>"011011000",
  17661=>"000000010",
  17662=>"000000111",
  17663=>"000000000",
  17664=>"000000000",
  17665=>"011111101",
  17666=>"111001000",
  17667=>"011000000",
  17668=>"011011111",
  17669=>"100000110",
  17670=>"000000000",
  17671=>"111001011",
  17672=>"011111111",
  17673=>"000000111",
  17674=>"000001111",
  17675=>"111111111",
  17676=>"001001111",
  17677=>"001000000",
  17678=>"101001101",
  17679=>"100010000",
  17680=>"000000111",
  17681=>"000000000",
  17682=>"111011000",
  17683=>"101111111",
  17684=>"011111111",
  17685=>"111111000",
  17686=>"110111110",
  17687=>"111111110",
  17688=>"111101000",
  17689=>"100111111",
  17690=>"111111000",
  17691=>"000000100",
  17692=>"000110111",
  17693=>"000000000",
  17694=>"010111111",
  17695=>"111111111",
  17696=>"110110000",
  17697=>"111011000",
  17698=>"100110110",
  17699=>"111111111",
  17700=>"101100000",
  17701=>"000000000",
  17702=>"000000000",
  17703=>"111111001",
  17704=>"000000000",
  17705=>"000001111",
  17706=>"000100000",
  17707=>"000111100",
  17708=>"000000000",
  17709=>"111111001",
  17710=>"000001001",
  17711=>"000000000",
  17712=>"000000111",
  17713=>"000000001",
  17714=>"000000100",
  17715=>"000000000",
  17716=>"000000110",
  17717=>"000111111",
  17718=>"111010111",
  17719=>"111111000",
  17720=>"000000000",
  17721=>"000000001",
  17722=>"111000000",
  17723=>"000010111",
  17724=>"111111111",
  17725=>"111111111",
  17726=>"110111110",
  17727=>"000000101",
  17728=>"111001000",
  17729=>"111111000",
  17730=>"010010011",
  17731=>"110110000",
  17732=>"000000000",
  17733=>"111110111",
  17734=>"011100110",
  17735=>"111111111",
  17736=>"011111111",
  17737=>"000000111",
  17738=>"000000000",
  17739=>"111111111",
  17740=>"000000001",
  17741=>"000000111",
  17742=>"110000100",
  17743=>"110111110",
  17744=>"110111110",
  17745=>"000000101",
  17746=>"110100000",
  17747=>"000111111",
  17748=>"000000000",
  17749=>"001000011",
  17750=>"111111111",
  17751=>"111101111",
  17752=>"111111111",
  17753=>"000000000",
  17754=>"111100000",
  17755=>"011111111",
  17756=>"111111101",
  17757=>"010000111",
  17758=>"111000010",
  17759=>"001011111",
  17760=>"111111111",
  17761=>"111111111",
  17762=>"010000111",
  17763=>"000000111",
  17764=>"100100110",
  17765=>"000000101",
  17766=>"111111111",
  17767=>"110110000",
  17768=>"111111111",
  17769=>"111111000",
  17770=>"000000110",
  17771=>"110000000",
  17772=>"000000111",
  17773=>"000000110",
  17774=>"111111111",
  17775=>"111111111",
  17776=>"000110111",
  17777=>"111110110",
  17778=>"100100111",
  17779=>"111001000",
  17780=>"000000000",
  17781=>"011011111",
  17782=>"110000000",
  17783=>"000000000",
  17784=>"000000000",
  17785=>"001000000",
  17786=>"110000000",
  17787=>"111101111",
  17788=>"000100011",
  17789=>"111111111",
  17790=>"111110100",
  17791=>"000000111",
  17792=>"110110110",
  17793=>"110111111",
  17794=>"111111111",
  17795=>"111111111",
  17796=>"100111111",
  17797=>"000001111",
  17798=>"000000000",
  17799=>"000110100",
  17800=>"000000001",
  17801=>"111111111",
  17802=>"000010000",
  17803=>"111111010",
  17804=>"111100111",
  17805=>"111100100",
  17806=>"110110111",
  17807=>"001111111",
  17808=>"000000000",
  17809=>"100000111",
  17810=>"101111111",
  17811=>"111111111",
  17812=>"000000000",
  17813=>"000000000",
  17814=>"111000100",
  17815=>"011001000",
  17816=>"111000000",
  17817=>"001001001",
  17818=>"000000011",
  17819=>"001101111",
  17820=>"111111111",
  17821=>"111111110",
  17822=>"000000000",
  17823=>"100111111",
  17824=>"000000111",
  17825=>"111011011",
  17826=>"011101100",
  17827=>"111111011",
  17828=>"111100111",
  17829=>"000000000",
  17830=>"000000111",
  17831=>"111111111",
  17832=>"100111111",
  17833=>"010111111",
  17834=>"111001001",
  17835=>"110000011",
  17836=>"000000000",
  17837=>"001011000",
  17838=>"111110100",
  17839=>"000000100",
  17840=>"111111001",
  17841=>"000000000",
  17842=>"000000000",
  17843=>"111111111",
  17844=>"000000000",
  17845=>"111000000",
  17846=>"111111111",
  17847=>"000000000",
  17848=>"111101100",
  17849=>"111111100",
  17850=>"100111100",
  17851=>"111011001",
  17852=>"000000000",
  17853=>"111111111",
  17854=>"000000000",
  17855=>"110111100",
  17856=>"111111111",
  17857=>"000000111",
  17858=>"000000111",
  17859=>"111111111",
  17860=>"000000111",
  17861=>"111001001",
  17862=>"111111110",
  17863=>"000000011",
  17864=>"011111111",
  17865=>"000000000",
  17866=>"111111111",
  17867=>"011111001",
  17868=>"111001001",
  17869=>"000101111",
  17870=>"111011000",
  17871=>"000000000",
  17872=>"101100001",
  17873=>"111001111",
  17874=>"000000000",
  17875=>"000000110",
  17876=>"100100110",
  17877=>"101111111",
  17878=>"111000000",
  17879=>"000001011",
  17880=>"101101000",
  17881=>"111000000",
  17882=>"000000110",
  17883=>"111111111",
  17884=>"011001011",
  17885=>"011000000",
  17886=>"000000011",
  17887=>"111111110",
  17888=>"000000001",
  17889=>"000000000",
  17890=>"000000000",
  17891=>"111111111",
  17892=>"111111111",
  17893=>"111111000",
  17894=>"000010000",
  17895=>"000000000",
  17896=>"011011001",
  17897=>"111111000",
  17898=>"100000000",
  17899=>"101111111",
  17900=>"000000111",
  17901=>"000000000",
  17902=>"101001000",
  17903=>"111111111",
  17904=>"000000000",
  17905=>"001000111",
  17906=>"111111011",
  17907=>"000010011",
  17908=>"111101001",
  17909=>"001000000",
  17910=>"000000000",
  17911=>"001101111",
  17912=>"000000000",
  17913=>"011111011",
  17914=>"111111111",
  17915=>"111111111",
  17916=>"000000000",
  17917=>"000001000",
  17918=>"111101101",
  17919=>"000111011",
  17920=>"111111111",
  17921=>"000000111",
  17922=>"001000001",
  17923=>"000000000",
  17924=>"011011000",
  17925=>"110100101",
  17926=>"001001000",
  17927=>"111111111",
  17928=>"010000111",
  17929=>"111111111",
  17930=>"001001001",
  17931=>"000000000",
  17932=>"010000011",
  17933=>"111000000",
  17934=>"111111011",
  17935=>"000110111",
  17936=>"000000000",
  17937=>"000000001",
  17938=>"000000100",
  17939=>"111111111",
  17940=>"111111111",
  17941=>"000111111",
  17942=>"000000000",
  17943=>"100100000",
  17944=>"000000000",
  17945=>"000000000",
  17946=>"100100100",
  17947=>"100110111",
  17948=>"000000000",
  17949=>"100101111",
  17950=>"000000000",
  17951=>"101111111",
  17952=>"111111101",
  17953=>"000000000",
  17954=>"001011111",
  17955=>"011111011",
  17956=>"110111111",
  17957=>"000110111",
  17958=>"111111110",
  17959=>"111111000",
  17960=>"000100000",
  17961=>"000000000",
  17962=>"000100111",
  17963=>"111000000",
  17964=>"011110110",
  17965=>"000000000",
  17966=>"011111111",
  17967=>"011111111",
  17968=>"100111111",
  17969=>"001001000",
  17970=>"111110100",
  17971=>"111111111",
  17972=>"110110000",
  17973=>"100100000",
  17974=>"011111111",
  17975=>"111111000",
  17976=>"101111111",
  17977=>"101111000",
  17978=>"111111111",
  17979=>"000011011",
  17980=>"000000000",
  17981=>"111111111",
  17982=>"111111111",
  17983=>"111111111",
  17984=>"111111110",
  17985=>"111011000",
  17986=>"000111110",
  17987=>"111111010",
  17988=>"111111011",
  17989=>"000000000",
  17990=>"100001111",
  17991=>"100000000",
  17992=>"011111100",
  17993=>"101000111",
  17994=>"011011111",
  17995=>"111111000",
  17996=>"011011011",
  17997=>"100111000",
  17998=>"000001001",
  17999=>"111111000",
  18000=>"100100000",
  18001=>"111111111",
  18002=>"000000000",
  18003=>"110100100",
  18004=>"001000001",
  18005=>"111111001",
  18006=>"000100000",
  18007=>"001000000",
  18008=>"000000100",
  18009=>"101000000",
  18010=>"111111011",
  18011=>"011011001",
  18012=>"111111111",
  18013=>"000000000",
  18014=>"011001000",
  18015=>"111111011",
  18016=>"001001111",
  18017=>"111100100",
  18018=>"001001100",
  18019=>"111111000",
  18020=>"110001001",
  18021=>"111111110",
  18022=>"111111111",
  18023=>"000000000",
  18024=>"111011011",
  18025=>"111111000",
  18026=>"110110000",
  18027=>"101001101",
  18028=>"111111011",
  18029=>"000000000",
  18030=>"000000000",
  18031=>"000000000",
  18032=>"111100111",
  18033=>"111001011",
  18034=>"011111100",
  18035=>"100100000",
  18036=>"111111000",
  18037=>"111011011",
  18038=>"001011111",
  18039=>"111000001",
  18040=>"111111111",
  18041=>"000000000",
  18042=>"111001001",
  18043=>"101111111",
  18044=>"111110100",
  18045=>"111111111",
  18046=>"111011111",
  18047=>"000100100",
  18048=>"000000011",
  18049=>"101000110",
  18050=>"000100111",
  18051=>"111111111",
  18052=>"000000000",
  18053=>"000000111",
  18054=>"110110110",
  18055=>"001011111",
  18056=>"010011111",
  18057=>"111000000",
  18058=>"011011110",
  18059=>"000000001",
  18060=>"111011001",
  18061=>"000000000",
  18062=>"000000100",
  18063=>"111111010",
  18064=>"000000000",
  18065=>"111001000",
  18066=>"000000000",
  18067=>"010010000",
  18068=>"000000000",
  18069=>"000001011",
  18070=>"000000000",
  18071=>"001000000",
  18072=>"000001001",
  18073=>"101100000",
  18074=>"001111000",
  18075=>"111111111",
  18076=>"100100001",
  18077=>"000000001",
  18078=>"110111111",
  18079=>"011010110",
  18080=>"000100111",
  18081=>"110111001",
  18082=>"000000001",
  18083=>"000000000",
  18084=>"000000011",
  18085=>"000001001",
  18086=>"111100111",
  18087=>"111011011",
  18088=>"111111010",
  18089=>"101111001",
  18090=>"011111110",
  18091=>"111111111",
  18092=>"101101101",
  18093=>"001000011",
  18094=>"011011011",
  18095=>"111111111",
  18096=>"111111010",
  18097=>"001011001",
  18098=>"111111111",
  18099=>"000000000",
  18100=>"100001001",
  18101=>"000000111",
  18102=>"000001011",
  18103=>"000000100",
  18104=>"001110000",
  18105=>"000111101",
  18106=>"000010000",
  18107=>"100100000",
  18108=>"111111111",
  18109=>"111111111",
  18110=>"111111111",
  18111=>"001001001",
  18112=>"111111111",
  18113=>"001001000",
  18114=>"111111111",
  18115=>"000000000",
  18116=>"100000101",
  18117=>"111111000",
  18118=>"111111000",
  18119=>"111111111",
  18120=>"000000000",
  18121=>"111111111",
  18122=>"011001101",
  18123=>"111111111",
  18124=>"110110000",
  18125=>"000000000",
  18126=>"000011011",
  18127=>"001101111",
  18128=>"111111111",
  18129=>"001111111",
  18130=>"001001111",
  18131=>"000000000",
  18132=>"000000111",
  18133=>"000000000",
  18134=>"001001100",
  18135=>"001000000",
  18136=>"110100111",
  18137=>"011001101",
  18138=>"100000111",
  18139=>"011111000",
  18140=>"001000000",
  18141=>"110000100",
  18142=>"000000000",
  18143=>"111111111",
  18144=>"000000001",
  18145=>"110110111",
  18146=>"111111111",
  18147=>"111111111",
  18148=>"111011001",
  18149=>"111111110",
  18150=>"111111111",
  18151=>"001111011",
  18152=>"000000011",
  18153=>"111111011",
  18154=>"111111011",
  18155=>"000000111",
  18156=>"000000000",
  18157=>"000000111",
  18158=>"000000110",
  18159=>"000000000",
  18160=>"100100010",
  18161=>"000000010",
  18162=>"110000000",
  18163=>"011001101",
  18164=>"111111111",
  18165=>"000111111",
  18166=>"000000011",
  18167=>"000000000",
  18168=>"011001000",
  18169=>"000000000",
  18170=>"001011011",
  18171=>"011001000",
  18172=>"111101000",
  18173=>"111000011",
  18174=>"000000000",
  18175=>"101111001",
  18176=>"001001001",
  18177=>"011011011",
  18178=>"110111111",
  18179=>"000000111",
  18180=>"001101111",
  18181=>"000000000",
  18182=>"000000000",
  18183=>"001011001",
  18184=>"111000000",
  18185=>"000000000",
  18186=>"111111000",
  18187=>"100110111",
  18188=>"111111100",
  18189=>"111111000",
  18190=>"000000000",
  18191=>"000000000",
  18192=>"000000000",
  18193=>"000001111",
  18194=>"111000000",
  18195=>"111111011",
  18196=>"000000001",
  18197=>"100111111",
  18198=>"000000000",
  18199=>"111111111",
  18200=>"110000000",
  18201=>"110111111",
  18202=>"101100111",
  18203=>"111111111",
  18204=>"100000000",
  18205=>"000000000",
  18206=>"100111111",
  18207=>"001111111",
  18208=>"000000000",
  18209=>"011111110",
  18210=>"100111111",
  18211=>"111111111",
  18212=>"011111111",
  18213=>"101000000",
  18214=>"000000001",
  18215=>"010000001",
  18216=>"111111111",
  18217=>"000000000",
  18218=>"000000000",
  18219=>"000111110",
  18220=>"000000011",
  18221=>"110100111",
  18222=>"010011111",
  18223=>"111111110",
  18224=>"000000000",
  18225=>"000000000",
  18226=>"111111111",
  18227=>"100111111",
  18228=>"001000000",
  18229=>"111111111",
  18230=>"000000000",
  18231=>"000000000",
  18232=>"001000000",
  18233=>"001000000",
  18234=>"111111011",
  18235=>"100111000",
  18236=>"011011011",
  18237=>"111111111",
  18238=>"010001011",
  18239=>"111001000",
  18240=>"100110000",
  18241=>"111111110",
  18242=>"111111111",
  18243=>"000011011",
  18244=>"001111101",
  18245=>"101001000",
  18246=>"000000111",
  18247=>"000000111",
  18248=>"000000000",
  18249=>"111111110",
  18250=>"000000111",
  18251=>"111111111",
  18252=>"111111111",
  18253=>"111000000",
  18254=>"011111111",
  18255=>"100100000",
  18256=>"011111111",
  18257=>"111001001",
  18258=>"000000000",
  18259=>"111111111",
  18260=>"111101111",
  18261=>"011011111",
  18262=>"000000000",
  18263=>"101111011",
  18264=>"001101110",
  18265=>"111111111",
  18266=>"000010000",
  18267=>"101111111",
  18268=>"000111111",
  18269=>"011011000",
  18270=>"000000101",
  18271=>"000000000",
  18272=>"000000000",
  18273=>"010011000",
  18274=>"011000000",
  18275=>"001000000",
  18276=>"000011001",
  18277=>"000000000",
  18278=>"111101000",
  18279=>"000001111",
  18280=>"001000100",
  18281=>"110111111",
  18282=>"111111111",
  18283=>"011111111",
  18284=>"111011011",
  18285=>"000000000",
  18286=>"000000000",
  18287=>"111011011",
  18288=>"000000000",
  18289=>"000000000",
  18290=>"110111111",
  18291=>"011001011",
  18292=>"000111110",
  18293=>"111111001",
  18294=>"111001000",
  18295=>"001111011",
  18296=>"111111111",
  18297=>"000000000",
  18298=>"000000100",
  18299=>"011111110",
  18300=>"110111111",
  18301=>"000001001",
  18302=>"001001111",
  18303=>"011111111",
  18304=>"011111111",
  18305=>"000111010",
  18306=>"000000001",
  18307=>"111111111",
  18308=>"100000001",
  18309=>"111111110",
  18310=>"000000000",
  18311=>"000000001",
  18312=>"000000000",
  18313=>"000110010",
  18314=>"001001000",
  18315=>"111111111",
  18316=>"101001111",
  18317=>"001101110",
  18318=>"001111001",
  18319=>"010111010",
  18320=>"000011011",
  18321=>"111001001",
  18322=>"110000101",
  18323=>"100110110",
  18324=>"111011000",
  18325=>"000010111",
  18326=>"001100100",
  18327=>"001000100",
  18328=>"000000000",
  18329=>"000100100",
  18330=>"100100100",
  18331=>"001111110",
  18332=>"000000011",
  18333=>"011011111",
  18334=>"000000000",
  18335=>"110111111",
  18336=>"000000001",
  18337=>"011110110",
  18338=>"000000001",
  18339=>"111000000",
  18340=>"111111111",
  18341=>"000001001",
  18342=>"001001000",
  18343=>"001111111",
  18344=>"000000000",
  18345=>"111100000",
  18346=>"000000000",
  18347=>"001000000",
  18348=>"000000000",
  18349=>"000110100",
  18350=>"111111101",
  18351=>"000000000",
  18352=>"000000000",
  18353=>"111111111",
  18354=>"001000111",
  18355=>"001001001",
  18356=>"100000100",
  18357=>"111111101",
  18358=>"001001001",
  18359=>"000111111",
  18360=>"000000111",
  18361=>"001000000",
  18362=>"000000110",
  18363=>"100001001",
  18364=>"000000000",
  18365=>"000000000",
  18366=>"000000000",
  18367=>"000010000",
  18368=>"111111111",
  18369=>"001001111",
  18370=>"111111111",
  18371=>"010011011",
  18372=>"110110111",
  18373=>"100100000",
  18374=>"111111111",
  18375=>"001001001",
  18376=>"001001001",
  18377=>"111111111",
  18378=>"001001000",
  18379=>"000000000",
  18380=>"000011000",
  18381=>"111111001",
  18382=>"000000000",
  18383=>"000111111",
  18384=>"000000000",
  18385=>"101111111",
  18386=>"111111111",
  18387=>"110111110",
  18388=>"111111111",
  18389=>"000000000",
  18390=>"000000000",
  18391=>"000000001",
  18392=>"111111111",
  18393=>"110111001",
  18394=>"111111111",
  18395=>"001100000",
  18396=>"010000100",
  18397=>"111111101",
  18398=>"000000000",
  18399=>"000000011",
  18400=>"000100110",
  18401=>"011000000",
  18402=>"000000000",
  18403=>"111111111",
  18404=>"000000000",
  18405=>"000101000",
  18406=>"111110100",
  18407=>"110110000",
  18408=>"001001111",
  18409=>"111111111",
  18410=>"000000001",
  18411=>"000000000",
  18412=>"111111111",
  18413=>"100100100",
  18414=>"000001111",
  18415=>"000000100",
  18416=>"000000000",
  18417=>"111111110",
  18418=>"011001001",
  18419=>"111111111",
  18420=>"000010000",
  18421=>"000000000",
  18422=>"111111111",
  18423=>"111111111",
  18424=>"101111101",
  18425=>"100111111",
  18426=>"001001101",
  18427=>"000000100",
  18428=>"111101111",
  18429=>"000000100",
  18430=>"000000111",
  18431=>"111111111",
  18432=>"000000011",
  18433=>"000001000",
  18434=>"110110110",
  18435=>"000000000",
  18436=>"011000110",
  18437=>"000000000",
  18438=>"000000000",
  18439=>"101000000",
  18440=>"000000000",
  18441=>"010000011",
  18442=>"000111111",
  18443=>"010000010",
  18444=>"000000000",
  18445=>"111111000",
  18446=>"111111101",
  18447=>"111111111",
  18448=>"001011011",
  18449=>"000001111",
  18450=>"111111111",
  18451=>"010000000",
  18452=>"000111111",
  18453=>"000000000",
  18454=>"000000000",
  18455=>"111110110",
  18456=>"000000000",
  18457=>"011111111",
  18458=>"001000001",
  18459=>"000111000",
  18460=>"111111111",
  18461=>"000111111",
  18462=>"101001101",
  18463=>"000111110",
  18464=>"011111111",
  18465=>"000101111",
  18466=>"000000001",
  18467=>"111111111",
  18468=>"111111111",
  18469=>"000000000",
  18470=>"111111111",
  18471=>"000000000",
  18472=>"000010111",
  18473=>"111110110",
  18474=>"110100000",
  18475=>"000000000",
  18476=>"000000000",
  18477=>"000000000",
  18478=>"111111111",
  18479=>"100100111",
  18480=>"111111000",
  18481=>"011000000",
  18482=>"001001111",
  18483=>"000000001",
  18484=>"000000000",
  18485=>"111111111",
  18486=>"000110111",
  18487=>"010000001",
  18488=>"000110110",
  18489=>"111111111",
  18490=>"000000000",
  18491=>"111111011",
  18492=>"011001101",
  18493=>"111111100",
  18494=>"111000000",
  18495=>"000000000",
  18496=>"111111000",
  18497=>"001000011",
  18498=>"000100111",
  18499=>"000000111",
  18500=>"000111110",
  18501=>"111000000",
  18502=>"101100000",
  18503=>"000000000",
  18504=>"000101000",
  18505=>"001000111",
  18506=>"000000000",
  18507=>"000001111",
  18508=>"101011011",
  18509=>"000000000",
  18510=>"000000000",
  18511=>"000000000",
  18512=>"111111111",
  18513=>"000000000",
  18514=>"000110110",
  18515=>"000000000",
  18516=>"111000001",
  18517=>"010000100",
  18518=>"000100110",
  18519=>"111100100",
  18520=>"000000000",
  18521=>"000000000",
  18522=>"001000100",
  18523=>"001001000",
  18524=>"111111111",
  18525=>"000000000",
  18526=>"011111000",
  18527=>"000011011",
  18528=>"001001000",
  18529=>"000100000",
  18530=>"111101000",
  18531=>"111111001",
  18532=>"111011111",
  18533=>"111111000",
  18534=>"111110011",
  18535=>"000000000",
  18536=>"111111000",
  18537=>"100100111",
  18538=>"111111000",
  18539=>"111111000",
  18540=>"011111111",
  18541=>"100000111",
  18542=>"111111111",
  18543=>"000000100",
  18544=>"111111111",
  18545=>"000001000",
  18546=>"010111111",
  18547=>"000001011",
  18548=>"100000000",
  18549=>"000111111",
  18550=>"111111111",
  18551=>"000000011",
  18552=>"001101000",
  18553=>"100101111",
  18554=>"000000100",
  18555=>"100100100",
  18556=>"011011111",
  18557=>"000000000",
  18558=>"000100100",
  18559=>"000000000",
  18560=>"111111010",
  18561=>"000000000",
  18562=>"000000111",
  18563=>"001000000",
  18564=>"000000111",
  18565=>"100100111",
  18566=>"011001001",
  18567=>"101111111",
  18568=>"000000010",
  18569=>"001001000",
  18570=>"000000000",
  18571=>"000110110",
  18572=>"111111001",
  18573=>"000000001",
  18574=>"011011001",
  18575=>"111111111",
  18576=>"000000000",
  18577=>"000110000",
  18578=>"011000010",
  18579=>"111100110",
  18580=>"101111000",
  18581=>"110000100",
  18582=>"001100100",
  18583=>"000000000",
  18584=>"000000001",
  18585=>"110111111",
  18586=>"111111111",
  18587=>"111100101",
  18588=>"000111011",
  18589=>"111011110",
  18590=>"000000011",
  18591=>"000000000",
  18592=>"111111111",
  18593=>"000000000",
  18594=>"111111111",
  18595=>"100110111",
  18596=>"001100111",
  18597=>"000001111",
  18598=>"101000000",
  18599=>"111111111",
  18600=>"000000000",
  18601=>"000000000",
  18602=>"000000000",
  18603=>"000000111",
  18604=>"000111111",
  18605=>"001001001",
  18606=>"011110111",
  18607=>"000000000",
  18608=>"111111111",
  18609=>"011011001",
  18610=>"110111111",
  18611=>"100100000",
  18612=>"100101101",
  18613=>"111111111",
  18614=>"000000000",
  18615=>"110111111",
  18616=>"011010000",
  18617=>"000000110",
  18618=>"000000000",
  18619=>"000000000",
  18620=>"000000000",
  18621=>"000011111",
  18622=>"111111111",
  18623=>"111001000",
  18624=>"000110000",
  18625=>"110000000",
  18626=>"111111110",
  18627=>"000000000",
  18628=>"001000001",
  18629=>"000000000",
  18630=>"100100111",
  18631=>"000110110",
  18632=>"111011100",
  18633=>"000000000",
  18634=>"010110111",
  18635=>"000000110",
  18636=>"000000000",
  18637=>"001111111",
  18638=>"101001101",
  18639=>"000000000",
  18640=>"111111111",
  18641=>"111111111",
  18642=>"111111111",
  18643=>"100100000",
  18644=>"001000001",
  18645=>"000000000",
  18646=>"000111111",
  18647=>"000110111",
  18648=>"111010010",
  18649=>"000000000",
  18650=>"001001111",
  18651=>"001000111",
  18652=>"011111111",
  18653=>"000111111",
  18654=>"100000100",
  18655=>"110110110",
  18656=>"001001001",
  18657=>"000000010",
  18658=>"001001011",
  18659=>"000000000",
  18660=>"001000000",
  18661=>"011001001",
  18662=>"000100111",
  18663=>"100101101",
  18664=>"101111111",
  18665=>"001000000",
  18666=>"111110010",
  18667=>"111100000",
  18668=>"011111010",
  18669=>"011000000",
  18670=>"000000000",
  18671=>"111111111",
  18672=>"111101111",
  18673=>"000000011",
  18674=>"111111111",
  18675=>"000000000",
  18676=>"000000011",
  18677=>"011000000",
  18678=>"100100111",
  18679=>"011111011",
  18680=>"001000000",
  18681=>"000000010",
  18682=>"111111111",
  18683=>"000000000",
  18684=>"110111011",
  18685=>"110000000",
  18686=>"111000000",
  18687=>"100110110",
  18688=>"000000000",
  18689=>"111101001",
  18690=>"111111111",
  18691=>"011111000",
  18692=>"011111110",
  18693=>"000000100",
  18694=>"111111110",
  18695=>"000000000",
  18696=>"111010111",
  18697=>"111100000",
  18698=>"111111111",
  18699=>"000000000",
  18700=>"111111111",
  18701=>"001001001",
  18702=>"000000100",
  18703=>"111111111",
  18704=>"111010111",
  18705=>"111111011",
  18706=>"000000000",
  18707=>"110011111",
  18708=>"000000000",
  18709=>"010011000",
  18710=>"101101001",
  18711=>"110110110",
  18712=>"111111111",
  18713=>"000000000",
  18714=>"101000111",
  18715=>"110011111",
  18716=>"111111111",
  18717=>"111111000",
  18718=>"000000000",
  18719=>"111010011",
  18720=>"100111001",
  18721=>"111111000",
  18722=>"110101111",
  18723=>"011011000",
  18724=>"000000000",
  18725=>"000100000",
  18726=>"000011000",
  18727=>"000000000",
  18728=>"111111100",
  18729=>"000000000",
  18730=>"000000000",
  18731=>"000000000",
  18732=>"000000000",
  18733=>"001001001",
  18734=>"011011111",
  18735=>"000000100",
  18736=>"000000000",
  18737=>"000000000",
  18738=>"000000000",
  18739=>"110111111",
  18740=>"001001000",
  18741=>"101111100",
  18742=>"000000000",
  18743=>"110100000",
  18744=>"000000000",
  18745=>"000000000",
  18746=>"111111111",
  18747=>"000000000",
  18748=>"100110110",
  18749=>"001110100",
  18750=>"110100100",
  18751=>"111111000",
  18752=>"000000000",
  18753=>"011001011",
  18754=>"011001001",
  18755=>"000000000",
  18756=>"010000000",
  18757=>"111111111",
  18758=>"000000111",
  18759=>"000000000",
  18760=>"000000100",
  18761=>"000011000",
  18762=>"000010100",
  18763=>"100100000",
  18764=>"110111000",
  18765=>"100100000",
  18766=>"111111111",
  18767=>"010010010",
  18768=>"000010011",
  18769=>"010111000",
  18770=>"111111111",
  18771=>"000000000",
  18772=>"000000100",
  18773=>"001011011",
  18774=>"000000001",
  18775=>"111111111",
  18776=>"111111111",
  18777=>"000100111",
  18778=>"111111111",
  18779=>"011111111",
  18780=>"101000000",
  18781=>"111111000",
  18782=>"000000000",
  18783=>"001001111",
  18784=>"111000111",
  18785=>"000000111",
  18786=>"000110000",
  18787=>"111001001",
  18788=>"110111011",
  18789=>"000011111",
  18790=>"001000100",
  18791=>"000000011",
  18792=>"001000000",
  18793=>"111000111",
  18794=>"000000111",
  18795=>"111111111",
  18796=>"111111111",
  18797=>"001111111",
  18798=>"000000000",
  18799=>"000000000",
  18800=>"000000000",
  18801=>"111111111",
  18802=>"111001001",
  18803=>"111111111",
  18804=>"100000000",
  18805=>"000100100",
  18806=>"001011011",
  18807=>"000000000",
  18808=>"000000111",
  18809=>"000000000",
  18810=>"000000000",
  18811=>"000000000",
  18812=>"011111111",
  18813=>"011001001",
  18814=>"110000000",
  18815=>"111111111",
  18816=>"000000000",
  18817=>"000000000",
  18818=>"000000000",
  18819=>"100000000",
  18820=>"110111111",
  18821=>"000000000",
  18822=>"111111111",
  18823=>"000011111",
  18824=>"111111001",
  18825=>"001000000",
  18826=>"111111101",
  18827=>"000000100",
  18828=>"011001000",
  18829=>"111011000",
  18830=>"110110111",
  18831=>"111111111",
  18832=>"111111111",
  18833=>"000000000",
  18834=>"000000010",
  18835=>"110001001",
  18836=>"000000100",
  18837=>"000001000",
  18838=>"000000000",
  18839=>"111111000",
  18840=>"000000000",
  18841=>"111100100",
  18842=>"100111111",
  18843=>"011111110",
  18844=>"000000111",
  18845=>"000100100",
  18846=>"110100111",
  18847=>"111111101",
  18848=>"110110000",
  18849=>"100100000",
  18850=>"000000000",
  18851=>"011011000",
  18852=>"000000000",
  18853=>"000000000",
  18854=>"000000111",
  18855=>"000000000",
  18856=>"111011000",
  18857=>"100000000",
  18858=>"000000000",
  18859=>"011111111",
  18860=>"000000000",
  18861=>"000000000",
  18862=>"001000000",
  18863=>"000000000",
  18864=>"111111101",
  18865=>"000000000",
  18866=>"110110000",
  18867=>"111011110",
  18868=>"110110110",
  18869=>"000110110",
  18870=>"000000100",
  18871=>"111111101",
  18872=>"000111111",
  18873=>"111000000",
  18874=>"001111000",
  18875=>"111111111",
  18876=>"001111000",
  18877=>"000000000",
  18878=>"100000000",
  18879=>"000000000",
  18880=>"111111111",
  18881=>"111111111",
  18882=>"000000000",
  18883=>"111111111",
  18884=>"000000100",
  18885=>"111111011",
  18886=>"000000000",
  18887=>"111000001",
  18888=>"000000011",
  18889=>"101110000",
  18890=>"000001001",
  18891=>"000000110",
  18892=>"110111001",
  18893=>"000000000",
  18894=>"000000110",
  18895=>"001001000",
  18896=>"111111111",
  18897=>"111111111",
  18898=>"111111111",
  18899=>"110100111",
  18900=>"100111111",
  18901=>"111111000",
  18902=>"111010000",
  18903=>"000000000",
  18904=>"001000000",
  18905=>"010000000",
  18906=>"110100110",
  18907=>"111111111",
  18908=>"110000000",
  18909=>"011011000",
  18910=>"000000000",
  18911=>"111111101",
  18912=>"111111111",
  18913=>"100000000",
  18914=>"000111011",
  18915=>"000000100",
  18916=>"000000000",
  18917=>"111100101",
  18918=>"000000000",
  18919=>"000011010",
  18920=>"011111111",
  18921=>"011111111",
  18922=>"111101101",
  18923=>"011111000",
  18924=>"000000010",
  18925=>"110110110",
  18926=>"111111111",
  18927=>"111111111",
  18928=>"000000000",
  18929=>"011011111",
  18930=>"111111111",
  18931=>"001101111",
  18932=>"111111011",
  18933=>"111111111",
  18934=>"100000000",
  18935=>"110010000",
  18936=>"111111111",
  18937=>"011001011",
  18938=>"101101100",
  18939=>"000110000",
  18940=>"011011000",
  18941=>"110111111",
  18942=>"111101111",
  18943=>"001001101",
  18944=>"000000000",
  18945=>"000000011",
  18946=>"101001101",
  18947=>"111100101",
  18948=>"000111111",
  18949=>"010000000",
  18950=>"111000000",
  18951=>"111111111",
  18952=>"111111000",
  18953=>"001000000",
  18954=>"000000111",
  18955=>"000000000",
  18956=>"110110100",
  18957=>"011000000",
  18958=>"011010000",
  18959=>"011101111",
  18960=>"000010011",
  18961=>"000000100",
  18962=>"000000001",
  18963=>"010000000",
  18964=>"000111110",
  18965=>"101101101",
  18966=>"000000111",
  18967=>"000111000",
  18968=>"000000000",
  18969=>"001000100",
  18970=>"111111111",
  18971=>"111111111",
  18972=>"100100100",
  18973=>"000110000",
  18974=>"001011001",
  18975=>"100011111",
  18976=>"000111111",
  18977=>"111111011",
  18978=>"000111011",
  18979=>"111111111",
  18980=>"000000001",
  18981=>"000111111",
  18982=>"000011011",
  18983=>"000000111",
  18984=>"000000000",
  18985=>"001101111",
  18986=>"000010111",
  18987=>"000000000",
  18988=>"011111011",
  18989=>"111011000",
  18990=>"111110000",
  18991=>"000000111",
  18992=>"001111001",
  18993=>"111111101",
  18994=>"100100100",
  18995=>"011000000",
  18996=>"000000000",
  18997=>"110000000",
  18998=>"000000000",
  18999=>"111011000",
  19000=>"110110110",
  19001=>"100111111",
  19002=>"111000011",
  19003=>"111111000",
  19004=>"111111101",
  19005=>"100000000",
  19006=>"111111000",
  19007=>"000000000",
  19008=>"111111011",
  19009=>"000000001",
  19010=>"000000000",
  19011=>"000000000",
  19012=>"000000000",
  19013=>"000100000",
  19014=>"111101111",
  19015=>"111111111",
  19016=>"000100111",
  19017=>"111111111",
  19018=>"000111111",
  19019=>"010111000",
  19020=>"000000111",
  19021=>"100000000",
  19022=>"000000000",
  19023=>"111111111",
  19024=>"000100000",
  19025=>"000011111",
  19026=>"000110110",
  19027=>"011001000",
  19028=>"100000000",
  19029=>"000000000",
  19030=>"000000011",
  19031=>"001000000",
  19032=>"000110111",
  19033=>"101000101",
  19034=>"111001000",
  19035=>"000101111",
  19036=>"001000100",
  19037=>"101111111",
  19038=>"111111111",
  19039=>"100000000",
  19040=>"111111111",
  19041=>"000011111",
  19042=>"000000000",
  19043=>"001011111",
  19044=>"101101000",
  19045=>"111011010",
  19046=>"000000000",
  19047=>"100101111",
  19048=>"111110000",
  19049=>"000000000",
  19050=>"000000000",
  19051=>"000110110",
  19052=>"111000001",
  19053=>"000000000",
  19054=>"100100111",
  19055=>"000011011",
  19056=>"001111111",
  19057=>"111000111",
  19058=>"111000000",
  19059=>"011011111",
  19060=>"111000000",
  19061=>"101001001",
  19062=>"000000000",
  19063=>"010111111",
  19064=>"011001000",
  19065=>"111111111",
  19066=>"111001000",
  19067=>"100110110",
  19068=>"010011111",
  19069=>"111111000",
  19070=>"000000011",
  19071=>"000011001",
  19072=>"000000000",
  19073=>"010011000",
  19074=>"111001000",
  19075=>"000000011",
  19076=>"001100111",
  19077=>"011000111",
  19078=>"001001001",
  19079=>"010000000",
  19080=>"000000000",
  19081=>"001110111",
  19082=>"000000000",
  19083=>"001000000",
  19084=>"000000000",
  19085=>"000000000",
  19086=>"000000000",
  19087=>"000000000",
  19088=>"111000000",
  19089=>"000010000",
  19090=>"000000111",
  19091=>"001000000",
  19092=>"011110000",
  19093=>"111111111",
  19094=>"000000101",
  19095=>"111011111",
  19096=>"111011011",
  19097=>"000000000",
  19098=>"111111011",
  19099=>"111111111",
  19100=>"000111111",
  19101=>"110110000",
  19102=>"010000000",
  19103=>"000000000",
  19104=>"111111110",
  19105=>"000000000",
  19106=>"000000001",
  19107=>"000000000",
  19108=>"111111000",
  19109=>"111111111",
  19110=>"000001000",
  19111=>"000000101",
  19112=>"000000000",
  19113=>"000001111",
  19114=>"000000000",
  19115=>"110111111",
  19116=>"001000000",
  19117=>"000000000",
  19118=>"111111111",
  19119=>"011111111",
  19120=>"000000000",
  19121=>"000000111",
  19122=>"111111111",
  19123=>"000000000",
  19124=>"000000000",
  19125=>"000000000",
  19126=>"010111101",
  19127=>"110000000",
  19128=>"110111111",
  19129=>"111001000",
  19130=>"111101000",
  19131=>"110111111",
  19132=>"101000111",
  19133=>"000000100",
  19134=>"110111111",
  19135=>"110000000",
  19136=>"111111111",
  19137=>"111111111",
  19138=>"111000000",
  19139=>"001000000",
  19140=>"000000000",
  19141=>"111000001",
  19142=>"000001000",
  19143=>"000000000",
  19144=>"000000011",
  19145=>"111111111",
  19146=>"000100111",
  19147=>"111111000",
  19148=>"000000100",
  19149=>"000011010",
  19150=>"011000000",
  19151=>"000000000",
  19152=>"011010010",
  19153=>"111111011",
  19154=>"111000000",
  19155=>"000000000",
  19156=>"111111100",
  19157=>"111101000",
  19158=>"111110110",
  19159=>"100000000",
  19160=>"100110011",
  19161=>"011111001",
  19162=>"000000000",
  19163=>"000000000",
  19164=>"000000000",
  19165=>"111111110",
  19166=>"000000000",
  19167=>"000000000",
  19168=>"000000000",
  19169=>"010000010",
  19170=>"111111011",
  19171=>"000001100",
  19172=>"110001011",
  19173=>"000011111",
  19174=>"000110111",
  19175=>"111100000",
  19176=>"000100111",
  19177=>"111111111",
  19178=>"101111111",
  19179=>"001111111",
  19180=>"010010010",
  19181=>"100000000",
  19182=>"000000001",
  19183=>"110000000",
  19184=>"010110011",
  19185=>"100111111",
  19186=>"111011011",
  19187=>"011101000",
  19188=>"000010111",
  19189=>"100000000",
  19190=>"111011001",
  19191=>"000000000",
  19192=>"000110111",
  19193=>"000011000",
  19194=>"111111111",
  19195=>"000011111",
  19196=>"000000001",
  19197=>"001001001",
  19198=>"000100100",
  19199=>"111111000",
  19200=>"011001000",
  19201=>"100100100",
  19202=>"011000000",
  19203=>"000111111",
  19204=>"000001000",
  19205=>"000010000",
  19206=>"010000000",
  19207=>"000101111",
  19208=>"001111111",
  19209=>"000000100",
  19210=>"111111111",
  19211=>"101000000",
  19212=>"111111111",
  19213=>"111111111",
  19214=>"000000000",
  19215=>"010000000",
  19216=>"110100000",
  19217=>"111001000",
  19218=>"000000000",
  19219=>"000000000",
  19220=>"111011000",
  19221=>"111111011",
  19222=>"100000000",
  19223=>"000000000",
  19224=>"110000110",
  19225=>"111111111",
  19226=>"000000011",
  19227=>"010011111",
  19228=>"110111100",
  19229=>"000000110",
  19230=>"111111111",
  19231=>"111111001",
  19232=>"110100000",
  19233=>"011111111",
  19234=>"111111111",
  19235=>"100100100",
  19236=>"100111001",
  19237=>"000001001",
  19238=>"000000000",
  19239=>"111111111",
  19240=>"111111111",
  19241=>"000101000",
  19242=>"011111111",
  19243=>"000000000",
  19244=>"000101000",
  19245=>"110110010",
  19246=>"000000000",
  19247=>"111111010",
  19248=>"100101111",
  19249=>"111111011",
  19250=>"000000000",
  19251=>"111111010",
  19252=>"111101001",
  19253=>"111110000",
  19254=>"000000001",
  19255=>"000011111",
  19256=>"000001001",
  19257=>"000000000",
  19258=>"111000010",
  19259=>"000011000",
  19260=>"000000000",
  19261=>"000001000",
  19262=>"100111111",
  19263=>"111111000",
  19264=>"111111011",
  19265=>"111111111",
  19266=>"101111111",
  19267=>"111000000",
  19268=>"000110000",
  19269=>"000000111",
  19270=>"111000000",
  19271=>"111111001",
  19272=>"111101110",
  19273=>"111000000",
  19274=>"100000011",
  19275=>"110100000",
  19276=>"111110111",
  19277=>"000000000",
  19278=>"110010000",
  19279=>"111111111",
  19280=>"111001001",
  19281=>"110001011",
  19282=>"001111011",
  19283=>"101000000",
  19284=>"000000000",
  19285=>"011011011",
  19286=>"111001000",
  19287=>"011001000",
  19288=>"111111111",
  19289=>"011111000",
  19290=>"111001000",
  19291=>"011001000",
  19292=>"111001101",
  19293=>"111001000",
  19294=>"111010011",
  19295=>"000000110",
  19296=>"011111011",
  19297=>"110111011",
  19298=>"110111111",
  19299=>"101101000",
  19300=>"110000000",
  19301=>"010000000",
  19302=>"110111111",
  19303=>"000000000",
  19304=>"000000001",
  19305=>"010010000",
  19306=>"111101111",
  19307=>"011110111",
  19308=>"100100110",
  19309=>"111111110",
  19310=>"000000000",
  19311=>"111100101",
  19312=>"100000000",
  19313=>"110110111",
  19314=>"000111111",
  19315=>"111111111",
  19316=>"101000000",
  19317=>"011011001",
  19318=>"110111111",
  19319=>"101100000",
  19320=>"000000011",
  19321=>"111111100",
  19322=>"111001000",
  19323=>"111111000",
  19324=>"111100100",
  19325=>"111111111",
  19326=>"110110000",
  19327=>"110110111",
  19328=>"000110010",
  19329=>"001111111",
  19330=>"001001000",
  19331=>"110111111",
  19332=>"001001001",
  19333=>"000000000",
  19334=>"000111111",
  19335=>"011100101",
  19336=>"011000000",
  19337=>"000000001",
  19338=>"000111011",
  19339=>"001111011",
  19340=>"101111111",
  19341=>"101110111",
  19342=>"110111111",
  19343=>"111111111",
  19344=>"000111111",
  19345=>"111111111",
  19346=>"111110000",
  19347=>"000000000",
  19348=>"111101000",
  19349=>"000000000",
  19350=>"011000000",
  19351=>"111111000",
  19352=>"000000001",
  19353=>"011111111",
  19354=>"111101111",
  19355=>"011000000",
  19356=>"000000000",
  19357=>"100000000",
  19358=>"000000000",
  19359=>"000100111",
  19360=>"111111011",
  19361=>"100000001",
  19362=>"001000000",
  19363=>"000111111",
  19364=>"001111111",
  19365=>"000000111",
  19366=>"100000111",
  19367=>"000000000",
  19368=>"011011010",
  19369=>"110000000",
  19370=>"000001011",
  19371=>"111011000",
  19372=>"010111000",
  19373=>"000100000",
  19374=>"000101111",
  19375=>"111111000",
  19376=>"000000000",
  19377=>"000000000",
  19378=>"000000111",
  19379=>"000000000",
  19380=>"000111111",
  19381=>"111111000",
  19382=>"000001000",
  19383=>"000100000",
  19384=>"000000100",
  19385=>"000000110",
  19386=>"111111111",
  19387=>"111110110",
  19388=>"000000101",
  19389=>"011000001",
  19390=>"000000111",
  19391=>"100000000",
  19392=>"000000000",
  19393=>"011010000",
  19394=>"111000000",
  19395=>"111111000",
  19396=>"110111111",
  19397=>"111101111",
  19398=>"000111011",
  19399=>"111011011",
  19400=>"011000000",
  19401=>"100111111",
  19402=>"011000000",
  19403=>"000000100",
  19404=>"000000000",
  19405=>"000100000",
  19406=>"001011001",
  19407=>"000111111",
  19408=>"100111111",
  19409=>"001000000",
  19410=>"111110110",
  19411=>"111111110",
  19412=>"000111111",
  19413=>"110111100",
  19414=>"000011000",
  19415=>"000000000",
  19416=>"001011000",
  19417=>"110010000",
  19418=>"110110110",
  19419=>"000011011",
  19420=>"110000000",
  19421=>"111111001",
  19422=>"000000000",
  19423=>"100100000",
  19424=>"001000011",
  19425=>"111011000",
  19426=>"111000000",
  19427=>"000000111",
  19428=>"011000000",
  19429=>"111111111",
  19430=>"111011000",
  19431=>"110111111",
  19432=>"111111000",
  19433=>"000111111",
  19434=>"000000111",
  19435=>"110111111",
  19436=>"000110100",
  19437=>"111001000",
  19438=>"001111111",
  19439=>"001001010",
  19440=>"111000100",
  19441=>"111010011",
  19442=>"111000000",
  19443=>"111000000",
  19444=>"000000000",
  19445=>"000000000",
  19446=>"000111111",
  19447=>"001111111",
  19448=>"111111000",
  19449=>"111101000",
  19450=>"000000000",
  19451=>"001000000",
  19452=>"110100101",
  19453=>"000100000",
  19454=>"001000000",
  19455=>"010000000",
  19456=>"100100000",
  19457=>"111111111",
  19458=>"000000000",
  19459=>"000000000",
  19460=>"011001011",
  19461=>"011011110",
  19462=>"101100101",
  19463=>"010111111",
  19464=>"101011011",
  19465=>"111111111",
  19466=>"111111001",
  19467=>"000000100",
  19468=>"001000000",
  19469=>"000010111",
  19470=>"111111111",
  19471=>"111111111",
  19472=>"000000000",
  19473=>"111000011",
  19474=>"110111111",
  19475=>"010000000",
  19476=>"110111000",
  19477=>"000000000",
  19478=>"100110111",
  19479=>"010001011",
  19480=>"110111111",
  19481=>"000011011",
  19482=>"110000100",
  19483=>"110111111",
  19484=>"000000000",
  19485=>"110111111",
  19486=>"100101001",
  19487=>"001000001",
  19488=>"000000000",
  19489=>"100111111",
  19490=>"000000000",
  19491=>"111111110",
  19492=>"111111111",
  19493=>"000111000",
  19494=>"111110000",
  19495=>"000000101",
  19496=>"011001000",
  19497=>"110000000",
  19498=>"111111111",
  19499=>"010011001",
  19500=>"001111111",
  19501=>"000000000",
  19502=>"001000001",
  19503=>"111111111",
  19504=>"110111111",
  19505=>"111111111",
  19506=>"000100100",
  19507=>"111111111",
  19508=>"000001111",
  19509=>"000000111",
  19510=>"001011000",
  19511=>"000000000",
  19512=>"001111000",
  19513=>"111100000",
  19514=>"111000000",
  19515=>"111001000",
  19516=>"000000000",
  19517=>"111111111",
  19518=>"001001001",
  19519=>"111111110",
  19520=>"001001001",
  19521=>"100000101",
  19522=>"000000000",
  19523=>"000001000",
  19524=>"000000100",
  19525=>"000001001",
  19526=>"100000000",
  19527=>"111111111",
  19528=>"000100100",
  19529=>"111111111",
  19530=>"111111111",
  19531=>"111111001",
  19532=>"111111110",
  19533=>"110010111",
  19534=>"011000000",
  19535=>"011111111",
  19536=>"110111111",
  19537=>"100101001",
  19538=>"001001001",
  19539=>"110111111",
  19540=>"001000001",
  19541=>"111010001",
  19542=>"000111111",
  19543=>"111111100",
  19544=>"111111111",
  19545=>"000000000",
  19546=>"111111111",
  19547=>"000110111",
  19548=>"100000000",
  19549=>"000000000",
  19550=>"000000000",
  19551=>"111111111",
  19552=>"000001001",
  19553=>"000000000",
  19554=>"100000011",
  19555=>"111111111",
  19556=>"000001111",
  19557=>"100111000",
  19558=>"100111111",
  19559=>"000000000",
  19560=>"000000000",
  19561=>"110111111",
  19562=>"000000000",
  19563=>"111000110",
  19564=>"110100000",
  19565=>"111111111",
  19566=>"000100111",
  19567=>"111111111",
  19568=>"111111111",
  19569=>"100111111",
  19570=>"001000000",
  19571=>"010000000",
  19572=>"000011111",
  19573=>"111111111",
  19574=>"000000000",
  19575=>"111011011",
  19576=>"000000000",
  19577=>"111111111",
  19578=>"111100111",
  19579=>"000000000",
  19580=>"000110000",
  19581=>"010011000",
  19582=>"000000000",
  19583=>"000000000",
  19584=>"100111111",
  19585=>"111111001",
  19586=>"100000000",
  19587=>"011111111",
  19588=>"111111111",
  19589=>"110111111",
  19590=>"001001001",
  19591=>"000000000",
  19592=>"111111111",
  19593=>"101000000",
  19594=>"111111111",
  19595=>"000000000",
  19596=>"101101001",
  19597=>"010010000",
  19598=>"110111000",
  19599=>"001000000",
  19600=>"011111010",
  19601=>"000000000",
  19602=>"111111101",
  19603=>"000000000",
  19604=>"111111111",
  19605=>"000110000",
  19606=>"000000000",
  19607=>"011101000",
  19608=>"000111000",
  19609=>"111101111",
  19610=>"111100100",
  19611=>"001000001",
  19612=>"111111010",
  19613=>"000010010",
  19614=>"111110100",
  19615=>"101101000",
  19616=>"111111111",
  19617=>"111111011",
  19618=>"001111111",
  19619=>"000111111",
  19620=>"111110110",
  19621=>"100111111",
  19622=>"000000000",
  19623=>"000000000",
  19624=>"000000000",
  19625=>"000000000",
  19626=>"000000000",
  19627=>"111111111",
  19628=>"111111110",
  19629=>"111111111",
  19630=>"000100000",
  19631=>"011011000",
  19632=>"010111111",
  19633=>"001001001",
  19634=>"110110110",
  19635=>"000000000",
  19636=>"000000111",
  19637=>"000111000",
  19638=>"111111000",
  19639=>"001001011",
  19640=>"101111111",
  19641=>"000111111",
  19642=>"101000111",
  19643=>"110111111",
  19644=>"000100000",
  19645=>"111111111",
  19646=>"111111111",
  19647=>"100111111",
  19648=>"111111000",
  19649=>"111111111",
  19650=>"111011111",
  19651=>"000000000",
  19652=>"110111111",
  19653=>"000000000",
  19654=>"110000011",
  19655=>"111111111",
  19656=>"000000011",
  19657=>"011000000",
  19658=>"111100111",
  19659=>"001001011",
  19660=>"110111111",
  19661=>"111000000",
  19662=>"111111111",
  19663=>"011011111",
  19664=>"000111000",
  19665=>"000111111",
  19666=>"000010011",
  19667=>"001000101",
  19668=>"011111111",
  19669=>"000000000",
  19670=>"000000000",
  19671=>"000000000",
  19672=>"111111111",
  19673=>"000000000",
  19674=>"000000000",
  19675=>"111111000",
  19676=>"000100000",
  19677=>"000000101",
  19678=>"000000000",
  19679=>"000000000",
  19680=>"111000000",
  19681=>"111011000",
  19682=>"111111110",
  19683=>"000000000",
  19684=>"111010111",
  19685=>"111111100",
  19686=>"100110111",
  19687=>"000000101",
  19688=>"111011001",
  19689=>"010000000",
  19690=>"111110000",
  19691=>"111101000",
  19692=>"000000000",
  19693=>"000000000",
  19694=>"000010000",
  19695=>"110110000",
  19696=>"111100101",
  19697=>"000111111",
  19698=>"011111111",
  19699=>"000000000",
  19700=>"111111111",
  19701=>"111111011",
  19702=>"011011001",
  19703=>"111111111",
  19704=>"111111111",
  19705=>"000000010",
  19706=>"000000000",
  19707=>"000000000",
  19708=>"110110000",
  19709=>"000000101",
  19710=>"000011010",
  19711=>"001000000",
  19712=>"110111111",
  19713=>"011011111",
  19714=>"111111111",
  19715=>"000001000",
  19716=>"100000000",
  19717=>"101001101",
  19718=>"000000000",
  19719=>"110100001",
  19720=>"000100000",
  19721=>"110110110",
  19722=>"000000000",
  19723=>"000000110",
  19724=>"100110110",
  19725=>"000010110",
  19726=>"000000000",
  19727=>"000000101",
  19728=>"110110110",
  19729=>"000000000",
  19730=>"000000000",
  19731=>"110010111",
  19732=>"101100100",
  19733=>"111000000",
  19734=>"000010000",
  19735=>"000100000",
  19736=>"111001001",
  19737=>"111111111",
  19738=>"000000000",
  19739=>"000000000",
  19740=>"001001001",
  19741=>"000001111",
  19742=>"000000000",
  19743=>"000001000",
  19744=>"001000000",
  19745=>"011011111",
  19746=>"000000100",
  19747=>"000000000",
  19748=>"000000011",
  19749=>"000110111",
  19750=>"000000000",
  19751=>"111111001",
  19752=>"000000111",
  19753=>"000000000",
  19754=>"000100000",
  19755=>"001000000",
  19756=>"000110000",
  19757=>"110010000",
  19758=>"111100100",
  19759=>"110110000",
  19760=>"000000000",
  19761=>"111000000",
  19762=>"111111111",
  19763=>"001000000",
  19764=>"000000000",
  19765=>"000100101",
  19766=>"000010000",
  19767=>"000100100",
  19768=>"000000000",
  19769=>"111100111",
  19770=>"101011001",
  19771=>"111100101",
  19772=>"000000000",
  19773=>"010000000",
  19774=>"000000000",
  19775=>"010000000",
  19776=>"001001000",
  19777=>"000000000",
  19778=>"010111001",
  19779=>"000000000",
  19780=>"111111111",
  19781=>"111111000",
  19782=>"110000110",
  19783=>"000011111",
  19784=>"000011000",
  19785=>"111101111",
  19786=>"111111110",
  19787=>"110111000",
  19788=>"100100010",
  19789=>"101001111",
  19790=>"111111000",
  19791=>"111111111",
  19792=>"001101001",
  19793=>"000011101",
  19794=>"000000000",
  19795=>"001000111",
  19796=>"111010110",
  19797=>"001001001",
  19798=>"000111110",
  19799=>"000000000",
  19800=>"000000000",
  19801=>"010011110",
  19802=>"000111111",
  19803=>"111011011",
  19804=>"000000111",
  19805=>"111111000",
  19806=>"100000000",
  19807=>"000010010",
  19808=>"111111001",
  19809=>"000000000",
  19810=>"000110100",
  19811=>"000000000",
  19812=>"011011111",
  19813=>"000000011",
  19814=>"000000000",
  19815=>"011001000",
  19816=>"011111000",
  19817=>"000100000",
  19818=>"000000001",
  19819=>"111111100",
  19820=>"111111011",
  19821=>"000010010",
  19822=>"111111111",
  19823=>"000110001",
  19824=>"000000000",
  19825=>"001111111",
  19826=>"111111111",
  19827=>"100110111",
  19828=>"100100000",
  19829=>"111111111",
  19830=>"000111111",
  19831=>"111111001",
  19832=>"000000000",
  19833=>"000000111",
  19834=>"110000110",
  19835=>"000010011",
  19836=>"110000010",
  19837=>"111100110",
  19838=>"000100110",
  19839=>"101000000",
  19840=>"000001011",
  19841=>"111010111",
  19842=>"000000000",
  19843=>"110100100",
  19844=>"000000000",
  19845=>"111110000",
  19846=>"110110000",
  19847=>"111111010",
  19848=>"000000000",
  19849=>"101001001",
  19850=>"111111000",
  19851=>"000000000",
  19852=>"000000000",
  19853=>"010010010",
  19854=>"000111111",
  19855=>"111111111",
  19856=>"000000000",
  19857=>"111111111",
  19858=>"111111101",
  19859=>"000000000",
  19860=>"000000000",
  19861=>"111101111",
  19862=>"100000010",
  19863=>"000000000",
  19864=>"000000000",
  19865=>"100111110",
  19866=>"111111111",
  19867=>"111111111",
  19868=>"000000000",
  19869=>"111111111",
  19870=>"000000110",
  19871=>"111111011",
  19872=>"011111111",
  19873=>"001001000",
  19874=>"000000001",
  19875=>"000000111",
  19876=>"111110000",
  19877=>"000000000",
  19878=>"110110000",
  19879=>"000000000",
  19880=>"000001101",
  19881=>"100111001",
  19882=>"000000000",
  19883=>"000000000",
  19884=>"000000000",
  19885=>"000001001",
  19886=>"000011000",
  19887=>"110100000",
  19888=>"111111100",
  19889=>"110000000",
  19890=>"001011111",
  19891=>"111111111",
  19892=>"101001000",
  19893=>"000001111",
  19894=>"111111111",
  19895=>"110100111",
  19896=>"011111100",
  19897=>"111111000",
  19898=>"001001111",
  19899=>"000111111",
  19900=>"111111111",
  19901=>"001000100",
  19902=>"001111100",
  19903=>"010010010",
  19904=>"000001111",
  19905=>"111111110",
  19906=>"111111111",
  19907=>"000000000",
  19908=>"110111111",
  19909=>"100110111",
  19910=>"011000000",
  19911=>"011111111",
  19912=>"000010000",
  19913=>"111000111",
  19914=>"000100000",
  19915=>"000000110",
  19916=>"000000000",
  19917=>"000000000",
  19918=>"111111011",
  19919=>"111111111",
  19920=>"001001001",
  19921=>"100110100",
  19922=>"111111110",
  19923=>"000000001",
  19924=>"011001000",
  19925=>"000111110",
  19926=>"010000000",
  19927=>"100100100",
  19928=>"000011011",
  19929=>"000110110",
  19930=>"000000000",
  19931=>"110111111",
  19932=>"000100101",
  19933=>"101000000",
  19934=>"001000000",
  19935=>"011011010",
  19936=>"000000100",
  19937=>"101000000",
  19938=>"111011111",
  19939=>"111111111",
  19940=>"110110000",
  19941=>"111111111",
  19942=>"000000000",
  19943=>"100111100",
  19944=>"111110101",
  19945=>"101000000",
  19946=>"000110100",
  19947=>"000000000",
  19948=>"111111111",
  19949=>"000001011",
  19950=>"100000000",
  19951=>"110011011",
  19952=>"001000111",
  19953=>"111111111",
  19954=>"111111111",
  19955=>"000000100",
  19956=>"001111000",
  19957=>"000010011",
  19958=>"010000000",
  19959=>"110110111",
  19960=>"011000110",
  19961=>"100110111",
  19962=>"111101000",
  19963=>"110100111",
  19964=>"001111111",
  19965=>"111111111",
  19966=>"111111111",
  19967=>"111111111",
  19968=>"110110111",
  19969=>"111110111",
  19970=>"011000010",
  19971=>"111111111",
  19972=>"000000000",
  19973=>"111011000",
  19974=>"000001000",
  19975=>"111111000",
  19976=>"000000001",
  19977=>"000111111",
  19978=>"111011111",
  19979=>"111000000",
  19980=>"011000000",
  19981=>"100111111",
  19982=>"100101100",
  19983=>"000000010",
  19984=>"000000000",
  19985=>"111111111",
  19986=>"000000000",
  19987=>"000000110",
  19988=>"000101101",
  19989=>"000000010",
  19990=>"111000100",
  19991=>"000001001",
  19992=>"111111111",
  19993=>"111111110",
  19994=>"111100110",
  19995=>"110000011",
  19996=>"000000111",
  19997=>"111111000",
  19998=>"001000110",
  19999=>"000000000",
  20000=>"110000000",
  20001=>"111111111",
  20002=>"111111111",
  20003=>"111111111",
  20004=>"000000000",
  20005=>"111111111",
  20006=>"111101100",
  20007=>"000001111",
  20008=>"000110111",
  20009=>"000000000",
  20010=>"000111110",
  20011=>"000111111",
  20012=>"000000111",
  20013=>"000000111",
  20014=>"000000011",
  20015=>"111111000",
  20016=>"111111111",
  20017=>"000111111",
  20018=>"100000000",
  20019=>"100000100",
  20020=>"000000000",
  20021=>"001001001",
  20022=>"000000000",
  20023=>"000000000",
  20024=>"000000000",
  20025=>"000000111",
  20026=>"000000000",
  20027=>"000000000",
  20028=>"000111111",
  20029=>"111100100",
  20030=>"010000101",
  20031=>"111111000",
  20032=>"000000101",
  20033=>"000000001",
  20034=>"000111111",
  20035=>"010000100",
  20036=>"000000111",
  20037=>"110111111",
  20038=>"000000000",
  20039=>"000000111",
  20040=>"011111111",
  20041=>"000000000",
  20042=>"000000111",
  20043=>"111111001",
  20044=>"111111111",
  20045=>"001000001",
  20046=>"000000000",
  20047=>"101111111",
  20048=>"010111111",
  20049=>"100101000",
  20050=>"000110011",
  20051=>"111101111",
  20052=>"000000000",
  20053=>"000000000",
  20054=>"110000000",
  20055=>"000000000",
  20056=>"000000110",
  20057=>"101000101",
  20058=>"100100000",
  20059=>"111110100",
  20060=>"000011111",
  20061=>"011011011",
  20062=>"100000000",
  20063=>"000000000",
  20064=>"000000000",
  20065=>"111110010",
  20066=>"100000000",
  20067=>"000100111",
  20068=>"000000000",
  20069=>"001000000",
  20070=>"111111000",
  20071=>"000000001",
  20072=>"000000000",
  20073=>"111000000",
  20074=>"111111111",
  20075=>"111011000",
  20076=>"111010100",
  20077=>"100111011",
  20078=>"111111110",
  20079=>"101110011",
  20080=>"011111111",
  20081=>"111111000",
  20082=>"001111010",
  20083=>"011011011",
  20084=>"111111111",
  20085=>"001001000",
  20086=>"001000000",
  20087=>"000000010",
  20088=>"110000000",
  20089=>"001000101",
  20090=>"001000000",
  20091=>"000010000",
  20092=>"000001000",
  20093=>"011011011",
  20094=>"000000001",
  20095=>"110010010",
  20096=>"111111111",
  20097=>"000000101",
  20098=>"011001100",
  20099=>"110000000",
  20100=>"111111111",
  20101=>"100000000",
  20102=>"111000001",
  20103=>"111111000",
  20104=>"100110111",
  20105=>"000000000",
  20106=>"111111111",
  20107=>"111111100",
  20108=>"110111010",
  20109=>"111111111",
  20110=>"110111100",
  20111=>"111111110",
  20112=>"000000001",
  20113=>"000000101",
  20114=>"000000000",
  20115=>"000000000",
  20116=>"011111111",
  20117=>"000000000",
  20118=>"000000011",
  20119=>"111111111",
  20120=>"000000000",
  20121=>"100001001",
  20122=>"111111111",
  20123=>"111111111",
  20124=>"000001000",
  20125=>"000000000",
  20126=>"111111111",
  20127=>"000000000",
  20128=>"111111011",
  20129=>"111111111",
  20130=>"000000010",
  20131=>"000000000",
  20132=>"111011111",
  20133=>"000000100",
  20134=>"110111000",
  20135=>"010100000",
  20136=>"000000100",
  20137=>"011000111",
  20138=>"001101110",
  20139=>"010111000",
  20140=>"000001001",
  20141=>"000000000",
  20142=>"110110111",
  20143=>"000000110",
  20144=>"111111000",
  20145=>"000000000",
  20146=>"111111110",
  20147=>"000011111",
  20148=>"000000001",
  20149=>"100000000",
  20150=>"111000000",
  20151=>"000011011",
  20152=>"110110100",
  20153=>"100100111",
  20154=>"111000101",
  20155=>"111110100",
  20156=>"000010000",
  20157=>"111100100",
  20158=>"000011111",
  20159=>"001001011",
  20160=>"000000001",
  20161=>"100100101",
  20162=>"000111011",
  20163=>"111011111",
  20164=>"000000001",
  20165=>"000000000",
  20166=>"000100111",
  20167=>"110111110",
  20168=>"100100111",
  20169=>"000010111",
  20170=>"000111110",
  20171=>"000111111",
  20172=>"000000111",
  20173=>"110010010",
  20174=>"000000111",
  20175=>"111110101",
  20176=>"101001000",
  20177=>"000000011",
  20178=>"111101000",
  20179=>"001001111",
  20180=>"000000000",
  20181=>"111010110",
  20182=>"111000000",
  20183=>"000000000",
  20184=>"000000000",
  20185=>"000110100",
  20186=>"000111000",
  20187=>"110000000",
  20188=>"110000000",
  20189=>"110000101",
  20190=>"010011010",
  20191=>"110100100",
  20192=>"000000000",
  20193=>"100000111",
  20194=>"000000000",
  20195=>"111011000",
  20196=>"001001110",
  20197=>"111101000",
  20198=>"111111100",
  20199=>"000000000",
  20200=>"000000110",
  20201=>"111100100",
  20202=>"011000100",
  20203=>"011000010",
  20204=>"000000111",
  20205=>"111111010",
  20206=>"111000110",
  20207=>"000100111",
  20208=>"111110100",
  20209=>"111110100",
  20210=>"000000111",
  20211=>"111011100",
  20212=>"111011001",
  20213=>"001000000",
  20214=>"011111011",
  20215=>"000000000",
  20216=>"000000111",
  20217=>"000001111",
  20218=>"100000110",
  20219=>"000111111",
  20220=>"111111111",
  20221=>"000111011",
  20222=>"111111110",
  20223=>"111001001",
  20224=>"000000000",
  20225=>"111011011",
  20226=>"000000011",
  20227=>"001010000",
  20228=>"000111101",
  20229=>"101000000",
  20230=>"000000111",
  20231=>"100101111",
  20232=>"111111000",
  20233=>"001000001",
  20234=>"000000000",
  20235=>"000111111",
  20236=>"000000111",
  20237=>"111111101",
  20238=>"111111111",
  20239=>"111111000",
  20240=>"101100100",
  20241=>"011110000",
  20242=>"110110000",
  20243=>"000000000",
  20244=>"111111111",
  20245=>"000000111",
  20246=>"000000001",
  20247=>"001001111",
  20248=>"111111011",
  20249=>"111001001",
  20250=>"000000000",
  20251=>"000000000",
  20252=>"011000001",
  20253=>"010010000",
  20254=>"000000000",
  20255=>"001000000",
  20256=>"001001000",
  20257=>"000000111",
  20258=>"110110111",
  20259=>"111111110",
  20260=>"101000100",
  20261=>"100111000",
  20262=>"111111110",
  20263=>"111111100",
  20264=>"111111111",
  20265=>"000010011",
  20266=>"000000000",
  20267=>"111101000",
  20268=>"101000000",
  20269=>"000000100",
  20270=>"111111111",
  20271=>"000001101",
  20272=>"111111111",
  20273=>"110111011",
  20274=>"000000000",
  20275=>"111000000",
  20276=>"111000000",
  20277=>"000010000",
  20278=>"111111000",
  20279=>"111111011",
  20280=>"000000010",
  20281=>"111001111",
  20282=>"011111111",
  20283=>"000000111",
  20284=>"110110110",
  20285=>"000000110",
  20286=>"101111111",
  20287=>"111110111",
  20288=>"011000000",
  20289=>"111111000",
  20290=>"111010000",
  20291=>"000000111",
  20292=>"110000100",
  20293=>"110110011",
  20294=>"110000000",
  20295=>"000010110",
  20296=>"000000000",
  20297=>"000000111",
  20298=>"111011001",
  20299=>"111000000",
  20300=>"111110111",
  20301=>"110111111",
  20302=>"110111000",
  20303=>"000001001",
  20304=>"000000000",
  20305=>"000000111",
  20306=>"110111100",
  20307=>"000000000",
  20308=>"111111000",
  20309=>"001000001",
  20310=>"111111111",
  20311=>"000000001",
  20312=>"001111111",
  20313=>"000111001",
  20314=>"011011111",
  20315=>"000000111",
  20316=>"011001110",
  20317=>"100111111",
  20318=>"100100110",
  20319=>"111111001",
  20320=>"111110000",
  20321=>"000011111",
  20322=>"000000000",
  20323=>"100000000",
  20324=>"111111000",
  20325=>"000000111",
  20326=>"111111000",
  20327=>"100111111",
  20328=>"111100000",
  20329=>"000001111",
  20330=>"000000010",
  20331=>"000000011",
  20332=>"111111010",
  20333=>"111100100",
  20334=>"001000000",
  20335=>"011011111",
  20336=>"000000000",
  20337=>"000001000",
  20338=>"010100100",
  20339=>"000111111",
  20340=>"000111111",
  20341=>"101101111",
  20342=>"001001111",
  20343=>"000000000",
  20344=>"111111010",
  20345=>"000000111",
  20346=>"011111111",
  20347=>"111111111",
  20348=>"111101000",
  20349=>"110000000",
  20350=>"000110110",
  20351=>"000000000",
  20352=>"111110111",
  20353=>"111111111",
  20354=>"000000110",
  20355=>"000000000",
  20356=>"110000111",
  20357=>"000100000",
  20358=>"100100100",
  20359=>"111000000",
  20360=>"000110000",
  20361=>"101111111",
  20362=>"001000000",
  20363=>"111001000",
  20364=>"111111111",
  20365=>"000100110",
  20366=>"000001000",
  20367=>"000000101",
  20368=>"001000000",
  20369=>"000100111",
  20370=>"010011000",
  20371=>"111001011",
  20372=>"100101000",
  20373=>"001011000",
  20374=>"111111111",
  20375=>"101000100",
  20376=>"111000001",
  20377=>"001000001",
  20378=>"110111111",
  20379=>"000000110",
  20380=>"011111111",
  20381=>"010111111",
  20382=>"111111101",
  20383=>"111111111",
  20384=>"001000000",
  20385=>"011111111",
  20386=>"110011000",
  20387=>"111100000",
  20388=>"100000100",
  20389=>"000111111",
  20390=>"000000000",
  20391=>"111111111",
  20392=>"110111111",
  20393=>"110110000",
  20394=>"100000000",
  20395=>"111111011",
  20396=>"000011011",
  20397=>"111011010",
  20398=>"111001111",
  20399=>"111111111",
  20400=>"000100111",
  20401=>"111111111",
  20402=>"100101110",
  20403=>"000000111",
  20404=>"000000000",
  20405=>"110000000",
  20406=>"111101101",
  20407=>"110010000",
  20408=>"000000000",
  20409=>"111011111",
  20410=>"000001000",
  20411=>"111111111",
  20412=>"000110111",
  20413=>"111101111",
  20414=>"000000111",
  20415=>"001001111",
  20416=>"011011010",
  20417=>"000000110",
  20418=>"000000000",
  20419=>"000000000",
  20420=>"100100111",
  20421=>"111111101",
  20422=>"111111001",
  20423=>"000000000",
  20424=>"111100110",
  20425=>"111111001",
  20426=>"000110000",
  20427=>"000000111",
  20428=>"010000110",
  20429=>"111000000",
  20430=>"000000000",
  20431=>"111111000",
  20432=>"010110111",
  20433=>"111111000",
  20434=>"000000101",
  20435=>"010111111",
  20436=>"101101000",
  20437=>"000111111",
  20438=>"000000000",
  20439=>"011000000",
  20440=>"010000001",
  20441=>"111111010",
  20442=>"000001000",
  20443=>"000100000",
  20444=>"101111111",
  20445=>"111111111",
  20446=>"110111111",
  20447=>"001000001",
  20448=>"111011111",
  20449=>"000000001",
  20450=>"000001111",
  20451=>"000000111",
  20452=>"011011111",
  20453=>"000011100",
  20454=>"000000100",
  20455=>"011110010",
  20456=>"000011010",
  20457=>"101111110",
  20458=>"000000000",
  20459=>"000000110",
  20460=>"000111000",
  20461=>"110000000",
  20462=>"000000111",
  20463=>"000000010",
  20464=>"101101101",
  20465=>"101001111",
  20466=>"111111110",
  20467=>"111011001",
  20468=>"000000000",
  20469=>"010000000",
  20470=>"111110110",
  20471=>"100111100",
  20472=>"111100000",
  20473=>"100100100",
  20474=>"000000000",
  20475=>"111110110",
  20476=>"111111111",
  20477=>"000000000",
  20478=>"110110111",
  20479=>"001111111",
  20480=>"000000000",
  20481=>"110111000",
  20482=>"100100000",
  20483=>"000000000",
  20484=>"111111010",
  20485=>"000000000",
  20486=>"111111111",
  20487=>"000001111",
  20488=>"100101111",
  20489=>"111110110",
  20490=>"000000000",
  20491=>"000000000",
  20492=>"111011011",
  20493=>"000000011",
  20494=>"111111110",
  20495=>"001011000",
  20496=>"111111111",
  20497=>"000111111",
  20498=>"100100111",
  20499=>"011011011",
  20500=>"111111111",
  20501=>"000000111",
  20502=>"110110110",
  20503=>"100110000",
  20504=>"111111000",
  20505=>"111111111",
  20506=>"111111000",
  20507=>"001111111",
  20508=>"110100000",
  20509=>"111111111",
  20510=>"110110010",
  20511=>"010111111",
  20512=>"000000000",
  20513=>"000100110",
  20514=>"000000000",
  20515=>"111111111",
  20516=>"110111100",
  20517=>"100110111",
  20518=>"000000000",
  20519=>"111111111",
  20520=>"100110000",
  20521=>"100000100",
  20522=>"001000000",
  20523=>"111111000",
  20524=>"111110000",
  20525=>"000000000",
  20526=>"111000101",
  20527=>"111110011",
  20528=>"000100100",
  20529=>"000000101",
  20530=>"010100000",
  20531=>"000100000",
  20532=>"011000000",
  20533=>"110110000",
  20534=>"110100000",
  20535=>"101101100",
  20536=>"111111111",
  20537=>"000110011",
  20538=>"000001111",
  20539=>"001011011",
  20540=>"000000000",
  20541=>"000000000",
  20542=>"111111111",
  20543=>"000000000",
  20544=>"011111000",
  20545=>"111100110",
  20546=>"110111111",
  20547=>"110000000",
  20548=>"000111111",
  20549=>"000000110",
  20550=>"110111001",
  20551=>"001000011",
  20552=>"111011110",
  20553=>"111101000",
  20554=>"010000111",
  20555=>"111111111",
  20556=>"111111000",
  20557=>"000110111",
  20558=>"111111111",
  20559=>"000111111",
  20560=>"000000111",
  20561=>"000000000",
  20562=>"000000001",
  20563=>"000100100",
  20564=>"111111000",
  20565=>"100100000",
  20566=>"001000000",
  20567=>"000000111",
  20568=>"111111000",
  20569=>"111101000",
  20570=>"011111110",
  20571=>"000011111",
  20572=>"010000000",
  20573=>"000000000",
  20574=>"110100000",
  20575=>"000000000",
  20576=>"111000000",
  20577=>"111111000",
  20578=>"111111111",
  20579=>"000000000",
  20580=>"111111000",
  20581=>"000000000",
  20582=>"110110011",
  20583=>"100111111",
  20584=>"111100000",
  20585=>"000000000",
  20586=>"111000000",
  20587=>"111000000",
  20588=>"111101011",
  20589=>"111111111",
  20590=>"000000000",
  20591=>"111111111",
  20592=>"111100000",
  20593=>"000000000",
  20594=>"000000011",
  20595=>"000000001",
  20596=>"000000000",
  20597=>"100111000",
  20598=>"110010000",
  20599=>"100100000",
  20600=>"111110110",
  20601=>"111111111",
  20602=>"000000001",
  20603=>"000011111",
  20604=>"100000011",
  20605=>"000000000",
  20606=>"111111111",
  20607=>"001001000",
  20608=>"000011111",
  20609=>"000000000",
  20610=>"000001111",
  20611=>"111110100",
  20612=>"000000100",
  20613=>"111101111",
  20614=>"000001111",
  20615=>"111111110",
  20616=>"001111111",
  20617=>"011111011",
  20618=>"111111111",
  20619=>"111111100",
  20620=>"001001001",
  20621=>"000000000",
  20622=>"111011111",
  20623=>"100000111",
  20624=>"111111111",
  20625=>"000000000",
  20626=>"110111111",
  20627=>"000000000",
  20628=>"010000000",
  20629=>"000100110",
  20630=>"111111111",
  20631=>"000000000",
  20632=>"101001000",
  20633=>"011001111",
  20634=>"000000000",
  20635=>"000000111",
  20636=>"111111000",
  20637=>"110101111",
  20638=>"111111110",
  20639=>"110011001",
  20640=>"100000111",
  20641=>"111111111",
  20642=>"000000000",
  20643=>"000111111",
  20644=>"111111111",
  20645=>"101101111",
  20646=>"001001111",
  20647=>"000001001",
  20648=>"101010111",
  20649=>"100111011",
  20650=>"111111111",
  20651=>"111000000",
  20652=>"000110111",
  20653=>"110111111",
  20654=>"111111000",
  20655=>"111111111",
  20656=>"111111111",
  20657=>"011111111",
  20658=>"110111111",
  20659=>"001000000",
  20660=>"110011011",
  20661=>"111111111",
  20662=>"011011111",
  20663=>"111111111",
  20664=>"000000100",
  20665=>"111111111",
  20666=>"000000000",
  20667=>"110110111",
  20668=>"000000000",
  20669=>"111111111",
  20670=>"111111111",
  20671=>"000100000",
  20672=>"111111111",
  20673=>"000001000",
  20674=>"111111111",
  20675=>"000000000",
  20676=>"111111111",
  20677=>"000000000",
  20678=>"111111111",
  20679=>"010000000",
  20680=>"000000000",
  20681=>"111001111",
  20682=>"000000001",
  20683=>"000011111",
  20684=>"000000000",
  20685=>"000000000",
  20686=>"000000000",
  20687=>"000000000",
  20688=>"010111111",
  20689=>"000110111",
  20690=>"000010010",
  20691=>"101000001",
  20692=>"000100000",
  20693=>"111111110",
  20694=>"000000010",
  20695=>"111111000",
  20696=>"111010000",
  20697=>"000000000",
  20698=>"111111111",
  20699=>"000011111",
  20700=>"100000000",
  20701=>"111111111",
  20702=>"000000000",
  20703=>"000000100",
  20704=>"111100100",
  20705=>"111111110",
  20706=>"111111101",
  20707=>"000000111",
  20708=>"111111111",
  20709=>"010011000",
  20710=>"111111111",
  20711=>"000000111",
  20712=>"111111111",
  20713=>"001001001",
  20714=>"110111011",
  20715=>"000000100",
  20716=>"000000101",
  20717=>"111111110",
  20718=>"111000000",
  20719=>"000000111",
  20720=>"001111111",
  20721=>"000000000",
  20722=>"111111111",
  20723=>"110110110",
  20724=>"001011111",
  20725=>"000000000",
  20726=>"000101000",
  20727=>"000001001",
  20728=>"111111111",
  20729=>"110000000",
  20730=>"111000000",
  20731=>"000000000",
  20732=>"110100110",
  20733=>"100111111",
  20734=>"000000111",
  20735=>"000000000",
  20736=>"011000000",
  20737=>"000000001",
  20738=>"001000010",
  20739=>"000000100",
  20740=>"001011111",
  20741=>"111001000",
  20742=>"000000000",
  20743=>"111000111",
  20744=>"100000000",
  20745=>"000000111",
  20746=>"110111011",
  20747=>"111111000",
  20748=>"000000000",
  20749=>"011011010",
  20750=>"111111000",
  20751=>"101111111",
  20752=>"111111110",
  20753=>"111111111",
  20754=>"000000000",
  20755=>"000010100",
  20756=>"101101101",
  20757=>"111111101",
  20758=>"000100000",
  20759=>"010000111",
  20760=>"000001000",
  20761=>"010111111",
  20762=>"111111110",
  20763=>"111111110",
  20764=>"100100000",
  20765=>"000000101",
  20766=>"100000100",
  20767=>"000000000",
  20768=>"000000000",
  20769=>"000000111",
  20770=>"000101111",
  20771=>"000000000",
  20772=>"101100000",
  20773=>"001000000",
  20774=>"000000010",
  20775=>"111000100",
  20776=>"000001001",
  20777=>"110111111",
  20778=>"000000001",
  20779=>"111110010",
  20780=>"000000000",
  20781=>"000010110",
  20782=>"000000000",
  20783=>"110000000",
  20784=>"000000101",
  20785=>"000000000",
  20786=>"110110110",
  20787=>"000000101",
  20788=>"000000000",
  20789=>"000000001",
  20790=>"000000100",
  20791=>"000000000",
  20792=>"000000000",
  20793=>"111111001",
  20794=>"011011011",
  20795=>"111111001",
  20796=>"000000001",
  20797=>"000000111",
  20798=>"000000000",
  20799=>"000000100",
  20800=>"111111111",
  20801=>"000000000",
  20802=>"001000000",
  20803=>"001101111",
  20804=>"100111111",
  20805=>"100110110",
  20806=>"111111111",
  20807=>"000000111",
  20808=>"011010011",
  20809=>"000111001",
  20810=>"000001000",
  20811=>"100011011",
  20812=>"101111011",
  20813=>"000000000",
  20814=>"001000000",
  20815=>"000110110",
  20816=>"110111111",
  20817=>"000110111",
  20818=>"010000000",
  20819=>"110110111",
  20820=>"101011000",
  20821=>"001011111",
  20822=>"000000111",
  20823=>"111111100",
  20824=>"111111111",
  20825=>"001011111",
  20826=>"000101111",
  20827=>"111111000",
  20828=>"100000000",
  20829=>"000000000",
  20830=>"011001011",
  20831=>"000000001",
  20832=>"111111111",
  20833=>"110000000",
  20834=>"001001011",
  20835=>"000000111",
  20836=>"111111111",
  20837=>"000000001",
  20838=>"011000000",
  20839=>"000000000",
  20840=>"011000011",
  20841=>"111111111",
  20842=>"000000000",
  20843=>"110110011",
  20844=>"011011001",
  20845=>"000110111",
  20846=>"111000000",
  20847=>"000000000",
  20848=>"000000000",
  20849=>"000000000",
  20850=>"111101111",
  20851=>"001000100",
  20852=>"000000111",
  20853=>"000000000",
  20854=>"000100110",
  20855=>"000100000",
  20856=>"111101111",
  20857=>"111111100",
  20858=>"111111111",
  20859=>"100110111",
  20860=>"111000000",
  20861=>"111111111",
  20862=>"010010000",
  20863=>"111111111",
  20864=>"111111001",
  20865=>"000000000",
  20866=>"000000111",
  20867=>"000000011",
  20868=>"000111010",
  20869=>"111111111",
  20870=>"100111000",
  20871=>"111011001",
  20872=>"011011000",
  20873=>"001011011",
  20874=>"011001001",
  20875=>"111101101",
  20876=>"101101111",
  20877=>"001001000",
  20878=>"110110000",
  20879=>"000001000",
  20880=>"111111111",
  20881=>"000000001",
  20882=>"111111001",
  20883=>"000000111",
  20884=>"111101100",
  20885=>"000100111",
  20886=>"001001001",
  20887=>"010000111",
  20888=>"111111111",
  20889=>"000000010",
  20890=>"110111111",
  20891=>"111111111",
  20892=>"001000110",
  20893=>"111000000",
  20894=>"010111000",
  20895=>"111111000",
  20896=>"000011110",
  20897=>"000000111",
  20898=>"111011000",
  20899=>"000111111",
  20900=>"000000000",
  20901=>"100101111",
  20902=>"001111111",
  20903=>"010000000",
  20904=>"111111000",
  20905=>"111110100",
  20906=>"111111111",
  20907=>"111110110",
  20908=>"000000000",
  20909=>"000000011",
  20910=>"000000000",
  20911=>"000000000",
  20912=>"110111111",
  20913=>"111110000",
  20914=>"111100100",
  20915=>"000000000",
  20916=>"001111111",
  20917=>"000000000",
  20918=>"001000110",
  20919=>"111111111",
  20920=>"111101000",
  20921=>"110110010",
  20922=>"001111111",
  20923=>"000000000",
  20924=>"000000000",
  20925=>"111111111",
  20926=>"111111111",
  20927=>"111111111",
  20928=>"110000111",
  20929=>"111111111",
  20930=>"111111010",
  20931=>"000000000",
  20932=>"111000001",
  20933=>"110110111",
  20934=>"110111111",
  20935=>"000010000",
  20936=>"000000000",
  20937=>"111001000",
  20938=>"000000111",
  20939=>"111100001",
  20940=>"111000000",
  20941=>"110110000",
  20942=>"010111100",
  20943=>"000111000",
  20944=>"111101111",
  20945=>"111111111",
  20946=>"110111111",
  20947=>"000000000",
  20948=>"011011111",
  20949=>"111111111",
  20950=>"000000000",
  20951=>"110110110",
  20952=>"011111111",
  20953=>"000000011",
  20954=>"000000000",
  20955=>"001000000",
  20956=>"110111111",
  20957=>"111000000",
  20958=>"000000001",
  20959=>"000000100",
  20960=>"100100110",
  20961=>"000000000",
  20962=>"000000100",
  20963=>"000000000",
  20964=>"000000000",
  20965=>"011010000",
  20966=>"111111111",
  20967=>"111000100",
  20968=>"111001100",
  20969=>"111111111",
  20970=>"011010000",
  20971=>"110000000",
  20972=>"111011101",
  20973=>"000000010",
  20974=>"000000000",
  20975=>"100111111",
  20976=>"111011111",
  20977=>"000000111",
  20978=>"111111100",
  20979=>"000011111",
  20980=>"111111111",
  20981=>"000010001",
  20982=>"001000000",
  20983=>"110110100",
  20984=>"111111011",
  20985=>"111111010",
  20986=>"001001111",
  20987=>"111111000",
  20988=>"000000000",
  20989=>"111110011",
  20990=>"001000000",
  20991=>"111111111",
  20992=>"111101000",
  20993=>"010111111",
  20994=>"000000000",
  20995=>"111111111",
  20996=>"110111111",
  20997=>"010110011",
  20998=>"000000000",
  20999=>"111111111",
  21000=>"110000010",
  21001=>"000000111",
  21002=>"000101111",
  21003=>"000000111",
  21004=>"000100000",
  21005=>"011000000",
  21006=>"100100100",
  21007=>"000110110",
  21008=>"000000000",
  21009=>"000000111",
  21010=>"111010000",
  21011=>"111100100",
  21012=>"010111111",
  21013=>"111111010",
  21014=>"010010000",
  21015=>"101101111",
  21016=>"000001111",
  21017=>"111111111",
  21018=>"111000000",
  21019=>"010110110",
  21020=>"111111001",
  21021=>"011011111",
  21022=>"000000001",
  21023=>"000000000",
  21024=>"111110000",
  21025=>"111111111",
  21026=>"111111100",
  21027=>"101001011",
  21028=>"100110100",
  21029=>"110111001",
  21030=>"000001111",
  21031=>"000000001",
  21032=>"000001001",
  21033=>"000000000",
  21034=>"111111111",
  21035=>"110110110",
  21036=>"111110110",
  21037=>"100100110",
  21038=>"000010011",
  21039=>"101000000",
  21040=>"111111111",
  21041=>"000000000",
  21042=>"000000000",
  21043=>"110100000",
  21044=>"111011000",
  21045=>"000000000",
  21046=>"000110100",
  21047=>"001111010",
  21048=>"111001011",
  21049=>"010110111",
  21050=>"111001000",
  21051=>"000001011",
  21052=>"111000000",
  21053=>"001111001",
  21054=>"111101000",
  21055=>"000000111",
  21056=>"001000000",
  21057=>"000000111",
  21058=>"000000000",
  21059=>"000000000",
  21060=>"000001000",
  21061=>"111111110",
  21062=>"000111101",
  21063=>"010000000",
  21064=>"000100000",
  21065=>"111000000",
  21066=>"111111111",
  21067=>"101011001",
  21068=>"000011011",
  21069=>"000000000",
  21070=>"000000001",
  21071=>"001111111",
  21072=>"010111110",
  21073=>"101111111",
  21074=>"111110000",
  21075=>"001001001",
  21076=>"110111111",
  21077=>"000001000",
  21078=>"111111100",
  21079=>"011111000",
  21080=>"001001001",
  21081=>"000000000",
  21082=>"100000000",
  21083=>"001111111",
  21084=>"000111110",
  21085=>"000000000",
  21086=>"111100000",
  21087=>"000111111",
  21088=>"001111111",
  21089=>"000011011",
  21090=>"000000001",
  21091=>"111111111",
  21092=>"111101100",
  21093=>"000000000",
  21094=>"000111101",
  21095=>"000000000",
  21096=>"000111111",
  21097=>"101100000",
  21098=>"000111111",
  21099=>"111010000",
  21100=>"100000100",
  21101=>"000000111",
  21102=>"011111111",
  21103=>"000110111",
  21104=>"000111011",
  21105=>"111111111",
  21106=>"100000000",
  21107=>"000000000",
  21108=>"110000000",
  21109=>"001000001",
  21110=>"110000000",
  21111=>"000000000",
  21112=>"110000000",
  21113=>"011000000",
  21114=>"000000001",
  21115=>"111000000",
  21116=>"001000000",
  21117=>"100110100",
  21118=>"000000000",
  21119=>"000000000",
  21120=>"000100111",
  21121=>"111111000",
  21122=>"000000110",
  21123=>"000100000",
  21124=>"110111000",
  21125=>"111000000",
  21126=>"111111111",
  21127=>"000000000",
  21128=>"111000000",
  21129=>"000110110",
  21130=>"000000000",
  21131=>"111110100",
  21132=>"000000001",
  21133=>"110111000",
  21134=>"000001111",
  21135=>"110110110",
  21136=>"001000000",
  21137=>"000000000",
  21138=>"011010000",
  21139=>"000111110",
  21140=>"000110111",
  21141=>"110100000",
  21142=>"101000000",
  21143=>"111111111",
  21144=>"000000000",
  21145=>"101101001",
  21146=>"011011111",
  21147=>"000000000",
  21148=>"000111110",
  21149=>"000000000",
  21150=>"111011000",
  21151=>"000110010",
  21152=>"110010000",
  21153=>"001000100",
  21154=>"011111111",
  21155=>"100111111",
  21156=>"000000001",
  21157=>"111111111",
  21158=>"101101111",
  21159=>"000001001",
  21160=>"000000100",
  21161=>"000000100",
  21162=>"111111111",
  21163=>"111111111",
  21164=>"111000000",
  21165=>"110110011",
  21166=>"111111111",
  21167=>"000001001",
  21168=>"111111000",
  21169=>"111111111",
  21170=>"111111111",
  21171=>"111111111",
  21172=>"110111111",
  21173=>"001000000",
  21174=>"000011111",
  21175=>"000000000",
  21176=>"110000000",
  21177=>"111111000",
  21178=>"000000000",
  21179=>"111000000",
  21180=>"000000111",
  21181=>"000101011",
  21182=>"111001010",
  21183=>"110100100",
  21184=>"111111111",
  21185=>"000000001",
  21186=>"000100100",
  21187=>"000000000",
  21188=>"001011110",
  21189=>"111111001",
  21190=>"001000000",
  21191=>"000011101",
  21192=>"100000010",
  21193=>"111111000",
  21194=>"111111111",
  21195=>"000010000",
  21196=>"111000000",
  21197=>"001111111",
  21198=>"110111111",
  21199=>"111111111",
  21200=>"110111111",
  21201=>"110111111",
  21202=>"101111111",
  21203=>"000000000",
  21204=>"000000110",
  21205=>"111000000",
  21206=>"100100100",
  21207=>"111000001",
  21208=>"000000000",
  21209=>"011110100",
  21210=>"001000001",
  21211=>"011000000",
  21212=>"111110111",
  21213=>"000000111",
  21214=>"011011111",
  21215=>"110001000",
  21216=>"000000100",
  21217=>"000001111",
  21218=>"111111111",
  21219=>"000000000",
  21220=>"000000000",
  21221=>"110110111",
  21222=>"111111111",
  21223=>"000000000",
  21224=>"000111111",
  21225=>"100111111",
  21226=>"011111111",
  21227=>"000000001",
  21228=>"000101111",
  21229=>"111001000",
  21230=>"110100110",
  21231=>"000000000",
  21232=>"000000000",
  21233=>"111111111",
  21234=>"110000000",
  21235=>"000001000",
  21236=>"000000000",
  21237=>"000111111",
  21238=>"111100011",
  21239=>"011000000",
  21240=>"000000000",
  21241=>"110011000",
  21242=>"000000000",
  21243=>"001000110",
  21244=>"100000000",
  21245=>"011001001",
  21246=>"000000000",
  21247=>"110100000",
  21248=>"000110100",
  21249=>"001000001",
  21250=>"000110111",
  21251=>"111111110",
  21252=>"111000111",
  21253=>"000000010",
  21254=>"111000111",
  21255=>"000100111",
  21256=>"000000000",
  21257=>"000000001",
  21258=>"000001011",
  21259=>"000000001",
  21260=>"111100000",
  21261=>"111111111",
  21262=>"111111111",
  21263=>"111111111",
  21264=>"000000000",
  21265=>"100100000",
  21266=>"101000000",
  21267=>"000100000",
  21268=>"000000000",
  21269=>"010001111",
  21270=>"001001001",
  21271=>"111111110",
  21272=>"001001111",
  21273=>"000000000",
  21274=>"000010111",
  21275=>"111110110",
  21276=>"110111111",
  21277=>"000111111",
  21278=>"000110110",
  21279=>"010110000",
  21280=>"110110000",
  21281=>"000001001",
  21282=>"111111111",
  21283=>"111100100",
  21284=>"000001000",
  21285=>"000000000",
  21286=>"111000000",
  21287=>"111111111",
  21288=>"110111111",
  21289=>"001111111",
  21290=>"111010011",
  21291=>"010000010",
  21292=>"000000000",
  21293=>"111011111",
  21294=>"000000111",
  21295=>"000001001",
  21296=>"110111111",
  21297=>"000000000",
  21298=>"111111111",
  21299=>"111000000",
  21300=>"000000000",
  21301=>"111010000",
  21302=>"010000000",
  21303=>"010110111",
  21304=>"001011000",
  21305=>"000000000",
  21306=>"110111111",
  21307=>"000111100",
  21308=>"111111000",
  21309=>"000000000",
  21310=>"110110110",
  21311=>"010111111",
  21312=>"101100101",
  21313=>"111111111",
  21314=>"000000000",
  21315=>"111000000",
  21316=>"000000000",
  21317=>"111111111",
  21318=>"000001011",
  21319=>"000000000",
  21320=>"000000000",
  21321=>"000110111",
  21322=>"110000001",
  21323=>"000000110",
  21324=>"110111111",
  21325=>"111111111",
  21326=>"000000000",
  21327=>"111000000",
  21328=>"000000000",
  21329=>"011111111",
  21330=>"111010000",
  21331=>"100000000",
  21332=>"000000000",
  21333=>"111001000",
  21334=>"111001010",
  21335=>"000000000",
  21336=>"111111111",
  21337=>"000000000",
  21338=>"111111111",
  21339=>"000101111",
  21340=>"111001001",
  21341=>"010111111",
  21342=>"000101111",
  21343=>"111111111",
  21344=>"111111111",
  21345=>"111000000",
  21346=>"000001101",
  21347=>"000010110",
  21348=>"111111000",
  21349=>"111100000",
  21350=>"111000000",
  21351=>"000000000",
  21352=>"100101011",
  21353=>"111011000",
  21354=>"000111111",
  21355=>"001111111",
  21356=>"000000000",
  21357=>"000111111",
  21358=>"100000100",
  21359=>"100100100",
  21360=>"000000111",
  21361=>"000100000",
  21362=>"000110010",
  21363=>"001011011",
  21364=>"000000000",
  21365=>"000000010",
  21366=>"000000000",
  21367=>"000000000",
  21368=>"000000000",
  21369=>"111011011",
  21370=>"111010000",
  21371=>"000000000",
  21372=>"000000111",
  21373=>"001001001",
  21374=>"000000000",
  21375=>"011111111",
  21376=>"000111111",
  21377=>"000000011",
  21378=>"111111111",
  21379=>"000000111",
  21380=>"000000000",
  21381=>"000000101",
  21382=>"111000000",
  21383=>"111000000",
  21384=>"000000001",
  21385=>"011011011",
  21386=>"000000000",
  21387=>"000111010",
  21388=>"111111111",
  21389=>"111111000",
  21390=>"111111000",
  21391=>"000000000",
  21392=>"010111110",
  21393=>"000000111",
  21394=>"111100000",
  21395=>"111110000",
  21396=>"111000000",
  21397=>"000000000",
  21398=>"111010000",
  21399=>"011111001",
  21400=>"001001000",
  21401=>"010111111",
  21402=>"111111111",
  21403=>"111110101",
  21404=>"101100100",
  21405=>"001000000",
  21406=>"111100000",
  21407=>"101000000",
  21408=>"010111111",
  21409=>"001110000",
  21410=>"011111111",
  21411=>"000000000",
  21412=>"111111101",
  21413=>"000110111",
  21414=>"000001111",
  21415=>"111010110",
  21416=>"110111111",
  21417=>"100000000",
  21418=>"111111010",
  21419=>"001000000",
  21420=>"000111111",
  21421=>"111100000",
  21422=>"000000000",
  21423=>"111110110",
  21424=>"111110111",
  21425=>"111111111",
  21426=>"111111111",
  21427=>"000011111",
  21428=>"000000000",
  21429=>"001001000",
  21430=>"110101000",
  21431=>"111000000",
  21432=>"111111000",
  21433=>"111111111",
  21434=>"111111110",
  21435=>"111111111",
  21436=>"111000000",
  21437=>"000110111",
  21438=>"000000000",
  21439=>"101100100",
  21440=>"000000000",
  21441=>"001000000",
  21442=>"000000001",
  21443=>"000000000",
  21444=>"111111110",
  21445=>"000001010",
  21446=>"111111111",
  21447=>"001000000",
  21448=>"000101101",
  21449=>"000000000",
  21450=>"100111011",
  21451=>"111011111",
  21452=>"101001101",
  21453=>"111111111",
  21454=>"101111111",
  21455=>"000000010",
  21456=>"101000010",
  21457=>"011011011",
  21458=>"111110110",
  21459=>"111000000",
  21460=>"001001111",
  21461=>"111000100",
  21462=>"111111110",
  21463=>"001011011",
  21464=>"111000000",
  21465=>"111111011",
  21466=>"000100111",
  21467=>"000000000",
  21468=>"100100000",
  21469=>"011111111",
  21470=>"110110111",
  21471=>"000000011",
  21472=>"111111111",
  21473=>"000000000",
  21474=>"000000000",
  21475=>"001111100",
  21476=>"111111111",
  21477=>"110000000",
  21478=>"000000000",
  21479=>"000000000",
  21480=>"011001000",
  21481=>"010011111",
  21482=>"111000000",
  21483=>"000000100",
  21484=>"100100100",
  21485=>"101111111",
  21486=>"111111111",
  21487=>"000011111",
  21488=>"010000000",
  21489=>"000000000",
  21490=>"111100100",
  21491=>"111111111",
  21492=>"111001000",
  21493=>"000011111",
  21494=>"000000000",
  21495=>"000001001",
  21496=>"000000010",
  21497=>"111111100",
  21498=>"110111111",
  21499=>"000000000",
  21500=>"110100101",
  21501=>"011011111",
  21502=>"110011000",
  21503=>"100000000",
  21504=>"111111110",
  21505=>"001000111",
  21506=>"111111111",
  21507=>"110111100",
  21508=>"001000100",
  21509=>"111111111",
  21510=>"000000000",
  21511=>"000000000",
  21512=>"000000000",
  21513=>"110110111",
  21514=>"000000000",
  21515=>"111111111",
  21516=>"000000110",
  21517=>"111000000",
  21518=>"000000000",
  21519=>"000000000",
  21520=>"001111111",
  21521=>"000000110",
  21522=>"000000101",
  21523=>"111111111",
  21524=>"111111111",
  21525=>"111111111",
  21526=>"111111111",
  21527=>"001000000",
  21528=>"111111110",
  21529=>"111111111",
  21530=>"100111111",
  21531=>"000000000",
  21532=>"111111111",
  21533=>"111001110",
  21534=>"011011011",
  21535=>"111111111",
  21536=>"111111111",
  21537=>"100111111",
  21538=>"111111110",
  21539=>"101100101",
  21540=>"111111111",
  21541=>"000000111",
  21542=>"111111111",
  21543=>"000000001",
  21544=>"111111111",
  21545=>"000000000",
  21546=>"000000000",
  21547=>"010000000",
  21548=>"001111111",
  21549=>"101110100",
  21550=>"001001101",
  21551=>"111110000",
  21552=>"001001101",
  21553=>"000000000",
  21554=>"100000100",
  21555=>"111010000",
  21556=>"111111001",
  21557=>"000000010",
  21558=>"000001111",
  21559=>"111110111",
  21560=>"000000111",
  21561=>"111111111",
  21562=>"000000000",
  21563=>"000000101",
  21564=>"100100111",
  21565=>"000010010",
  21566=>"100000010",
  21567=>"000000111",
  21568=>"111111000",
  21569=>"011111001",
  21570=>"111100100",
  21571=>"111111111",
  21572=>"000010111",
  21573=>"000000000",
  21574=>"111000000",
  21575=>"111111011",
  21576=>"011111111",
  21577=>"000000000",
  21578=>"111111111",
  21579=>"000001000",
  21580=>"000000101",
  21581=>"100000000",
  21582=>"000000001",
  21583=>"000000000",
  21584=>"000000000",
  21585=>"100010000",
  21586=>"000000000",
  21587=>"110110100",
  21588=>"000000000",
  21589=>"001001111",
  21590=>"001000000",
  21591=>"000000101",
  21592=>"001001001",
  21593=>"001000000",
  21594=>"000101111",
  21595=>"000000000",
  21596=>"011000100",
  21597=>"111111111",
  21598=>"000000000",
  21599=>"100000000",
  21600=>"001001001",
  21601=>"001110110",
  21602=>"010010111",
  21603=>"111111000",
  21604=>"111111000",
  21605=>"111111111",
  21606=>"110100100",
  21607=>"000000001",
  21608=>"111000101",
  21609=>"000000111",
  21610=>"100000000",
  21611=>"000000000",
  21612=>"001001001",
  21613=>"111011000",
  21614=>"000000000",
  21615=>"000110011",
  21616=>"000000100",
  21617=>"000000100",
  21618=>"101101101",
  21619=>"000000101",
  21620=>"000000000",
  21621=>"111111000",
  21622=>"001101101",
  21623=>"000000000",
  21624=>"010000000",
  21625=>"000000000",
  21626=>"001000000",
  21627=>"111111111",
  21628=>"100110100",
  21629=>"111101001",
  21630=>"111001000",
  21631=>"111111111",
  21632=>"001111000",
  21633=>"000000000",
  21634=>"111111000",
  21635=>"011011011",
  21636=>"000000000",
  21637=>"111111111",
  21638=>"111111110",
  21639=>"000101111",
  21640=>"100110011",
  21641=>"101111111",
  21642=>"100111111",
  21643=>"000000001",
  21644=>"000000000",
  21645=>"111011000",
  21646=>"100111111",
  21647=>"011000000",
  21648=>"111101111",
  21649=>"000000000",
  21650=>"000000000",
  21651=>"110010100",
  21652=>"101000000",
  21653=>"000000000",
  21654=>"000000000",
  21655=>"001101111",
  21656=>"000000000",
  21657=>"100000100",
  21658=>"001111111",
  21659=>"000000000",
  21660=>"111111111",
  21661=>"000000100",
  21662=>"010010000",
  21663=>"111111111",
  21664=>"000000000",
  21665=>"001001111",
  21666=>"101101111",
  21667=>"111111001",
  21668=>"011000000",
  21669=>"010000000",
  21670=>"111111111",
  21671=>"000011011",
  21672=>"000000100",
  21673=>"001111111",
  21674=>"111100000",
  21675=>"000000000",
  21676=>"000000001",
  21677=>"011111110",
  21678=>"111111111",
  21679=>"111111111",
  21680=>"011001101",
  21681=>"011000010",
  21682=>"111111111",
  21683=>"001000000",
  21684=>"111000000",
  21685=>"000011111",
  21686=>"101000000",
  21687=>"111001000",
  21688=>"111101000",
  21689=>"000000000",
  21690=>"111101000",
  21691=>"000000000",
  21692=>"111000000",
  21693=>"000000000",
  21694=>"111111100",
  21695=>"111111111",
  21696=>"110111111",
  21697=>"000000000",
  21698=>"100111111",
  21699=>"000001111",
  21700=>"000000000",
  21701=>"111111111",
  21702=>"110100101",
  21703=>"000000000",
  21704=>"000111111",
  21705=>"111111111",
  21706=>"011011000",
  21707=>"011000011",
  21708=>"000111111",
  21709=>"000000000",
  21710=>"101000001",
  21711=>"110110110",
  21712=>"000000000",
  21713=>"011111111",
  21714=>"101011111",
  21715=>"111111111",
  21716=>"111111001",
  21717=>"000000010",
  21718=>"000000111",
  21719=>"100110111",
  21720=>"111111111",
  21721=>"111111101",
  21722=>"000000000",
  21723=>"111111111",
  21724=>"111111001",
  21725=>"001001001",
  21726=>"000000000",
  21727=>"111111111",
  21728=>"000000100",
  21729=>"111111011",
  21730=>"111000000",
  21731=>"010111111",
  21732=>"000000000",
  21733=>"000000000",
  21734=>"110100000",
  21735=>"111111111",
  21736=>"000000000",
  21737=>"000000111",
  21738=>"111000110",
  21739=>"000000111",
  21740=>"111111111",
  21741=>"111111111",
  21742=>"000000100",
  21743=>"111001000",
  21744=>"111111111",
  21745=>"100100000",
  21746=>"111111111",
  21747=>"000000001",
  21748=>"000101111",
  21749=>"111011000",
  21750=>"011111111",
  21751=>"101000101",
  21752=>"111000000",
  21753=>"111111111",
  21754=>"000000011",
  21755=>"111111111",
  21756=>"000000111",
  21757=>"111111111",
  21758=>"111111000",
  21759=>"110111111",
  21760=>"000000000",
  21761=>"101000100",
  21762=>"110110110",
  21763=>"111111110",
  21764=>"001000000",
  21765=>"000000000",
  21766=>"001001000",
  21767=>"001001001",
  21768=>"000000000",
  21769=>"101000000",
  21770=>"000000000",
  21771=>"000000100",
  21772=>"101000001",
  21773=>"000000000",
  21774=>"000000000",
  21775=>"111110000",
  21776=>"111111111",
  21777=>"000000111",
  21778=>"000001111",
  21779=>"111011011",
  21780=>"111111011",
  21781=>"111011111",
  21782=>"111111100",
  21783=>"111111111",
  21784=>"001111011",
  21785=>"101001001",
  21786=>"000000000",
  21787=>"111111100",
  21788=>"001001001",
  21789=>"001011111",
  21790=>"000001001",
  21791=>"101101111",
  21792=>"110111111",
  21793=>"000000111",
  21794=>"010010001",
  21795=>"010011111",
  21796=>"000000000",
  21797=>"111111111",
  21798=>"010011011",
  21799=>"110101101",
  21800=>"101000000",
  21801=>"000000000",
  21802=>"000011011",
  21803=>"000110000",
  21804=>"000000000",
  21805=>"111000111",
  21806=>"000000110",
  21807=>"000000000",
  21808=>"110110110",
  21809=>"000000000",
  21810=>"111000000",
  21811=>"000000000",
  21812=>"111111111",
  21813=>"111111111",
  21814=>"101000111",
  21815=>"001000000",
  21816=>"001000001",
  21817=>"011000111",
  21818=>"000000000",
  21819=>"111000110",
  21820=>"111111111",
  21821=>"000001101",
  21822=>"100110111",
  21823=>"111111011",
  21824=>"000000111",
  21825=>"111111100",
  21826=>"000000100",
  21827=>"000110111",
  21828=>"111111111",
  21829=>"111111111",
  21830=>"110110111",
  21831=>"000000000",
  21832=>"000000000",
  21833=>"000000111",
  21834=>"111001000",
  21835=>"001111111",
  21836=>"001000011",
  21837=>"111011111",
  21838=>"000000000",
  21839=>"110110110",
  21840=>"011111000",
  21841=>"000000000",
  21842=>"010110000",
  21843=>"000000111",
  21844=>"111100000",
  21845=>"011011001",
  21846=>"111111001",
  21847=>"000000111",
  21848=>"000000111",
  21849=>"111001000",
  21850=>"000000000",
  21851=>"111111111",
  21852=>"000000001",
  21853=>"111111100",
  21854=>"001000001",
  21855=>"001001000",
  21856=>"000000111",
  21857=>"001101111",
  21858=>"100000000",
  21859=>"111111111",
  21860=>"011011011",
  21861=>"000000111",
  21862=>"111111111",
  21863=>"000000000",
  21864=>"000110111",
  21865=>"000000111",
  21866=>"000001111",
  21867=>"111101011",
  21868=>"000100110",
  21869=>"000000000",
  21870=>"111100000",
  21871=>"001000000",
  21872=>"000000111",
  21873=>"000000000",
  21874=>"111111111",
  21875=>"000000000",
  21876=>"000000000",
  21877=>"001111111",
  21878=>"111111111",
  21879=>"000000000",
  21880=>"000111111",
  21881=>"000000110",
  21882=>"001000001",
  21883=>"110110010",
  21884=>"101111111",
  21885=>"000000000",
  21886=>"111111111",
  21887=>"100000111",
  21888=>"000000000",
  21889=>"000000000",
  21890=>"000000000",
  21891=>"001001101",
  21892=>"111110000",
  21893=>"000000110",
  21894=>"000000100",
  21895=>"110110111",
  21896=>"000000101",
  21897=>"111111111",
  21898=>"000000000",
  21899=>"001111111",
  21900=>"101111111",
  21901=>"111111111",
  21902=>"111111000",
  21903=>"000000000",
  21904=>"000000000",
  21905=>"100000100",
  21906=>"111001101",
  21907=>"111111111",
  21908=>"000101101",
  21909=>"111110010",
  21910=>"000000001",
  21911=>"001000100",
  21912=>"111111111",
  21913=>"000001110",
  21914=>"000000000",
  21915=>"111111111",
  21916=>"111111111",
  21917=>"111111111",
  21918=>"000000001",
  21919=>"000000000",
  21920=>"010111000",
  21921=>"000000001",
  21922=>"111111001",
  21923=>"000000000",
  21924=>"100110000",
  21925=>"001111111",
  21926=>"001111111",
  21927=>"000000000",
  21928=>"000000000",
  21929=>"000001000",
  21930=>"101111111",
  21931=>"001000000",
  21932=>"011000000",
  21933=>"000100000",
  21934=>"111111001",
  21935=>"111111101",
  21936=>"101000111",
  21937=>"110110111",
  21938=>"000000000",
  21939=>"000000011",
  21940=>"101001001",
  21941=>"111111111",
  21942=>"111111111",
  21943=>"000000000",
  21944=>"000000111",
  21945=>"000000100",
  21946=>"100000100",
  21947=>"001001111",
  21948=>"000000101",
  21949=>"100000001",
  21950=>"000000000",
  21951=>"011011000",
  21952=>"000000100",
  21953=>"111111111",
  21954=>"011000010",
  21955=>"000000110",
  21956=>"000100101",
  21957=>"010000000",
  21958=>"111000000",
  21959=>"000000100",
  21960=>"001000001",
  21961=>"111111111",
  21962=>"111111111",
  21963=>"100100111",
  21964=>"101000000",
  21965=>"100111111",
  21966=>"000000000",
  21967=>"011011001",
  21968=>"000010000",
  21969=>"101000011",
  21970=>"111111001",
  21971=>"101001001",
  21972=>"110111110",
  21973=>"111001001",
  21974=>"000000011",
  21975=>"000001001",
  21976=>"001000111",
  21977=>"111111111",
  21978=>"111100101",
  21979=>"111111111",
  21980=>"111111111",
  21981=>"111111001",
  21982=>"111111011",
  21983=>"000000000",
  21984=>"000000001",
  21985=>"010000000",
  21986=>"000000000",
  21987=>"101100111",
  21988=>"000110011",
  21989=>"111111111",
  21990=>"111101111",
  21991=>"000000000",
  21992=>"000000000",
  21993=>"110111111",
  21994=>"000000000",
  21995=>"011011000",
  21996=>"001111111",
  21997=>"110110111",
  21998=>"000110111",
  21999=>"000000000",
  22000=>"000000000",
  22001=>"001111111",
  22002=>"000000001",
  22003=>"000110100",
  22004=>"101101111",
  22005=>"111111111",
  22006=>"010000000",
  22007=>"110011011",
  22008=>"000000100",
  22009=>"110110010",
  22010=>"011011011",
  22011=>"000000111",
  22012=>"000000100",
  22013=>"111111111",
  22014=>"100100111",
  22015=>"100100100",
  22016=>"010111111",
  22017=>"111111111",
  22018=>"000001111",
  22019=>"101111100",
  22020=>"010010010",
  22021=>"001011111",
  22022=>"000000000",
  22023=>"111111111",
  22024=>"111111111",
  22025=>"100100100",
  22026=>"111111111",
  22027=>"100110111",
  22028=>"010000110",
  22029=>"001001000",
  22030=>"000000000",
  22031=>"111111111",
  22032=>"101001001",
  22033=>"000001000",
  22034=>"000001000",
  22035=>"000000000",
  22036=>"111111111",
  22037=>"000000000",
  22038=>"111111111",
  22039=>"011011000",
  22040=>"110110111",
  22041=>"000000000",
  22042=>"001000011",
  22043=>"000000000",
  22044=>"010000000",
  22045=>"000000100",
  22046=>"000100000",
  22047=>"000010000",
  22048=>"111111111",
  22049=>"101101111",
  22050=>"110000000",
  22051=>"111111111",
  22052=>"001001001",
  22053=>"001000000",
  22054=>"111111111",
  22055=>"000000000",
  22056=>"111111111",
  22057=>"111111011",
  22058=>"000000001",
  22059=>"011010110",
  22060=>"111111000",
  22061=>"000110100",
  22062=>"011011011",
  22063=>"111001001",
  22064=>"001000010",
  22065=>"000010000",
  22066=>"000000000",
  22067=>"001001111",
  22068=>"110001000",
  22069=>"011011011",
  22070=>"110111111",
  22071=>"111011011",
  22072=>"000000000",
  22073=>"001000110",
  22074=>"000000000",
  22075=>"000011111",
  22076=>"111111111",
  22077=>"011000000",
  22078=>"011011111",
  22079=>"011000010",
  22080=>"011001001",
  22081=>"000000000",
  22082=>"000000001",
  22083=>"100000000",
  22084=>"000000000",
  22085=>"000000000",
  22086=>"000000011",
  22087=>"000100111",
  22088=>"000000010",
  22089=>"100100111",
  22090=>"000000111",
  22091=>"111011001",
  22092=>"000000111",
  22093=>"101000111",
  22094=>"000110111",
  22095=>"111111100",
  22096=>"111111111",
  22097=>"000000000",
  22098=>"000000000",
  22099=>"001111100",
  22100=>"011010010",
  22101=>"000010011",
  22102=>"111011011",
  22103=>"111111111",
  22104=>"110100100",
  22105=>"001000000",
  22106=>"000000001",
  22107=>"000000000",
  22108=>"000000010",
  22109=>"000000001",
  22110=>"000000000",
  22111=>"011100100",
  22112=>"000111111",
  22113=>"001111100",
  22114=>"000000000",
  22115=>"000000111",
  22116=>"000000000",
  22117=>"000000000",
  22118=>"000000000",
  22119=>"011011111",
  22120=>"111111111",
  22121=>"101000100",
  22122=>"110111111",
  22123=>"000000000",
  22124=>"100100000",
  22125=>"111111000",
  22126=>"101111111",
  22127=>"000001001",
  22128=>"111000111",
  22129=>"000000000",
  22130=>"010010110",
  22131=>"111111110",
  22132=>"001000000",
  22133=>"000000000",
  22134=>"000000111",
  22135=>"111101001",
  22136=>"100110100",
  22137=>"011000000",
  22138=>"001011001",
  22139=>"010110000",
  22140=>"000100111",
  22141=>"011010011",
  22142=>"111011001",
  22143=>"111111111",
  22144=>"111010010",
  22145=>"111111111",
  22146=>"111111111",
  22147=>"000001011",
  22148=>"001001000",
  22149=>"000000000",
  22150=>"001011000",
  22151=>"011011111",
  22152=>"111111111",
  22153=>"110001000",
  22154=>"110110110",
  22155=>"111111110",
  22156=>"000000000",
  22157=>"000100000",
  22158=>"000111111",
  22159=>"000000000",
  22160=>"111111111",
  22161=>"010111111",
  22162=>"011010011",
  22163=>"000001011",
  22164=>"011000000",
  22165=>"100111010",
  22166=>"010000000",
  22167=>"111111111",
  22168=>"111110111",
  22169=>"011010000",
  22170=>"001001000",
  22171=>"010000000",
  22172=>"111111111",
  22173=>"010011111",
  22174=>"111111001",
  22175=>"100100100",
  22176=>"000000111",
  22177=>"000111111",
  22178=>"000000010",
  22179=>"101101111",
  22180=>"001000000",
  22181=>"000000000",
  22182=>"111111111",
  22183=>"100100100",
  22184=>"100111111",
  22185=>"011111111",
  22186=>"111000000",
  22187=>"111110111",
  22188=>"000001011",
  22189=>"000000000",
  22190=>"101100000",
  22191=>"101101000",
  22192=>"111111111",
  22193=>"110100100",
  22194=>"111101111",
  22195=>"111101100",
  22196=>"111000000",
  22197=>"011000000",
  22198=>"001000000",
  22199=>"100100100",
  22200=>"100000000",
  22201=>"011111001",
  22202=>"011000000",
  22203=>"111011011",
  22204=>"000000000",
  22205=>"111111001",
  22206=>"101111111",
  22207=>"101001001",
  22208=>"011001000",
  22209=>"110010000",
  22210=>"110111111",
  22211=>"101001111",
  22212=>"001011011",
  22213=>"111111111",
  22214=>"111111111",
  22215=>"111000001",
  22216=>"111101111",
  22217=>"000000011",
  22218=>"000010111",
  22219=>"111111111",
  22220=>"000000111",
  22221=>"000000001",
  22222=>"101111100",
  22223=>"001000000",
  22224=>"000000000",
  22225=>"000000000",
  22226=>"000000000",
  22227=>"000000000",
  22228=>"010000000",
  22229=>"110110111",
  22230=>"000000010",
  22231=>"110110110",
  22232=>"011010000",
  22233=>"001000000",
  22234=>"000000000",
  22235=>"000000000",
  22236=>"111111000",
  22237=>"000000110",
  22238=>"000000000",
  22239=>"011000010",
  22240=>"110000000",
  22241=>"110111111",
  22242=>"000000000",
  22243=>"111111111",
  22244=>"001001000",
  22245=>"100001111",
  22246=>"000101111",
  22247=>"001000000",
  22248=>"000000111",
  22249=>"100100110",
  22250=>"000000110",
  22251=>"100100011",
  22252=>"000000111",
  22253=>"010111111",
  22254=>"110110111",
  22255=>"101111111",
  22256=>"111101111",
  22257=>"000000001",
  22258=>"000000000",
  22259=>"000000111",
  22260=>"001011111",
  22261=>"000000011",
  22262=>"000000000",
  22263=>"111111111",
  22264=>"111111111",
  22265=>"111011011",
  22266=>"000000111",
  22267=>"111011010",
  22268=>"001000000",
  22269=>"000000000",
  22270=>"000011000",
  22271=>"000011000",
  22272=>"010000110",
  22273=>"110110100",
  22274=>"000000111",
  22275=>"010000000",
  22276=>"110100010",
  22277=>"110111011",
  22278=>"101100000",
  22279=>"111111111",
  22280=>"111111111",
  22281=>"110010000",
  22282=>"000001000",
  22283=>"010010000",
  22284=>"001001111",
  22285=>"111000001",
  22286=>"111000011",
  22287=>"111111111",
  22288=>"000000011",
  22289=>"111111111",
  22290=>"000000000",
  22291=>"111011010",
  22292=>"111111111",
  22293=>"001001001",
  22294=>"000000000",
  22295=>"111111111",
  22296=>"101101100",
  22297=>"010110100",
  22298=>"000000000",
  22299=>"000001000",
  22300=>"100000000",
  22301=>"001011011",
  22302=>"000011011",
  22303=>"111111111",
  22304=>"000000010",
  22305=>"110000000",
  22306=>"000001001",
  22307=>"111111110",
  22308=>"000000000",
  22309=>"000000001",
  22310=>"101001011",
  22311=>"000011011",
  22312=>"111111010",
  22313=>"000000000",
  22314=>"111101111",
  22315=>"111111111",
  22316=>"000000100",
  22317=>"100100000",
  22318=>"000110100",
  22319=>"111111111",
  22320=>"111000011",
  22321=>"111000111",
  22322=>"111111111",
  22323=>"000000000",
  22324=>"111001111",
  22325=>"110011011",
  22326=>"111011011",
  22327=>"000000001",
  22328=>"110110111",
  22329=>"010000000",
  22330=>"111111111",
  22331=>"111100010",
  22332=>"100100000",
  22333=>"111000000",
  22334=>"011111111",
  22335=>"111111111",
  22336=>"000000000",
  22337=>"111101000",
  22338=>"001000111",
  22339=>"010011010",
  22340=>"111111111",
  22341=>"111111111",
  22342=>"111111111",
  22343=>"001101101",
  22344=>"000001001",
  22345=>"011111000",
  22346=>"001001011",
  22347=>"001001000",
  22348=>"000000000",
  22349=>"000000000",
  22350=>"001001111",
  22351=>"001001011",
  22352=>"000000001",
  22353=>"000000000",
  22354=>"111001111",
  22355=>"001001001",
  22356=>"000000000",
  22357=>"011111011",
  22358=>"000000000",
  22359=>"110110100",
  22360=>"001001000",
  22361=>"110100110",
  22362=>"000110111",
  22363=>"111111110",
  22364=>"000000000",
  22365=>"011111010",
  22366=>"111111101",
  22367=>"001001000",
  22368=>"000000000",
  22369=>"000000000",
  22370=>"000000000",
  22371=>"000000111",
  22372=>"001001000",
  22373=>"000000000",
  22374=>"000000000",
  22375=>"000010010",
  22376=>"000000000",
  22377=>"111100001",
  22378=>"000010110",
  22379=>"111111011",
  22380=>"000000000",
  22381=>"111111110",
  22382=>"010010110",
  22383=>"110100111",
  22384=>"001001011",
  22385=>"000000000",
  22386=>"111100100",
  22387=>"001001000",
  22388=>"000000000",
  22389=>"100111111",
  22390=>"010111111",
  22391=>"111111111",
  22392=>"000000001",
  22393=>"011111111",
  22394=>"000000001",
  22395=>"001011000",
  22396=>"100000000",
  22397=>"101001000",
  22398=>"000001000",
  22399=>"111001001",
  22400=>"111000000",
  22401=>"111011011",
  22402=>"001000000",
  22403=>"110100100",
  22404=>"010011011",
  22405=>"111111111",
  22406=>"000000111",
  22407=>"000000111",
  22408=>"111111101",
  22409=>"000110000",
  22410=>"101000000",
  22411=>"111111111",
  22412=>"111001001",
  22413=>"001000001",
  22414=>"001001001",
  22415=>"110000000",
  22416=>"000001111",
  22417=>"111110100",
  22418=>"011001111",
  22419=>"001001011",
  22420=>"111011010",
  22421=>"000110111",
  22422=>"000000000",
  22423=>"000000000",
  22424=>"111111111",
  22425=>"011011011",
  22426=>"111000000",
  22427=>"110111111",
  22428=>"001000000",
  22429=>"001001010",
  22430=>"111111111",
  22431=>"000000000",
  22432=>"000010111",
  22433=>"000000111",
  22434=>"101111000",
  22435=>"011011011",
  22436=>"101101000",
  22437=>"000000000",
  22438=>"100111111",
  22439=>"011000001",
  22440=>"110111110",
  22441=>"111111110",
  22442=>"000100111",
  22443=>"111111111",
  22444=>"000000011",
  22445=>"000000000",
  22446=>"000011001",
  22447=>"111111000",
  22448=>"000000001",
  22449=>"111111111",
  22450=>"011011110",
  22451=>"110010000",
  22452=>"111100111",
  22453=>"100100000",
  22454=>"010111110",
  22455=>"010110100",
  22456=>"000000100",
  22457=>"111111011",
  22458=>"001000000",
  22459=>"101001000",
  22460=>"111111111",
  22461=>"111111111",
  22462=>"111111111",
  22463=>"101000000",
  22464=>"111111011",
  22465=>"100000100",
  22466=>"001000010",
  22467=>"111111111",
  22468=>"000000000",
  22469=>"001011011",
  22470=>"000000011",
  22471=>"111111111",
  22472=>"101000111",
  22473=>"001000011",
  22474=>"011010111",
  22475=>"000000000",
  22476=>"000001100",
  22477=>"111111111",
  22478=>"001000000",
  22479=>"010000000",
  22480=>"111111111",
  22481=>"101101101",
  22482=>"000000000",
  22483=>"011111111",
  22484=>"000110000",
  22485=>"110110100",
  22486=>"001000000",
  22487=>"110110101",
  22488=>"000000000",
  22489=>"111111110",
  22490=>"000001001",
  22491=>"000000010",
  22492=>"001111111",
  22493=>"111011111",
  22494=>"111111111",
  22495=>"000100100",
  22496=>"110110100",
  22497=>"001011110",
  22498=>"111111111",
  22499=>"111111000",
  22500=>"001000000",
  22501=>"111111001",
  22502=>"110111111",
  22503=>"000000000",
  22504=>"000000010",
  22505=>"001001111",
  22506=>"000000000",
  22507=>"111111111",
  22508=>"000000000",
  22509=>"001001000",
  22510=>"110110110",
  22511=>"000000000",
  22512=>"111011111",
  22513=>"111001111",
  22514=>"000010000",
  22515=>"111111111",
  22516=>"001101111",
  22517=>"000000000",
  22518=>"000001000",
  22519=>"000000000",
  22520=>"111111011",
  22521=>"000001011",
  22522=>"010111110",
  22523=>"111111111",
  22524=>"000110110",
  22525=>"000000000",
  22526=>"001011010",
  22527=>"000000110",
  22528=>"001001000",
  22529=>"100110000",
  22530=>"000000000",
  22531=>"001000100",
  22532=>"000000111",
  22533=>"110111111",
  22534=>"111111111",
  22535=>"100000101",
  22536=>"000010111",
  22537=>"111111111",
  22538=>"111111000",
  22539=>"000000000",
  22540=>"110111010",
  22541=>"111100111",
  22542=>"111111111",
  22543=>"110111111",
  22544=>"010000000",
  22545=>"000111111",
  22546=>"000001111",
  22547=>"111100000",
  22548=>"111000100",
  22549=>"111010010",
  22550=>"000000000",
  22551=>"011011000",
  22552=>"111111111",
  22553=>"110101111",
  22554=>"111111111",
  22555=>"111011111",
  22556=>"000000000",
  22557=>"011111111",
  22558=>"000000101",
  22559=>"111111001",
  22560=>"000001001",
  22561=>"111111010",
  22562=>"110110111",
  22563=>"001001111",
  22564=>"000100111",
  22565=>"110101111",
  22566=>"000111111",
  22567=>"111100000",
  22568=>"111111111",
  22569=>"001000000",
  22570=>"111011000",
  22571=>"111111111",
  22572=>"000000000",
  22573=>"000110110",
  22574=>"001011001",
  22575=>"000000000",
  22576=>"000000000",
  22577=>"111001111",
  22578=>"000000000",
  22579=>"111011100",
  22580=>"001001011",
  22581=>"111111111",
  22582=>"001000000",
  22583=>"111111111",
  22584=>"000000000",
  22585=>"110000111",
  22586=>"110110111",
  22587=>"000010011",
  22588=>"000000001",
  22589=>"000000000",
  22590=>"101111111",
  22591=>"110110000",
  22592=>"111111111",
  22593=>"101101100",
  22594=>"010111111",
  22595=>"000000000",
  22596=>"100000000",
  22597=>"000000000",
  22598=>"011010110",
  22599=>"111111011",
  22600=>"111111000",
  22601=>"000000111",
  22602=>"000000000",
  22603=>"001111011",
  22604=>"000000001",
  22605=>"101100111",
  22606=>"000111011",
  22607=>"001001000",
  22608=>"000000000",
  22609=>"000000110",
  22610=>"000000000",
  22611=>"001001001",
  22612=>"000000000",
  22613=>"100101111",
  22614=>"000111111",
  22615=>"000111111",
  22616=>"001000111",
  22617=>"101000000",
  22618=>"010010000",
  22619=>"011011111",
  22620=>"011111001",
  22621=>"000001001",
  22622=>"000001101",
  22623=>"111111100",
  22624=>"000000111",
  22625=>"111111011",
  22626=>"000000000",
  22627=>"100111111",
  22628=>"111110110",
  22629=>"111111111",
  22630=>"000010011",
  22631=>"111001101",
  22632=>"000111011",
  22633=>"101001101",
  22634=>"111111111",
  22635=>"000000000",
  22636=>"110110111",
  22637=>"111111111",
  22638=>"000000000",
  22639=>"000000111",
  22640=>"111111000",
  22641=>"001000111",
  22642=>"101101111",
  22643=>"010011000",
  22644=>"111111111",
  22645=>"111111100",
  22646=>"000000000",
  22647=>"011000110",
  22648=>"100000000",
  22649=>"000000000",
  22650=>"111001100",
  22651=>"000000000",
  22652=>"110111101",
  22653=>"111001111",
  22654=>"000000000",
  22655=>"000000000",
  22656=>"100000100",
  22657=>"110010000",
  22658=>"101111101",
  22659=>"001001101",
  22660=>"100100111",
  22661=>"111011011",
  22662=>"111111111",
  22663=>"000000001",
  22664=>"111111111",
  22665=>"111000000",
  22666=>"111111111",
  22667=>"111111110",
  22668=>"001000000",
  22669=>"000100101",
  22670=>"000000000",
  22671=>"110111111",
  22672=>"000000000",
  22673=>"000000000",
  22674=>"100000000",
  22675=>"111111000",
  22676=>"101001101",
  22677=>"000000000",
  22678=>"011111011",
  22679=>"110111101",
  22680=>"101001001",
  22681=>"000101111",
  22682=>"001000100",
  22683=>"000000000",
  22684=>"011000001",
  22685=>"100000000",
  22686=>"000110011",
  22687=>"111111111",
  22688=>"000111111",
  22689=>"111110000",
  22690=>"000111011",
  22691=>"000000100",
  22692=>"001001000",
  22693=>"111111111",
  22694=>"000000101",
  22695=>"000011111",
  22696=>"001111101",
  22697=>"000000000",
  22698=>"000000000",
  22699=>"000000000",
  22700=>"111111000",
  22701=>"111111011",
  22702=>"000001111",
  22703=>"001101001",
  22704=>"011111111",
  22705=>"111111101",
  22706=>"011111010",
  22707=>"101000000",
  22708=>"101100000",
  22709=>"000000100",
  22710=>"000000101",
  22711=>"000000000",
  22712=>"001000000",
  22713=>"111111111",
  22714=>"001111111",
  22715=>"000010110",
  22716=>"000000010",
  22717=>"010010000",
  22718=>"111110110",
  22719=>"000110110",
  22720=>"111111111",
  22721=>"111111111",
  22722=>"001000000",
  22723=>"111111101",
  22724=>"111111000",
  22725=>"000000000",
  22726=>"111110110",
  22727=>"000000000",
  22728=>"100111111",
  22729=>"000000000",
  22730=>"000000000",
  22731=>"111111111",
  22732=>"000000000",
  22733=>"111111111",
  22734=>"000000100",
  22735=>"001000000",
  22736=>"111111100",
  22737=>"111111111",
  22738=>"010110111",
  22739=>"111111110",
  22740=>"100101101",
  22741=>"000000110",
  22742=>"100000100",
  22743=>"000001001",
  22744=>"111111111",
  22745=>"000111000",
  22746=>"111111111",
  22747=>"111111110",
  22748=>"000110100",
  22749=>"011110110",
  22750=>"000110111",
  22751=>"000010001",
  22752=>"111110000",
  22753=>"000000110",
  22754=>"000000000",
  22755=>"011111000",
  22756=>"110101000",
  22757=>"100111011",
  22758=>"000000000",
  22759=>"110111010",
  22760=>"111111011",
  22761=>"100000000",
  22762=>"000000000",
  22763=>"000000000",
  22764=>"000000000",
  22765=>"111111110",
  22766=>"000000110",
  22767=>"111111000",
  22768=>"001001111",
  22769=>"000000000",
  22770=>"000000000",
  22771=>"111111111",
  22772=>"101000001",
  22773=>"111111111",
  22774=>"000000000",
  22775=>"011011011",
  22776=>"111111111",
  22777=>"111111111",
  22778=>"000000111",
  22779=>"101110110",
  22780=>"000000000",
  22781=>"010111010",
  22782=>"000000000",
  22783=>"101100100",
  22784=>"111111000",
  22785=>"011011000",
  22786=>"000100110",
  22787=>"011111011",
  22788=>"000000000",
  22789=>"101101111",
  22790=>"110111111",
  22791=>"111111101",
  22792=>"110111111",
  22793=>"000000000",
  22794=>"110110110",
  22795=>"000101101",
  22796=>"001111111",
  22797=>"000000100",
  22798=>"000000000",
  22799=>"111110000",
  22800=>"000000000",
  22801=>"111000000",
  22802=>"111001000",
  22803=>"000111100",
  22804=>"000000111",
  22805=>"111011110",
  22806=>"101101100",
  22807=>"000000000",
  22808=>"110110111",
  22809=>"101000111",
  22810=>"000000011",
  22811=>"010011011",
  22812=>"011011000",
  22813=>"000000110",
  22814=>"111101111",
  22815=>"000001000",
  22816=>"000000000",
  22817=>"000010010",
  22818=>"111111111",
  22819=>"111101000",
  22820=>"000000111",
  22821=>"010000100",
  22822=>"111111111",
  22823=>"000000000",
  22824=>"110111111",
  22825=>"000000010",
  22826=>"111110000",
  22827=>"000000000",
  22828=>"000001111",
  22829=>"000000000",
  22830=>"000000100",
  22831=>"000001111",
  22832=>"110110110",
  22833=>"000000000",
  22834=>"111111111",
  22835=>"100000000",
  22836=>"111000110",
  22837=>"001000101",
  22838=>"111111001",
  22839=>"000000000",
  22840=>"110110110",
  22841=>"111001101",
  22842=>"111111001",
  22843=>"011000011",
  22844=>"000000101",
  22845=>"000000000",
  22846=>"000000100",
  22847=>"100000000",
  22848=>"111111110",
  22849=>"111111111",
  22850=>"000011000",
  22851=>"111111111",
  22852=>"111111111",
  22853=>"000100100",
  22854=>"111000000",
  22855=>"100110111",
  22856=>"000000001",
  22857=>"000100000",
  22858=>"100000000",
  22859=>"111100000",
  22860=>"100000100",
  22861=>"111001011",
  22862=>"000000000",
  22863=>"000000000",
  22864=>"110111111",
  22865=>"000000111",
  22866=>"111111111",
  22867=>"000110111",
  22868=>"011000011",
  22869=>"001011011",
  22870=>"000000000",
  22871=>"011110000",
  22872=>"100000111",
  22873=>"111111000",
  22874=>"000000000",
  22875=>"000000111",
  22876=>"000000100",
  22877=>"111111111",
  22878=>"111111111",
  22879=>"000000000",
  22880=>"111110000",
  22881=>"000011001",
  22882=>"010010010",
  22883=>"000000000",
  22884=>"010111111",
  22885=>"000000001",
  22886=>"100010011",
  22887=>"000000000",
  22888=>"111111001",
  22889=>"110100100",
  22890=>"111001000",
  22891=>"111000000",
  22892=>"000000100",
  22893=>"011011011",
  22894=>"000000000",
  22895=>"010110000",
  22896=>"000000101",
  22897=>"000000000",
  22898=>"011010000",
  22899=>"000101111",
  22900=>"100110110",
  22901=>"000000111",
  22902=>"000000111",
  22903=>"100000000",
  22904=>"100000000",
  22905=>"000101100",
  22906=>"000000000",
  22907=>"111111111",
  22908=>"000110110",
  22909=>"000000001",
  22910=>"000000000",
  22911=>"000000000",
  22912=>"000000011",
  22913=>"111111011",
  22914=>"000000000",
  22915=>"111111111",
  22916=>"100101110",
  22917=>"000110111",
  22918=>"000000000",
  22919=>"110111111",
  22920=>"111111111",
  22921=>"110101100",
  22922=>"000000010",
  22923=>"100100100",
  22924=>"111001000",
  22925=>"111111100",
  22926=>"111111111",
  22927=>"111111111",
  22928=>"000100101",
  22929=>"000001001",
  22930=>"000000111",
  22931=>"000000000",
  22932=>"000110111",
  22933=>"000000010",
  22934=>"000000000",
  22935=>"000000000",
  22936=>"111111101",
  22937=>"000000100",
  22938=>"000000011",
  22939=>"000000001",
  22940=>"000000000",
  22941=>"000001111",
  22942=>"001100101",
  22943=>"101111111",
  22944=>"000111111",
  22945=>"001000000",
  22946=>"000000111",
  22947=>"001000110",
  22948=>"111101101",
  22949=>"101111111",
  22950=>"000000000",
  22951=>"000000000",
  22952=>"011110000",
  22953=>"011011011",
  22954=>"000000011",
  22955=>"010100001",
  22956=>"111111111",
  22957=>"001101111",
  22958=>"000000000",
  22959=>"000000100",
  22960=>"001101111",
  22961=>"000100000",
  22962=>"100100111",
  22963=>"000110010",
  22964=>"000111111",
  22965=>"000101011",
  22966=>"001101111",
  22967=>"111111111",
  22968=>"000000001",
  22969=>"000000000",
  22970=>"000001011",
  22971=>"001101101",
  22972=>"000000000",
  22973=>"111111111",
  22974=>"011111011",
  22975=>"111111101",
  22976=>"000000000",
  22977=>"000000000",
  22978=>"000000000",
  22979=>"111111000",
  22980=>"000100111",
  22981=>"110111010",
  22982=>"000000000",
  22983=>"011000000",
  22984=>"101111111",
  22985=>"101101111",
  22986=>"000000000",
  22987=>"111111111",
  22988=>"001000111",
  22989=>"111011000",
  22990=>"110111111",
  22991=>"000011111",
  22992=>"000110000",
  22993=>"001111111",
  22994=>"100100001",
  22995=>"000000000",
  22996=>"110110000",
  22997=>"001111110",
  22998=>"000000000",
  22999=>"111111100",
  23000=>"000101101",
  23001=>"000000110",
  23002=>"000000000",
  23003=>"000000001",
  23004=>"111111011",
  23005=>"011010001",
  23006=>"011011011",
  23007=>"000000111",
  23008=>"000000000",
  23009=>"111111111",
  23010=>"000000000",
  23011=>"110111101",
  23012=>"010000000",
  23013=>"000000111",
  23014=>"111111001",
  23015=>"000000100",
  23016=>"111111111",
  23017=>"011000000",
  23018=>"110110101",
  23019=>"111111100",
  23020=>"110000001",
  23021=>"000000010",
  23022=>"101101111",
  23023=>"111111111",
  23024=>"001000101",
  23025=>"111111001",
  23026=>"111111111",
  23027=>"111100010",
  23028=>"000001001",
  23029=>"001001000",
  23030=>"000000111",
  23031=>"000000000",
  23032=>"000011111",
  23033=>"010011011",
  23034=>"110010100",
  23035=>"100000001",
  23036=>"110111111",
  23037=>"100000111",
  23038=>"001111110",
  23039=>"001001001",
  23040=>"001001001",
  23041=>"000000001",
  23042=>"111111111",
  23043=>"111111111",
  23044=>"000000001",
  23045=>"000111111",
  23046=>"000000000",
  23047=>"111111111",
  23048=>"111000110",
  23049=>"100000100",
  23050=>"011111111",
  23051=>"000010111",
  23052=>"000110110",
  23053=>"111111001",
  23054=>"000101111",
  23055=>"000001000",
  23056=>"000000000",
  23057=>"011001111",
  23058=>"111001000",
  23059=>"000111110",
  23060=>"000000000",
  23061=>"111111000",
  23062=>"111011000",
  23063=>"001011011",
  23064=>"011001011",
  23065=>"111001000",
  23066=>"010011011",
  23067=>"001111111",
  23068=>"100000000",
  23069=>"111111101",
  23070=>"111110100",
  23071=>"000111111",
  23072=>"000000000",
  23073=>"000110111",
  23074=>"111000000",
  23075=>"111001011",
  23076=>"000010000",
  23077=>"111000000",
  23078=>"000000111",
  23079=>"000000000",
  23080=>"011000001",
  23081=>"000000000",
  23082=>"001011111",
  23083=>"111111100",
  23084=>"111011000",
  23085=>"011101000",
  23086=>"000000000",
  23087=>"111000000",
  23088=>"111111001",
  23089=>"111111000",
  23090=>"000001011",
  23091=>"000000101",
  23092=>"111001000",
  23093=>"111011001",
  23094=>"110100101",
  23095=>"100000000",
  23096=>"000010000",
  23097=>"111111110",
  23098=>"000000000",
  23099=>"010000001",
  23100=>"000000000",
  23101=>"000000000",
  23102=>"111110110",
  23103=>"111000000",
  23104=>"011001000",
  23105=>"000000000",
  23106=>"001111111",
  23107=>"000000001",
  23108=>"100000000",
  23109=>"001000000",
  23110=>"000111111",
  23111=>"111100000",
  23112=>"110111000",
  23113=>"000000101",
  23114=>"010111111",
  23115=>"011011001",
  23116=>"000000011",
  23117=>"001000000",
  23118=>"000000100",
  23119=>"000000000",
  23120=>"000000000",
  23121=>"111000000",
  23122=>"100011001",
  23123=>"010000000",
  23124=>"111111000",
  23125=>"000001111",
  23126=>"000000001",
  23127=>"111111111",
  23128=>"011001000",
  23129=>"000000000",
  23130=>"100000110",
  23131=>"000011111",
  23132=>"000010111",
  23133=>"111000010",
  23134=>"011111111",
  23135=>"100000000",
  23136=>"110000111",
  23137=>"000000110",
  23138=>"000000000",
  23139=>"111000000",
  23140=>"110010111",
  23141=>"111101001",
  23142=>"010000000",
  23143=>"111000001",
  23144=>"111111101",
  23145=>"111101111",
  23146=>"000111111",
  23147=>"000011011",
  23148=>"011011111",
  23149=>"000000000",
  23150=>"111111111",
  23151=>"000101111",
  23152=>"010000111",
  23153=>"011001000",
  23154=>"110100001",
  23155=>"100111111",
  23156=>"111000000",
  23157=>"111111000",
  23158=>"111100000",
  23159=>"000000000",
  23160=>"000101111",
  23161=>"111111111",
  23162=>"000011011",
  23163=>"111100000",
  23164=>"011001000",
  23165=>"111111111",
  23166=>"010000000",
  23167=>"000000000",
  23168=>"000000000",
  23169=>"001111111",
  23170=>"000000111",
  23171=>"101111111",
  23172=>"010111111",
  23173=>"111000111",
  23174=>"110000000",
  23175=>"111000000",
  23176=>"000000000",
  23177=>"000000001",
  23178=>"000000000",
  23179=>"111000000",
  23180=>"110110100",
  23181=>"000110010",
  23182=>"111011011",
  23183=>"110010000",
  23184=>"111001000",
  23185=>"110111110",
  23186=>"010100111",
  23187=>"110000000",
  23188=>"001001111",
  23189=>"000111110",
  23190=>"101111111",
  23191=>"111111111",
  23192=>"000000000",
  23193=>"001111111",
  23194=>"000001010",
  23195=>"111011001",
  23196=>"000000000",
  23197=>"001111001",
  23198=>"111111100",
  23199=>"001000000",
  23200=>"000000000",
  23201=>"011011001",
  23202=>"111111000",
  23203=>"000011000",
  23204=>"111000001",
  23205=>"111000111",
  23206=>"111111000",
  23207=>"111111000",
  23208=>"001000101",
  23209=>"111001000",
  23210=>"111011000",
  23211=>"111111111",
  23212=>"000000000",
  23213=>"100110100",
  23214=>"000001111",
  23215=>"101000000",
  23216=>"000000000",
  23217=>"100100000",
  23218=>"011111111",
  23219=>"111101000",
  23220=>"000000111",
  23221=>"000000000",
  23222=>"000111111",
  23223=>"001001111",
  23224=>"111000000",
  23225=>"111001001",
  23226=>"001000011",
  23227=>"101110100",
  23228=>"111000000",
  23229=>"000000000",
  23230=>"011000000",
  23231=>"111011011",
  23232=>"000000000",
  23233=>"000110111",
  23234=>"110110110",
  23235=>"101111000",
  23236=>"001001001",
  23237=>"100111111",
  23238=>"000000000",
  23239=>"100101110",
  23240=>"111111111",
  23241=>"011011011",
  23242=>"000111111",
  23243=>"001001000",
  23244=>"111111111",
  23245=>"000000000",
  23246=>"000000001",
  23247=>"000000000",
  23248=>"101111111",
  23249=>"111001001",
  23250=>"000011111",
  23251=>"000000000",
  23252=>"100000000",
  23253=>"110000000",
  23254=>"100100111",
  23255=>"111111111",
  23256=>"111111111",
  23257=>"000100111",
  23258=>"111000000",
  23259=>"001101111",
  23260=>"000110111",
  23261=>"111110111",
  23262=>"000000000",
  23263=>"011001000",
  23264=>"100110111",
  23265=>"001000000",
  23266=>"111001001",
  23267=>"000000000",
  23268=>"101101000",
  23269=>"100110111",
  23270=>"100010011",
  23271=>"111001111",
  23272=>"111111111",
  23273=>"001001001",
  23274=>"111111000",
  23275=>"111111111",
  23276=>"101000000",
  23277=>"000000100",
  23278=>"111001101",
  23279=>"111000000",
  23280=>"111111111",
  23281=>"000000000",
  23282=>"001000000",
  23283=>"000000100",
  23284=>"000000000",
  23285=>"111011000",
  23286=>"000100111",
  23287=>"001001110",
  23288=>"001000000",
  23289=>"111111101",
  23290=>"000000000",
  23291=>"111111111",
  23292=>"110111111",
  23293=>"110000001",
  23294=>"110100111",
  23295=>"000000000",
  23296=>"000000000",
  23297=>"100110110",
  23298=>"111111001",
  23299=>"011111000",
  23300=>"000111111",
  23301=>"110000000",
  23302=>"111111010",
  23303=>"000000001",
  23304=>"010010011",
  23305=>"101110100",
  23306=>"001101111",
  23307=>"001000000",
  23308=>"110100100",
  23309=>"111010100",
  23310=>"000111111",
  23311=>"111111001",
  23312=>"111111110",
  23313=>"000000000",
  23314=>"100100110",
  23315=>"000000111",
  23316=>"000000000",
  23317=>"011111001",
  23318=>"100000000",
  23319=>"000101111",
  23320=>"111111111",
  23321=>"100111000",
  23322=>"000000111",
  23323=>"000000010",
  23324=>"110000000",
  23325=>"111101111",
  23326=>"011011011",
  23327=>"000111111",
  23328=>"010111111",
  23329=>"110111101",
  23330=>"111111111",
  23331=>"111000001",
  23332=>"000000000",
  23333=>"000000100",
  23334=>"000000000",
  23335=>"000001100",
  23336=>"110000011",
  23337=>"010110111",
  23338=>"000010000",
  23339=>"001111000",
  23340=>"000011111",
  23341=>"100110110",
  23342=>"000000111",
  23343=>"010010000",
  23344=>"111011111",
  23345=>"010000000",
  23346=>"110110000",
  23347=>"110000110",
  23348=>"110101111",
  23349=>"111101111",
  23350=>"001000000",
  23351=>"111111110",
  23352=>"000111000",
  23353=>"111000000",
  23354=>"111110000",
  23355=>"001001011",
  23356=>"000000000",
  23357=>"000000110",
  23358=>"111000001",
  23359=>"111111111",
  23360=>"011111111",
  23361=>"111111101",
  23362=>"000000000",
  23363=>"111000111",
  23364=>"101001111",
  23365=>"111111110",
  23366=>"111101000",
  23367=>"100110011",
  23368=>"111000000",
  23369=>"110111111",
  23370=>"111000000",
  23371=>"001000000",
  23372=>"000010010",
  23373=>"000000011",
  23374=>"010011111",
  23375=>"000011011",
  23376=>"000001001",
  23377=>"001001111",
  23378=>"001000000",
  23379=>"111000000",
  23380=>"001001000",
  23381=>"001011111",
  23382=>"111011111",
  23383=>"000000000",
  23384=>"011001001",
  23385=>"101000101",
  23386=>"111000001",
  23387=>"011111111",
  23388=>"111000000",
  23389=>"111100000",
  23390=>"001000001",
  23391=>"111111110",
  23392=>"100000111",
  23393=>"110100100",
  23394=>"100111001",
  23395=>"000000111",
  23396=>"100000000",
  23397=>"000111100",
  23398=>"000001111",
  23399=>"000001000",
  23400=>"111000001",
  23401=>"000110111",
  23402=>"011011111",
  23403=>"111000000",
  23404=>"000111111",
  23405=>"000111111",
  23406=>"110010000",
  23407=>"111000010",
  23408=>"000000011",
  23409=>"000001110",
  23410=>"000000101",
  23411=>"101110000",
  23412=>"000000000",
  23413=>"000000110",
  23414=>"110000100",
  23415=>"000000111",
  23416=>"000000000",
  23417=>"101111001",
  23418=>"000110111",
  23419=>"100000000",
  23420=>"000100000",
  23421=>"111111111",
  23422=>"001001000",
  23423=>"111001000",
  23424=>"001001111",
  23425=>"111101001",
  23426=>"100000000",
  23427=>"000011110",
  23428=>"000000001",
  23429=>"000100111",
  23430=>"010110110",
  23431=>"100000111",
  23432=>"000000111",
  23433=>"000000001",
  23434=>"011111111",
  23435=>"000001000",
  23436=>"000000001",
  23437=>"111101100",
  23438=>"100111111",
  23439=>"101111111",
  23440=>"000100100",
  23441=>"110100000",
  23442=>"111110111",
  23443=>"110000000",
  23444=>"011001100",
  23445=>"011001000",
  23446=>"101011011",
  23447=>"110110000",
  23448=>"111100011",
  23449=>"101101111",
  23450=>"111000000",
  23451=>"111011000",
  23452=>"111111111",
  23453=>"111001001",
  23454=>"111001000",
  23455=>"000000100",
  23456=>"000000111",
  23457=>"001011011",
  23458=>"010001101",
  23459=>"000000000",
  23460=>"001001111",
  23461=>"111111100",
  23462=>"101100111",
  23463=>"111111111",
  23464=>"111001000",
  23465=>"011000000",
  23466=>"111110000",
  23467=>"111001000",
  23468=>"101000000",
  23469=>"111000001",
  23470=>"011000000",
  23471=>"000001001",
  23472=>"001001001",
  23473=>"111000000",
  23474=>"111001000",
  23475=>"000000100",
  23476=>"111111100",
  23477=>"011001000",
  23478=>"011111111",
  23479=>"000000110",
  23480=>"111010001",
  23481=>"000111111",
  23482=>"100000010",
  23483=>"111111011",
  23484=>"011111110",
  23485=>"000011011",
  23486=>"000000000",
  23487=>"111110110",
  23488=>"011000000",
  23489=>"111000000",
  23490=>"111111111",
  23491=>"111000000",
  23492=>"011110111",
  23493=>"011011111",
  23494=>"001001101",
  23495=>"111111111",
  23496=>"000011111",
  23497=>"000101111",
  23498=>"000000001",
  23499=>"111001000",
  23500=>"111111111",
  23501=>"110111011",
  23502=>"001000000",
  23503=>"111111110",
  23504=>"001001111",
  23505=>"100000000",
  23506=>"111111000",
  23507=>"101111111",
  23508=>"111111011",
  23509=>"011111111",
  23510=>"001111111",
  23511=>"000000001",
  23512=>"101111111",
  23513=>"111101000",
  23514=>"111000000",
  23515=>"000001111",
  23516=>"111111011",
  23517=>"000000000",
  23518=>"100100111",
  23519=>"110000110",
  23520=>"011000000",
  23521=>"101000000",
  23522=>"100000000",
  23523=>"100000000",
  23524=>"111110111",
  23525=>"111111011",
  23526=>"000000000",
  23527=>"000000111",
  23528=>"010100000",
  23529=>"111000000",
  23530=>"000000010",
  23531=>"000000000",
  23532=>"111001001",
  23533=>"001011001",
  23534=>"001000000",
  23535=>"111111111",
  23536=>"111111000",
  23537=>"010001011",
  23538=>"111111111",
  23539=>"000000000",
  23540=>"001000000",
  23541=>"111101000",
  23542=>"100000111",
  23543=>"000000100",
  23544=>"111111110",
  23545=>"111111000",
  23546=>"100110111",
  23547=>"000111000",
  23548=>"011111111",
  23549=>"000000000",
  23550=>"000000000",
  23551=>"111000100",
  23552=>"111100000",
  23553=>"011111000",
  23554=>"111000000",
  23555=>"000011111",
  23556=>"111101001",
  23557=>"111111000",
  23558=>"000101100",
  23559=>"000000100",
  23560=>"000000111",
  23561=>"100000101",
  23562=>"111111000",
  23563=>"001101101",
  23564=>"001001000",
  23565=>"000000001",
  23566=>"110100000",
  23567=>"000100000",
  23568=>"000001101",
  23569=>"000000000",
  23570=>"000000110",
  23571=>"111101101",
  23572=>"010000000",
  23573=>"110110111",
  23574=>"000001111",
  23575=>"001000001",
  23576=>"111011001",
  23577=>"000000101",
  23578=>"111111111",
  23579=>"000000000",
  23580=>"111101100",
  23581=>"000000000",
  23582=>"100011000",
  23583=>"000000100",
  23584=>"000000011",
  23585=>"110100000",
  23586=>"111111111",
  23587=>"000000001",
  23588=>"001000111",
  23589=>"000000110",
  23590=>"110111110",
  23591=>"111111000",
  23592=>"001111111",
  23593=>"111111000",
  23594=>"111101101",
  23595=>"001000000",
  23596=>"001001111",
  23597=>"111111011",
  23598=>"111111011",
  23599=>"000010000",
  23600=>"111111000",
  23601=>"000101111",
  23602=>"001000000",
  23603=>"110010010",
  23604=>"111000000",
  23605=>"001001000",
  23606=>"001000110",
  23607=>"001001000",
  23608=>"000000000",
  23609=>"110110000",
  23610=>"001001001",
  23611=>"000000000",
  23612=>"111000001",
  23613=>"000000101",
  23614=>"111100100",
  23615=>"001000000",
  23616=>"001000000",
  23617=>"010010000",
  23618=>"101001111",
  23619=>"000011000",
  23620=>"000001011",
  23621=>"111001011",
  23622=>"001000000",
  23623=>"001100000",
  23624=>"110000000",
  23625=>"000000011",
  23626=>"000001000",
  23627=>"000100101",
  23628=>"000100001",
  23629=>"000000111",
  23630=>"111000000",
  23631=>"000001111",
  23632=>"000000000",
  23633=>"101000111",
  23634=>"111111110",
  23635=>"000000100",
  23636=>"000000000",
  23637=>"100110111",
  23638=>"000000000",
  23639=>"001001001",
  23640=>"101001110",
  23641=>"100000000",
  23642=>"111110000",
  23643=>"001010010",
  23644=>"111100110",
  23645=>"111011010",
  23646=>"001001111",
  23647=>"000000111",
  23648=>"000000010",
  23649=>"000000111",
  23650=>"111101111",
  23651=>"110100111",
  23652=>"000000001",
  23653=>"000000001",
  23654=>"100011001",
  23655=>"000001111",
  23656=>"001000000",
  23657=>"111111111",
  23658=>"110111000",
  23659=>"111111011",
  23660=>"010011001",
  23661=>"111111110",
  23662=>"110100110",
  23663=>"000000011",
  23664=>"000111111",
  23665=>"010011000",
  23666=>"000000000",
  23667=>"000000111",
  23668=>"111000011",
  23669=>"011111111",
  23670=>"100111111",
  23671=>"000100101",
  23672=>"000000000",
  23673=>"111101000",
  23674=>"001101111",
  23675=>"000000111",
  23676=>"000000001",
  23677=>"001011001",
  23678=>"101110111",
  23679=>"001111111",
  23680=>"000000000",
  23681=>"001001111",
  23682=>"000100111",
  23683=>"000001011",
  23684=>"011011000",
  23685=>"111111000",
  23686=>"111110000",
  23687=>"000000000",
  23688=>"000100000",
  23689=>"011111000",
  23690=>"100000000",
  23691=>"011000011",
  23692=>"001001101",
  23693=>"000000001",
  23694=>"110111111",
  23695=>"000000000",
  23696=>"111101111",
  23697=>"100000100",
  23698=>"000000000",
  23699=>"011000000",
  23700=>"111111111",
  23701=>"101111100",
  23702=>"111100010",
  23703=>"000000000",
  23704=>"000000111",
  23705=>"111111110",
  23706=>"001111111",
  23707=>"111111000",
  23708=>"000000111",
  23709=>"000000111",
  23710=>"100000011",
  23711=>"011000000",
  23712=>"000000000",
  23713=>"111000000",
  23714=>"000111111",
  23715=>"111000101",
  23716=>"001001001",
  23717=>"010111111",
  23718=>"110111111",
  23719=>"001001001",
  23720=>"111111101",
  23721=>"000001000",
  23722=>"000000000",
  23723=>"110100111",
  23724=>"001000101",
  23725=>"110010000",
  23726=>"111110110",
  23727=>"111000000",
  23728=>"000001111",
  23729=>"000011011",
  23730=>"010111111",
  23731=>"100111111",
  23732=>"001111110",
  23733=>"000000000",
  23734=>"111111000",
  23735=>"111110000",
  23736=>"000000000",
  23737=>"000111011",
  23738=>"001001001",
  23739=>"000001111",
  23740=>"111000000",
  23741=>"001000000",
  23742=>"110000110",
  23743=>"111100100",
  23744=>"111110100",
  23745=>"000110000",
  23746=>"111111110",
  23747=>"111111111",
  23748=>"000000010",
  23749=>"000111111",
  23750=>"001001101",
  23751=>"000110000",
  23752=>"011111010",
  23753=>"000000000",
  23754=>"111111111",
  23755=>"111100000",
  23756=>"010010000",
  23757=>"010011000",
  23758=>"110111011",
  23759=>"100000111",
  23760=>"101101000",
  23761=>"011111010",
  23762=>"101111000",
  23763=>"000100101",
  23764=>"000001111",
  23765=>"000000001",
  23766=>"011010010",
  23767=>"001111111",
  23768=>"000000111",
  23769=>"001000000",
  23770=>"000100111",
  23771=>"010010111",
  23772=>"000000000",
  23773=>"000001000",
  23774=>"001001100",
  23775=>"000011000",
  23776=>"111110111",
  23777=>"011111101",
  23778=>"111000000",
  23779=>"000100111",
  23780=>"111111111",
  23781=>"100100000",
  23782=>"111111000",
  23783=>"000000000",
  23784=>"111101110",
  23785=>"000111111",
  23786=>"111111111",
  23787=>"000000000",
  23788=>"111001000",
  23789=>"111010000",
  23790=>"111111000",
  23791=>"111111111",
  23792=>"000001001",
  23793=>"000000000",
  23794=>"111111111",
  23795=>"111111110",
  23796=>"101111111",
  23797=>"000110010",
  23798=>"111111001",
  23799=>"111111111",
  23800=>"111111111",
  23801=>"011001000",
  23802=>"000011011",
  23803=>"000001000",
  23804=>"000000010",
  23805=>"111000001",
  23806=>"110000001",
  23807=>"001011111",
  23808=>"001000001",
  23809=>"100111100",
  23810=>"111111000",
  23811=>"000001000",
  23812=>"100100111",
  23813=>"111111000",
  23814=>"111101000",
  23815=>"010010011",
  23816=>"011111011",
  23817=>"111111111",
  23818=>"111101100",
  23819=>"000111111",
  23820=>"111111111",
  23821=>"000000100",
  23822=>"111111111",
  23823=>"111111000",
  23824=>"000000000",
  23825=>"000111111",
  23826=>"000000000",
  23827=>"111101101",
  23828=>"000000000",
  23829=>"110100111",
  23830=>"110110100",
  23831=>"000101111",
  23832=>"001001111",
  23833=>"001000000",
  23834=>"111101010",
  23835=>"010110110",
  23836=>"110110100",
  23837=>"011001000",
  23838=>"100110111",
  23839=>"000011111",
  23840=>"001100100",
  23841=>"001001011",
  23842=>"011011111",
  23843=>"000000111",
  23844=>"010111110",
  23845=>"001000001",
  23846=>"101111100",
  23847=>"011000101",
  23848=>"111000000",
  23849=>"000000000",
  23850=>"111101000",
  23851=>"000000000",
  23852=>"000000000",
  23853=>"001001001",
  23854=>"001111111",
  23855=>"000000000",
  23856=>"000100100",
  23857=>"011000000",
  23858=>"001001000",
  23859=>"111110110",
  23860=>"000101000",
  23861=>"111111110",
  23862=>"000000010",
  23863=>"011001111",
  23864=>"000001111",
  23865=>"101000000",
  23866=>"000000011",
  23867=>"111111000",
  23868=>"111111000",
  23869=>"000000111",
  23870=>"001000000",
  23871=>"000000111",
  23872=>"011101100",
  23873=>"101101111",
  23874=>"001000000",
  23875=>"101001101",
  23876=>"000000000",
  23877=>"000000111",
  23878=>"000000000",
  23879=>"001011011",
  23880=>"110111000",
  23881=>"011111000",
  23882=>"000011111",
  23883=>"100110111",
  23884=>"111111001",
  23885=>"000000111",
  23886=>"111111111",
  23887=>"001011001",
  23888=>"000100101",
  23889=>"111111111",
  23890=>"111011111",
  23891=>"000000000",
  23892=>"111111111",
  23893=>"011011011",
  23894=>"111110000",
  23895=>"110000011",
  23896=>"111111111",
  23897=>"010001000",
  23898=>"001000000",
  23899=>"100111111",
  23900=>"000110011",
  23901=>"000000000",
  23902=>"111010000",
  23903=>"000001011",
  23904=>"001001001",
  23905=>"000000000",
  23906=>"001100111",
  23907=>"111111111",
  23908=>"110010111",
  23909=>"001000000",
  23910=>"111111111",
  23911=>"001001111",
  23912=>"000000000",
  23913=>"101010111",
  23914=>"100000000",
  23915=>"000000000",
  23916=>"001001001",
  23917=>"111111111",
  23918=>"011010000",
  23919=>"000000000",
  23920=>"000001000",
  23921=>"000000101",
  23922=>"001011000",
  23923=>"111111000",
  23924=>"111000111",
  23925=>"111100000",
  23926=>"000000111",
  23927=>"001001000",
  23928=>"000000000",
  23929=>"010111111",
  23930=>"010010010",
  23931=>"000111010",
  23932=>"101101000",
  23933=>"111001000",
  23934=>"100111111",
  23935=>"111100101",
  23936=>"011000000",
  23937=>"000000000",
  23938=>"001000110",
  23939=>"111111111",
  23940=>"111111000",
  23941=>"111111111",
  23942=>"000000000",
  23943=>"000111110",
  23944=>"110000000",
  23945=>"000000101",
  23946=>"001000111",
  23947=>"000101001",
  23948=>"111111111",
  23949=>"000000001",
  23950=>"111100100",
  23951=>"000000000",
  23952=>"010110000",
  23953=>"111111100",
  23954=>"100000000",
  23955=>"110111011",
  23956=>"000000000",
  23957=>"000000010",
  23958=>"000000100",
  23959=>"011010010",
  23960=>"001001001",
  23961=>"000001111",
  23962=>"011111010",
  23963=>"111111000",
  23964=>"111111111",
  23965=>"000000000",
  23966=>"111000000",
  23967=>"001001101",
  23968=>"000000011",
  23969=>"100110100",
  23970=>"000000100",
  23971=>"000111100",
  23972=>"001011111",
  23973=>"001011011",
  23974=>"111111111",
  23975=>"111001000",
  23976=>"110110000",
  23977=>"010000011",
  23978=>"000100111",
  23979=>"000010010",
  23980=>"000110000",
  23981=>"110110000",
  23982=>"111000000",
  23983=>"111111000",
  23984=>"010011111",
  23985=>"000000000",
  23986=>"000000000",
  23987=>"000001011",
  23988=>"111001001",
  23989=>"100000111",
  23990=>"000000000",
  23991=>"111001000",
  23992=>"001000000",
  23993=>"111110110",
  23994=>"000000101",
  23995=>"000000000",
  23996=>"000001111",
  23997=>"110110010",
  23998=>"111000000",
  23999=>"001001011",
  24000=>"111111011",
  24001=>"001001101",
  24002=>"101111111",
  24003=>"000000000",
  24004=>"111111111",
  24005=>"111111000",
  24006=>"111010000",
  24007=>"001000000",
  24008=>"100110111",
  24009=>"000000000",
  24010=>"000011000",
  24011=>"000000100",
  24012=>"000000111",
  24013=>"000000000",
  24014=>"001001000",
  24015=>"000100111",
  24016=>"000010000",
  24017=>"111111111",
  24018=>"111111111",
  24019=>"111111111",
  24020=>"011111111",
  24021=>"111001101",
  24022=>"000011111",
  24023=>"000100000",
  24024=>"111111110",
  24025=>"110111111",
  24026=>"011111111",
  24027=>"111001111",
  24028=>"101000000",
  24029=>"000110110",
  24030=>"001001000",
  24031=>"110100001",
  24032=>"110111111",
  24033=>"111100111",
  24034=>"101000111",
  24035=>"000010111",
  24036=>"000000010",
  24037=>"000000010",
  24038=>"000010111",
  24039=>"000000111",
  24040=>"111111001",
  24041=>"111000100",
  24042=>"000111111",
  24043=>"111100111",
  24044=>"010000000",
  24045=>"111110000",
  24046=>"001000000",
  24047=>"001001111",
  24048=>"000111111",
  24049=>"111111111",
  24050=>"111001001",
  24051=>"000110010",
  24052=>"111111111",
  24053=>"000101100",
  24054=>"000000000",
  24055=>"110000110",
  24056=>"111111001",
  24057=>"000100100",
  24058=>"111111111",
  24059=>"000001111",
  24060=>"000000000",
  24061=>"110110100",
  24062=>"110011000",
  24063=>"000111111",
  24064=>"000000000",
  24065=>"000000000",
  24066=>"000111111",
  24067=>"111011001",
  24068=>"110110100",
  24069=>"001000000",
  24070=>"000000000",
  24071=>"111111111",
  24072=>"011000000",
  24073=>"000000000",
  24074=>"011000000",
  24075=>"000000000",
  24076=>"110100100",
  24077=>"101111111",
  24078=>"000001000",
  24079=>"111111111",
  24080=>"111110111",
  24081=>"000000000",
  24082=>"101000000",
  24083=>"001001000",
  24084=>"011110110",
  24085=>"000000111",
  24086=>"111111111",
  24087=>"001101011",
  24088=>"110100001",
  24089=>"011011011",
  24090=>"001000000",
  24091=>"000000010",
  24092=>"010111010",
  24093=>"000000000",
  24094=>"001011111",
  24095=>"001001001",
  24096=>"111111011",
  24097=>"110110100",
  24098=>"001000110",
  24099=>"111000101",
  24100=>"111010000",
  24101=>"111111011",
  24102=>"111111000",
  24103=>"100000000",
  24104=>"111111011",
  24105=>"000000000",
  24106=>"000111111",
  24107=>"000000000",
  24108=>"111111111",
  24109=>"111111111",
  24110=>"000000101",
  24111=>"111111001",
  24112=>"000000001",
  24113=>"000000000",
  24114=>"111100010",
  24115=>"111111000",
  24116=>"011111111",
  24117=>"000000111",
  24118=>"001000001",
  24119=>"101011111",
  24120=>"001111100",
  24121=>"101111111",
  24122=>"000000000",
  24123=>"000000000",
  24124=>"111000000",
  24125=>"001001001",
  24126=>"010000111",
  24127=>"111001000",
  24128=>"001000000",
  24129=>"111111000",
  24130=>"000000000",
  24131=>"111111101",
  24132=>"000000000",
  24133=>"111111111",
  24134=>"000000111",
  24135=>"111111111",
  24136=>"100100000",
  24137=>"010000000",
  24138=>"000000000",
  24139=>"000000111",
  24140=>"111011111",
  24141=>"000010000",
  24142=>"000000001",
  24143=>"111111111",
  24144=>"000000001",
  24145=>"000001111",
  24146=>"111001111",
  24147=>"011011011",
  24148=>"000000111",
  24149=>"111111111",
  24150=>"000000000",
  24151=>"111110111",
  24152=>"100100100",
  24153=>"111100101",
  24154=>"000011111",
  24155=>"111111001",
  24156=>"000111111",
  24157=>"111101101",
  24158=>"111111101",
  24159=>"001000110",
  24160=>"000110111",
  24161=>"111111111",
  24162=>"000000000",
  24163=>"000000000",
  24164=>"010000011",
  24165=>"000000000",
  24166=>"111100111",
  24167=>"000000000",
  24168=>"111111111",
  24169=>"011000000",
  24170=>"001011111",
  24171=>"001000111",
  24172=>"000000000",
  24173=>"000000011",
  24174=>"111111000",
  24175=>"000000000",
  24176=>"000000111",
  24177=>"000010010",
  24178=>"011000000",
  24179=>"100101111",
  24180=>"111000110",
  24181=>"110110100",
  24182=>"111011000",
  24183=>"000000000",
  24184=>"111110111",
  24185=>"111111101",
  24186=>"111111110",
  24187=>"111111111",
  24188=>"100010110",
  24189=>"111111111",
  24190=>"000000000",
  24191=>"000000000",
  24192=>"000000000",
  24193=>"111111111",
  24194=>"010110110",
  24195=>"001001000",
  24196=>"111111111",
  24197=>"011000101",
  24198=>"010010010",
  24199=>"000000100",
  24200=>"111111010",
  24201=>"101000000",
  24202=>"000000000",
  24203=>"111111111",
  24204=>"111111111",
  24205=>"000000000",
  24206=>"001000000",
  24207=>"110111111",
  24208=>"111111111",
  24209=>"000111111",
  24210=>"000100111",
  24211=>"111111111",
  24212=>"101111111",
  24213=>"110111101",
  24214=>"111111000",
  24215=>"111111111",
  24216=>"001001111",
  24217=>"100000100",
  24218=>"000000000",
  24219=>"111111111",
  24220=>"111111011",
  24221=>"000000000",
  24222=>"111111111",
  24223=>"111111111",
  24224=>"000000000",
  24225=>"000010001",
  24226=>"111111111",
  24227=>"111111011",
  24228=>"000000000",
  24229=>"111100000",
  24230=>"111001001",
  24231=>"000010111",
  24232=>"111111111",
  24233=>"000001011",
  24234=>"111111011",
  24235=>"111111111",
  24236=>"001011011",
  24237=>"100000000",
  24238=>"111101011",
  24239=>"000000000",
  24240=>"000110111",
  24241=>"111111111",
  24242=>"110110000",
  24243=>"111000000",
  24244=>"011011111",
  24245=>"100000000",
  24246=>"000000000",
  24247=>"111111111",
  24248=>"111111111",
  24249=>"000000000",
  24250=>"000000000",
  24251=>"000111011",
  24252=>"101100101",
  24253=>"111110000",
  24254=>"000001001",
  24255=>"111111111",
  24256=>"111111111",
  24257=>"111011001",
  24258=>"000000011",
  24259=>"000111011",
  24260=>"000000000",
  24261=>"111111111",
  24262=>"111111100",
  24263=>"100101011",
  24264=>"011000000",
  24265=>"000000000",
  24266=>"111110010",
  24267=>"000000000",
  24268=>"111011011",
  24269=>"011111111",
  24270=>"111111111",
  24271=>"000000000",
  24272=>"000000001",
  24273=>"000010000",
  24274=>"000000000",
  24275=>"000000000",
  24276=>"100100011",
  24277=>"111111111",
  24278=>"111111111",
  24279=>"011011111",
  24280=>"000000000",
  24281=>"111111111",
  24282=>"000000000",
  24283=>"000000000",
  24284=>"111110001",
  24285=>"110100001",
  24286=>"000001001",
  24287=>"000000000",
  24288=>"111111110",
  24289=>"110111000",
  24290=>"111111000",
  24291=>"110110111",
  24292=>"111111111",
  24293=>"111111110",
  24294=>"110111111",
  24295=>"110000100",
  24296=>"000000000",
  24297=>"000000000",
  24298=>"111111111",
  24299=>"000000111",
  24300=>"000000000",
  24301=>"000110111",
  24302=>"000100101",
  24303=>"000000000",
  24304=>"110011010",
  24305=>"111100111",
  24306=>"000000000",
  24307=>"000001000",
  24308=>"000110100",
  24309=>"000100010",
  24310=>"001011011",
  24311=>"111111111",
  24312=>"110111111",
  24313=>"000000000",
  24314=>"000111111",
  24315=>"000100000",
  24316=>"111111111",
  24317=>"100000001",
  24318=>"111111111",
  24319=>"111111111",
  24320=>"001001011",
  24321=>"001000000",
  24322=>"000000000",
  24323=>"111111010",
  24324=>"111111111",
  24325=>"100111101",
  24326=>"000101111",
  24327=>"100000110",
  24328=>"111111011",
  24329=>"001000000",
  24330=>"111100101",
  24331=>"001000000",
  24332=>"000111111",
  24333=>"000000110",
  24334=>"111110110",
  24335=>"111101000",
  24336=>"111111111",
  24337=>"000000000",
  24338=>"111110110",
  24339=>"011001000",
  24340=>"001001000",
  24341=>"101000111",
  24342=>"111111001",
  24343=>"110111111",
  24344=>"100000000",
  24345=>"111101111",
  24346=>"100000001",
  24347=>"111111111",
  24348=>"111111001",
  24349=>"000111000",
  24350=>"010011000",
  24351=>"000001111",
  24352=>"001000000",
  24353=>"100111111",
  24354=>"000000000",
  24355=>"000001001",
  24356=>"110100110",
  24357=>"111111111",
  24358=>"011011001",
  24359=>"000000000",
  24360=>"111111111",
  24361=>"011111111",
  24362=>"101111111",
  24363=>"000000000",
  24364=>"111110111",
  24365=>"110110110",
  24366=>"001111000",
  24367=>"000100101",
  24368=>"110011111",
  24369=>"111111111",
  24370=>"000000100",
  24371=>"111010111",
  24372=>"000000000",
  24373=>"110000000",
  24374=>"000001111",
  24375=>"100000100",
  24376=>"000000000",
  24377=>"111111110",
  24378=>"111111111",
  24379=>"111111111",
  24380=>"101101011",
  24381=>"000000000",
  24382=>"000000000",
  24383=>"001000000",
  24384=>"000011000",
  24385=>"000000011",
  24386=>"110000000",
  24387=>"111110110",
  24388=>"000110111",
  24389=>"111111111",
  24390=>"000000000",
  24391=>"000001001",
  24392=>"000110111",
  24393=>"000000000",
  24394=>"101111111",
  24395=>"000000010",
  24396=>"000000100",
  24397=>"101111000",
  24398=>"111111111",
  24399=>"011011011",
  24400=>"011011001",
  24401=>"111011111",
  24402=>"001011111",
  24403=>"100100111",
  24404=>"111111110",
  24405=>"011101011",
  24406=>"000011101",
  24407=>"111111111",
  24408=>"111000000",
  24409=>"000000000",
  24410=>"100000000",
  24411=>"000000000",
  24412=>"000000000",
  24413=>"111111111",
  24414=>"000000000",
  24415=>"100000111",
  24416=>"111111111",
  24417=>"000000000",
  24418=>"011011011",
  24419=>"111111111",
  24420=>"000000000",
  24421=>"111100100",
  24422=>"000000001",
  24423=>"111111111",
  24424=>"001000000",
  24425=>"000000000",
  24426=>"111111110",
  24427=>"111000000",
  24428=>"000000000",
  24429=>"000011111",
  24430=>"100100000",
  24431=>"111111011",
  24432=>"000000000",
  24433=>"100100101",
  24434=>"000000000",
  24435=>"011001000",
  24436=>"010000000",
  24437=>"010000000",
  24438=>"111111111",
  24439=>"000000000",
  24440=>"011001000",
  24441=>"000000000",
  24442=>"110110111",
  24443=>"111101001",
  24444=>"110111110",
  24445=>"110100111",
  24446=>"111111111",
  24447=>"111111111",
  24448=>"000010010",
  24449=>"100110111",
  24450=>"110110000",
  24451=>"000000000",
  24452=>"000000000",
  24453=>"000000000",
  24454=>"111111111",
  24455=>"000000000",
  24456=>"000111111",
  24457=>"000001000",
  24458=>"111110100",
  24459=>"111111111",
  24460=>"111111111",
  24461=>"000000000",
  24462=>"111111111",
  24463=>"111111111",
  24464=>"111111111",
  24465=>"111110111",
  24466=>"111111111",
  24467=>"100010000",
  24468=>"000000000",
  24469=>"000000110",
  24470=>"000000000",
  24471=>"000000000",
  24472=>"111111101",
  24473=>"111111111",
  24474=>"111111111",
  24475=>"110110000",
  24476=>"101111111",
  24477=>"111111111",
  24478=>"001000101",
  24479=>"000000100",
  24480=>"100100111",
  24481=>"011000011",
  24482=>"000100100",
  24483=>"000000000",
  24484=>"101011111",
  24485=>"111111111",
  24486=>"000000000",
  24487=>"100100001",
  24488=>"000000000",
  24489=>"111111111",
  24490=>"001111111",
  24491=>"001000000",
  24492=>"000000000",
  24493=>"011010001",
  24494=>"000010011",
  24495=>"000000000",
  24496=>"101111111",
  24497=>"011011011",
  24498=>"001111111",
  24499=>"000101000",
  24500=>"000000000",
  24501=>"111111111",
  24502=>"111000000",
  24503=>"001000000",
  24504=>"111111010",
  24505=>"000000000",
  24506=>"000000100",
  24507=>"111111111",
  24508=>"111111110",
  24509=>"111111111",
  24510=>"000111001",
  24511=>"001001001",
  24512=>"111111111",
  24513=>"000000000",
  24514=>"000000000",
  24515=>"000000000",
  24516=>"000000000",
  24517=>"001000000",
  24518=>"011111001",
  24519=>"000000000",
  24520=>"001001000",
  24521=>"100000000",
  24522=>"010111111",
  24523=>"011011111",
  24524=>"000000000",
  24525=>"111111111",
  24526=>"000001001",
  24527=>"000000110",
  24528=>"000111011",
  24529=>"111111111",
  24530=>"111001001",
  24531=>"000000000",
  24532=>"001000000",
  24533=>"000100110",
  24534=>"111111111",
  24535=>"000001000",
  24536=>"000100011",
  24537=>"000000100",
  24538=>"000000000",
  24539=>"000000000",
  24540=>"000000000",
  24541=>"111111111",
  24542=>"001100111",
  24543=>"000000000",
  24544=>"000000000",
  24545=>"000100101",
  24546=>"111111111",
  24547=>"001000111",
  24548=>"111111111",
  24549=>"111001001",
  24550=>"001001110",
  24551=>"110111111",
  24552=>"100111111",
  24553=>"000000000",
  24554=>"010000000",
  24555=>"111111111",
  24556=>"011011111",
  24557=>"011000000",
  24558=>"111111011",
  24559=>"111111111",
  24560=>"100100101",
  24561=>"111111111",
  24562=>"000000000",
  24563=>"000000111",
  24564=>"000000000",
  24565=>"111111111",
  24566=>"000000000",
  24567=>"100111111",
  24568=>"111100110",
  24569=>"110010110",
  24570=>"111111011",
  24571=>"000111001",
  24572=>"111100100",
  24573=>"111111111",
  24574=>"111111011",
  24575=>"000000000",
  24576=>"111111111",
  24577=>"100000000",
  24578=>"101001100",
  24579=>"111101100",
  24580=>"100100110",
  24581=>"100000001",
  24582=>"010000000",
  24583=>"001111111",
  24584=>"111110000",
  24585=>"110111111",
  24586=>"000000000",
  24587=>"000000011",
  24588=>"000100100",
  24589=>"111111111",
  24590=>"000100110",
  24591=>"111111111",
  24592=>"011001000",
  24593=>"000110111",
  24594=>"011011000",
  24595=>"100100111",
  24596=>"000000000",
  24597=>"001001000",
  24598=>"000000000",
  24599=>"011011011",
  24600=>"110110110",
  24601=>"101101001",
  24602=>"000110000",
  24603=>"110100101",
  24604=>"000000000",
  24605=>"111111111",
  24606=>"100000000",
  24607=>"000011000",
  24608=>"111111111",
  24609=>"110000000",
  24610=>"111111100",
  24611=>"011010000",
  24612=>"000000000",
  24613=>"100000111",
  24614=>"111110100",
  24615=>"000000000",
  24616=>"001011001",
  24617=>"000100110",
  24618=>"000000000",
  24619=>"011111111",
  24620=>"111111111",
  24621=>"000000000",
  24622=>"000110110",
  24623=>"000000000",
  24624=>"111111111",
  24625=>"000000000",
  24626=>"000000000",
  24627=>"111111111",
  24628=>"001111111",
  24629=>"001111011",
  24630=>"111110110",
  24631=>"011100100",
  24632=>"011111100",
  24633=>"110110000",
  24634=>"111001111",
  24635=>"100100001",
  24636=>"111111111",
  24637=>"111010010",
  24638=>"001001001",
  24639=>"111001111",
  24640=>"110111000",
  24641=>"011111111",
  24642=>"000000000",
  24643=>"000000011",
  24644=>"101101000",
  24645=>"110100110",
  24646=>"000000010",
  24647=>"111111111",
  24648=>"101000001",
  24649=>"111111111",
  24650=>"001001010",
  24651=>"000111111",
  24652=>"011011011",
  24653=>"111100000",
  24654=>"111111111",
  24655=>"011111111",
  24656=>"111010000",
  24657=>"101101000",
  24658=>"100000000",
  24659=>"001100111",
  24660=>"111111111",
  24661=>"000000000",
  24662=>"100000110",
  24663=>"111111111",
  24664=>"000000000",
  24665=>"111100111",
  24666=>"000010010",
  24667=>"111111111",
  24668=>"000110000",
  24669=>"111111111",
  24670=>"100001001",
  24671=>"111110111",
  24672=>"001000000",
  24673=>"110100000",
  24674=>"000000000",
  24675=>"000000000",
  24676=>"110000000",
  24677=>"010000001",
  24678=>"000000111",
  24679=>"010111101",
  24680=>"000110111",
  24681=>"000000000",
  24682=>"000000000",
  24683=>"000000000",
  24684=>"011111100",
  24685=>"111111111",
  24686=>"111111000",
  24687=>"000001000",
  24688=>"000110111",
  24689=>"000000111",
  24690=>"101111111",
  24691=>"000000001",
  24692=>"111101001",
  24693=>"000000000",
  24694=>"000000100",
  24695=>"000000000",
  24696=>"111111111",
  24697=>"111111101",
  24698=>"011000000",
  24699=>"111111111",
  24700=>"000000100",
  24701=>"110111011",
  24702=>"000000000",
  24703=>"000000000",
  24704=>"011111111",
  24705=>"111011000",
  24706=>"001000000",
  24707=>"000000001",
  24708=>"111110111",
  24709=>"111111111",
  24710=>"001000000",
  24711=>"000000000",
  24712=>"100100000",
  24713=>"001001001",
  24714=>"001001000",
  24715=>"000000110",
  24716=>"101100100",
  24717=>"000011001",
  24718=>"111111111",
  24719=>"111110111",
  24720=>"100001011",
  24721=>"000111111",
  24722=>"000001001",
  24723=>"100110110",
  24724=>"110110000",
  24725=>"110100110",
  24726=>"011110011",
  24727=>"011000000",
  24728=>"111000100",
  24729=>"000000000",
  24730=>"111111111",
  24731=>"000011000",
  24732=>"101000000",
  24733=>"100011111",
  24734=>"111011010",
  24735=>"000000000",
  24736=>"010010110",
  24737=>"011001000",
  24738=>"111111101",
  24739=>"111011001",
  24740=>"000100000",
  24741=>"111100100",
  24742=>"000110110",
  24743=>"111001001",
  24744=>"110011111",
  24745=>"111111111",
  24746=>"000000110",
  24747=>"111101110",
  24748=>"011001111",
  24749=>"000111011",
  24750=>"110000000",
  24751=>"101101001",
  24752=>"001000000",
  24753=>"001101001",
  24754=>"100101100",
  24755=>"111111000",
  24756=>"111111110",
  24757=>"000000100",
  24758=>"111111110",
  24759=>"111000001",
  24760=>"111111111",
  24761=>"000001001",
  24762=>"000111111",
  24763=>"000001111",
  24764=>"000111111",
  24765=>"000001111",
  24766=>"111111111",
  24767=>"111111111",
  24768=>"111110011",
  24769=>"111111111",
  24770=>"000001110",
  24771=>"000000000",
  24772=>"111111001",
  24773=>"000001111",
  24774=>"000000000",
  24775=>"110111100",
  24776=>"111011011",
  24777=>"111111100",
  24778=>"001001111",
  24779=>"000000000",
  24780=>"111111100",
  24781=>"111111111",
  24782=>"000000000",
  24783=>"000011000",
  24784=>"100100100",
  24785=>"010111111",
  24786=>"100100000",
  24787=>"000000000",
  24788=>"001001001",
  24789=>"111111110",
  24790=>"000000000",
  24791=>"111100100",
  24792=>"111111111",
  24793=>"111001101",
  24794=>"000000000",
  24795=>"000100111",
  24796=>"000000000",
  24797=>"000000011",
  24798=>"000000000",
  24799=>"100111100",
  24800=>"000000000",
  24801=>"110110100",
  24802=>"000000000",
  24803=>"110111111",
  24804=>"111100111",
  24805=>"111111100",
  24806=>"000011011",
  24807=>"110110001",
  24808=>"111100000",
  24809=>"101110010",
  24810=>"011000100",
  24811=>"110110011",
  24812=>"001001000",
  24813=>"000011111",
  24814=>"000000100",
  24815=>"110000000",
  24816=>"111000000",
  24817=>"011111111",
  24818=>"111111111",
  24819=>"000001100",
  24820=>"110110110",
  24821=>"110111101",
  24822=>"000011010",
  24823=>"111111011",
  24824=>"000000000",
  24825=>"010000000",
  24826=>"111111111",
  24827=>"110100000",
  24828=>"000111111",
  24829=>"101000000",
  24830=>"110100000",
  24831=>"110000000",
  24832=>"010010100",
  24833=>"100010010",
  24834=>"110000111",
  24835=>"111111111",
  24836=>"011011000",
  24837=>"111001000",
  24838=>"000000011",
  24839=>"110110111",
  24840=>"111111111",
  24841=>"000000010",
  24842=>"111111100",
  24843=>"111111100",
  24844=>"100000000",
  24845=>"111000000",
  24846=>"111111100",
  24847=>"000000001",
  24848=>"111000000",
  24849=>"111111111",
  24850=>"111110110",
  24851=>"111111111",
  24852=>"000000000",
  24853=>"111111000",
  24854=>"000000000",
  24855=>"111101101",
  24856=>"001101110",
  24857=>"000111011",
  24858=>"111111010",
  24859=>"000000000",
  24860=>"000000000",
  24861=>"111111111",
  24862=>"010110111",
  24863=>"001000110",
  24864=>"000000011",
  24865=>"000000000",
  24866=>"111111111",
  24867=>"100111111",
  24868=>"011011011",
  24869=>"111111110",
  24870=>"000001000",
  24871=>"111111000",
  24872=>"011000101",
  24873=>"000000010",
  24874=>"010000000",
  24875=>"110111111",
  24876=>"011011111",
  24877=>"111111101",
  24878=>"000000000",
  24879=>"111011000",
  24880=>"111111111",
  24881=>"111011011",
  24882=>"000000000",
  24883=>"011111001",
  24884=>"111111111",
  24885=>"100111111",
  24886=>"111000111",
  24887=>"111110111",
  24888=>"011111000",
  24889=>"000000000",
  24890=>"000001011",
  24891=>"111111111",
  24892=>"000000000",
  24893=>"001001111",
  24894=>"100000000",
  24895=>"111111000",
  24896=>"000000100",
  24897=>"000000000",
  24898=>"100000000",
  24899=>"001001001",
  24900=>"111110010",
  24901=>"100100111",
  24902=>"000110000",
  24903=>"000110110",
  24904=>"111111111",
  24905=>"000000110",
  24906=>"110111111",
  24907=>"111111111",
  24908=>"100000110",
  24909=>"000100101",
  24910=>"111111100",
  24911=>"011111110",
  24912=>"011001001",
  24913=>"110000000",
  24914=>"000000001",
  24915=>"111111000",
  24916=>"000000000",
  24917=>"001001011",
  24918=>"000010000",
  24919=>"111101101",
  24920=>"111111111",
  24921=>"111111000",
  24922=>"000000000",
  24923=>"111111100",
  24924=>"000000000",
  24925=>"001001000",
  24926=>"111011111",
  24927=>"000000000",
  24928=>"111111110",
  24929=>"111110000",
  24930=>"000100111",
  24931=>"111111111",
  24932=>"001111111",
  24933=>"101111011",
  24934=>"100111111",
  24935=>"111111111",
  24936=>"110110111",
  24937=>"000011011",
  24938=>"001000000",
  24939=>"111001011",
  24940=>"000000100",
  24941=>"000111111",
  24942=>"010111001",
  24943=>"011000010",
  24944=>"000000000",
  24945=>"000000000",
  24946=>"111111001",
  24947=>"100000011",
  24948=>"000110110",
  24949=>"010000000",
  24950=>"000000000",
  24951=>"111111111",
  24952=>"000101111",
  24953=>"000000000",
  24954=>"000000000",
  24955=>"110000000",
  24956=>"011011111",
  24957=>"011000000",
  24958=>"101000000",
  24959=>"111111000",
  24960=>"111101100",
  24961=>"111010101",
  24962=>"111011001",
  24963=>"000000000",
  24964=>"110111111",
  24965=>"000000100",
  24966=>"110000100",
  24967=>"111111111",
  24968=>"101000000",
  24969=>"000000000",
  24970=>"101111111",
  24971=>"000000000",
  24972=>"111100111",
  24973=>"100110000",
  24974=>"111111111",
  24975=>"000000000",
  24976=>"000000000",
  24977=>"011111111",
  24978=>"100000000",
  24979=>"111001000",
  24980=>"001001000",
  24981=>"000000001",
  24982=>"000000000",
  24983=>"000000100",
  24984=>"000100110",
  24985=>"110111111",
  24986=>"000100100",
  24987=>"111111111",
  24988=>"100000111",
  24989=>"111100110",
  24990=>"101111111",
  24991=>"000000000",
  24992=>"110111111",
  24993=>"111000000",
  24994=>"111111111",
  24995=>"000001000",
  24996=>"111111111",
  24997=>"011001001",
  24998=>"100000000",
  24999=>"000000000",
  25000=>"010100000",
  25001=>"111111111",
  25002=>"010000000",
  25003=>"000000000",
  25004=>"100110111",
  25005=>"111111111",
  25006=>"111111111",
  25007=>"101000000",
  25008=>"110110011",
  25009=>"111111111",
  25010=>"110111111",
  25011=>"000011011",
  25012=>"011111111",
  25013=>"001011111",
  25014=>"111010100",
  25015=>"100000000",
  25016=>"000001101",
  25017=>"000000000",
  25018=>"111111111",
  25019=>"100000000",
  25020=>"000100110",
  25021=>"001001111",
  25022=>"101100111",
  25023=>"000010010",
  25024=>"000000101",
  25025=>"111111000",
  25026=>"111111111",
  25027=>"001111111",
  25028=>"000000000",
  25029=>"110110100",
  25030=>"000010110",
  25031=>"000010110",
  25032=>"011010000",
  25033=>"110110000",
  25034=>"111100111",
  25035=>"111111111",
  25036=>"111111111",
  25037=>"000000000",
  25038=>"100111001",
  25039=>"011111111",
  25040=>"000000000",
  25041=>"010010010",
  25042=>"000000001",
  25043=>"111111111",
  25044=>"111100000",
  25045=>"110010000",
  25046=>"100100111",
  25047=>"000010111",
  25048=>"100000000",
  25049=>"111111111",
  25050=>"000000000",
  25051=>"000000100",
  25052=>"111110010",
  25053=>"000001000",
  25054=>"111111111",
  25055=>"000000000",
  25056=>"111011000",
  25057=>"111111011",
  25058=>"000011111",
  25059=>"111111111",
  25060=>"100011111",
  25061=>"111111111",
  25062=>"111111111",
  25063=>"001001000",
  25064=>"111111111",
  25065=>"110110111",
  25066=>"010000000",
  25067=>"000000000",
  25068=>"110111011",
  25069=>"000000100",
  25070=>"001001001",
  25071=>"000000000",
  25072=>"000000000",
  25073=>"010111111",
  25074=>"111111111",
  25075=>"000000000",
  25076=>"000000000",
  25077=>"111111111",
  25078=>"111111111",
  25079=>"000100110",
  25080=>"000010010",
  25081=>"001001001",
  25082=>"000000000",
  25083=>"100111111",
  25084=>"011000000",
  25085=>"101101101",
  25086=>"000000000",
  25087=>"000000000",
  25088=>"000000000",
  25089=>"101000011",
  25090=>"000000011",
  25091=>"111011001",
  25092=>"101000100",
  25093=>"111111111",
  25094=>"000101111",
  25095=>"000010011",
  25096=>"001000110",
  25097=>"000000000",
  25098=>"111111111",
  25099=>"110111111",
  25100=>"111111111",
  25101=>"000001001",
  25102=>"000000000",
  25103=>"111111111",
  25104=>"011111111",
  25105=>"110001111",
  25106=>"000000000",
  25107=>"111111000",
  25108=>"111111001",
  25109=>"000111111",
  25110=>"100100100",
  25111=>"000111100",
  25112=>"000000000",
  25113=>"110100100",
  25114=>"000000000",
  25115=>"110110100",
  25116=>"001001001",
  25117=>"010111000",
  25118=>"000000011",
  25119=>"100000100",
  25120=>"111111111",
  25121=>"111111111",
  25122=>"011111111",
  25123=>"001001111",
  25124=>"101111111",
  25125=>"111111111",
  25126=>"110111111",
  25127=>"001000000",
  25128=>"111111111",
  25129=>"000000000",
  25130=>"000000000",
  25131=>"000100111",
  25132=>"000111101",
  25133=>"000000000",
  25134=>"000000000",
  25135=>"000100000",
  25136=>"000110110",
  25137=>"111111111",
  25138=>"100110111",
  25139=>"000000100",
  25140=>"111111111",
  25141=>"111111111",
  25142=>"000000011",
  25143=>"000001000",
  25144=>"111111111",
  25145=>"111111111",
  25146=>"000000000",
  25147=>"100000111",
  25148=>"111111111",
  25149=>"100100100",
  25150=>"111100111",
  25151=>"000000000",
  25152=>"111111111",
  25153=>"111111111",
  25154=>"111100110",
  25155=>"011000000",
  25156=>"000000000",
  25157=>"110100000",
  25158=>"111000010",
  25159=>"111111000",
  25160=>"111011011",
  25161=>"111111000",
  25162=>"111111111",
  25163=>"000000000",
  25164=>"111100100",
  25165=>"111000000",
  25166=>"000000000",
  25167=>"111111000",
  25168=>"001111001",
  25169=>"000000000",
  25170=>"010100000",
  25171=>"100100100",
  25172=>"000000000",
  25173=>"000000000",
  25174=>"100110000",
  25175=>"111000000",
  25176=>"000000100",
  25177=>"111111111",
  25178=>"000110111",
  25179=>"011000100",
  25180=>"000000111",
  25181=>"010111011",
  25182=>"001001011",
  25183=>"100100100",
  25184=>"000000000",
  25185=>"111111000",
  25186=>"111101111",
  25187=>"111001000",
  25188=>"000000001",
  25189=>"000111111",
  25190=>"000000000",
  25191=>"100000000",
  25192=>"000000000",
  25193=>"111111111",
  25194=>"001011011",
  25195=>"000000100",
  25196=>"001100111",
  25197=>"110111000",
  25198=>"000000000",
  25199=>"111111010",
  25200=>"110111000",
  25201=>"000000000",
  25202=>"011111011",
  25203=>"000100000",
  25204=>"000000000",
  25205=>"001001101",
  25206=>"111001000",
  25207=>"111111111",
  25208=>"000000000",
  25209=>"000000000",
  25210=>"101100000",
  25211=>"011010010",
  25212=>"111111111",
  25213=>"010110000",
  25214=>"100101000",
  25215=>"000000010",
  25216=>"000010000",
  25217=>"111111110",
  25218=>"100101000",
  25219=>"011110110",
  25220=>"111111111",
  25221=>"111111000",
  25222=>"100110100",
  25223=>"111111110",
  25224=>"000000111",
  25225=>"000111111",
  25226=>"000000000",
  25227=>"111111000",
  25228=>"001000000",
  25229=>"100100111",
  25230=>"111111111",
  25231=>"111111111",
  25232=>"000000000",
  25233=>"000000000",
  25234=>"011111111",
  25235=>"000000000",
  25236=>"110000000",
  25237=>"001011111",
  25238=>"000000001",
  25239=>"000000000",
  25240=>"101000110",
  25241=>"000001011",
  25242=>"000000000",
  25243=>"000000000",
  25244=>"111111111",
  25245=>"000000101",
  25246=>"111111111",
  25247=>"000000000",
  25248=>"100100111",
  25249=>"000000010",
  25250=>"111111000",
  25251=>"111100111",
  25252=>"111011111",
  25253=>"011001000",
  25254=>"110111111",
  25255=>"111111111",
  25256=>"001011111",
  25257=>"000000011",
  25258=>"000000000",
  25259=>"000000000",
  25260=>"001011111",
  25261=>"011011111",
  25262=>"111111111",
  25263=>"111011111",
  25264=>"111110000",
  25265=>"111011001",
  25266=>"111111110",
  25267=>"111111111",
  25268=>"111100100",
  25269=>"111111111",
  25270=>"111111111",
  25271=>"111110110",
  25272=>"111100111",
  25273=>"111111111",
  25274=>"000000000",
  25275=>"011000000",
  25276=>"000000000",
  25277=>"111000001",
  25278=>"111111111",
  25279=>"111111111",
  25280=>"010010010",
  25281=>"000000000",
  25282=>"001000000",
  25283=>"011111111",
  25284=>"000000000",
  25285=>"010111111",
  25286=>"111111111",
  25287=>"000000000",
  25288=>"000011001",
  25289=>"111111001",
  25290=>"001000111",
  25291=>"011011000",
  25292=>"000000000",
  25293=>"100111111",
  25294=>"110000000",
  25295=>"111111111",
  25296=>"111111001",
  25297=>"000100101",
  25298=>"111011111",
  25299=>"111111010",
  25300=>"001111000",
  25301=>"011000000",
  25302=>"000000000",
  25303=>"100000000",
  25304=>"000000000",
  25305=>"100100110",
  25306=>"110010000",
  25307=>"000001111",
  25308=>"111011111",
  25309=>"110110010",
  25310=>"111111111",
  25311=>"011111111",
  25312=>"000000000",
  25313=>"011000011",
  25314=>"000000000",
  25315=>"000000000",
  25316=>"111100100",
  25317=>"000001011",
  25318=>"000000000",
  25319=>"111111111",
  25320=>"000000000",
  25321=>"000000000",
  25322=>"000000111",
  25323=>"011001000",
  25324=>"000010000",
  25325=>"000111011",
  25326=>"000000000",
  25327=>"111111111",
  25328=>"111111000",
  25329=>"111111111",
  25330=>"000000000",
  25331=>"000000000",
  25332=>"111011011",
  25333=>"111111111",
  25334=>"101001000",
  25335=>"000000100",
  25336=>"100000000",
  25337=>"000010100",
  25338=>"111111111",
  25339=>"000000000",
  25340=>"000000000",
  25341=>"101111111",
  25342=>"011011011",
  25343=>"000000111",
  25344=>"111100100",
  25345=>"000000011",
  25346=>"100000100",
  25347=>"000000000",
  25348=>"011011110",
  25349=>"111111111",
  25350=>"000000000",
  25351=>"011001111",
  25352=>"000000000",
  25353=>"111000000",
  25354=>"110111111",
  25355=>"011010111",
  25356=>"111111100",
  25357=>"000000000",
  25358=>"001000000",
  25359=>"110000000",
  25360=>"111111111",
  25361=>"000000000",
  25362=>"000000000",
  25363=>"000101111",
  25364=>"110000100",
  25365=>"000000110",
  25366=>"001011111",
  25367=>"111111111",
  25368=>"000010000",
  25369=>"111111000",
  25370=>"100000000",
  25371=>"111111111",
  25372=>"001001100",
  25373=>"111111110",
  25374=>"000110111",
  25375=>"111111111",
  25376=>"111001000",
  25377=>"001001011",
  25378=>"111111111",
  25379=>"000000000",
  25380=>"001001001",
  25381=>"010010001",
  25382=>"111111111",
  25383=>"000000011",
  25384=>"101001000",
  25385=>"000010000",
  25386=>"011111000",
  25387=>"110111111",
  25388=>"011000000",
  25389=>"000000000",
  25390=>"111000111",
  25391=>"111111001",
  25392=>"001110111",
  25393=>"100110000",
  25394=>"100101100",
  25395=>"000000000",
  25396=>"111111111",
  25397=>"111100111",
  25398=>"111111111",
  25399=>"011001111",
  25400=>"000000000",
  25401=>"110000111",
  25402=>"000000000",
  25403=>"110010011",
  25404=>"000000000",
  25405=>"111111110",
  25406=>"111111101",
  25407=>"111111111",
  25408=>"000000000",
  25409=>"000000000",
  25410=>"111111111",
  25411=>"000001101",
  25412=>"000000001",
  25413=>"010011011",
  25414=>"111111111",
  25415=>"110110111",
  25416=>"111110111",
  25417=>"001101111",
  25418=>"111111011",
  25419=>"100101011",
  25420=>"000111111",
  25421=>"011011111",
  25422=>"000001111",
  25423=>"000100110",
  25424=>"100110110",
  25425=>"000010110",
  25426=>"110111011",
  25427=>"111111111",
  25428=>"100000000",
  25429=>"011011011",
  25430=>"111111111",
  25431=>"110110000",
  25432=>"000000000",
  25433=>"011111111",
  25434=>"111110000",
  25435=>"101111111",
  25436=>"000000000",
  25437=>"111001000",
  25438=>"000000000",
  25439=>"000000000",
  25440=>"000000100",
  25441=>"000000000",
  25442=>"000000110",
  25443=>"111111111",
  25444=>"111111110",
  25445=>"000000000",
  25446=>"111111111",
  25447=>"111000111",
  25448=>"101111011",
  25449=>"000000000",
  25450=>"000000000",
  25451=>"000000000",
  25452=>"000000000",
  25453=>"101001000",
  25454=>"000000000",
  25455=>"111111000",
  25456=>"110110000",
  25457=>"000000000",
  25458=>"111111111",
  25459=>"111111110",
  25460=>"100100100",
  25461=>"001000010",
  25462=>"011000110",
  25463=>"111111111",
  25464=>"000000000",
  25465=>"000000100",
  25466=>"001011000",
  25467=>"111111111",
  25468=>"111111111",
  25469=>"000001000",
  25470=>"000000000",
  25471=>"000011000",
  25472=>"010000000",
  25473=>"001011111",
  25474=>"111100000",
  25475=>"111011000",
  25476=>"100111111",
  25477=>"110110111",
  25478=>"000011000",
  25479=>"000100110",
  25480=>"100110000",
  25481=>"100110111",
  25482=>"000000000",
  25483=>"110111111",
  25484=>"111111111",
  25485=>"111111111",
  25486=>"111111111",
  25487=>"000000000",
  25488=>"110000000",
  25489=>"111001000",
  25490=>"010111111",
  25491=>"001000000",
  25492=>"000000111",
  25493=>"000001011",
  25494=>"111100100",
  25495=>"000111100",
  25496=>"111000000",
  25497=>"011001110",
  25498=>"000000000",
  25499=>"110111111",
  25500=>"111110000",
  25501=>"001011000",
  25502=>"111001000",
  25503=>"111111111",
  25504=>"000000000",
  25505=>"011011001",
  25506=>"100110110",
  25507=>"011110000",
  25508=>"000000100",
  25509=>"000111111",
  25510=>"000000111",
  25511=>"000000011",
  25512=>"111111010",
  25513=>"111111110",
  25514=>"000000000",
  25515=>"011011011",
  25516=>"000000001",
  25517=>"001000000",
  25518=>"000010000",
  25519=>"111011000",
  25520=>"011011000",
  25521=>"000000000",
  25522=>"110110111",
  25523=>"000000000",
  25524=>"111111111",
  25525=>"101100101",
  25526=>"101001000",
  25527=>"110000110",
  25528=>"111111000",
  25529=>"110111111",
  25530=>"111101000",
  25531=>"000000000",
  25532=>"100100111",
  25533=>"101111111",
  25534=>"011000000",
  25535=>"111110000",
  25536=>"011011111",
  25537=>"000000100",
  25538=>"111111111",
  25539=>"110010111",
  25540=>"011111001",
  25541=>"000000000",
  25542=>"111111001",
  25543=>"111001000",
  25544=>"111100111",
  25545=>"011111111",
  25546=>"000000000",
  25547=>"000000010",
  25548=>"000000000",
  25549=>"111111111",
  25550=>"111111111",
  25551=>"000000000",
  25552=>"000000000",
  25553=>"000000000",
  25554=>"111001001",
  25555=>"111111111",
  25556=>"001000000",
  25557=>"000000011",
  25558=>"000000111",
  25559=>"110000000",
  25560=>"000011010",
  25561=>"000000000",
  25562=>"000000000",
  25563=>"111111111",
  25564=>"111111111",
  25565=>"111111111",
  25566=>"111000100",
  25567=>"011000001",
  25568=>"000000000",
  25569=>"101111111",
  25570=>"000100100",
  25571=>"010111111",
  25572=>"000000000",
  25573=>"000000001",
  25574=>"000000010",
  25575=>"000000000",
  25576=>"000000000",
  25577=>"011110110",
  25578=>"000000000",
  25579=>"111111111",
  25580=>"000000111",
  25581=>"100110110",
  25582=>"111111011",
  25583=>"000000010",
  25584=>"111111000",
  25585=>"110000000",
  25586=>"111111111",
  25587=>"110100000",
  25588=>"001001101",
  25589=>"111111111",
  25590=>"000000000",
  25591=>"000000000",
  25592=>"111110000",
  25593=>"000100100",
  25594=>"010000101",
  25595=>"111111111",
  25596=>"011011000",
  25597=>"111111011",
  25598=>"000000000",
  25599=>"111011000",
  25600=>"011111111",
  25601=>"000000001",
  25602=>"000010010",
  25603=>"111111111",
  25604=>"000000010",
  25605=>"011000100",
  25606=>"101000000",
  25607=>"110100100",
  25608=>"000000001",
  25609=>"101101111",
  25610=>"000000000",
  25611=>"000111011",
  25612=>"111111011",
  25613=>"000001000",
  25614=>"000000111",
  25615=>"000000000",
  25616=>"111000000",
  25617=>"000000100",
  25618=>"100000000",
  25619=>"111111000",
  25620=>"000000100",
  25621=>"000111000",
  25622=>"000000000",
  25623=>"110111110",
  25624=>"001111010",
  25625=>"001000000",
  25626=>"000000000",
  25627=>"000000000",
  25628=>"111100100",
  25629=>"011011111",
  25630=>"011111110",
  25631=>"111111111",
  25632=>"000100000",
  25633=>"111111111",
  25634=>"000000011",
  25635=>"000110111",
  25636=>"000000000",
  25637=>"111111011",
  25638=>"000000100",
  25639=>"100100101",
  25640=>"000000000",
  25641=>"000000000",
  25642=>"000001000",
  25643=>"111011000",
  25644=>"011000000",
  25645=>"111000100",
  25646=>"001111111",
  25647=>"110000000",
  25648=>"110111111",
  25649=>"111101101",
  25650=>"100100100",
  25651=>"100100100",
  25652=>"100101001",
  25653=>"001001001",
  25654=>"000000100",
  25655=>"000000010",
  25656=>"001000000",
  25657=>"111111111",
  25658=>"000100110",
  25659=>"111111000",
  25660=>"000000000",
  25661=>"111111100",
  25662=>"111111011",
  25663=>"000000000",
  25664=>"010000000",
  25665=>"111111110",
  25666=>"111111111",
  25667=>"011011000",
  25668=>"111111111",
  25669=>"110110111",
  25670=>"000011000",
  25671=>"000000000",
  25672=>"011011001",
  25673=>"000000000",
  25674=>"111111010",
  25675=>"011001000",
  25676=>"100110111",
  25677=>"011011000",
  25678=>"110111010",
  25679=>"000111101",
  25680=>"001001000",
  25681=>"111000000",
  25682=>"000000000",
  25683=>"111111111",
  25684=>"101000000",
  25685=>"000000000",
  25686=>"100000100",
  25687=>"111110011",
  25688=>"000000000",
  25689=>"000000000",
  25690=>"001001111",
  25691=>"001000000",
  25692=>"000000000",
  25693=>"100111011",
  25694=>"111111111",
  25695=>"000000000",
  25696=>"000000000",
  25697=>"111111111",
  25698=>"000000000",
  25699=>"100100100",
  25700=>"000000000",
  25701=>"111000000",
  25702=>"001000000",
  25703=>"000000000",
  25704=>"111111111",
  25705=>"000000001",
  25706=>"111111111",
  25707=>"010011000",
  25708=>"011010000",
  25709=>"000000000",
  25710=>"111111010",
  25711=>"000000000",
  25712=>"000000000",
  25713=>"110000000",
  25714=>"111000001",
  25715=>"111111100",
  25716=>"111111110",
  25717=>"111111001",
  25718=>"111000011",
  25719=>"000011111",
  25720=>"001000000",
  25721=>"010111111",
  25722=>"101000001",
  25723=>"011000000",
  25724=>"000000000",
  25725=>"100111111",
  25726=>"111111001",
  25727=>"011011000",
  25728=>"000000000",
  25729=>"111111111",
  25730=>"000000000",
  25731=>"101101001",
  25732=>"000000111",
  25733=>"000000000",
  25734=>"110111111",
  25735=>"111111111",
  25736=>"110110110",
  25737=>"000010010",
  25738=>"111111110",
  25739=>"000000000",
  25740=>"111111111",
  25741=>"000000000",
  25742=>"111111111",
  25743=>"000111111",
  25744=>"000000000",
  25745=>"101101100",
  25746=>"111111010",
  25747=>"000000000",
  25748=>"111111111",
  25749=>"000000110",
  25750=>"000000000",
  25751=>"111111111",
  25752=>"111000100",
  25753=>"000101111",
  25754=>"000000100",
  25755=>"111111000",
  25756=>"000001010",
  25757=>"000000000",
  25758=>"101000000",
  25759=>"111111111",
  25760=>"000000000",
  25761=>"100111110",
  25762=>"111000000",
  25763=>"111000000",
  25764=>"001101001",
  25765=>"111000010",
  25766=>"111111111",
  25767=>"000000000",
  25768=>"001111111",
  25769=>"000000000",
  25770=>"000111111",
  25771=>"110111111",
  25772=>"000000000",
  25773=>"011011001",
  25774=>"100100111",
  25775=>"000111010",
  25776=>"111111111",
  25777=>"010111111",
  25778=>"101111010",
  25779=>"000101010",
  25780=>"101100100",
  25781=>"000000000",
  25782=>"000000000",
  25783=>"001011111",
  25784=>"111011111",
  25785=>"111111111",
  25786=>"000100100",
  25787=>"101100110",
  25788=>"011011001",
  25789=>"111101000",
  25790=>"111111010",
  25791=>"000011011",
  25792=>"001101101",
  25793=>"000000000",
  25794=>"111111111",
  25795=>"111111111",
  25796=>"000000000",
  25797=>"000011001",
  25798=>"111100000",
  25799=>"111110101",
  25800=>"111011111",
  25801=>"000000000",
  25802=>"000000000",
  25803=>"101111111",
  25804=>"100111110",
  25805=>"001111010",
  25806=>"000000000",
  25807=>"111111111",
  25808=>"000000000",
  25809=>"000000101",
  25810=>"111111010",
  25811=>"000000000",
  25812=>"000100110",
  25813=>"001110100",
  25814=>"000001000",
  25815=>"110111011",
  25816=>"000000000",
  25817=>"111101100",
  25818=>"000111000",
  25819=>"000000011",
  25820=>"111111111",
  25821=>"011001001",
  25822=>"011011011",
  25823=>"111111011",
  25824=>"001101111",
  25825=>"000000111",
  25826=>"000000000",
  25827=>"111111111",
  25828=>"000000000",
  25829=>"101111000",
  25830=>"110111111",
  25831=>"000111111",
  25832=>"000000010",
  25833=>"000000000",
  25834=>"000100101",
  25835=>"000010011",
  25836=>"000000000",
  25837=>"000000010",
  25838=>"110111111",
  25839=>"000000000",
  25840=>"001000000",
  25841=>"111111000",
  25842=>"000000000",
  25843=>"011101101",
  25844=>"101101111",
  25845=>"000000000",
  25846=>"011111011",
  25847=>"001000000",
  25848=>"000010000",
  25849=>"111111110",
  25850=>"111111111",
  25851=>"111111000",
  25852=>"011011011",
  25853=>"001000000",
  25854=>"000010011",
  25855=>"000000001",
  25856=>"111111000",
  25857=>"001111000",
  25858=>"111010000",
  25859=>"111111010",
  25860=>"001001111",
  25861=>"111111001",
  25862=>"000101111",
  25863=>"110110111",
  25864=>"011010000",
  25865=>"000000000",
  25866=>"111110110",
  25867=>"111111111",
  25868=>"001001001",
  25869=>"111011000",
  25870=>"111111000",
  25871=>"000011011",
  25872=>"000000000",
  25873=>"000101101",
  25874=>"011111011",
  25875=>"001010010",
  25876=>"111111011",
  25877=>"100000100",
  25878=>"011011001",
  25879=>"111111111",
  25880=>"111101011",
  25881=>"001001000",
  25882=>"000000000",
  25883=>"000111010",
  25884=>"000000000",
  25885=>"000000011",
  25886=>"001111111",
  25887=>"000111111",
  25888=>"011011001",
  25889=>"000000000",
  25890=>"111000000",
  25891=>"000000000",
  25892=>"000000110",
  25893=>"111011001",
  25894=>"000111111",
  25895=>"001000000",
  25896=>"110110010",
  25897=>"110111110",
  25898=>"000011110",
  25899=>"000000111",
  25900=>"010000000",
  25901=>"111111100",
  25902=>"110010111",
  25903=>"000000000",
  25904=>"110110110",
  25905=>"001001001",
  25906=>"000000010",
  25907=>"000000000",
  25908=>"110100111",
  25909=>"000111111",
  25910=>"100110011",
  25911=>"000000000",
  25912=>"000000111",
  25913=>"000001001",
  25914=>"000001001",
  25915=>"101000000",
  25916=>"000000100",
  25917=>"111110100",
  25918=>"100110110",
  25919=>"111111101",
  25920=>"000000000",
  25921=>"111110010",
  25922=>"011000000",
  25923=>"001000101",
  25924=>"111111111",
  25925=>"010011111",
  25926=>"111111111",
  25927=>"000000000",
  25928=>"000001001",
  25929=>"100000000",
  25930=>"000010000",
  25931=>"010110000",
  25932=>"011010000",
  25933=>"111111010",
  25934=>"000000000",
  25935=>"000110110",
  25936=>"100110100",
  25937=>"001000000",
  25938=>"111011000",
  25939=>"000000001",
  25940=>"101101001",
  25941=>"011011011",
  25942=>"110110010",
  25943=>"111110110",
  25944=>"001000000",
  25945=>"000011000",
  25946=>"111110110",
  25947=>"000000101",
  25948=>"111000000",
  25949=>"000000000",
  25950=>"000000000",
  25951=>"000111000",
  25952=>"000000000",
  25953=>"011011011",
  25954=>"010111111",
  25955=>"000011011",
  25956=>"110111111",
  25957=>"000000000",
  25958=>"111111111",
  25959=>"011011111",
  25960=>"111010000",
  25961=>"101001001",
  25962=>"000000001",
  25963=>"111101100",
  25964=>"110100100",
  25965=>"001011000",
  25966=>"000111111",
  25967=>"111110110",
  25968=>"000000000",
  25969=>"111010010",
  25970=>"111111000",
  25971=>"110110111",
  25972=>"011001001",
  25973=>"000000101",
  25974=>"101111111",
  25975=>"000000000",
  25976=>"000000000",
  25977=>"000010010",
  25978=>"010111111",
  25979=>"101001001",
  25980=>"111111111",
  25981=>"011111111",
  25982=>"000001111",
  25983=>"001001000",
  25984=>"111110110",
  25985=>"000010000",
  25986=>"000010110",
  25987=>"111101100",
  25988=>"000111000",
  25989=>"000000110",
  25990=>"000000000",
  25991=>"000000101",
  25992=>"010111111",
  25993=>"111101000",
  25994=>"000000000",
  25995=>"101101100",
  25996=>"000000000",
  25997=>"001001001",
  25998=>"111110110",
  25999=>"101000000",
  26000=>"111110110",
  26001=>"010111111",
  26002=>"011011010",
  26003=>"001011111",
  26004=>"000000000",
  26005=>"000000000",
  26006=>"111011000",
  26007=>"001001000",
  26008=>"100111111",
  26009=>"001000000",
  26010=>"001101001",
  26011=>"000000000",
  26012=>"110010010",
  26013=>"111101111",
  26014=>"101001011",
  26015=>"000000000",
  26016=>"001000101",
  26017=>"001001001",
  26018=>"111001000",
  26019=>"011011000",
  26020=>"011000000",
  26021=>"111111111",
  26022=>"000000000",
  26023=>"111111111",
  26024=>"100100110",
  26025=>"001100111",
  26026=>"111111111",
  26027=>"000100101",
  26028=>"111111001",
  26029=>"100000011",
  26030=>"000000000",
  26031=>"111111000",
  26032=>"111000000",
  26033=>"111111111",
  26034=>"000111111",
  26035=>"000000000",
  26036=>"011111111",
  26037=>"111001111",
  26038=>"001001111",
  26039=>"111001000",
  26040=>"111010010",
  26041=>"111111011",
  26042=>"111010000",
  26043=>"101111110",
  26044=>"000000101",
  26045=>"100000000",
  26046=>"101001111",
  26047=>"011011011",
  26048=>"000000111",
  26049=>"010010110",
  26050=>"000001001",
  26051=>"101011000",
  26052=>"111000000",
  26053=>"110111011",
  26054=>"000000000",
  26055=>"111001000",
  26056=>"111000100",
  26057=>"000010000",
  26058=>"001000000",
  26059=>"111111111",
  26060=>"111000000",
  26061=>"000110010",
  26062=>"000000000",
  26063=>"000000000",
  26064=>"110000000",
  26065=>"111111011",
  26066=>"111111111",
  26067=>"000101011",
  26068=>"111111111",
  26069=>"111011000",
  26070=>"111100100",
  26071=>"111100111",
  26072=>"000100101",
  26073=>"111101000",
  26074=>"001001000",
  26075=>"000111111",
  26076=>"111111100",
  26077=>"000100100",
  26078=>"000000001",
  26079=>"001111111",
  26080=>"111100111",
  26081=>"111111111",
  26082=>"101101101",
  26083=>"111100000",
  26084=>"111110000",
  26085=>"000000100",
  26086=>"011111111",
  26087=>"000000000",
  26088=>"000000000",
  26089=>"111111111",
  26090=>"000000101",
  26091=>"010011000",
  26092=>"000101111",
  26093=>"100100111",
  26094=>"100000100",
  26095=>"000000000",
  26096=>"100100001",
  26097=>"001001111",
  26098=>"111110100",
  26099=>"001000001",
  26100=>"001000001",
  26101=>"000000000",
  26102=>"110111110",
  26103=>"100111110",
  26104=>"110110000",
  26105=>"000001011",
  26106=>"101101111",
  26107=>"111111111",
  26108=>"000100111",
  26109=>"111111110",
  26110=>"111111111",
  26111=>"000000111",
  26112=>"110111011",
  26113=>"010000000",
  26114=>"111000100",
  26115=>"000000000",
  26116=>"111111001",
  26117=>"000000000",
  26118=>"000111111",
  26119=>"110000000",
  26120=>"111111111",
  26121=>"110111111",
  26122=>"000000000",
  26123=>"100100100",
  26124=>"000111111",
  26125=>"011111000",
  26126=>"000100011",
  26127=>"011010000",
  26128=>"110000000",
  26129=>"010111111",
  26130=>"000101110",
  26131=>"000000110",
  26132=>"111111111",
  26133=>"000000000",
  26134=>"000000000",
  26135=>"111000000",
  26136=>"000000000",
  26137=>"111111111",
  26138=>"111000100",
  26139=>"100011000",
  26140=>"111111111",
  26141=>"000000111",
  26142=>"100011001",
  26143=>"111111110",
  26144=>"011011000",
  26145=>"111111111",
  26146=>"000110110",
  26147=>"111111111",
  26148=>"111000001",
  26149=>"110110110",
  26150=>"011011000",
  26151=>"111000111",
  26152=>"100100100",
  26153=>"000110000",
  26154=>"000000100",
  26155=>"000000000",
  26156=>"000000110",
  26157=>"000000000",
  26158=>"000000111",
  26159=>"000001111",
  26160=>"111111001",
  26161=>"000001111",
  26162=>"000111111",
  26163=>"111111001",
  26164=>"110100000",
  26165=>"010000000",
  26166=>"000000001",
  26167=>"101000000",
  26168=>"000000000",
  26169=>"011110000",
  26170=>"000000000",
  26171=>"001101111",
  26172=>"111111101",
  26173=>"001011111",
  26174=>"010101111",
  26175=>"010010111",
  26176=>"100101111",
  26177=>"000110111",
  26178=>"100000001",
  26179=>"111111110",
  26180=>"000110111",
  26181=>"001100100",
  26182=>"111110000",
  26183=>"000000000",
  26184=>"001011101",
  26185=>"000000111",
  26186=>"111001101",
  26187=>"100110000",
  26188=>"111111111",
  26189=>"000000000",
  26190=>"000000000",
  26191=>"111111111",
  26192=>"000111110",
  26193=>"100110000",
  26194=>"000101010",
  26195=>"111100111",
  26196=>"000000110",
  26197=>"111111110",
  26198=>"111101110",
  26199=>"000001111",
  26200=>"111111100",
  26201=>"000000111",
  26202=>"111111111",
  26203=>"110111001",
  26204=>"111111001",
  26205=>"011111111",
  26206=>"000000011",
  26207=>"000000000",
  26208=>"001000010",
  26209=>"101101101",
  26210=>"111111111",
  26211=>"000100111",
  26212=>"111000000",
  26213=>"000000000",
  26214=>"000000000",
  26215=>"111111111",
  26216=>"111111111",
  26217=>"010000000",
  26218=>"001011111",
  26219=>"111111110",
  26220=>"011011111",
  26221=>"000000010",
  26222=>"000000000",
  26223=>"010111111",
  26224=>"101100111",
  26225=>"001000101",
  26226=>"000000011",
  26227=>"110000000",
  26228=>"000001000",
  26229=>"000000000",
  26230=>"000100000",
  26231=>"000000000",
  26232=>"000001111",
  26233=>"111100000",
  26234=>"100000000",
  26235=>"000111110",
  26236=>"001000001",
  26237=>"000000000",
  26238=>"000000000",
  26239=>"000101111",
  26240=>"110011011",
  26241=>"000000111",
  26242=>"110110111",
  26243=>"100001011",
  26244=>"000001111",
  26245=>"110000000",
  26246=>"001011000",
  26247=>"110111100",
  26248=>"111111111",
  26249=>"011000001",
  26250=>"000111111",
  26251=>"011001000",
  26252=>"111101111",
  26253=>"111111110",
  26254=>"110100110",
  26255=>"000111111",
  26256=>"001101111",
  26257=>"000000000",
  26258=>"111100111",
  26259=>"001000011",
  26260=>"100100101",
  26261=>"000010000",
  26262=>"110000000",
  26263=>"000000000",
  26264=>"100000000",
  26265=>"111111010",
  26266=>"000111111",
  26267=>"111111111",
  26268=>"111111110",
  26269=>"111110111",
  26270=>"111111111",
  26271=>"001001000",
  26272=>"111110110",
  26273=>"011110110",
  26274=>"000111111",
  26275=>"000000111",
  26276=>"111001001",
  26277=>"010000000",
  26278=>"111111111",
  26279=>"000011100",
  26280=>"000011010",
  26281=>"001100111",
  26282=>"000010111",
  26283=>"110110111",
  26284=>"000111111",
  26285=>"100100111",
  26286=>"000000111",
  26287=>"000000000",
  26288=>"000011111",
  26289=>"010011011",
  26290=>"011111011",
  26291=>"111000111",
  26292=>"110010000",
  26293=>"000100000",
  26294=>"011111111",
  26295=>"000000000",
  26296=>"000000000",
  26297=>"000111011",
  26298=>"111001000",
  26299=>"000000001",
  26300=>"000000000",
  26301=>"000111111",
  26302=>"100000000",
  26303=>"000000000",
  26304=>"000101011",
  26305=>"000110110",
  26306=>"110100100",
  26307=>"011111010",
  26308=>"000000111",
  26309=>"000000000",
  26310=>"110010000",
  26311=>"000101111",
  26312=>"010111011",
  26313=>"111111101",
  26314=>"111111100",
  26315=>"000000000",
  26316=>"000000000",
  26317=>"011111101",
  26318=>"111111111",
  26319=>"111111111",
  26320=>"000000111",
  26321=>"000000111",
  26322=>"111000001",
  26323=>"000000111",
  26324=>"100101001",
  26325=>"001011110",
  26326=>"000000000",
  26327=>"000000110",
  26328=>"000000000",
  26329=>"000000000",
  26330=>"000000110",
  26331=>"111111000",
  26332=>"111111111",
  26333=>"001001000",
  26334=>"111111001",
  26335=>"000000000",
  26336=>"000000111",
  26337=>"000000000",
  26338=>"011001011",
  26339=>"000000010",
  26340=>"000010111",
  26341=>"011111111",
  26342=>"010110111",
  26343=>"110111110",
  26344=>"111111111",
  26345=>"001101111",
  26346=>"111111100",
  26347=>"000000111",
  26348=>"001000000",
  26349=>"011000110",
  26350=>"111000000",
  26351=>"110000000",
  26352=>"011110010",
  26353=>"111000001",
  26354=>"111111111",
  26355=>"111111111",
  26356=>"111111111",
  26357=>"000100000",
  26358=>"011011011",
  26359=>"000000000",
  26360=>"000001111",
  26361=>"000011001",
  26362=>"000000010",
  26363=>"001111111",
  26364=>"001001001",
  26365=>"111111111",
  26366=>"001111100",
  26367=>"000001001",
  26368=>"101100000",
  26369=>"001000100",
  26370=>"111011001",
  26371=>"000000000",
  26372=>"000100110",
  26373=>"001000010",
  26374=>"000111111",
  26375=>"000000000",
  26376=>"000000000",
  26377=>"111111000",
  26378=>"111000000",
  26379=>"001001110",
  26380=>"000001001",
  26381=>"100101101",
  26382=>"111111000",
  26383=>"111110000",
  26384=>"000000000",
  26385=>"000000000",
  26386=>"000000000",
  26387=>"000000000",
  26388=>"000011111",
  26389=>"000111111",
  26390=>"011111001",
  26391=>"000000101",
  26392=>"001000100",
  26393=>"111111000",
  26394=>"111000000",
  26395=>"011011000",
  26396=>"000001011",
  26397=>"111111000",
  26398=>"000000000",
  26399=>"111101110",
  26400=>"110000100",
  26401=>"001011111",
  26402=>"000000000",
  26403=>"000000110",
  26404=>"110110111",
  26405=>"111111111",
  26406=>"101101111",
  26407=>"100000000",
  26408=>"000000000",
  26409=>"001111111",
  26410=>"100000100",
  26411=>"110110101",
  26412=>"000110000",
  26413=>"001001111",
  26414=>"000110011",
  26415=>"000000000",
  26416=>"111110110",
  26417=>"000000000",
  26418=>"000000011",
  26419=>"000110010",
  26420=>"111000000",
  26421=>"111010011",
  26422=>"111111010",
  26423=>"111111011",
  26424=>"000000000",
  26425=>"101001101",
  26426=>"000000000",
  26427=>"111111111",
  26428=>"110110111",
  26429=>"000110110",
  26430=>"001001000",
  26431=>"000111111",
  26432=>"111000000",
  26433=>"011011010",
  26434=>"111111111",
  26435=>"000000000",
  26436=>"000000111",
  26437=>"000010010",
  26438=>"000010000",
  26439=>"001001000",
  26440=>"111111111",
  26441=>"111010000",
  26442=>"111111111",
  26443=>"001001011",
  26444=>"111000000",
  26445=>"111111000",
  26446=>"111111111",
  26447=>"000001000",
  26448=>"000000000",
  26449=>"111111000",
  26450=>"001000111",
  26451=>"000001011",
  26452=>"000011111",
  26453=>"001001001",
  26454=>"111111011",
  26455=>"000000000",
  26456=>"010000011",
  26457=>"111001011",
  26458=>"001001000",
  26459=>"000000111",
  26460=>"110111111",
  26461=>"111000000",
  26462=>"111000111",
  26463=>"000100000",
  26464=>"000000000",
  26465=>"110000000",
  26466=>"001001111",
  26467=>"100000000",
  26468=>"000001011",
  26469=>"000000001",
  26470=>"010000000",
  26471=>"110100000",
  26472=>"001100111",
  26473=>"000011000",
  26474=>"000000000",
  26475=>"100000001",
  26476=>"001111111",
  26477=>"111010111",
  26478=>"000010000",
  26479=>"000000000",
  26480=>"000001111",
  26481=>"111111100",
  26482=>"111000001",
  26483=>"111111001",
  26484=>"000010111",
  26485=>"000000000",
  26486=>"110110100",
  26487=>"111111110",
  26488=>"000000111",
  26489=>"000000000",
  26490=>"011001011",
  26491=>"000011111",
  26492=>"000100111",
  26493=>"000100100",
  26494=>"000000000",
  26495=>"101000000",
  26496=>"111011001",
  26497=>"110111111",
  26498=>"010011001",
  26499=>"111110100",
  26500=>"111010111",
  26501=>"000000000",
  26502=>"100110111",
  26503=>"000000111",
  26504=>"000000001",
  26505=>"000000000",
  26506=>"111111000",
  26507=>"000110111",
  26508=>"111111111",
  26509=>"001000000",
  26510=>"110111111",
  26511=>"010111111",
  26512=>"110110010",
  26513=>"110000100",
  26514=>"011000000",
  26515=>"111111101",
  26516=>"111100000",
  26517=>"010000000",
  26518=>"111111111",
  26519=>"000000011",
  26520=>"111111111",
  26521=>"111111011",
  26522=>"000000000",
  26523=>"101111111",
  26524=>"011011110",
  26525=>"011101110",
  26526=>"111011101",
  26527=>"110111110",
  26528=>"111111000",
  26529=>"001000010",
  26530=>"000000100",
  26531=>"000000000",
  26532=>"110101111",
  26533=>"100000111",
  26534=>"001001101",
  26535=>"111111110",
  26536=>"111111111",
  26537=>"111111111",
  26538=>"111111111",
  26539=>"111111101",
  26540=>"000000000",
  26541=>"100111111",
  26542=>"111111111",
  26543=>"010011111",
  26544=>"100000000",
  26545=>"100111111",
  26546=>"000000000",
  26547=>"000100000",
  26548=>"000100100",
  26549=>"111000111",
  26550=>"000000000",
  26551=>"111111111",
  26552=>"110111111",
  26553=>"111111010",
  26554=>"000000000",
  26555=>"000010000",
  26556=>"001111111",
  26557=>"000110000",
  26558=>"000000000",
  26559=>"000000000",
  26560=>"001000000",
  26561=>"000000000",
  26562=>"000000001",
  26563=>"100000000",
  26564=>"001001111",
  26565=>"011111111",
  26566=>"111111110",
  26567=>"000000000",
  26568=>"001000000",
  26569=>"111110111",
  26570=>"000000100",
  26571=>"000000111",
  26572=>"110000000",
  26573=>"001000000",
  26574=>"111100111",
  26575=>"111000000",
  26576=>"100111111",
  26577=>"101101001",
  26578=>"010010000",
  26579=>"111111111",
  26580=>"000000111",
  26581=>"111000100",
  26582=>"111111111",
  26583=>"001111111",
  26584=>"000001111",
  26585=>"000000111",
  26586=>"000000110",
  26587=>"111101111",
  26588=>"111000000",
  26589=>"001000000",
  26590=>"111111111",
  26591=>"000011010",
  26592=>"110100110",
  26593=>"000000000",
  26594=>"111111111",
  26595=>"011011000",
  26596=>"111111001",
  26597=>"000111111",
  26598=>"011010010",
  26599=>"111010010",
  26600=>"001111111",
  26601=>"111111011",
  26602=>"000011111",
  26603=>"111111111",
  26604=>"111001011",
  26605=>"001000001",
  26606=>"101101001",
  26607=>"110001000",
  26608=>"100000000",
  26609=>"111111111",
  26610=>"100111111",
  26611=>"101000000",
  26612=>"100110111",
  26613=>"011000000",
  26614=>"100111111",
  26615=>"011010000",
  26616=>"000000111",
  26617=>"011011011",
  26618=>"000111111",
  26619=>"111100000",
  26620=>"111000111",
  26621=>"000111111",
  26622=>"000000011",
  26623=>"000000000",
  26624=>"110111111",
  26625=>"111010100",
  26626=>"001001111",
  26627=>"000000000",
  26628=>"111111111",
  26629=>"110110000",
  26630=>"101101001",
  26631=>"000000000",
  26632=>"100110100",
  26633=>"111011001",
  26634=>"111111111",
  26635=>"000000000",
  26636=>"011011011",
  26637=>"000000111",
  26638=>"111010010",
  26639=>"111111011",
  26640=>"000000000",
  26641=>"000000001",
  26642=>"111111111",
  26643=>"111111000",
  26644=>"111111111",
  26645=>"110111011",
  26646=>"000000000",
  26647=>"101000000",
  26648=>"000000000",
  26649=>"001001011",
  26650=>"000001001",
  26651=>"111011000",
  26652=>"111001111",
  26653=>"111001111",
  26654=>"001010100",
  26655=>"000010110",
  26656=>"001000111",
  26657=>"110111110",
  26658=>"111111111",
  26659=>"100100100",
  26660=>"011111111",
  26661=>"111111111",
  26662=>"000000000",
  26663=>"100100000",
  26664=>"111111111",
  26665=>"111111111",
  26666=>"111111111",
  26667=>"111111111",
  26668=>"000000000",
  26669=>"000011111",
  26670=>"111011011",
  26671=>"111111111",
  26672=>"000000111",
  26673=>"000000101",
  26674=>"100100000",
  26675=>"100001000",
  26676=>"000000000",
  26677=>"000000000",
  26678=>"100001000",
  26679=>"111111111",
  26680=>"101000010",
  26681=>"111111111",
  26682=>"111111111",
  26683=>"000000000",
  26684=>"000000000",
  26685=>"111111111",
  26686=>"010000001",
  26687=>"011011011",
  26688=>"010111010",
  26689=>"000111111",
  26690=>"011011111",
  26691=>"100000100",
  26692=>"000000000",
  26693=>"111011001",
  26694=>"001000000",
  26695=>"111100000",
  26696=>"000000001",
  26697=>"111111111",
  26698=>"111000000",
  26699=>"100110111",
  26700=>"000110100",
  26701=>"000000000",
  26702=>"000000000",
  26703=>"000111011",
  26704=>"111100000",
  26705=>"000000000",
  26706=>"000000000",
  26707=>"011011110",
  26708=>"000000001",
  26709=>"110111100",
  26710=>"111110110",
  26711=>"111111011",
  26712=>"100000000",
  26713=>"110110000",
  26714=>"111111110",
  26715=>"000111110",
  26716=>"111101111",
  26717=>"111111111",
  26718=>"101111111",
  26719=>"100000000",
  26720=>"100000100",
  26721=>"000001001",
  26722=>"011110000",
  26723=>"111111111",
  26724=>"101000000",
  26725=>"100100100",
  26726=>"000011011",
  26727=>"001000000",
  26728=>"000000000",
  26729=>"111111010",
  26730=>"101000000",
  26731=>"001001010",
  26732=>"110000010",
  26733=>"111111111",
  26734=>"000000000",
  26735=>"111111000",
  26736=>"000000000",
  26737=>"111111001",
  26738=>"011011011",
  26739=>"001000000",
  26740=>"111111111",
  26741=>"001111111",
  26742=>"010011011",
  26743=>"111011011",
  26744=>"001111111",
  26745=>"111111001",
  26746=>"000000000",
  26747=>"000001011",
  26748=>"000000000",
  26749=>"111111111",
  26750=>"100000000",
  26751=>"001001001",
  26752=>"110110111",
  26753=>"110100000",
  26754=>"000000000",
  26755=>"000000001",
  26756=>"111100100",
  26757=>"100000000",
  26758=>"000000000",
  26759=>"000000000",
  26760=>"000000000",
  26761=>"000000000",
  26762=>"111101101",
  26763=>"000000011",
  26764=>"000000000",
  26765=>"000000000",
  26766=>"110000111",
  26767=>"011110110",
  26768=>"000010111",
  26769=>"101111011",
  26770=>"000000001",
  26771=>"000000000",
  26772=>"111111111",
  26773=>"000001011",
  26774=>"111000000",
  26775=>"111011000",
  26776=>"111111011",
  26777=>"110100000",
  26778=>"111111111",
  26779=>"000000000",
  26780=>"101000000",
  26781=>"100100100",
  26782=>"000001101",
  26783=>"110000000",
  26784=>"111101110",
  26785=>"000000000",
  26786=>"111111111",
  26787=>"000000000",
  26788=>"100100111",
  26789=>"111101111",
  26790=>"111100111",
  26791=>"000001001",
  26792=>"100111111",
  26793=>"011011111",
  26794=>"101111000",
  26795=>"000001000",
  26796=>"111111000",
  26797=>"000011011",
  26798=>"111111101",
  26799=>"100000000",
  26800=>"111111000",
  26801=>"110111111",
  26802=>"111100100",
  26803=>"000000000",
  26804=>"001000000",
  26805=>"001001001",
  26806=>"111111011",
  26807=>"000000100",
  26808=>"000000001",
  26809=>"111111000",
  26810=>"110100100",
  26811=>"111100111",
  26812=>"111111111",
  26813=>"000000000",
  26814=>"111111111",
  26815=>"111111111",
  26816=>"111111111",
  26817=>"101000000",
  26818=>"000000000",
  26819=>"111111111",
  26820=>"000000000",
  26821=>"011110111",
  26822=>"111011010",
  26823=>"000000000",
  26824=>"000000000",
  26825=>"111111111",
  26826=>"100001001",
  26827=>"110111110",
  26828=>"111011011",
  26829=>"000110011",
  26830=>"000000000",
  26831=>"000000000",
  26832=>"111111001",
  26833=>"111110110",
  26834=>"000000111",
  26835=>"001111111",
  26836=>"110000000",
  26837=>"111111100",
  26838=>"011111111",
  26839=>"110000000",
  26840=>"000000000",
  26841=>"111000011",
  26842=>"000000000",
  26843=>"000000100",
  26844=>"100100111",
  26845=>"001111111",
  26846=>"001001011",
  26847=>"111111010",
  26848=>"000000000",
  26849=>"011111111",
  26850=>"111000000",
  26851=>"110000000",
  26852=>"001001001",
  26853=>"110110111",
  26854=>"000000100",
  26855=>"000000000",
  26856=>"000000000",
  26857=>"001001001",
  26858=>"000001111",
  26859=>"001000100",
  26860=>"000000000",
  26861=>"100111110",
  26862=>"000000111",
  26863=>"000000111",
  26864=>"111110000",
  26865=>"011011011",
  26866=>"100100000",
  26867=>"011101101",
  26868=>"110000001",
  26869=>"000000000",
  26870=>"000000101",
  26871=>"000000000",
  26872=>"000000001",
  26873=>"000000000",
  26874=>"100000101",
  26875=>"000000000",
  26876=>"001001111",
  26877=>"001001100",
  26878=>"000000000",
  26879=>"001011000",
  26880=>"000000000",
  26881=>"001011000",
  26882=>"111111110",
  26883=>"111001011",
  26884=>"101111101",
  26885=>"111100000",
  26886=>"110100000",
  26887=>"000000111",
  26888=>"111111111",
  26889=>"110110100",
  26890=>"001000011",
  26891=>"100000001",
  26892=>"000000000",
  26893=>"000000001",
  26894=>"000000000",
  26895=>"000111111",
  26896=>"000000011",
  26897=>"111111111",
  26898=>"111011011",
  26899=>"000000000",
  26900=>"000000000",
  26901=>"000000000",
  26902=>"000011011",
  26903=>"111111111",
  26904=>"101000000",
  26905=>"111111100",
  26906=>"111001011",
  26907=>"100100111",
  26908=>"000000011",
  26909=>"100000001",
  26910=>"111111111",
  26911=>"011101111",
  26912=>"000000000",
  26913=>"111100000",
  26914=>"111111000",
  26915=>"000000111",
  26916=>"110010011",
  26917=>"001000011",
  26918=>"001110111",
  26919=>"111111101",
  26920=>"011011010",
  26921=>"001101111",
  26922=>"001000000",
  26923=>"000000010",
  26924=>"000000000",
  26925=>"111111111",
  26926=>"000000000",
  26927=>"000000000",
  26928=>"110100111",
  26929=>"000110111",
  26930=>"110110000",
  26931=>"000000001",
  26932=>"000000000",
  26933=>"000001001",
  26934=>"110100001",
  26935=>"100101001",
  26936=>"111000000",
  26937=>"111000111",
  26938=>"110111111",
  26939=>"111111111",
  26940=>"111001001",
  26941=>"000000000",
  26942=>"000001001",
  26943=>"000000000",
  26944=>"111111111",
  26945=>"000000000",
  26946=>"111001001",
  26947=>"111111111",
  26948=>"100000001",
  26949=>"111111111",
  26950=>"111000000",
  26951=>"001001001",
  26952=>"110000000",
  26953=>"111111111",
  26954=>"111111111",
  26955=>"110110100",
  26956=>"000000000",
  26957=>"100000000",
  26958=>"000100101",
  26959=>"111101101",
  26960=>"000000000",
  26961=>"101100010",
  26962=>"100000001",
  26963=>"111100100",
  26964=>"000000000",
  26965=>"011011011",
  26966=>"000000000",
  26967=>"101001111",
  26968=>"111111011",
  26969=>"101111111",
  26970=>"000000000",
  26971=>"111110000",
  26972=>"110111111",
  26973=>"111111111",
  26974=>"111001101",
  26975=>"000010000",
  26976=>"111111111",
  26977=>"111011011",
  26978=>"011001000",
  26979=>"111111111",
  26980=>"101111111",
  26981=>"111111111",
  26982=>"111111111",
  26983=>"001001001",
  26984=>"001001000",
  26985=>"000100111",
  26986=>"111111111",
  26987=>"000000000",
  26988=>"110000000",
  26989=>"101000000",
  26990=>"000111111",
  26991=>"000100000",
  26992=>"000000000",
  26993=>"000010000",
  26994=>"000000000",
  26995=>"111000000",
  26996=>"110010100",
  26997=>"111001000",
  26998=>"000010010",
  26999=>"001001001",
  27000=>"111111111",
  27001=>"101000100",
  27002=>"111111111",
  27003=>"011111011",
  27004=>"000111111",
  27005=>"111111111",
  27006=>"011001011",
  27007=>"111111111",
  27008=>"000000000",
  27009=>"000000000",
  27010=>"100111111",
  27011=>"111111111",
  27012=>"000000000",
  27013=>"010010000",
  27014=>"000100100",
  27015=>"111000000",
  27016=>"000000000",
  27017=>"000000000",
  27018=>"000000000",
  27019=>"001011111",
  27020=>"111111111",
  27021=>"000010010",
  27022=>"111111000",
  27023=>"111111111",
  27024=>"110111111",
  27025=>"110111011",
  27026=>"000000000",
  27027=>"100101111",
  27028=>"000000000",
  27029=>"000000000",
  27030=>"111100000",
  27031=>"010000110",
  27032=>"111111111",
  27033=>"000000000",
  27034=>"000000000",
  27035=>"111001001",
  27036=>"010000000",
  27037=>"000000000",
  27038=>"001100000",
  27039=>"111111111",
  27040=>"100100000",
  27041=>"000000011",
  27042=>"110100011",
  27043=>"111111111",
  27044=>"111111111",
  27045=>"010110110",
  27046=>"000000000",
  27047=>"000000111",
  27048=>"000000000",
  27049=>"110101111",
  27050=>"000000111",
  27051=>"000000001",
  27052=>"100110000",
  27053=>"110111111",
  27054=>"000000000",
  27055=>"111111111",
  27056=>"000000000",
  27057=>"011011011",
  27058=>"100101011",
  27059=>"101111101",
  27060=>"111111100",
  27061=>"100110000",
  27062=>"111111000",
  27063=>"000000000",
  27064=>"111111010",
  27065=>"000000000",
  27066=>"111011001",
  27067=>"111111111",
  27068=>"111111111",
  27069=>"000000000",
  27070=>"111100000",
  27071=>"001011010",
  27072=>"000000001",
  27073=>"000000110",
  27074=>"011111111",
  27075=>"111000000",
  27076=>"111100101",
  27077=>"111100000",
  27078=>"111111111",
  27079=>"000010010",
  27080=>"111111000",
  27081=>"111100000",
  27082=>"111011011",
  27083=>"111111100",
  27084=>"000000000",
  27085=>"111000000",
  27086=>"111111111",
  27087=>"111111111",
  27088=>"000000000",
  27089=>"111010111",
  27090=>"100100111",
  27091=>"111111111",
  27092=>"010000000",
  27093=>"010110111",
  27094=>"000000000",
  27095=>"111111111",
  27096=>"000000000",
  27097=>"000001011",
  27098=>"100111111",
  27099=>"111111110",
  27100=>"000111011",
  27101=>"100000001",
  27102=>"111011001",
  27103=>"000011111",
  27104=>"011000100",
  27105=>"000110000",
  27106=>"111111110",
  27107=>"111100111",
  27108=>"111101111",
  27109=>"111111100",
  27110=>"011011011",
  27111=>"111111111",
  27112=>"101101101",
  27113=>"000000000",
  27114=>"111101111",
  27115=>"101110111",
  27116=>"111111111",
  27117=>"111110111",
  27118=>"111110111",
  27119=>"010000000",
  27120=>"000100110",
  27121=>"000000000",
  27122=>"000000000",
  27123=>"000000000",
  27124=>"001011101",
  27125=>"110110100",
  27126=>"111001001",
  27127=>"000011010",
  27128=>"000000000",
  27129=>"111110000",
  27130=>"001011001",
  27131=>"000000000",
  27132=>"010110110",
  27133=>"000000100",
  27134=>"110111111",
  27135=>"111000000",
  27136=>"000110110",
  27137=>"110000000",
  27138=>"111111110",
  27139=>"000100101",
  27140=>"001101100",
  27141=>"000000111",
  27142=>"111000000",
  27143=>"111111111",
  27144=>"100000000",
  27145=>"111111000",
  27146=>"000000000",
  27147=>"111000010",
  27148=>"111000100",
  27149=>"000010110",
  27150=>"000110110",
  27151=>"000011111",
  27152=>"111001011",
  27153=>"111000001",
  27154=>"111011111",
  27155=>"000000000",
  27156=>"001100100",
  27157=>"000110000",
  27158=>"000000000",
  27159=>"000001001",
  27160=>"000101000",
  27161=>"110111111",
  27162=>"111110111",
  27163=>"111111111",
  27164=>"000000000",
  27165=>"001000000",
  27166=>"100111111",
  27167=>"000011111",
  27168=>"011011000",
  27169=>"111111001",
  27170=>"000000011",
  27171=>"000000000",
  27172=>"000000000",
  27173=>"000001111",
  27174=>"001000100",
  27175=>"111011111",
  27176=>"101101001",
  27177=>"110000000",
  27178=>"000000000",
  27179=>"001001111",
  27180=>"111111111",
  27181=>"111111000",
  27182=>"111111110",
  27183=>"001000000",
  27184=>"111001000",
  27185=>"001001111",
  27186=>"110110011",
  27187=>"000000000",
  27188=>"000000000",
  27189=>"110010000",
  27190=>"101100001",
  27191=>"000000000",
  27192=>"001010110",
  27193=>"100000000",
  27194=>"000000000",
  27195=>"000000110",
  27196=>"111000000",
  27197=>"111000000",
  27198=>"110000001",
  27199=>"111001101",
  27200=>"100100111",
  27201=>"000000100",
  27202=>"000110111",
  27203=>"001001111",
  27204=>"000100110",
  27205=>"101101101",
  27206=>"111111101",
  27207=>"111111111",
  27208=>"001001000",
  27209=>"111001111",
  27210=>"111110010",
  27211=>"110000000",
  27212=>"000111111",
  27213=>"110110111",
  27214=>"100111111",
  27215=>"000000000",
  27216=>"000000000",
  27217=>"000001000",
  27218=>"100100111",
  27219=>"000111111",
  27220=>"110101000",
  27221=>"111111111",
  27222=>"101000000",
  27223=>"000000001",
  27224=>"000000000",
  27225=>"111111111",
  27226=>"001101101",
  27227=>"100110000",
  27228=>"000111111",
  27229=>"001111111",
  27230=>"111111001",
  27231=>"100111111",
  27232=>"111111111",
  27233=>"001111110",
  27234=>"111110110",
  27235=>"000000000",
  27236=>"000000000",
  27237=>"000000110",
  27238=>"101000000",
  27239=>"000010010",
  27240=>"000000110",
  27241=>"111111111",
  27242=>"111000000",
  27243=>"000000111",
  27244=>"111011001",
  27245=>"000000000",
  27246=>"101000111",
  27247=>"001000010",
  27248=>"001000011",
  27249=>"011011000",
  27250=>"111111000",
  27251=>"100111010",
  27252=>"111001000",
  27253=>"111111100",
  27254=>"000001000",
  27255=>"111000000",
  27256=>"011011011",
  27257=>"111000000",
  27258=>"111110000",
  27259=>"010001000",
  27260=>"110111111",
  27261=>"100111111",
  27262=>"111111111",
  27263=>"000000000",
  27264=>"111011000",
  27265=>"011010000",
  27266=>"111011111",
  27267=>"000011100",
  27268=>"111111000",
  27269=>"011000000",
  27270=>"111111001",
  27271=>"000000000",
  27272=>"000000101",
  27273=>"111111011",
  27274=>"000000100",
  27275=>"111101000",
  27276=>"111111111",
  27277=>"000011011",
  27278=>"001001111",
  27279=>"000000000",
  27280=>"100111111",
  27281=>"000000000",
  27282=>"001000111",
  27283=>"001011011",
  27284=>"000000111",
  27285=>"000100111",
  27286=>"000000000",
  27287=>"111000000",
  27288=>"110000000",
  27289=>"111000000",
  27290=>"101101000",
  27291=>"000010000",
  27292=>"111111000",
  27293=>"100110011",
  27294=>"001111000",
  27295=>"110010111",
  27296=>"101001001",
  27297=>"100111111",
  27298=>"000000000",
  27299=>"111100001",
  27300=>"111001000",
  27301=>"110000000",
  27302=>"000000111",
  27303=>"111101001",
  27304=>"111111110",
  27305=>"000000100",
  27306=>"000010000",
  27307=>"000000110",
  27308=>"111110111",
  27309=>"000111111",
  27310=>"011000000",
  27311=>"101111111",
  27312=>"110111111",
  27313=>"101101111",
  27314=>"111011010",
  27315=>"100101111",
  27316=>"101101111",
  27317=>"000000000",
  27318=>"000000000",
  27319=>"011111111",
  27320=>"101000000",
  27321=>"111000000",
  27322=>"111110110",
  27323=>"000010111",
  27324=>"000000111",
  27325=>"000111111",
  27326=>"111111111",
  27327=>"100111111",
  27328=>"111111111",
  27329=>"001001111",
  27330=>"000110000",
  27331=>"100100111",
  27332=>"000010000",
  27333=>"111111110",
  27334=>"110010000",
  27335=>"000011111",
  27336=>"000000000",
  27337=>"101111111",
  27338=>"101000000",
  27339=>"011011000",
  27340=>"111011111",
  27341=>"100001001",
  27342=>"001001001",
  27343=>"111111001",
  27344=>"110000010",
  27345=>"111000000",
  27346=>"001101100",
  27347=>"011011000",
  27348=>"111111000",
  27349=>"100110110",
  27350=>"111111000",
  27351=>"100100100",
  27352=>"111111001",
  27353=>"000111111",
  27354=>"111111000",
  27355=>"000001111",
  27356=>"000100111",
  27357=>"110111111",
  27358=>"111000000",
  27359=>"001000000",
  27360=>"000000000",
  27361=>"000000000",
  27362=>"011000111",
  27363=>"111111001",
  27364=>"100000011",
  27365=>"011011011",
  27366=>"111111111",
  27367=>"101111010",
  27368=>"000000000",
  27369=>"111111111",
  27370=>"000001000",
  27371=>"000001110",
  27372=>"000000000",
  27373=>"101100111",
  27374=>"000000110",
  27375=>"011000000",
  27376=>"000000000",
  27377=>"100000001",
  27378=>"001001001",
  27379=>"011011000",
  27380=>"000000111",
  27381=>"000101101",
  27382=>"110111111",
  27383=>"111010011",
  27384=>"111111111",
  27385=>"110000000",
  27386=>"100000100",
  27387=>"000111111",
  27388=>"100111101",
  27389=>"111100100",
  27390=>"111100000",
  27391=>"001111111",
  27392=>"111000000",
  27393=>"001111011",
  27394=>"111111011",
  27395=>"000111111",
  27396=>"000000100",
  27397=>"110111100",
  27398=>"110000000",
  27399=>"111111111",
  27400=>"101101011",
  27401=>"000000000",
  27402=>"000000111",
  27403=>"111000100",
  27404=>"111111111",
  27405=>"000000000",
  27406=>"100111111",
  27407=>"111111111",
  27408=>"110110110",
  27409=>"111011001",
  27410=>"111001001",
  27411=>"111000111",
  27412=>"000111001",
  27413=>"111111111",
  27414=>"100100100",
  27415=>"111111111",
  27416=>"100100101",
  27417=>"100100111",
  27418=>"111101001",
  27419=>"000000000",
  27420=>"000100100",
  27421=>"111111111",
  27422=>"111111111",
  27423=>"000010111",
  27424=>"111111000",
  27425=>"000000000",
  27426=>"111111111",
  27427=>"000101101",
  27428=>"100001001",
  27429=>"111111111",
  27430=>"000000000",
  27431=>"111110000",
  27432=>"000000000",
  27433=>"101111000",
  27434=>"000011100",
  27435=>"000111111",
  27436=>"011010000",
  27437=>"110100000",
  27438=>"000000111",
  27439=>"000000011",
  27440=>"000001001",
  27441=>"000000001",
  27442=>"111111111",
  27443=>"010000000",
  27444=>"111111000",
  27445=>"111011010",
  27446=>"100100111",
  27447=>"111000000",
  27448=>"000110110",
  27449=>"111000000",
  27450=>"111111111",
  27451=>"111111000",
  27452=>"111100101",
  27453=>"000000111",
  27454=>"000100111",
  27455=>"011011111",
  27456=>"000000100",
  27457=>"110100111",
  27458=>"100111101",
  27459=>"111110000",
  27460=>"000000000",
  27461=>"000100111",
  27462=>"111001111",
  27463=>"111001000",
  27464=>"010000111",
  27465=>"000000000",
  27466=>"001110111",
  27467=>"001110110",
  27468=>"011111111",
  27469=>"000000111",
  27470=>"100000000",
  27471=>"000000110",
  27472=>"000000001",
  27473=>"000000000",
  27474=>"001111111",
  27475=>"100111111",
  27476=>"000000000",
  27477=>"010111111",
  27478=>"000000000",
  27479=>"101111111",
  27480=>"110111111",
  27481=>"000000011",
  27482=>"000000110",
  27483=>"010000000",
  27484=>"000000100",
  27485=>"101111000",
  27486=>"000111110",
  27487=>"001100101",
  27488=>"001111111",
  27489=>"100111111",
  27490=>"101111111",
  27491=>"111000010",
  27492=>"000000000",
  27493=>"101111111",
  27494=>"111000000",
  27495=>"000000000",
  27496=>"100110111",
  27497=>"011111110",
  27498=>"011111111",
  27499=>"000001101",
  27500=>"001101111",
  27501=>"111000100",
  27502=>"001111111",
  27503=>"000101111",
  27504=>"110111011",
  27505=>"100000010",
  27506=>"111000111",
  27507=>"011111111",
  27508=>"000111111",
  27509=>"101100100",
  27510=>"000100111",
  27511=>"000000101",
  27512=>"111000000",
  27513=>"111111000",
  27514=>"111111001",
  27515=>"111001000",
  27516=>"111001001",
  27517=>"011000000",
  27518=>"111101000",
  27519=>"100111001",
  27520=>"001111111",
  27521=>"000000000",
  27522=>"101111111",
  27523=>"000000111",
  27524=>"011000110",
  27525=>"010111000",
  27526=>"011111100",
  27527=>"100100000",
  27528=>"100000111",
  27529=>"111000000",
  27530=>"000100000",
  27531=>"000000000",
  27532=>"001111100",
  27533=>"000111111",
  27534=>"000000111",
  27535=>"000000000",
  27536=>"000101100",
  27537=>"111111111",
  27538=>"000010010",
  27539=>"111100110",
  27540=>"000011011",
  27541=>"000000000",
  27542=>"100000000",
  27543=>"110110110",
  27544=>"111111111",
  27545=>"001100100",
  27546=>"111000000",
  27547=>"111111111",
  27548=>"111011000",
  27549=>"000010000",
  27550=>"000011011",
  27551=>"111111000",
  27552=>"111011000",
  27553=>"000111111",
  27554=>"100100100",
  27555=>"111111111",
  27556=>"111010100",
  27557=>"000000000",
  27558=>"111000000",
  27559=>"000000000",
  27560=>"100111100",
  27561=>"110100101",
  27562=>"001011111",
  27563=>"000011111",
  27564=>"000000000",
  27565=>"000000111",
  27566=>"000111111",
  27567=>"110111111",
  27568=>"110100111",
  27569=>"111000000",
  27570=>"000110000",
  27571=>"000111111",
  27572=>"111111000",
  27573=>"111000000",
  27574=>"111111111",
  27575=>"111110000",
  27576=>"000000011",
  27577=>"000011011",
  27578=>"001101111",
  27579=>"000101111",
  27580=>"111001000",
  27581=>"001001101",
  27582=>"111111110",
  27583=>"110101001",
  27584=>"111011000",
  27585=>"100000110",
  27586=>"000000011",
  27587=>"101111001",
  27588=>"100000000",
  27589=>"111011010",
  27590=>"000000000",
  27591=>"111111110",
  27592=>"111000000",
  27593=>"111101000",
  27594=>"000000000",
  27595=>"001001111",
  27596=>"000000010",
  27597=>"011011111",
  27598=>"011111010",
  27599=>"101000100",
  27600=>"000000000",
  27601=>"001111011",
  27602=>"111111111",
  27603=>"001000000",
  27604=>"001001000",
  27605=>"111111000",
  27606=>"000000001",
  27607=>"100000000",
  27608=>"101011000",
  27609=>"000111010",
  27610=>"000010011",
  27611=>"011000000",
  27612=>"101111111",
  27613=>"001010111",
  27614=>"000011011",
  27615=>"000100100",
  27616=>"011111011",
  27617=>"011001111",
  27618=>"110111111",
  27619=>"110000000",
  27620=>"000000001",
  27621=>"101001111",
  27622=>"111100000",
  27623=>"000000000",
  27624=>"011111111",
  27625=>"000000100",
  27626=>"001000010",
  27627=>"100110100",
  27628=>"000110111",
  27629=>"000011011",
  27630=>"000000000",
  27631=>"000000001",
  27632=>"111111111",
  27633=>"111111001",
  27634=>"100000000",
  27635=>"110000000",
  27636=>"001111111",
  27637=>"101001111",
  27638=>"100100000",
  27639=>"000000100",
  27640=>"111111001",
  27641=>"001111111",
  27642=>"011111110",
  27643=>"111111111",
  27644=>"111111000",
  27645=>"001100100",
  27646=>"000000000",
  27647=>"110011011",
  27648=>"111111111",
  27649=>"101001001",
  27650=>"101101101",
  27651=>"000000111",
  27652=>"100110111",
  27653=>"010000000",
  27654=>"111111111",
  27655=>"000000001",
  27656=>"010110111",
  27657=>"011111110",
  27658=>"111010011",
  27659=>"110111111",
  27660=>"001001101",
  27661=>"110000001",
  27662=>"111111001",
  27663=>"101100000",
  27664=>"111111111",
  27665=>"011110111",
  27666=>"000000000",
  27667=>"000000001",
  27668=>"111111111",
  27669=>"000000101",
  27670=>"110110100",
  27671=>"000000000",
  27672=>"101001111",
  27673=>"111111100",
  27674=>"000000000",
  27675=>"100000000",
  27676=>"111011111",
  27677=>"110011010",
  27678=>"000100100",
  27679=>"111111111",
  27680=>"000000110",
  27681=>"110000000",
  27682=>"111111110",
  27683=>"111111111",
  27684=>"111111111",
  27685=>"000010000",
  27686=>"111111111",
  27687=>"011000000",
  27688=>"100110111",
  27689=>"000011111",
  27690=>"111101111",
  27691=>"111110111",
  27692=>"111011011",
  27693=>"000000000",
  27694=>"111111111",
  27695=>"101001001",
  27696=>"111111011",
  27697=>"000000000",
  27698=>"000000000",
  27699=>"111111111",
  27700=>"110010110",
  27701=>"000000000",
  27702=>"100110110",
  27703=>"101100111",
  27704=>"000001000",
  27705=>"000000000",
  27706=>"111111111",
  27707=>"000000000",
  27708=>"111111111",
  27709=>"100000000",
  27710=>"111111111",
  27711=>"111111111",
  27712=>"000000000",
  27713=>"010011111",
  27714=>"111110110",
  27715=>"111111111",
  27716=>"111111111",
  27717=>"100100100",
  27718=>"011111101",
  27719=>"111111011",
  27720=>"010000000",
  27721=>"111111111",
  27722=>"000000011",
  27723=>"111110111",
  27724=>"110000110",
  27725=>"110100111",
  27726=>"111111100",
  27727=>"000011000",
  27728=>"111111111",
  27729=>"000000000",
  27730=>"011011000",
  27731=>"111111001",
  27732=>"111111111",
  27733=>"000010000",
  27734=>"111011011",
  27735=>"101111111",
  27736=>"111011111",
  27737=>"000000111",
  27738=>"000000010",
  27739=>"111111111",
  27740=>"000000011",
  27741=>"111111111",
  27742=>"111111001",
  27743=>"111111111",
  27744=>"111111100",
  27745=>"000000000",
  27746=>"000000101",
  27747=>"000000000",
  27748=>"111111111",
  27749=>"111101110",
  27750=>"000000000",
  27751=>"010110000",
  27752=>"000000001",
  27753=>"010010011",
  27754=>"011010000",
  27755=>"110000001",
  27756=>"111111110",
  27757=>"001001111",
  27758=>"000000110",
  27759=>"000111111",
  27760=>"111000000",
  27761=>"000000110",
  27762=>"000000001",
  27763=>"000000001",
  27764=>"000000000",
  27765=>"001101111",
  27766=>"000000000",
  27767=>"111111111",
  27768=>"101001111",
  27769=>"111100000",
  27770=>"111111000",
  27771=>"011011000",
  27772=>"100000000",
  27773=>"000000000",
  27774=>"000000000",
  27775=>"000000000",
  27776=>"000000101",
  27777=>"111111111",
  27778=>"000000000",
  27779=>"001001000",
  27780=>"000000000",
  27781=>"111111111",
  27782=>"001000110",
  27783=>"000000000",
  27784=>"011011111",
  27785=>"000000000",
  27786=>"011111111",
  27787=>"000000000",
  27788=>"000000111",
  27789=>"111111110",
  27790=>"000000111",
  27791=>"111100111",
  27792=>"000000000",
  27793=>"000000000",
  27794=>"111111101",
  27795=>"001000000",
  27796=>"000000110",
  27797=>"111111011",
  27798=>"000000011",
  27799=>"001000000",
  27800=>"100111111",
  27801=>"111111111",
  27802=>"111111111",
  27803=>"000000001",
  27804=>"111100000",
  27805=>"100000000",
  27806=>"100000000",
  27807=>"111111111",
  27808=>"111000000",
  27809=>"110000100",
  27810=>"000000000",
  27811=>"000000110",
  27812=>"100100111",
  27813=>"111000000",
  27814=>"110000000",
  27815=>"000000000",
  27816=>"110100111",
  27817=>"000000000",
  27818=>"001000100",
  27819=>"000000001",
  27820=>"001001111",
  27821=>"100110111",
  27822=>"100111111",
  27823=>"000011011",
  27824=>"111111111",
  27825=>"111110111",
  27826=>"110110010",
  27827=>"001000000",
  27828=>"111111001",
  27829=>"111111111",
  27830=>"000000000",
  27831=>"000001001",
  27832=>"000110110",
  27833=>"000000000",
  27834=>"100100100",
  27835=>"100100000",
  27836=>"000110110",
  27837=>"000000000",
  27838=>"111111111",
  27839=>"000110111",
  27840=>"011011011",
  27841=>"000000000",
  27842=>"000000000",
  27843=>"110000000",
  27844=>"111111010",
  27845=>"011111111",
  27846=>"111111111",
  27847=>"011011111",
  27848=>"111111111",
  27849=>"000000000",
  27850=>"100001111",
  27851=>"000000001",
  27852=>"000000100",
  27853=>"000011011",
  27854=>"111111111",
  27855=>"000000000",
  27856=>"111111111",
  27857=>"000111111",
  27858=>"000011111",
  27859=>"001101111",
  27860=>"111111111",
  27861=>"111111111",
  27862=>"000000011",
  27863=>"111111111",
  27864=>"000000000",
  27865=>"000000000",
  27866=>"000000000",
  27867=>"110010000",
  27868=>"100100000",
  27869=>"000000000",
  27870=>"000000011",
  27871=>"001101100",
  27872=>"010010000",
  27873=>"000110111",
  27874=>"110010111",
  27875=>"000000000",
  27876=>"000000000",
  27877=>"111111111",
  27878=>"000000000",
  27879=>"111111111",
  27880=>"000100000",
  27881=>"010000000",
  27882=>"010011010",
  27883=>"000000100",
  27884=>"111111111",
  27885=>"111011011",
  27886=>"001001111",
  27887=>"000000000",
  27888=>"100111111",
  27889=>"111111111",
  27890=>"000001001",
  27891=>"000111111",
  27892=>"000000000",
  27893=>"110110110",
  27894=>"001001001",
  27895=>"111111111",
  27896=>"011011111",
  27897=>"111111110",
  27898=>"000100000",
  27899=>"110110110",
  27900=>"001011011",
  27901=>"110110111",
  27902=>"111000111",
  27903=>"000111111",
  27904=>"100111111",
  27905=>"111111111",
  27906=>"000000000",
  27907=>"000000000",
  27908=>"111111111",
  27909=>"000000000",
  27910=>"001001000",
  27911=>"001001001",
  27912=>"111110110",
  27913=>"000000000",
  27914=>"111111111",
  27915=>"000011111",
  27916=>"100100100",
  27917=>"111111111",
  27918=>"001001000",
  27919=>"000100100",
  27920=>"001000101",
  27921=>"000000000",
  27922=>"011000000",
  27923=>"111100111",
  27924=>"000100111",
  27925=>"001000000",
  27926=>"000000000",
  27927=>"111111111",
  27928=>"000000000",
  27929=>"000000001",
  27930=>"000000000",
  27931=>"000000110",
  27932=>"111000000",
  27933=>"000000001",
  27934=>"000010111",
  27935=>"000011011",
  27936=>"001011001",
  27937=>"111111111",
  27938=>"001011011",
  27939=>"000000000",
  27940=>"111000000",
  27941=>"000000011",
  27942=>"111010100",
  27943=>"001100111",
  27944=>"111110101",
  27945=>"000000000",
  27946=>"000000011",
  27947=>"000000000",
  27948=>"111111111",
  27949=>"110110110",
  27950=>"000000000",
  27951=>"000000000",
  27952=>"000000000",
  27953=>"000000000",
  27954=>"111111110",
  27955=>"011011000",
  27956=>"110111110",
  27957=>"001011001",
  27958=>"010010111",
  27959=>"111111111",
  27960=>"001000000",
  27961=>"000000000",
  27962=>"000000100",
  27963=>"111111111",
  27964=>"100101001",
  27965=>"100000000",
  27966=>"000000000",
  27967=>"001000000",
  27968=>"000000001",
  27969=>"000000000",
  27970=>"111111111",
  27971=>"111111111",
  27972=>"011000000",
  27973=>"100100110",
  27974=>"111001000",
  27975=>"000000000",
  27976=>"000000000",
  27977=>"000111111",
  27978=>"111111111",
  27979=>"001001000",
  27980=>"000110111",
  27981=>"000111000",
  27982=>"111000111",
  27983=>"000000000",
  27984=>"000111100",
  27985=>"000000000",
  27986=>"000000000",
  27987=>"001000000",
  27988=>"000000000",
  27989=>"001001001",
  27990=>"100000000",
  27991=>"000000110",
  27992=>"101111111",
  27993=>"001111000",
  27994=>"001000010",
  27995=>"001011011",
  27996=>"000000000",
  27997=>"011000111",
  27998=>"000000000",
  27999=>"110111110",
  28000=>"111000000",
  28001=>"010111111",
  28002=>"000000000",
  28003=>"000000000",
  28004=>"100110110",
  28005=>"100000000",
  28006=>"000000000",
  28007=>"100100100",
  28008=>"011011111",
  28009=>"000000000",
  28010=>"111111111",
  28011=>"101001111",
  28012=>"100110100",
  28013=>"100100101",
  28014=>"000000000",
  28015=>"011001011",
  28016=>"000110011",
  28017=>"001011111",
  28018=>"000100111",
  28019=>"101100000",
  28020=>"000111111",
  28021=>"100000100",
  28022=>"111001011",
  28023=>"000100100",
  28024=>"111101101",
  28025=>"111000000",
  28026=>"110110100",
  28027=>"000000000",
  28028=>"111111111",
  28029=>"111111111",
  28030=>"111111111",
  28031=>"000000100",
  28032=>"100100111",
  28033=>"000000100",
  28034=>"111111111",
  28035=>"111101111",
  28036=>"000000000",
  28037=>"000000000",
  28038=>"000000011",
  28039=>"001111111",
  28040=>"110110000",
  28041=>"111111100",
  28042=>"001000000",
  28043=>"000000111",
  28044=>"111111111",
  28045=>"111111111",
  28046=>"000000000",
  28047=>"111111111",
  28048=>"010000010",
  28049=>"000000000",
  28050=>"110011111",
  28051=>"111001111",
  28052=>"010111111",
  28053=>"000010000",
  28054=>"000000010",
  28055=>"111111111",
  28056=>"001000000",
  28057=>"111111111",
  28058=>"001000000",
  28059=>"110000111",
  28060=>"000000111",
  28061=>"111000000",
  28062=>"000000000",
  28063=>"000000000",
  28064=>"110111000",
  28065=>"001000001",
  28066=>"100000101",
  28067=>"000000000",
  28068=>"110111111",
  28069=>"111111000",
  28070=>"111111111",
  28071=>"000000000",
  28072=>"000011011",
  28073=>"000100111",
  28074=>"110111111",
  28075=>"000000000",
  28076=>"111111000",
  28077=>"000000000",
  28078=>"000000000",
  28079=>"110110100",
  28080=>"111111111",
  28081=>"000000000",
  28082=>"000000000",
  28083=>"111111111",
  28084=>"000000000",
  28085=>"000000000",
  28086=>"110110110",
  28087=>"111110000",
  28088=>"111001000",
  28089=>"111111011",
  28090=>"001101111",
  28091=>"110110000",
  28092=>"000000011",
  28093=>"100000101",
  28094=>"000000100",
  28095=>"101111111",
  28096=>"111111111",
  28097=>"000000000",
  28098=>"000010111",
  28099=>"101111111",
  28100=>"011011111",
  28101=>"110000100",
  28102=>"000000000",
  28103=>"000000000",
  28104=>"000000000",
  28105=>"000000000",
  28106=>"001000100",
  28107=>"000000000",
  28108=>"110000000",
  28109=>"111111111",
  28110=>"000000000",
  28111=>"111111011",
  28112=>"000101001",
  28113=>"100000001",
  28114=>"000000000",
  28115=>"000010000",
  28116=>"111111111",
  28117=>"011110000",
  28118=>"000000111",
  28119=>"010011001",
  28120=>"111011000",
  28121=>"000110000",
  28122=>"000000000",
  28123=>"000000000",
  28124=>"100000110",
  28125=>"111110111",
  28126=>"111111111",
  28127=>"100011111",
  28128=>"000000000",
  28129=>"111101011",
  28130=>"000001001",
  28131=>"000000000",
  28132=>"000000000",
  28133=>"111111111",
  28134=>"000000000",
  28135=>"011000111",
  28136=>"111111111",
  28137=>"100000000",
  28138=>"000011010",
  28139=>"111111011",
  28140=>"000000000",
  28141=>"111110110",
  28142=>"000000010",
  28143=>"000000000",
  28144=>"010111111",
  28145=>"000000000",
  28146=>"111000000",
  28147=>"111111111",
  28148=>"000001000",
  28149=>"000000011",
  28150=>"111111001",
  28151=>"110110000",
  28152=>"000000001",
  28153=>"000110110",
  28154=>"011000001",
  28155=>"111111111",
  28156=>"000111111",
  28157=>"111111111",
  28158=>"111111111",
  28159=>"111111111",
  28160=>"111111100",
  28161=>"100111111",
  28162=>"000000000",
  28163=>"000100100",
  28164=>"110110000",
  28165=>"000000000",
  28166=>"011000011",
  28167=>"111111111",
  28168=>"000000010",
  28169=>"011111001",
  28170=>"000111111",
  28171=>"111111111",
  28172=>"000000000",
  28173=>"111111000",
  28174=>"001111111",
  28175=>"111101100",
  28176=>"011011111",
  28177=>"111011000",
  28178=>"000000000",
  28179=>"000000000",
  28180=>"000000000",
  28181=>"111001111",
  28182=>"000001001",
  28183=>"101000100",
  28184=>"111111111",
  28185=>"100111111",
  28186=>"111110000",
  28187=>"000110111",
  28188=>"000000000",
  28189=>"100100000",
  28190=>"110000001",
  28191=>"111000010",
  28192=>"110100100",
  28193=>"010100110",
  28194=>"000000000",
  28195=>"111111111",
  28196=>"100111000",
  28197=>"000000010",
  28198=>"000000000",
  28199=>"000011110",
  28200=>"000000000",
  28201=>"000000000",
  28202=>"111111100",
  28203=>"000000000",
  28204=>"111000000",
  28205=>"111111000",
  28206=>"111001001",
  28207=>"000000000",
  28208=>"111101101",
  28209=>"111111000",
  28210=>"111111000",
  28211=>"011110000",
  28212=>"111011000",
  28213=>"111000000",
  28214=>"111111001",
  28215=>"000000000",
  28216=>"010010001",
  28217=>"000000000",
  28218=>"001111111",
  28219=>"000000111",
  28220=>"111111111",
  28221=>"100000000",
  28222=>"000110110",
  28223=>"111001101",
  28224=>"010000100",
  28225=>"011000011",
  28226=>"111000000",
  28227=>"010110111",
  28228=>"111001001",
  28229=>"111110100",
  28230=>"000011111",
  28231=>"111111111",
  28232=>"101101000",
  28233=>"000000001",
  28234=>"011111110",
  28235=>"111111111",
  28236=>"001011011",
  28237=>"000000000",
  28238=>"111000000",
  28239=>"000000110",
  28240=>"000000000",
  28241=>"100000000",
  28242=>"000101111",
  28243=>"000001111",
  28244=>"000000000",
  28245=>"111110000",
  28246=>"111111101",
  28247=>"000101000",
  28248=>"001000000",
  28249=>"000001111",
  28250=>"111111111",
  28251=>"000000000",
  28252=>"000000010",
  28253=>"111111111",
  28254=>"000000000",
  28255=>"001101100",
  28256=>"000111111",
  28257=>"001101101",
  28258=>"111111001",
  28259=>"000000000",
  28260=>"000000000",
  28261=>"110000000",
  28262=>"111111100",
  28263=>"000000010",
  28264=>"111111111",
  28265=>"111111111",
  28266=>"000110000",
  28267=>"001001000",
  28268=>"000111111",
  28269=>"000000000",
  28270=>"000010111",
  28271=>"100111111",
  28272=>"111110110",
  28273=>"000000000",
  28274=>"111111001",
  28275=>"101111111",
  28276=>"000100011",
  28277=>"000000111",
  28278=>"000000000",
  28279=>"010000000",
  28280=>"111000000",
  28281=>"001000000",
  28282=>"000111111",
  28283=>"000000000",
  28284=>"111111111",
  28285=>"011111111",
  28286=>"111111110",
  28287=>"011000111",
  28288=>"111111111",
  28289=>"000000001",
  28290=>"111111111",
  28291=>"110110000",
  28292=>"111111110",
  28293=>"111100111",
  28294=>"111111111",
  28295=>"000000111",
  28296=>"111001000",
  28297=>"000000101",
  28298=>"000010000",
  28299=>"000000000",
  28300=>"000100111",
  28301=>"000000000",
  28302=>"100111111",
  28303=>"111111100",
  28304=>"001000000",
  28305=>"011000000",
  28306=>"111111000",
  28307=>"000111110",
  28308=>"110110100",
  28309=>"111111111",
  28310=>"111111100",
  28311=>"111111000",
  28312=>"000000000",
  28313=>"100000111",
  28314=>"111000000",
  28315=>"000000000",
  28316=>"111101101",
  28317=>"110111111",
  28318=>"001111111",
  28319=>"111010111",
  28320=>"111111111",
  28321=>"001111001",
  28322=>"000110010",
  28323=>"011111011",
  28324=>"000110000",
  28325=>"011010110",
  28326=>"000000000",
  28327=>"111100000",
  28328=>"000000000",
  28329=>"111110111",
  28330=>"001000000",
  28331=>"000111111",
  28332=>"111111111",
  28333=>"100111111",
  28334=>"111111001",
  28335=>"000010111",
  28336=>"000000111",
  28337=>"001000011",
  28338=>"110111110",
  28339=>"000000000",
  28340=>"000000000",
  28341=>"111111111",
  28342=>"111111111",
  28343=>"000011010",
  28344=>"100000001",
  28345=>"000000001",
  28346=>"000000111",
  28347=>"000111111",
  28348=>"000000000",
  28349=>"000000100",
  28350=>"111000000",
  28351=>"111111111",
  28352=>"000000000",
  28353=>"000000000",
  28354=>"011011011",
  28355=>"100000000",
  28356=>"000111111",
  28357=>"110110100",
  28358=>"101111000",
  28359=>"110000000",
  28360=>"110101111",
  28361=>"000000010",
  28362=>"101000000",
  28363=>"000010011",
  28364=>"000111111",
  28365=>"101000111",
  28366=>"111111110",
  28367=>"011111100",
  28368=>"100100111",
  28369=>"000111111",
  28370=>"000111111",
  28371=>"111111111",
  28372=>"000000010",
  28373=>"001111111",
  28374=>"111111110",
  28375=>"111111000",
  28376=>"110000000",
  28377=>"110110111",
  28378=>"000000000",
  28379=>"000000000",
  28380=>"010111111",
  28381=>"001000000",
  28382=>"000111111",
  28383=>"000000000",
  28384=>"000011111",
  28385=>"000010000",
  28386=>"111111111",
  28387=>"000000000",
  28388=>"111001000",
  28389=>"001000000",
  28390=>"100100111",
  28391=>"011110111",
  28392=>"000001000",
  28393=>"000000101",
  28394=>"111111110",
  28395=>"111111111",
  28396=>"111111111",
  28397=>"111000111",
  28398=>"110111111",
  28399=>"101000111",
  28400=>"010100001",
  28401=>"100000000",
  28402=>"000111111",
  28403=>"000000000",
  28404=>"111111111",
  28405=>"100000000",
  28406=>"001111001",
  28407=>"111000011",
  28408=>"000011111",
  28409=>"111000000",
  28410=>"000000000",
  28411=>"000101111",
  28412=>"011111010",
  28413=>"011111000",
  28414=>"111111001",
  28415=>"111111111",
  28416=>"000000000",
  28417=>"111011001",
  28418=>"000000000",
  28419=>"000000000",
  28420=>"000000100",
  28421=>"101000000",
  28422=>"000000000",
  28423=>"000010110",
  28424=>"110101101",
  28425=>"000111111",
  28426=>"001100110",
  28427=>"000010011",
  28428=>"000000000",
  28429=>"000000000",
  28430=>"111111111",
  28431=>"000111111",
  28432=>"110111111",
  28433=>"001111111",
  28434=>"111000000",
  28435=>"000111111",
  28436=>"001111111",
  28437=>"001000001",
  28438=>"100100111",
  28439=>"111111111",
  28440=>"111111000",
  28441=>"111100000",
  28442=>"011111010",
  28443=>"100000000",
  28444=>"011011010",
  28445=>"010000000",
  28446=>"000000000",
  28447=>"000111111",
  28448=>"101110111",
  28449=>"011000000",
  28450=>"000000110",
  28451=>"001101101",
  28452=>"111000000",
  28453=>"111111111",
  28454=>"000011111",
  28455=>"000000100",
  28456=>"110110000",
  28457=>"000000111",
  28458=>"000110111",
  28459=>"001000000",
  28460=>"000001000",
  28461=>"010111001",
  28462=>"111110000",
  28463=>"000000000",
  28464=>"010000111",
  28465=>"000001001",
  28466=>"110111111",
  28467=>"101111111",
  28468=>"000000011",
  28469=>"111000011",
  28470=>"111110000",
  28471=>"000000000",
  28472=>"110111110",
  28473=>"111101000",
  28474=>"000000000",
  28475=>"110011111",
  28476=>"111111000",
  28477=>"010000000",
  28478=>"000000000",
  28479=>"000000000",
  28480=>"000000000",
  28481=>"111111000",
  28482=>"000111001",
  28483=>"111111000",
  28484=>"111001111",
  28485=>"001001000",
  28486=>"111100000",
  28487=>"000000000",
  28488=>"000000000",
  28489=>"000111111",
  28490=>"111111111",
  28491=>"000011011",
  28492=>"001000101",
  28493=>"000000000",
  28494=>"011000111",
  28495=>"000000000",
  28496=>"001000000",
  28497=>"110010000",
  28498=>"000000000",
  28499=>"011011111",
  28500=>"010110000",
  28501=>"001001111",
  28502=>"010011000",
  28503=>"111111111",
  28504=>"011111110",
  28505=>"111100000",
  28506=>"100111111",
  28507=>"111100100",
  28508=>"000000000",
  28509=>"000000111",
  28510=>"000000000",
  28511=>"110100110",
  28512=>"000000000",
  28513=>"111111001",
  28514=>"011010000",
  28515=>"000000000",
  28516=>"111111000",
  28517=>"000000000",
  28518=>"000000000",
  28519=>"000000110",
  28520=>"100100000",
  28521=>"001111111",
  28522=>"001001000",
  28523=>"011011001",
  28524=>"110111110",
  28525=>"111111000",
  28526=>"000111010",
  28527=>"000011000",
  28528=>"110111111",
  28529=>"111010000",
  28530=>"111000000",
  28531=>"000111111",
  28532=>"111111111",
  28533=>"111111101",
  28534=>"000000000",
  28535=>"000000000",
  28536=>"111101000",
  28537=>"000000000",
  28538=>"000000000",
  28539=>"111111110",
  28540=>"000000000",
  28541=>"001000000",
  28542=>"110111000",
  28543=>"000000000",
  28544=>"001001000",
  28545=>"110110110",
  28546=>"111011000",
  28547=>"000000111",
  28548=>"100011111",
  28549=>"111000000",
  28550=>"100010000",
  28551=>"101000000",
  28552=>"000001000",
  28553=>"111111000",
  28554=>"100000100",
  28555=>"000111111",
  28556=>"111111111",
  28557=>"101100000",
  28558=>"000100000",
  28559=>"000000000",
  28560=>"000010000",
  28561=>"000000000",
  28562=>"011111111",
  28563=>"011011000",
  28564=>"000000111",
  28565=>"000000000",
  28566=>"101111111",
  28567=>"111111100",
  28568=>"110000000",
  28569=>"000111111",
  28570=>"000000000",
  28571=>"101111111",
  28572=>"001001110",
  28573=>"000111100",
  28574=>"111101000",
  28575=>"111000000",
  28576=>"111111000",
  28577=>"111101001",
  28578=>"011111100",
  28579=>"000000000",
  28580=>"111100000",
  28581=>"010000011",
  28582=>"000000001",
  28583=>"000000000",
  28584=>"000000011",
  28585=>"100000000",
  28586=>"001000000",
  28587=>"000000111",
  28588=>"000000000",
  28589=>"011111100",
  28590=>"000000000",
  28591=>"001111000",
  28592=>"011001001",
  28593=>"110010001",
  28594=>"000001111",
  28595=>"010010000",
  28596=>"110100100",
  28597=>"000111111",
  28598=>"111111101",
  28599=>"111111001",
  28600=>"000000000",
  28601=>"111111100",
  28602=>"111100000",
  28603=>"111011011",
  28604=>"111111111",
  28605=>"000000000",
  28606=>"111111000",
  28607=>"101100001",
  28608=>"101111110",
  28609=>"000001000",
  28610=>"000110111",
  28611=>"000000111",
  28612=>"000000000",
  28613=>"100110000",
  28614=>"010000000",
  28615=>"111100000",
  28616=>"111110000",
  28617=>"000010010",
  28618=>"011011111",
  28619=>"000111000",
  28620=>"000000000",
  28621=>"000100110",
  28622=>"000110110",
  28623=>"101101110",
  28624=>"000010110",
  28625=>"000010110",
  28626=>"000000101",
  28627=>"111111111",
  28628=>"000000000",
  28629=>"000101001",
  28630=>"000000010",
  28631=>"000000000",
  28632=>"111000000",
  28633=>"001011000",
  28634=>"000100111",
  28635=>"111111000",
  28636=>"100100101",
  28637=>"010111110",
  28638=>"111100001",
  28639=>"010011001",
  28640=>"000010000",
  28641=>"000000000",
  28642=>"000000000",
  28643=>"000000000",
  28644=>"111111000",
  28645=>"111111111",
  28646=>"001001111",
  28647=>"000000000",
  28648=>"010111010",
  28649=>"111111111",
  28650=>"000000000",
  28651=>"111111000",
  28652=>"100000111",
  28653=>"011011110",
  28654=>"111111011",
  28655=>"000000001",
  28656=>"000000010",
  28657=>"000110111",
  28658=>"000110100",
  28659=>"110110110",
  28660=>"010111000",
  28661=>"111011101",
  28662=>"111111000",
  28663=>"111000001",
  28664=>"000011011",
  28665=>"010111010",
  28666=>"110100000",
  28667=>"111111000",
  28668=>"000100111",
  28669=>"111101101",
  28670=>"000000000",
  28671=>"111011000",
  28672=>"000000000",
  28673=>"110110000",
  28674=>"100000000",
  28675=>"000000000",
  28676=>"000000000",
  28677=>"110110000",
  28678=>"000000000",
  28679=>"111110110",
  28680=>"000000001",
  28681=>"000000101",
  28682=>"001111111",
  28683=>"000111100",
  28684=>"000000000",
  28685=>"111111111",
  28686=>"000000010",
  28687=>"111111000",
  28688=>"000101000",
  28689=>"000110110",
  28690=>"000011001",
  28691=>"100100100",
  28692=>"111111000",
  28693=>"010000000",
  28694=>"111111000",
  28695=>"011000001",
  28696=>"011000001",
  28697=>"111111001",
  28698=>"000000100",
  28699=>"011111000",
  28700=>"111111111",
  28701=>"011000000",
  28702=>"111111110",
  28703=>"111111000",
  28704=>"001001000",
  28705=>"111111011",
  28706=>"110111110",
  28707=>"010011111",
  28708=>"000101000",
  28709=>"111111000",
  28710=>"000000000",
  28711=>"000101111",
  28712=>"000001111",
  28713=>"000000000",
  28714=>"011111111",
  28715=>"010111111",
  28716=>"110110111",
  28717=>"110010000",
  28718=>"111111110",
  28719=>"000000000",
  28720=>"111110111",
  28721=>"111000000",
  28722=>"100100100",
  28723=>"111001000",
  28724=>"111111000",
  28725=>"111011001",
  28726=>"011111111",
  28727=>"111011111",
  28728=>"111111111",
  28729=>"111001000",
  28730=>"000000000",
  28731=>"111110111",
  28732=>"100000000",
  28733=>"000000100",
  28734=>"000000011",
  28735=>"000000000",
  28736=>"000000000",
  28737=>"000000111",
  28738=>"000101111",
  28739=>"110111111",
  28740=>"000000000",
  28741=>"110110000",
  28742=>"000111001",
  28743=>"110000100",
  28744=>"110010010",
  28745=>"000000111",
  28746=>"111100100",
  28747=>"001100001",
  28748=>"111000111",
  28749=>"000000001",
  28750=>"000000110",
  28751=>"000111101",
  28752=>"111111000",
  28753=>"011000100",
  28754=>"111111111",
  28755=>"000000000",
  28756=>"000000001",
  28757=>"000000000",
  28758=>"011011101",
  28759=>"000000000",
  28760=>"000000000",
  28761=>"101111111",
  28762=>"111111000",
  28763=>"011011000",
  28764=>"001000111",
  28765=>"001000000",
  28766=>"111111000",
  28767=>"101101111",
  28768=>"000100000",
  28769=>"111111111",
  28770=>"011111111",
  28771=>"000111011",
  28772=>"001001000",
  28773=>"100000111",
  28774=>"000000111",
  28775=>"000000000",
  28776=>"000000000",
  28777=>"000000000",
  28778=>"000101101",
  28779=>"000000000",
  28780=>"000000000",
  28781=>"001000011",
  28782=>"111001001",
  28783=>"000000000",
  28784=>"000000000",
  28785=>"111111111",
  28786=>"101111111",
  28787=>"111011000",
  28788=>"111111111",
  28789=>"000110111",
  28790=>"111100111",
  28791=>"000111110",
  28792=>"000000000",
  28793=>"000000101",
  28794=>"000111001",
  28795=>"000110111",
  28796=>"111111011",
  28797=>"000000000",
  28798=>"000001111",
  28799=>"110110000",
  28800=>"111111111",
  28801=>"010110110",
  28802=>"000000011",
  28803=>"000000011",
  28804=>"000000000",
  28805=>"000000100",
  28806=>"000101000",
  28807=>"010011111",
  28808=>"111010000",
  28809=>"100000101",
  28810=>"001000000",
  28811=>"111110110",
  28812=>"011000001",
  28813=>"001010000",
  28814=>"111111111",
  28815=>"111111111",
  28816=>"110111001",
  28817=>"011010000",
  28818=>"100000000",
  28819=>"101101000",
  28820=>"000000000",
  28821=>"000000000",
  28822=>"111110111",
  28823=>"111100000",
  28824=>"000000000",
  28825=>"111111101",
  28826=>"000000000",
  28827=>"111000111",
  28828=>"000000001",
  28829=>"000000101",
  28830=>"111001001",
  28831=>"111111111",
  28832=>"000000000",
  28833=>"000000000",
  28834=>"100000000",
  28835=>"111111111",
  28836=>"001001001",
  28837=>"111100000",
  28838=>"111111010",
  28839=>"111111110",
  28840=>"000111110",
  28841=>"110111111",
  28842=>"111001111",
  28843=>"000111111",
  28844=>"111111001",
  28845=>"001001110",
  28846=>"000000111",
  28847=>"000111000",
  28848=>"110111111",
  28849=>"111100000",
  28850=>"111011011",
  28851=>"111111001",
  28852=>"111000000",
  28853=>"000000111",
  28854=>"011111101",
  28855=>"000000001",
  28856=>"111111000",
  28857=>"000000000",
  28858=>"001000000",
  28859=>"111001000",
  28860=>"000000011",
  28861=>"111111111",
  28862=>"000111111",
  28863=>"001111101",
  28864=>"111111100",
  28865=>"111111101",
  28866=>"110111111",
  28867=>"100110111",
  28868=>"101111111",
  28869=>"111111011",
  28870=>"000000111",
  28871=>"000001000",
  28872=>"111000001",
  28873=>"111001000",
  28874=>"100000001",
  28875=>"001000000",
  28876=>"000101111",
  28877=>"111110000",
  28878=>"000000001",
  28879=>"001000000",
  28880=>"111010000",
  28881=>"111000000",
  28882=>"111010000",
  28883=>"111000000",
  28884=>"111000000",
  28885=>"111111111",
  28886=>"101000000",
  28887=>"000101001",
  28888=>"000000001",
  28889=>"101101101",
  28890=>"000000111",
  28891=>"000000000",
  28892=>"111111111",
  28893=>"000000000",
  28894=>"010010000",
  28895=>"000000111",
  28896=>"000000000",
  28897=>"110111000",
  28898=>"111011000",
  28899=>"111111101",
  28900=>"000000000",
  28901=>"100100000",
  28902=>"000111011",
  28903=>"000101111",
  28904=>"111111011",
  28905=>"111111111",
  28906=>"000111111",
  28907=>"000000000",
  28908=>"111111100",
  28909=>"000000000",
  28910=>"111001001",
  28911=>"101001111",
  28912=>"111111111",
  28913=>"110100111",
  28914=>"111111111",
  28915=>"000000111",
  28916=>"000000000",
  28917=>"001000111",
  28918=>"000001011",
  28919=>"000000000",
  28920=>"000110111",
  28921=>"111110000",
  28922=>"000000011",
  28923=>"000110111",
  28924=>"111111000",
  28925=>"001000111",
  28926=>"110000110",
  28927=>"000000001",
  28928=>"111111101",
  28929=>"011001000",
  28930=>"111110100",
  28931=>"000000111",
  28932=>"111111001",
  28933=>"000101111",
  28934=>"000000000",
  28935=>"111110101",
  28936=>"110111100",
  28937=>"000000000",
  28938=>"110100000",
  28939=>"000000000",
  28940=>"111100111",
  28941=>"011011011",
  28942=>"101111111",
  28943=>"111000000",
  28944=>"000000111",
  28945=>"000000000",
  28946=>"000000111",
  28947=>"111111000",
  28948=>"001000000",
  28949=>"001001101",
  28950=>"011000100",
  28951=>"000000000",
  28952=>"111111111",
  28953=>"101101001",
  28954=>"110110111",
  28955=>"000000000",
  28956=>"011011011",
  28957=>"001000000",
  28958=>"111111111",
  28959=>"010010000",
  28960=>"000000000",
  28961=>"111111111",
  28962=>"000110111",
  28963=>"001001101",
  28964=>"000010111",
  28965=>"000000000",
  28966=>"000000000",
  28967=>"001111000",
  28968=>"111110111",
  28969=>"000000000",
  28970=>"010111111",
  28971=>"000000111",
  28972=>"000000000",
  28973=>"000000000",
  28974=>"010111111",
  28975=>"000000001",
  28976=>"000000100",
  28977=>"000000111",
  28978=>"010000000",
  28979=>"111000000",
  28980=>"000000010",
  28981=>"000000010",
  28982=>"010000010",
  28983=>"001000001",
  28984=>"000010010",
  28985=>"000000111",
  28986=>"111100000",
  28987=>"000100000",
  28988=>"110111111",
  28989=>"000001001",
  28990=>"111111111",
  28991=>"111111001",
  28992=>"111000000",
  28993=>"011000000",
  28994=>"001001000",
  28995=>"000000010",
  28996=>"011001111",
  28997=>"001111111",
  28998=>"010010010",
  28999=>"000000000",
  29000=>"111111001",
  29001=>"111100100",
  29002=>"111000000",
  29003=>"011111001",
  29004=>"000011111",
  29005=>"000000000",
  29006=>"000000001",
  29007=>"000000111",
  29008=>"100101001",
  29009=>"000001111",
  29010=>"001001000",
  29011=>"000000000",
  29012=>"011000000",
  29013=>"000010000",
  29014=>"111111111",
  29015=>"000000111",
  29016=>"000001111",
  29017=>"001000000",
  29018=>"010000000",
  29019=>"111111111",
  29020=>"000001111",
  29021=>"000000010",
  29022=>"011000111",
  29023=>"001001000",
  29024=>"110001000",
  29025=>"010110111",
  29026=>"111111011",
  29027=>"111110100",
  29028=>"001000000",
  29029=>"000011000",
  29030=>"100001111",
  29031=>"001001111",
  29032=>"110110100",
  29033=>"000000101",
  29034=>"011111110",
  29035=>"101001000",
  29036=>"010110000",
  29037=>"000001111",
  29038=>"000000111",
  29039=>"111111010",
  29040=>"111111111",
  29041=>"111001000",
  29042=>"000110111",
  29043=>"111100000",
  29044=>"000000000",
  29045=>"111111111",
  29046=>"101100111",
  29047=>"000000000",
  29048=>"111111111",
  29049=>"000001111",
  29050=>"111111111",
  29051=>"111000010",
  29052=>"100101111",
  29053=>"110111111",
  29054=>"000000000",
  29055=>"111111111",
  29056=>"000100111",
  29057=>"110111111",
  29058=>"111111000",
  29059=>"000100100",
  29060=>"000000000",
  29061=>"000000000",
  29062=>"101101111",
  29063=>"000000000",
  29064=>"110111111",
  29065=>"011011011",
  29066=>"111000000",
  29067=>"101101001",
  29068=>"111111111",
  29069=>"110110110",
  29070=>"000011111",
  29071=>"111111111",
  29072=>"011011111",
  29073=>"000000111",
  29074=>"010110010",
  29075=>"111111100",
  29076=>"000101000",
  29077=>"000000000",
  29078=>"001011111",
  29079=>"000110111",
  29080=>"101000011",
  29081=>"111000110",
  29082=>"111111111",
  29083=>"000111111",
  29084=>"000000111",
  29085=>"000000001",
  29086=>"000000001",
  29087=>"110000010",
  29088=>"001000011",
  29089=>"100100110",
  29090=>"001111111",
  29091=>"100100111",
  29092=>"111111111",
  29093=>"111111010",
  29094=>"100110111",
  29095=>"000000000",
  29096=>"111000000",
  29097=>"110000000",
  29098=>"101111111",
  29099=>"000000000",
  29100=>"000000000",
  29101=>"000000111",
  29102=>"100101111",
  29103=>"111100101",
  29104=>"100101101",
  29105=>"000110111",
  29106=>"000101111",
  29107=>"111111100",
  29108=>"110111101",
  29109=>"111111101",
  29110=>"111101111",
  29111=>"101111000",
  29112=>"000000110",
  29113=>"000000111",
  29114=>"111111110",
  29115=>"101111111",
  29116=>"101111111",
  29117=>"111111111",
  29118=>"000010000",
  29119=>"111110111",
  29120=>"000000011",
  29121=>"111111100",
  29122=>"111111111",
  29123=>"110111001",
  29124=>"110101111",
  29125=>"111001001",
  29126=>"010000000",
  29127=>"100000011",
  29128=>"001000000",
  29129=>"010111111",
  29130=>"001000111",
  29131=>"000000000",
  29132=>"011000000",
  29133=>"011111000",
  29134=>"111000010",
  29135=>"111111111",
  29136=>"101111111",
  29137=>"111100100",
  29138=>"000000000",
  29139=>"011011000",
  29140=>"000000000",
  29141=>"001000001",
  29142=>"111000000",
  29143=>"000011010",
  29144=>"101100100",
  29145=>"000000000",
  29146=>"111100000",
  29147=>"111111111",
  29148=>"111101101",
  29149=>"111101001",
  29150=>"000000111",
  29151=>"001000001",
  29152=>"001001001",
  29153=>"111010000",
  29154=>"001111111",
  29155=>"111000000",
  29156=>"111110000",
  29157=>"011111111",
  29158=>"011000000",
  29159=>"000000111",
  29160=>"001001101",
  29161=>"000000111",
  29162=>"000000000",
  29163=>"110111101",
  29164=>"100100101",
  29165=>"000101111",
  29166=>"001000000",
  29167=>"000110111",
  29168=>"111100000",
  29169=>"100111111",
  29170=>"011000000",
  29171=>"101000000",
  29172=>"000000000",
  29173=>"000001001",
  29174=>"110110111",
  29175=>"001000000",
  29176=>"000000000",
  29177=>"101100111",
  29178=>"100000101",
  29179=>"110000000",
  29180=>"000100011",
  29181=>"000000000",
  29182=>"101001000",
  29183=>"000000000",
  29184=>"000001001",
  29185=>"111111111",
  29186=>"111101111",
  29187=>"100000000",
  29188=>"111110111",
  29189=>"101000111",
  29190=>"011011010",
  29191=>"111111111",
  29192=>"000000000",
  29193=>"111011001",
  29194=>"111111111",
  29195=>"111111101",
  29196=>"100100100",
  29197=>"111111111",
  29198=>"110110010",
  29199=>"000101000",
  29200=>"111100000",
  29201=>"011000000",
  29202=>"111111111",
  29203=>"111101111",
  29204=>"000000000",
  29205=>"000000011",
  29206=>"111000000",
  29207=>"001000110",
  29208=>"100000101",
  29209=>"001000000",
  29210=>"111111111",
  29211=>"111111110",
  29212=>"100000000",
  29213=>"100101111",
  29214=>"110111000",
  29215=>"111111100",
  29216=>"110000000",
  29217=>"111111110",
  29218=>"110111110",
  29219=>"101000111",
  29220=>"111101100",
  29221=>"110110100",
  29222=>"111000000",
  29223=>"010001001",
  29224=>"101000101",
  29225=>"000000000",
  29226=>"111111111",
  29227=>"111111111",
  29228=>"000000000",
  29229=>"110000000",
  29230=>"000100100",
  29231=>"111001011",
  29232=>"111111111",
  29233=>"111111000",
  29234=>"011001000",
  29235=>"111010011",
  29236=>"110100000",
  29237=>"110111110",
  29238=>"001000000",
  29239=>"110011011",
  29240=>"111111111",
  29241=>"111111111",
  29242=>"000011111",
  29243=>"111111111",
  29244=>"100000000",
  29245=>"111010011",
  29246=>"111111111",
  29247=>"111000000",
  29248=>"000010001",
  29249=>"111001000",
  29250=>"101111111",
  29251=>"111010001",
  29252=>"110111111",
  29253=>"011000000",
  29254=>"000000000",
  29255=>"111111111",
  29256=>"111111011",
  29257=>"111111111",
  29258=>"110111111",
  29259=>"111011001",
  29260=>"000000001",
  29261=>"001101111",
  29262=>"111000110",
  29263=>"010110110",
  29264=>"010000111",
  29265=>"111101111",
  29266=>"111111000",
  29267=>"000000000",
  29268=>"000101001",
  29269=>"111111001",
  29270=>"000000010",
  29271=>"100101000",
  29272=>"000000000",
  29273=>"111001101",
  29274=>"111001000",
  29275=>"110110000",
  29276=>"110110110",
  29277=>"101000000",
  29278=>"100111111",
  29279=>"111011000",
  29280=>"100111111",
  29281=>"010010000",
  29282=>"000000000",
  29283=>"000000000",
  29284=>"110110010",
  29285=>"001001111",
  29286=>"111101111",
  29287=>"000000000",
  29288=>"011011010",
  29289=>"000001010",
  29290=>"011101111",
  29291=>"111111111",
  29292=>"111000001",
  29293=>"000110000",
  29294=>"001101101",
  29295=>"001001000",
  29296=>"000000000",
  29297=>"110010001",
  29298=>"110100000",
  29299=>"011111111",
  29300=>"000111111",
  29301=>"111111100",
  29302=>"111011111",
  29303=>"111111111",
  29304=>"000000010",
  29305=>"111110110",
  29306=>"000000000",
  29307=>"001111111",
  29308=>"000000000",
  29309=>"111111111",
  29310=>"000000000",
  29311=>"011011001",
  29312=>"011000000",
  29313=>"001000111",
  29314=>"011000100",
  29315=>"000000001",
  29316=>"110000000",
  29317=>"000000101",
  29318=>"000000110",
  29319=>"000000000",
  29320=>"011001000",
  29321=>"011001000",
  29322=>"110110110",
  29323=>"111011011",
  29324=>"000000100",
  29325=>"100000000",
  29326=>"111111101",
  29327=>"000000111",
  29328=>"111001000",
  29329=>"000000011",
  29330=>"000000000",
  29331=>"111111111",
  29332=>"110111111",
  29333=>"001000100",
  29334=>"011011001",
  29335=>"000000100",
  29336=>"111101111",
  29337=>"111111111",
  29338=>"000000000",
  29339=>"001111001",
  29340=>"111111111",
  29341=>"101111111",
  29342=>"110110111",
  29343=>"111111111",
  29344=>"011010111",
  29345=>"110111111",
  29346=>"111111111",
  29347=>"010010100",
  29348=>"001000000",
  29349=>"111110100",
  29350=>"111111010",
  29351=>"111110000",
  29352=>"000000000",
  29353=>"011001000",
  29354=>"000000000",
  29355=>"000001001",
  29356=>"111111111",
  29357=>"000001111",
  29358=>"111111111",
  29359=>"011111101",
  29360=>"111111111",
  29361=>"000000000",
  29362=>"011111010",
  29363=>"111111101",
  29364=>"111110110",
  29365=>"000000001",
  29366=>"001001001",
  29367=>"111111111",
  29368=>"111000000",
  29369=>"111111111",
  29370=>"111000000",
  29371=>"100000000",
  29372=>"001001111",
  29373=>"000000000",
  29374=>"000001111",
  29375=>"000000000",
  29376=>"000000001",
  29377=>"111111010",
  29378=>"000000000",
  29379=>"111111001",
  29380=>"111111000",
  29381=>"000000011",
  29382=>"111011001",
  29383=>"110011001",
  29384=>"001001000",
  29385=>"100100111",
  29386=>"010111100",
  29387=>"000000110",
  29388=>"111111111",
  29389=>"111111111",
  29390=>"111111110",
  29391=>"011000000",
  29392=>"011001011",
  29393=>"011000000",
  29394=>"111000100",
  29395=>"010000010",
  29396=>"001000000",
  29397=>"100100110",
  29398=>"000000001",
  29399=>"011101111",
  29400=>"111101110",
  29401=>"111110110",
  29402=>"001001000",
  29403=>"010010000",
  29404=>"000000000",
  29405=>"001000000",
  29406=>"000000110",
  29407=>"111111111",
  29408=>"001000000",
  29409=>"000001011",
  29410=>"000000000",
  29411=>"111110000",
  29412=>"000000000",
  29413=>"001101101",
  29414=>"010000000",
  29415=>"110010010",
  29416=>"101101111",
  29417=>"000000000",
  29418=>"111111111",
  29419=>"111010010",
  29420=>"000011010",
  29421=>"000000000",
  29422=>"111000001",
  29423=>"010000100",
  29424=>"011011011",
  29425=>"111110111",
  29426=>"011000000",
  29427=>"110000001",
  29428=>"011001110",
  29429=>"111110000",
  29430=>"000000100",
  29431=>"101111111",
  29432=>"000000000",
  29433=>"011111111",
  29434=>"001000000",
  29435=>"111001111",
  29436=>"100100111",
  29437=>"111111111",
  29438=>"011110110",
  29439=>"110110000",
  29440=>"111111110",
  29441=>"111111000",
  29442=>"111111000",
  29443=>"111101100",
  29444=>"000000000",
  29445=>"001000000",
  29446=>"101101111",
  29447=>"110010011",
  29448=>"111111111",
  29449=>"111111111",
  29450=>"000000001",
  29451=>"000000000",
  29452=>"000000101",
  29453=>"100100000",
  29454=>"111111111",
  29455=>"000100000",
  29456=>"000000000",
  29457=>"001110111",
  29458=>"000000000",
  29459=>"111011111",
  29460=>"111101111",
  29461=>"010110111",
  29462=>"100000000",
  29463=>"111111111",
  29464=>"011011010",
  29465=>"000000000",
  29466=>"111111111",
  29467=>"110110110",
  29468=>"110100000",
  29469=>"000000010",
  29470=>"011111000",
  29471=>"000111110",
  29472=>"010111111",
  29473=>"111110000",
  29474=>"111111010",
  29475=>"011000000",
  29476=>"001101101",
  29477=>"000100111",
  29478=>"000000000",
  29479=>"110110111",
  29480=>"111100100",
  29481=>"111111111",
  29482=>"000110110",
  29483=>"000000000",
  29484=>"000000111",
  29485=>"001011101",
  29486=>"111101111",
  29487=>"111111111",
  29488=>"000000000",
  29489=>"000011110",
  29490=>"010011111",
  29491=>"000000000",
  29492=>"011001000",
  29493=>"111110111",
  29494=>"110110110",
  29495=>"000001001",
  29496=>"111111000",
  29497=>"001101111",
  29498=>"001000001",
  29499=>"011010010",
  29500=>"110000000",
  29501=>"101101111",
  29502=>"100100100",
  29503=>"100010111",
  29504=>"100000100",
  29505=>"111111111",
  29506=>"000000001",
  29507=>"000000000",
  29508=>"000000000",
  29509=>"111100110",
  29510=>"011001011",
  29511=>"000000100",
  29512=>"111111111",
  29513=>"000001111",
  29514=>"000000000",
  29515=>"000000100",
  29516=>"000000001",
  29517=>"000000000",
  29518=>"111110110",
  29519=>"000000000",
  29520=>"011001000",
  29521=>"110000000",
  29522=>"000000001",
  29523=>"000000000",
  29524=>"111111000",
  29525=>"000000001",
  29526=>"111111111",
  29527=>"000000000",
  29528=>"111111111",
  29529=>"000001000",
  29530=>"110100100",
  29531=>"011000101",
  29532=>"011001001",
  29533=>"010110110",
  29534=>"111100000",
  29535=>"111000000",
  29536=>"111011111",
  29537=>"111011000",
  29538=>"100100100",
  29539=>"000000111",
  29540=>"000000000",
  29541=>"111111111",
  29542=>"000111111",
  29543=>"100100001",
  29544=>"001100100",
  29545=>"011000000",
  29546=>"000000000",
  29547=>"111100100",
  29548=>"111001000",
  29549=>"111000000",
  29550=>"111111111",
  29551=>"100000000",
  29552=>"100000000",
  29553=>"111111110",
  29554=>"000010111",
  29555=>"010111000",
  29556=>"111010000",
  29557=>"110110110",
  29558=>"111001001",
  29559=>"001001100",
  29560=>"100000000",
  29561=>"000000000",
  29562=>"111111111",
  29563=>"110100100",
  29564=>"111101001",
  29565=>"111111111",
  29566=>"000000010",
  29567=>"000101000",
  29568=>"000000100",
  29569=>"110010001",
  29570=>"011011000",
  29571=>"000000011",
  29572=>"001000111",
  29573=>"111111111",
  29574=>"001001111",
  29575=>"101100100",
  29576=>"110111111",
  29577=>"111111111",
  29578=>"010110111",
  29579=>"000000000",
  29580=>"000000101",
  29581=>"111010011",
  29582=>"000000000",
  29583=>"001001011",
  29584=>"000100111",
  29585=>"111111111",
  29586=>"111010110",
  29587=>"011011000",
  29588=>"111111111",
  29589=>"000000000",
  29590=>"111000011",
  29591=>"001001100",
  29592=>"011111111",
  29593=>"111111111",
  29594=>"000000000",
  29595=>"000000101",
  29596=>"000000000",
  29597=>"100000000",
  29598=>"100000000",
  29599=>"011111111",
  29600=>"001001000",
  29601=>"001000001",
  29602=>"111111011",
  29603=>"001001000",
  29604=>"101100101",
  29605=>"111110010",
  29606=>"001001001",
  29607=>"111010000",
  29608=>"101101101",
  29609=>"110000111",
  29610=>"111111000",
  29611=>"110111111",
  29612=>"110000000",
  29613=>"000001000",
  29614=>"010111111",
  29615=>"000000000",
  29616=>"011001111",
  29617=>"010110000",
  29618=>"111111101",
  29619=>"001111111",
  29620=>"110010000",
  29621=>"000010111",
  29622=>"111111111",
  29623=>"000000011",
  29624=>"000000000",
  29625=>"000000000",
  29626=>"111101000",
  29627=>"111111111",
  29628=>"000000000",
  29629=>"000000111",
  29630=>"000000010",
  29631=>"110110100",
  29632=>"111111011",
  29633=>"111000000",
  29634=>"000110000",
  29635=>"111111100",
  29636=>"000111111",
  29637=>"111011111",
  29638=>"111011011",
  29639=>"111001001",
  29640=>"001000000",
  29641=>"000000000",
  29642=>"011011100",
  29643=>"111101010",
  29644=>"111111111",
  29645=>"111111111",
  29646=>"000000000",
  29647=>"111000000",
  29648=>"110110110",
  29649=>"111111111",
  29650=>"110110000",
  29651=>"011001001",
  29652=>"000000000",
  29653=>"110100000",
  29654=>"111111111",
  29655=>"011011011",
  29656=>"000000000",
  29657=>"000110110",
  29658=>"111110000",
  29659=>"001011111",
  29660=>"001000000",
  29661=>"000100111",
  29662=>"000011111",
  29663=>"111111011",
  29664=>"011010000",
  29665=>"111111011",
  29666=>"011111111",
  29667=>"111111111",
  29668=>"111000001",
  29669=>"111111111",
  29670=>"110111111",
  29671=>"011000000",
  29672=>"111111111",
  29673=>"100010111",
  29674=>"000110010",
  29675=>"000000100",
  29676=>"111111111",
  29677=>"011010110",
  29678=>"110111111",
  29679=>"001000000",
  29680=>"000011010",
  29681=>"011111111",
  29682=>"000011111",
  29683=>"111111111",
  29684=>"001001011",
  29685=>"000000000",
  29686=>"111111110",
  29687=>"110000100",
  29688=>"001000001",
  29689=>"001001001",
  29690=>"111111110",
  29691=>"000000111",
  29692=>"111111111",
  29693=>"100110111",
  29694=>"111100100",
  29695=>"000001001",
  29696=>"000000000",
  29697=>"111111000",
  29698=>"000000000",
  29699=>"111111000",
  29700=>"100110111",
  29701=>"000111011",
  29702=>"111011011",
  29703=>"111111111",
  29704=>"111111000",
  29705=>"100111010",
  29706=>"111000100",
  29707=>"001000110",
  29708=>"000000000",
  29709=>"111111000",
  29710=>"111000000",
  29711=>"000000000",
  29712=>"000000011",
  29713=>"111111110",
  29714=>"000000100",
  29715=>"011000100",
  29716=>"111110111",
  29717=>"000000000",
  29718=>"000000000",
  29719=>"101001001",
  29720=>"111100000",
  29721=>"001001001",
  29722=>"111001101",
  29723=>"001011011",
  29724=>"000000000",
  29725=>"110100111",
  29726=>"111111011",
  29727=>"000000111",
  29728=>"001000000",
  29729=>"110110101",
  29730=>"011001001",
  29731=>"111110110",
  29732=>"110110111",
  29733=>"111111111",
  29734=>"000000000",
  29735=>"111011111",
  29736=>"111111111",
  29737=>"000111111",
  29738=>"111111111",
  29739=>"000000000",
  29740=>"001111001",
  29741=>"011111111",
  29742=>"000000101",
  29743=>"001101111",
  29744=>"000000111",
  29745=>"011111111",
  29746=>"001100111",
  29747=>"100000000",
  29748=>"000000000",
  29749=>"000000111",
  29750=>"011000011",
  29751=>"110111111",
  29752=>"111111111",
  29753=>"111111101",
  29754=>"001000000",
  29755=>"000100000",
  29756=>"011011000",
  29757=>"000000000",
  29758=>"110110110",
  29759=>"001000000",
  29760=>"111000000",
  29761=>"000110110",
  29762=>"111111010",
  29763=>"011111010",
  29764=>"111111000",
  29765=>"101001001",
  29766=>"111110000",
  29767=>"111110110",
  29768=>"111111111",
  29769=>"100110110",
  29770=>"111011011",
  29771=>"111111111",
  29772=>"000100100",
  29773=>"001001000",
  29774=>"000000000",
  29775=>"111111111",
  29776=>"111000000",
  29777=>"000000111",
  29778=>"111101111",
  29779=>"000001111",
  29780=>"001001111",
  29781=>"111111110",
  29782=>"101100111",
  29783=>"000001011",
  29784=>"000110111",
  29785=>"000000000",
  29786=>"111111000",
  29787=>"110110110",
  29788=>"110100000",
  29789=>"000000000",
  29790=>"111111111",
  29791=>"011111101",
  29792=>"000111111",
  29793=>"000001111",
  29794=>"110110100",
  29795=>"000011011",
  29796=>"001111111",
  29797=>"001011000",
  29798=>"110111111",
  29799=>"101011011",
  29800=>"000000000",
  29801=>"100000100",
  29802=>"111111000",
  29803=>"111111000",
  29804=>"011011011",
  29805=>"100110111",
  29806=>"000110000",
  29807=>"111111111",
  29808=>"000011100",
  29809=>"000100111",
  29810=>"001000000",
  29811=>"110001001",
  29812=>"111111111",
  29813=>"000000000",
  29814=>"000000000",
  29815=>"111111001",
  29816=>"010011111",
  29817=>"110111111",
  29818=>"011011111",
  29819=>"000000010",
  29820=>"000011001",
  29821=>"001000111",
  29822=>"111111001",
  29823=>"001011111",
  29824=>"100110100",
  29825=>"000000001",
  29826=>"111100100",
  29827=>"000111111",
  29828=>"111000000",
  29829=>"000000000",
  29830=>"111100000",
  29831=>"000111010",
  29832=>"000000000",
  29833=>"000100110",
  29834=>"111111100",
  29835=>"000000000",
  29836=>"000000000",
  29837=>"111101100",
  29838=>"011111111",
  29839=>"111000000",
  29840=>"111111111",
  29841=>"111111111",
  29842=>"001000001",
  29843=>"000000000",
  29844=>"111111111",
  29845=>"001000110",
  29846=>"111111111",
  29847=>"111111000",
  29848=>"110100001",
  29849=>"000000000",
  29850=>"000000000",
  29851=>"000000000",
  29852=>"111000000",
  29853=>"111000000",
  29854=>"011011011",
  29855=>"000000000",
  29856=>"111111011",
  29857=>"111111010",
  29858=>"111001000",
  29859=>"111111111",
  29860=>"110110111",
  29861=>"111100110",
  29862=>"111111111",
  29863=>"000001110",
  29864=>"111101111",
  29865=>"000000000",
  29866=>"000111111",
  29867=>"000111111",
  29868=>"111111001",
  29869=>"000000000",
  29870=>"001001111",
  29871=>"000000000",
  29872=>"000111011",
  29873=>"000000111",
  29874=>"100111000",
  29875=>"000000000",
  29876=>"000000000",
  29877=>"000000101",
  29878=>"111000001",
  29879=>"111111111",
  29880=>"111111000",
  29881=>"000100001",
  29882=>"001000000",
  29883=>"000000000",
  29884=>"000100100",
  29885=>"000000000",
  29886=>"110111111",
  29887=>"110000000",
  29888=>"000000000",
  29889=>"110100100",
  29890=>"011000000",
  29891=>"000000000",
  29892=>"111111000",
  29893=>"111111111",
  29894=>"010010010",
  29895=>"001001111",
  29896=>"000001011",
  29897=>"000111111",
  29898=>"000011011",
  29899=>"000000000",
  29900=>"011011000",
  29901=>"110111011",
  29902=>"111111111",
  29903=>"101000000",
  29904=>"000000111",
  29905=>"000000000",
  29906=>"110110110",
  29907=>"000000011",
  29908=>"001101000",
  29909=>"111000000",
  29910=>"000000111",
  29911=>"000001000",
  29912=>"000000001",
  29913=>"110110000",
  29914=>"010000000",
  29915=>"001111100",
  29916=>"110111111",
  29917=>"000000000",
  29918=>"000010010",
  29919=>"001001000",
  29920=>"000111110",
  29921=>"000111100",
  29922=>"111011000",
  29923=>"111000000",
  29924=>"111011110",
  29925=>"111111111",
  29926=>"111000000",
  29927=>"111111111",
  29928=>"110110000",
  29929=>"111111111",
  29930=>"111110000",
  29931=>"000001111",
  29932=>"000110000",
  29933=>"111000110",
  29934=>"111000110",
  29935=>"000000000",
  29936=>"101111111",
  29937=>"111001011",
  29938=>"111011000",
  29939=>"001000111",
  29940=>"000111111",
  29941=>"010000000",
  29942=>"000000000",
  29943=>"000000111",
  29944=>"000000000",
  29945=>"000000000",
  29946=>"000000001",
  29947=>"111111100",
  29948=>"110110111",
  29949=>"100000011",
  29950=>"111111001",
  29951=>"111111111",
  29952=>"000000000",
  29953=>"000001011",
  29954=>"001000111",
  29955=>"111111111",
  29956=>"110111111",
  29957=>"111111110",
  29958=>"111111111",
  29959=>"001000000",
  29960=>"000101111",
  29961=>"111111111",
  29962=>"010000000",
  29963=>"000000001",
  29964=>"000000000",
  29965=>"000000100",
  29966=>"111111111",
  29967=>"011111111",
  29968=>"000111011",
  29969=>"101000000",
  29970=>"000000000",
  29971=>"000000000",
  29972=>"111111000",
  29973=>"111000000",
  29974=>"000000000",
  29975=>"001000001",
  29976=>"001111001",
  29977=>"111111111",
  29978=>"000000001",
  29979=>"100100100",
  29980=>"110100101",
  29981=>"100000000",
  29982=>"111000000",
  29983=>"111111100",
  29984=>"100111111",
  29985=>"111111111",
  29986=>"000100111",
  29987=>"000001001",
  29988=>"110010001",
  29989=>"011011011",
  29990=>"000000000",
  29991=>"111111111",
  29992=>"011111000",
  29993=>"000000000",
  29994=>"001011111",
  29995=>"101100111",
  29996=>"111111111",
  29997=>"000100110",
  29998=>"000100000",
  29999=>"000001001",
  30000=>"100100100",
  30001=>"001001111",
  30002=>"000000000",
  30003=>"111100100",
  30004=>"000000000",
  30005=>"000000000",
  30006=>"111001011",
  30007=>"111111111",
  30008=>"000000111",
  30009=>"111100111",
  30010=>"000001101",
  30011=>"111111110",
  30012=>"111111111",
  30013=>"111111000",
  30014=>"111111111",
  30015=>"011001001",
  30016=>"111000000",
  30017=>"011000101",
  30018=>"001001111",
  30019=>"000000001",
  30020=>"000000000",
  30021=>"000110110",
  30022=>"111111000",
  30023=>"111000000",
  30024=>"000000111",
  30025=>"100110110",
  30026=>"001001000",
  30027=>"000000001",
  30028=>"011110010",
  30029=>"000000000",
  30030=>"111111111",
  30031=>"110111111",
  30032=>"001001011",
  30033=>"100110111",
  30034=>"001000000",
  30035=>"111111111",
  30036=>"111111111",
  30037=>"001111111",
  30038=>"001110111",
  30039=>"110110011",
  30040=>"011111111",
  30041=>"000000000",
  30042=>"001011001",
  30043=>"110110110",
  30044=>"000000000",
  30045=>"111111100",
  30046=>"111111111",
  30047=>"111111110",
  30048=>"111100100",
  30049=>"111110000",
  30050=>"000000100",
  30051=>"000111111",
  30052=>"000000000",
  30053=>"001101111",
  30054=>"111101111",
  30055=>"011000111",
  30056=>"000001001",
  30057=>"000000010",
  30058=>"001000000",
  30059=>"000011011",
  30060=>"100110111",
  30061=>"001000000",
  30062=>"000000111",
  30063=>"111111111",
  30064=>"000011111",
  30065=>"110000000",
  30066=>"000000000",
  30067=>"001101000",
  30068=>"000000000",
  30069=>"111111111",
  30070=>"111100011",
  30071=>"111101101",
  30072=>"000000000",
  30073=>"111101000",
  30074=>"000000011",
  30075=>"111111111",
  30076=>"111111111",
  30077=>"010000000",
  30078=>"001000100",
  30079=>"110110100",
  30080=>"000000010",
  30081=>"001011010",
  30082=>"110111101",
  30083=>"110111111",
  30084=>"000000111",
  30085=>"000000111",
  30086=>"010111001",
  30087=>"000000000",
  30088=>"000000000",
  30089=>"111111111",
  30090=>"000100011",
  30091=>"111111111",
  30092=>"111111111",
  30093=>"000010000",
  30094=>"000000011",
  30095=>"111111111",
  30096=>"110110100",
  30097=>"111111111",
  30098=>"011010000",
  30099=>"111111111",
  30100=>"000000111",
  30101=>"000010000",
  30102=>"010111111",
  30103=>"000001001",
  30104=>"000000100",
  30105=>"100110001",
  30106=>"001000100",
  30107=>"000000111",
  30108=>"111111111",
  30109=>"111111111",
  30110=>"101101111",
  30111=>"000000000",
  30112=>"100000000",
  30113=>"001000000",
  30114=>"001000110",
  30115=>"111111111",
  30116=>"000000000",
  30117=>"000100100",
  30118=>"100111101",
  30119=>"000000000",
  30120=>"111111100",
  30121=>"000000101",
  30122=>"001000000",
  30123=>"001000000",
  30124=>"110010111",
  30125=>"111101111",
  30126=>"011000001",
  30127=>"111100000",
  30128=>"111000000",
  30129=>"000010000",
  30130=>"111000000",
  30131=>"111001000",
  30132=>"111101011",
  30133=>"001000111",
  30134=>"110111000",
  30135=>"111101111",
  30136=>"111111111",
  30137=>"111011111",
  30138=>"000000001",
  30139=>"100100111",
  30140=>"001001011",
  30141=>"011100110",
  30142=>"000000000",
  30143=>"000000000",
  30144=>"100100000",
  30145=>"000011011",
  30146=>"111111111",
  30147=>"111111011",
  30148=>"001100111",
  30149=>"001111111",
  30150=>"001000001",
  30151=>"100111111",
  30152=>"011100111",
  30153=>"111111100",
  30154=>"000000101",
  30155=>"000010111",
  30156=>"000100000",
  30157=>"111111000",
  30158=>"000000000",
  30159=>"111111111",
  30160=>"111000111",
  30161=>"000000011",
  30162=>"100100111",
  30163=>"011111111",
  30164=>"110010000",
  30165=>"011010000",
  30166=>"100000000",
  30167=>"001000011",
  30168=>"111111111",
  30169=>"011011111",
  30170=>"000111111",
  30171=>"111011111",
  30172=>"001011011",
  30173=>"001001000",
  30174=>"001011000",
  30175=>"000000000",
  30176=>"000000000",
  30177=>"000000111",
  30178=>"010001011",
  30179=>"111111111",
  30180=>"001000111",
  30181=>"111111111",
  30182=>"000111111",
  30183=>"100100110",
  30184=>"010000000",
  30185=>"111001001",
  30186=>"000000001",
  30187=>"111000000",
  30188=>"111100000",
  30189=>"001000100",
  30190=>"000000111",
  30191=>"011000000",
  30192=>"111111111",
  30193=>"010011111",
  30194=>"101011011",
  30195=>"111011111",
  30196=>"111110111",
  30197=>"000000111",
  30198=>"111011000",
  30199=>"010110110",
  30200=>"000000000",
  30201=>"001101001",
  30202=>"111111111",
  30203=>"000000000",
  30204=>"111011010",
  30205=>"011011111",
  30206=>"000001000",
  30207=>"000000000",
  30208=>"111111100",
  30209=>"111000000",
  30210=>"111000000",
  30211=>"100000000",
  30212=>"000000000",
  30213=>"111111100",
  30214=>"011000000",
  30215=>"111111111",
  30216=>"000000000",
  30217=>"000000111",
  30218=>"111001000",
  30219=>"111011111",
  30220=>"111000100",
  30221=>"111111111",
  30222=>"111000000",
  30223=>"000111111",
  30224=>"000101111",
  30225=>"000000111",
  30226=>"111111111",
  30227=>"000111111",
  30228=>"111110000",
  30229=>"111111111",
  30230=>"000000000",
  30231=>"011111111",
  30232=>"111111110",
  30233=>"111111111",
  30234=>"000000111",
  30235=>"000000000",
  30236=>"000001001",
  30237=>"111111010",
  30238=>"001001100",
  30239=>"000000111",
  30240=>"000100000",
  30241=>"111100111",
  30242=>"000110111",
  30243=>"000001001",
  30244=>"000000000",
  30245=>"111000000",
  30246=>"000000000",
  30247=>"111000000",
  30248=>"100111011",
  30249=>"111110100",
  30250=>"111111011",
  30251=>"000000111",
  30252=>"000101111",
  30253=>"111111000",
  30254=>"000100000",
  30255=>"111111111",
  30256=>"001111011",
  30257=>"100111111",
  30258=>"000000000",
  30259=>"111000111",
  30260=>"000000101",
  30261=>"110111011",
  30262=>"000000000",
  30263=>"111110111",
  30264=>"001111111",
  30265=>"000000110",
  30266=>"000000001",
  30267=>"011111000",
  30268=>"110000000",
  30269=>"011111011",
  30270=>"111110111",
  30271=>"011011001",
  30272=>"011111110",
  30273=>"100100101",
  30274=>"000000001",
  30275=>"111111111",
  30276=>"111111111",
  30277=>"011011111",
  30278=>"111000000",
  30279=>"111111111",
  30280=>"011111100",
  30281=>"000000000",
  30282=>"111111000",
  30283=>"011110111",
  30284=>"110111111",
  30285=>"111111000",
  30286=>"111010110",
  30287=>"000110110",
  30288=>"110110000",
  30289=>"100111111",
  30290=>"111111000",
  30291=>"100000001",
  30292=>"111111111",
  30293=>"111111111",
  30294=>"111100111",
  30295=>"000000100",
  30296=>"001000001",
  30297=>"101000111",
  30298=>"111000000",
  30299=>"000100111",
  30300=>"111000100",
  30301=>"000000111",
  30302=>"111111000",
  30303=>"000110000",
  30304=>"111101001",
  30305=>"111111111",
  30306=>"111000000",
  30307=>"000000000",
  30308=>"001000000",
  30309=>"001111111",
  30310=>"000110110",
  30311=>"000000110",
  30312=>"111100111",
  30313=>"111000000",
  30314=>"110111110",
  30315=>"000000110",
  30316=>"111111000",
  30317=>"111111111",
  30318=>"100111110",
  30319=>"000000000",
  30320=>"111110111",
  30321=>"100111001",
  30322=>"000000100",
  30323=>"000000000",
  30324=>"000001000",
  30325=>"111111000",
  30326=>"111111000",
  30327=>"001111111",
  30328=>"111000011",
  30329=>"011111001",
  30330=>"111100000",
  30331=>"000111111",
  30332=>"110110110",
  30333=>"111000000",
  30334=>"111011001",
  30335=>"000000110",
  30336=>"000100000",
  30337=>"000111101",
  30338=>"000100111",
  30339=>"000000000",
  30340=>"000110111",
  30341=>"000000100",
  30342=>"111001000",
  30343=>"111111000",
  30344=>"001000100",
  30345=>"001111111",
  30346=>"000000111",
  30347=>"000011001",
  30348=>"110111111",
  30349=>"000000000",
  30350=>"111111000",
  30351=>"111111001",
  30352=>"000000011",
  30353=>"000000101",
  30354=>"000101111",
  30355=>"111000100",
  30356=>"000000100",
  30357=>"011000000",
  30358=>"111111111",
  30359=>"000000111",
  30360=>"010000000",
  30361=>"000100111",
  30362=>"000000111",
  30363=>"000000000",
  30364=>"110111111",
  30365=>"000000110",
  30366=>"111111111",
  30367=>"000000000",
  30368=>"011000000",
  30369=>"111100100",
  30370=>"101000000",
  30371=>"111000000",
  30372=>"011000000",
  30373=>"111111111",
  30374=>"000000000",
  30375=>"010110110",
  30376=>"001000000",
  30377=>"000000111",
  30378=>"000000100",
  30379=>"110010000",
  30380=>"010011011",
  30381=>"001011011",
  30382=>"111111000",
  30383=>"111111100",
  30384=>"111111000",
  30385=>"011000000",
  30386=>"011111010",
  30387=>"000000000",
  30388=>"010110110",
  30389=>"110000000",
  30390=>"000000010",
  30391=>"000010010",
  30392=>"000000001",
  30393=>"000000000",
  30394=>"000000000",
  30395=>"010111011",
  30396=>"111000000",
  30397=>"110110000",
  30398=>"101100111",
  30399=>"000000100",
  30400=>"000000000",
  30401=>"111000000",
  30402=>"111111111",
  30403=>"000000000",
  30404=>"001000000",
  30405=>"111011000",
  30406=>"100000000",
  30407=>"111111111",
  30408=>"010010111",
  30409=>"000111100",
  30410=>"000000000",
  30411=>"000100111",
  30412=>"111100000",
  30413=>"011000000",
  30414=>"111000001",
  30415=>"111000111",
  30416=>"000000000",
  30417=>"000111111",
  30418=>"000000001",
  30419=>"000000000",
  30420=>"111101000",
  30421=>"111111111",
  30422=>"111111101",
  30423=>"100001100",
  30424=>"111111011",
  30425=>"111110111",
  30426=>"000001111",
  30427=>"000001000",
  30428=>"111000000",
  30429=>"000000111",
  30430=>"111011010",
  30431=>"000100100",
  30432=>"100000000",
  30433=>"111111111",
  30434=>"000000111",
  30435=>"000000000",
  30436=>"111111111",
  30437=>"100100111",
  30438=>"000010000",
  30439=>"111001000",
  30440=>"110111111",
  30441=>"001100001",
  30442=>"111010000",
  30443=>"111000101",
  30444=>"000100100",
  30445=>"111110000",
  30446=>"000110110",
  30447=>"111111001",
  30448=>"111000000",
  30449=>"011000000",
  30450=>"111000000",
  30451=>"000100000",
  30452=>"000110111",
  30453=>"000100100",
  30454=>"010000011",
  30455=>"000000000",
  30456=>"111111101",
  30457=>"000000111",
  30458=>"111111011",
  30459=>"011011000",
  30460=>"000000010",
  30461=>"000010010",
  30462=>"010011011",
  30463=>"111111111",
  30464=>"111111000",
  30465=>"011000000",
  30466=>"110111111",
  30467=>"111110000",
  30468=>"000110111",
  30469=>"111110000",
  30470=>"100000101",
  30471=>"000000111",
  30472=>"000000000",
  30473=>"100000000",
  30474=>"000111111",
  30475=>"111111111",
  30476=>"000000001",
  30477=>"111111110",
  30478=>"111111001",
  30479=>"111111000",
  30480=>"000000100",
  30481=>"000000000",
  30482=>"011001000",
  30483=>"000000000",
  30484=>"000110110",
  30485=>"000000000",
  30486=>"110000000",
  30487=>"100101111",
  30488=>"000000000",
  30489=>"110000100",
  30490=>"000000110",
  30491=>"011111111",
  30492=>"001111001",
  30493=>"111111111",
  30494=>"000000111",
  30495=>"111010000",
  30496=>"000010000",
  30497=>"000000100",
  30498=>"000000111",
  30499=>"111010000",
  30500=>"111111110",
  30501=>"111101111",
  30502=>"001011111",
  30503=>"001111100",
  30504=>"000000011",
  30505=>"000000000",
  30506=>"111111111",
  30507=>"000000010",
  30508=>"000111001",
  30509=>"000000100",
  30510=>"000010111",
  30511=>"000000000",
  30512=>"110110110",
  30513=>"111111000",
  30514=>"110111010",
  30515=>"111111111",
  30516=>"111000000",
  30517=>"111100100",
  30518=>"000110111",
  30519=>"000101000",
  30520=>"101111111",
  30521=>"000000000",
  30522=>"000000000",
  30523=>"111000100",
  30524=>"110000110",
  30525=>"000000001",
  30526=>"000111111",
  30527=>"000000000",
  30528=>"000101000",
  30529=>"110111111",
  30530=>"000011001",
  30531=>"000000111",
  30532=>"000111000",
  30533=>"001111111",
  30534=>"100100000",
  30535=>"111000010",
  30536=>"000111011",
  30537=>"000000000",
  30538=>"000000000",
  30539=>"100100111",
  30540=>"000000111",
  30541=>"000000011",
  30542=>"010111111",
  30543=>"110000100",
  30544=>"001001011",
  30545=>"000100101",
  30546=>"100110101",
  30547=>"000100111",
  30548=>"000000011",
  30549=>"111010000",
  30550=>"000001001",
  30551=>"000101111",
  30552=>"111100111",
  30553=>"000000000",
  30554=>"000001011",
  30555=>"000000011",
  30556=>"111000000",
  30557=>"001011000",
  30558=>"111101111",
  30559=>"000000000",
  30560=>"111111000",
  30561=>"010000111",
  30562=>"000110011",
  30563=>"000000000",
  30564=>"100100011",
  30565=>"000000110",
  30566=>"100000001",
  30567=>"000000000",
  30568=>"111010010",
  30569=>"111111111",
  30570=>"000111111",
  30571=>"000001111",
  30572=>"000000000",
  30573=>"000000000",
  30574=>"000000000",
  30575=>"000000000",
  30576=>"011000111",
  30577=>"010111011",
  30578=>"000000100",
  30579=>"111111111",
  30580=>"000000000",
  30581=>"000111111",
  30582=>"000000000",
  30583=>"000000000",
  30584=>"111110111",
  30585=>"111111000",
  30586=>"011000000",
  30587=>"111000000",
  30588=>"000000111",
  30589=>"001100000",
  30590=>"000000101",
  30591=>"111000111",
  30592=>"000000010",
  30593=>"111000000",
  30594=>"100000001",
  30595=>"000000000",
  30596=>"001101000",
  30597=>"000111000",
  30598=>"010110011",
  30599=>"111000100",
  30600=>"101111111",
  30601=>"101111111",
  30602=>"111111111",
  30603=>"000100000",
  30604=>"011001001",
  30605=>"111111000",
  30606=>"010011000",
  30607=>"000000000",
  30608=>"000000111",
  30609=>"000000000",
  30610=>"000000111",
  30611=>"001000001",
  30612=>"000111111",
  30613=>"010010011",
  30614=>"000000001",
  30615=>"110110000",
  30616=>"011010000",
  30617=>"000001011",
  30618=>"111100001",
  30619=>"000001111",
  30620=>"111100100",
  30621=>"111111000",
  30622=>"000110111",
  30623=>"000000000",
  30624=>"111001000",
  30625=>"000010111",
  30626=>"110110111",
  30627=>"110111111",
  30628=>"000100111",
  30629=>"000000000",
  30630=>"001111111",
  30631=>"100111111",
  30632=>"100000001",
  30633=>"000000000",
  30634=>"000100011",
  30635=>"111111000",
  30636=>"000000000",
  30637=>"111111111",
  30638=>"001000000",
  30639=>"111111011",
  30640=>"011000000",
  30641=>"111111111",
  30642=>"111111111",
  30643=>"111011111",
  30644=>"001110111",
  30645=>"111000100",
  30646=>"000101111",
  30647=>"111111100",
  30648=>"101100100",
  30649=>"000111111",
  30650=>"000011111",
  30651=>"001000001",
  30652=>"011001000",
  30653=>"111110000",
  30654=>"101100111",
  30655=>"010000010",
  30656=>"111111111",
  30657=>"000000001",
  30658=>"111111011",
  30659=>"000000000",
  30660=>"000110011",
  30661=>"111001111",
  30662=>"101000010",
  30663=>"000000001",
  30664=>"111011010",
  30665=>"000100011",
  30666=>"000000000",
  30667=>"011000000",
  30668=>"111001000",
  30669=>"000101011",
  30670=>"111101000",
  30671=>"111111111",
  30672=>"111010000",
  30673=>"111111111",
  30674=>"000100110",
  30675=>"111111001",
  30676=>"000111000",
  30677=>"000000111",
  30678=>"111111101",
  30679=>"111111011",
  30680=>"111000000",
  30681=>"110111111",
  30682=>"000000111",
  30683=>"000000001",
  30684=>"000111110",
  30685=>"000111111",
  30686=>"111001111",
  30687=>"000000110",
  30688=>"011111111",
  30689=>"000000000",
  30690=>"011111111",
  30691=>"111111100",
  30692=>"000111111",
  30693=>"101000011",
  30694=>"000000000",
  30695=>"111111111",
  30696=>"111100111",
  30697=>"000111111",
  30698=>"111110100",
  30699=>"000000000",
  30700=>"111000100",
  30701=>"001111100",
  30702=>"000000000",
  30703=>"111111111",
  30704=>"000000111",
  30705=>"000000000",
  30706=>"011111011",
  30707=>"111000100",
  30708=>"111111000",
  30709=>"111111111",
  30710=>"000111111",
  30711=>"111011111",
  30712=>"111000000",
  30713=>"001000000",
  30714=>"000000010",
  30715=>"011000000",
  30716=>"000000000",
  30717=>"110110110",
  30718=>"011000010",
  30719=>"001001011",
  30720=>"111111111",
  30721=>"000110111",
  30722=>"111001111",
  30723=>"100100110",
  30724=>"101111111",
  30725=>"111000000",
  30726=>"100101111",
  30727=>"111011011",
  30728=>"100001111",
  30729=>"111110110",
  30730=>"111111000",
  30731=>"111111110",
  30732=>"101101100",
  30733=>"110000000",
  30734=>"000110111",
  30735=>"000011111",
  30736=>"111100110",
  30737=>"000000000",
  30738=>"111111111",
  30739=>"111111001",
  30740=>"111111000",
  30741=>"000000110",
  30742=>"000000100",
  30743=>"001001001",
  30744=>"111111100",
  30745=>"000011111",
  30746=>"000000111",
  30747=>"110111000",
  30748=>"000000111",
  30749=>"000001000",
  30750=>"000001001",
  30751=>"000000000",
  30752=>"110110110",
  30753=>"000010111",
  30754=>"111000000",
  30755=>"000000000",
  30756=>"111111010",
  30757=>"001100111",
  30758=>"000111110",
  30759=>"101000011",
  30760=>"111111111",
  30761=>"000000000",
  30762=>"101000111",
  30763=>"000000000",
  30764=>"001001111",
  30765=>"111000000",
  30766=>"001000000",
  30767=>"001111110",
  30768=>"000011111",
  30769=>"001000000",
  30770=>"001001001",
  30771=>"000100111",
  30772=>"000000000",
  30773=>"111111111",
  30774=>"000111010",
  30775=>"001000011",
  30776=>"000000000",
  30777=>"000000111",
  30778=>"101001000",
  30779=>"110110000",
  30780=>"111001001",
  30781=>"000001000",
  30782=>"010010010",
  30783=>"111100111",
  30784=>"001101000",
  30785=>"000000000",
  30786=>"101100111",
  30787=>"101111111",
  30788=>"111111100",
  30789=>"111111011",
  30790=>"000000111",
  30791=>"111111111",
  30792=>"001001001",
  30793=>"111101111",
  30794=>"000010010",
  30795=>"111111000",
  30796=>"111110110",
  30797=>"011111111",
  30798=>"001111110",
  30799=>"000000111",
  30800=>"000000000",
  30801=>"110110111",
  30802=>"000000000",
  30803=>"001111111",
  30804=>"000000001",
  30805=>"000000000",
  30806=>"011011111",
  30807=>"111111000",
  30808=>"011010010",
  30809=>"111001000",
  30810=>"111111000",
  30811=>"000000001",
  30812=>"111000000",
  30813=>"000110111",
  30814=>"111001001",
  30815=>"000000000",
  30816=>"000010000",
  30817=>"111001111",
  30818=>"000110111",
  30819=>"111111000",
  30820=>"111111111",
  30821=>"110000000",
  30822=>"000000001",
  30823=>"000000000",
  30824=>"000000000",
  30825=>"011000000",
  30826=>"001000000",
  30827=>"111111001",
  30828=>"111111111",
  30829=>"000000000",
  30830=>"101000001",
  30831=>"000000000",
  30832=>"000000100",
  30833=>"001101111",
  30834=>"111111010",
  30835=>"111111111",
  30836=>"000010111",
  30837=>"001001011",
  30838=>"111100000",
  30839=>"111000001",
  30840=>"111111110",
  30841=>"111010010",
  30842=>"111101001",
  30843=>"111101101",
  30844=>"110111101",
  30845=>"000000000",
  30846=>"110111001",
  30847=>"000000000",
  30848=>"010111111",
  30849=>"110100110",
  30850=>"000000000",
  30851=>"111111111",
  30852=>"000000000",
  30853=>"101100111",
  30854=>"111110000",
  30855=>"001001111",
  30856=>"111111110",
  30857=>"111111111",
  30858=>"111111101",
  30859=>"011000011",
  30860=>"111111111",
  30861=>"111110100",
  30862=>"000001101",
  30863=>"000001000",
  30864=>"000000100",
  30865=>"001001001",
  30866=>"110110100",
  30867=>"101111101",
  30868=>"000000111",
  30869=>"001101100",
  30870=>"111110111",
  30871=>"011000000",
  30872=>"001011111",
  30873=>"011011001",
  30874=>"000000010",
  30875=>"111000100",
  30876=>"110010010",
  30877=>"111110110",
  30878=>"000000110",
  30879=>"000000111",
  30880=>"000000111",
  30881=>"011111110",
  30882=>"001001001",
  30883=>"111111111",
  30884=>"001001001",
  30885=>"100100111",
  30886=>"011111111",
  30887=>"110110110",
  30888=>"001000000",
  30889=>"000000111",
  30890=>"111111111",
  30891=>"111101111",
  30892=>"111111010",
  30893=>"001001001",
  30894=>"000000000",
  30895=>"111111110",
  30896=>"111111111",
  30897=>"001111011",
  30898=>"011010011",
  30899=>"000000001",
  30900=>"000110100",
  30901=>"000000000",
  30902=>"000000000",
  30903=>"111110111",
  30904=>"010011111",
  30905=>"001000000",
  30906=>"000000000",
  30907=>"000000000",
  30908=>"000111111",
  30909=>"001001001",
  30910=>"110010000",
  30911=>"111110110",
  30912=>"100100000",
  30913=>"010111111",
  30914=>"110100111",
  30915=>"000010010",
  30916=>"111000000",
  30917=>"110010000",
  30918=>"000000000",
  30919=>"111111010",
  30920=>"000000010",
  30921=>"000000011",
  30922=>"111000101",
  30923=>"111110000",
  30924=>"100100111",
  30925=>"000001111",
  30926=>"000111111",
  30927=>"001001101",
  30928=>"011000000",
  30929=>"000000111",
  30930=>"101101000",
  30931=>"010111111",
  30932=>"111111111",
  30933=>"000000100",
  30934=>"000000010",
  30935=>"100000011",
  30936=>"111110000",
  30937=>"111111011",
  30938=>"111000100",
  30939=>"000111111",
  30940=>"010111110",
  30941=>"011001100",
  30942=>"001111111",
  30943=>"000000000",
  30944=>"001000111",
  30945=>"000000000",
  30946=>"101000000",
  30947=>"000000000",
  30948=>"111001001",
  30949=>"000001000",
  30950=>"101110010",
  30951=>"011111111",
  30952=>"110100100",
  30953=>"111110110",
  30954=>"111111111",
  30955=>"000000111",
  30956=>"100110000",
  30957=>"000000011",
  30958=>"000000010",
  30959=>"000110110",
  30960=>"111101111",
  30961=>"000111111",
  30962=>"001101000",
  30963=>"000000000",
  30964=>"010010111",
  30965=>"000100000",
  30966=>"111111110",
  30967=>"001001000",
  30968=>"011000000",
  30969=>"000000000",
  30970=>"011011011",
  30971=>"010011000",
  30972=>"001011111",
  30973=>"000000011",
  30974=>"000000000",
  30975=>"000001111",
  30976=>"111111111",
  30977=>"001000000",
  30978=>"000110111",
  30979=>"111110000",
  30980=>"100011011",
  30981=>"110110000",
  30982=>"110110111",
  30983=>"111010000",
  30984=>"011001000",
  30985=>"000001111",
  30986=>"001111111",
  30987=>"000000000",
  30988=>"111100000",
  30989=>"100110100",
  30990=>"000111111",
  30991=>"000000110",
  30992=>"000000101",
  30993=>"111111111",
  30994=>"001001001",
  30995=>"000001111",
  30996=>"111011000",
  30997=>"111111000",
  30998=>"011001101",
  30999=>"111111111",
  31000=>"011000000",
  31001=>"111111111",
  31002=>"000001001",
  31003=>"111000000",
  31004=>"100101111",
  31005=>"111111010",
  31006=>"000000000",
  31007=>"111101011",
  31008=>"001110111",
  31009=>"110111110",
  31010=>"001000000",
  31011=>"110111111",
  31012=>"001000010",
  31013=>"111111111",
  31014=>"100000001",
  31015=>"111111000",
  31016=>"001111010",
  31017=>"000010010",
  31018=>"010000000",
  31019=>"111010000",
  31020=>"001000000",
  31021=>"111111111",
  31022=>"100100000",
  31023=>"110111010",
  31024=>"001001001",
  31025=>"000111111",
  31026=>"011000000",
  31027=>"011010111",
  31028=>"111111100",
  31029=>"110110111",
  31030=>"000000100",
  31031=>"111111111",
  31032=>"001011010",
  31033=>"111101111",
  31034=>"000001111",
  31035=>"111011011",
  31036=>"111111010",
  31037=>"001111101",
  31038=>"000000001",
  31039=>"111110010",
  31040=>"000000000",
  31041=>"100110111",
  31042=>"000000110",
  31043=>"100111101",
  31044=>"111001000",
  31045=>"001000100",
  31046=>"000000100",
  31047=>"000000000",
  31048=>"000000000",
  31049=>"111101000",
  31050=>"010010110",
  31051=>"000000000",
  31052=>"000000000",
  31053=>"111111111",
  31054=>"001000101",
  31055=>"110110100",
  31056=>"000001001",
  31057=>"000101111",
  31058=>"000000000",
  31059=>"000111110",
  31060=>"000010111",
  31061=>"111011011",
  31062=>"010011000",
  31063=>"111101111",
  31064=>"111111001",
  31065=>"000000000",
  31066=>"000000010",
  31067=>"101010000",
  31068=>"100110110",
  31069=>"111011100",
  31070=>"000000101",
  31071=>"001011111",
  31072=>"010111110",
  31073=>"000000001",
  31074=>"000000101",
  31075=>"101001000",
  31076=>"111111111",
  31077=>"000000011",
  31078=>"110110010",
  31079=>"011111111",
  31080=>"000000000",
  31081=>"000000000",
  31082=>"010110000",
  31083=>"001111111",
  31084=>"000101111",
  31085=>"000011110",
  31086=>"000000000",
  31087=>"001001000",
  31088=>"000000000",
  31089=>"000010111",
  31090=>"000000101",
  31091=>"100100100",
  31092=>"000000000",
  31093=>"000111111",
  31094=>"000000101",
  31095=>"000000000",
  31096=>"000000000",
  31097=>"111001000",
  31098=>"001000001",
  31099=>"000000000",
  31100=>"100000001",
  31101=>"111111000",
  31102=>"000111111",
  31103=>"101101111",
  31104=>"011111111",
  31105=>"000100100",
  31106=>"111111110",
  31107=>"001000000",
  31108=>"110100000",
  31109=>"000001001",
  31110=>"000000111",
  31111=>"011111111",
  31112=>"000000000",
  31113=>"000000000",
  31114=>"100100100",
  31115=>"111101000",
  31116=>"111101111",
  31117=>"100100100",
  31118=>"111011000",
  31119=>"000000000",
  31120=>"000001111",
  31121=>"010110111",
  31122=>"111111000",
  31123=>"011110110",
  31124=>"111111111",
  31125=>"110111111",
  31126=>"100000000",
  31127=>"001001001",
  31128=>"011011011",
  31129=>"000001001",
  31130=>"010011011",
  31131=>"111111000",
  31132=>"010111111",
  31133=>"100000000",
  31134=>"000000000",
  31135=>"100111111",
  31136=>"010111111",
  31137=>"111011011",
  31138=>"111111100",
  31139=>"111101111",
  31140=>"010010111",
  31141=>"010000000",
  31142=>"111101101",
  31143=>"111000000",
  31144=>"100000000",
  31145=>"000011000",
  31146=>"000000110",
  31147=>"011001000",
  31148=>"000000000",
  31149=>"000000100",
  31150=>"000010110",
  31151=>"111111101",
  31152=>"111111110",
  31153=>"101000110",
  31154=>"011001000",
  31155=>"001111111",
  31156=>"111111111",
  31157=>"111111111",
  31158=>"011111111",
  31159=>"000000000",
  31160=>"000111111",
  31161=>"000110111",
  31162=>"111111111",
  31163=>"000000110",
  31164=>"011000111",
  31165=>"000000110",
  31166=>"000000000",
  31167=>"000000000",
  31168=>"111011111",
  31169=>"000000111",
  31170=>"000000011",
  31171=>"000000000",
  31172=>"000000001",
  31173=>"000001111",
  31174=>"010110100",
  31175=>"011001000",
  31176=>"000001000",
  31177=>"000000000",
  31178=>"000000000",
  31179=>"001001000",
  31180=>"111000001",
  31181=>"111111010",
  31182=>"001001000",
  31183=>"010111110",
  31184=>"110000000",
  31185=>"101000000",
  31186=>"110110110",
  31187=>"111011001",
  31188=>"111011011",
  31189=>"001000000",
  31190=>"001001001",
  31191=>"000000000",
  31192=>"000000000",
  31193=>"101101001",
  31194=>"011011000",
  31195=>"011000010",
  31196=>"110110110",
  31197=>"111111000",
  31198=>"111110111",
  31199=>"000000001",
  31200=>"001000111",
  31201=>"100111110",
  31202=>"000011010",
  31203=>"111000000",
  31204=>"000000000",
  31205=>"110110110",
  31206=>"111011111",
  31207=>"110111111",
  31208=>"000000000",
  31209=>"100100110",
  31210=>"000000000",
  31211=>"100110000",
  31212=>"011011011",
  31213=>"100100111",
  31214=>"000101110",
  31215=>"110111011",
  31216=>"000000101",
  31217=>"000110111",
  31218=>"000000101",
  31219=>"111111011",
  31220=>"010000000",
  31221=>"111111111",
  31222=>"001000001",
  31223=>"110110110",
  31224=>"000001011",
  31225=>"100000001",
  31226=>"000010110",
  31227=>"111111111",
  31228=>"010000111",
  31229=>"000001001",
  31230=>"000000000",
  31231=>"000000001",
  31232=>"011000000",
  31233=>"110111110",
  31234=>"000000000",
  31235=>"111111111",
  31236=>"111111011",
  31237=>"110110000",
  31238=>"111111110",
  31239=>"001000000",
  31240=>"011011011",
  31241=>"110111111",
  31242=>"111111111",
  31243=>"000110111",
  31244=>"000110000",
  31245=>"111111111",
  31246=>"001001000",
  31247=>"000000000",
  31248=>"110000000",
  31249=>"111111111",
  31250=>"000000000",
  31251=>"000000000",
  31252=>"000000000",
  31253=>"010110111",
  31254=>"110110110",
  31255=>"011111101",
  31256=>"100000100",
  31257=>"111111000",
  31258=>"111000000",
  31259=>"000101111",
  31260=>"111011011",
  31261=>"011001001",
  31262=>"000100110",
  31263=>"001011000",
  31264=>"000000111",
  31265=>"000000100",
  31266=>"011000000",
  31267=>"000000000",
  31268=>"100110111",
  31269=>"111111101",
  31270=>"111111000",
  31271=>"011011111",
  31272=>"000100100",
  31273=>"000000100",
  31274=>"000000000",
  31275=>"100000111",
  31276=>"111111110",
  31277=>"010111100",
  31278=>"000000000",
  31279=>"000100100",
  31280=>"111111110",
  31281=>"000000100",
  31282=>"000000000",
  31283=>"001001001",
  31284=>"000011000",
  31285=>"001000000",
  31286=>"111111001",
  31287=>"000000000",
  31288=>"000010111",
  31289=>"101000000",
  31290=>"000001111",
  31291=>"111111111",
  31292=>"001001111",
  31293=>"011111100",
  31294=>"111111111",
  31295=>"111111111",
  31296=>"111111100",
  31297=>"011010000",
  31298=>"111111110",
  31299=>"000000101",
  31300=>"000001000",
  31301=>"101111111",
  31302=>"000000110",
  31303=>"000111111",
  31304=>"011111001",
  31305=>"111001001",
  31306=>"111000000",
  31307=>"000000000",
  31308=>"010000111",
  31309=>"100101000",
  31310=>"111111111",
  31311=>"000000111",
  31312=>"001100000",
  31313=>"011111111",
  31314=>"000000000",
  31315=>"000000000",
  31316=>"111111111",
  31317=>"111111110",
  31318=>"001001111",
  31319=>"100110111",
  31320=>"111111110",
  31321=>"001000111",
  31322=>"111111000",
  31323=>"110110111",
  31324=>"111111000",
  31325=>"111111010",
  31326=>"111000000",
  31327=>"100011011",
  31328=>"111001111",
  31329=>"011010011",
  31330=>"100100000",
  31331=>"111001000",
  31332=>"110110000",
  31333=>"001000000",
  31334=>"000001111",
  31335=>"111111011",
  31336=>"111111000",
  31337=>"111011011",
  31338=>"110111111",
  31339=>"000000010",
  31340=>"111111011",
  31341=>"110010000",
  31342=>"101000111",
  31343=>"000100111",
  31344=>"000000100",
  31345=>"000000000",
  31346=>"000000010",
  31347=>"111111111",
  31348=>"111000000",
  31349=>"000010110",
  31350=>"110111111",
  31351=>"000000000",
  31352=>"001000000",
  31353=>"000101111",
  31354=>"101100000",
  31355=>"110101111",
  31356=>"000000000",
  31357=>"000000000",
  31358=>"111111111",
  31359=>"111110110",
  31360=>"000000000",
  31361=>"101101001",
  31362=>"110011000",
  31363=>"111111111",
  31364=>"000001000",
  31365=>"000111111",
  31366=>"111111111",
  31367=>"100100110",
  31368=>"100000000",
  31369=>"000111111",
  31370=>"001001000",
  31371=>"110011010",
  31372=>"000000011",
  31373=>"000001111",
  31374=>"111111111",
  31375=>"000000000",
  31376=>"000000001",
  31377=>"111110000",
  31378=>"110111110",
  31379=>"000000100",
  31380=>"111111111",
  31381=>"000100000",
  31382=>"000000100",
  31383=>"111011111",
  31384=>"001000000",
  31385=>"000000000",
  31386=>"100011111",
  31387=>"111001000",
  31388=>"111110110",
  31389=>"110000000",
  31390=>"001000000",
  31391=>"000000000",
  31392=>"000100100",
  31393=>"000110110",
  31394=>"000000000",
  31395=>"111111010",
  31396=>"111111111",
  31397=>"111111111",
  31398=>"000100111",
  31399=>"101011001",
  31400=>"110011101",
  31401=>"000000100",
  31402=>"000000000",
  31403=>"001111111",
  31404=>"001101001",
  31405=>"100100110",
  31406=>"111111110",
  31407=>"111110100",
  31408=>"011111111",
  31409=>"111110101",
  31410=>"001011011",
  31411=>"010000000",
  31412=>"000011000",
  31413=>"000000000",
  31414=>"101111111",
  31415=>"111111011",
  31416=>"011111111",
  31417=>"000000000",
  31418=>"111100000",
  31419=>"111101000",
  31420=>"001000000",
  31421=>"001001011",
  31422=>"111110111",
  31423=>"110110111",
  31424=>"111100111",
  31425=>"001011111",
  31426=>"000000110",
  31427=>"111111111",
  31428=>"111111000",
  31429=>"000111110",
  31430=>"000110110",
  31431=>"001000000",
  31432=>"000111111",
  31433=>"011000000",
  31434=>"100100110",
  31435=>"000000000",
  31436=>"111101111",
  31437=>"010110110",
  31438=>"000000000",
  31439=>"000000000",
  31440=>"000000000",
  31441=>"000101111",
  31442=>"111110000",
  31443=>"000000000",
  31444=>"101101011",
  31445=>"000001111",
  31446=>"111011000",
  31447=>"110111111",
  31448=>"111111111",
  31449=>"111111111",
  31450=>"111111110",
  31451=>"011001011",
  31452=>"000000111",
  31453=>"011111111",
  31454=>"000000000",
  31455=>"001111111",
  31456=>"000000111",
  31457=>"010010110",
  31458=>"000111111",
  31459=>"111110000",
  31460=>"000000100",
  31461=>"011000000",
  31462=>"110110111",
  31463=>"111001110",
  31464=>"111111000",
  31465=>"100111111",
  31466=>"000011111",
  31467=>"111111111",
  31468=>"000000000",
  31469=>"000000000",
  31470=>"111111111",
  31471=>"000000000",
  31472=>"111111110",
  31473=>"000100000",
  31474=>"000100111",
  31475=>"000000000",
  31476=>"111111111",
  31477=>"100000000",
  31478=>"101110110",
  31479=>"011000000",
  31480=>"111111000",
  31481=>"010000000",
  31482=>"111001100",
  31483=>"000100111",
  31484=>"111111111",
  31485=>"000101111",
  31486=>"111111110",
  31487=>"011111111",
  31488=>"000000001",
  31489=>"000000000",
  31490=>"000000001",
  31491=>"111111110",
  31492=>"110111111",
  31493=>"000111111",
  31494=>"001000000",
  31495=>"000000000",
  31496=>"110011000",
  31497=>"011111111",
  31498=>"111111111",
  31499=>"111001001",
  31500=>"000000000",
  31501=>"111011111",
  31502=>"111110010",
  31503=>"111011111",
  31504=>"000000000",
  31505=>"000110110",
  31506=>"111101001",
  31507=>"111111111",
  31508=>"111111111",
  31509=>"000011111",
  31510=>"000011100",
  31511=>"001000001",
  31512=>"011111110",
  31513=>"111110110",
  31514=>"111111000",
  31515=>"000000100",
  31516=>"001011011",
  31517=>"000000000",
  31518=>"000000000",
  31519=>"011111010",
  31520=>"111111111",
  31521=>"011000100",
  31522=>"111110000",
  31523=>"000000000",
  31524=>"000010011",
  31525=>"000100100",
  31526=>"011001011",
  31527=>"100000000",
  31528=>"000000011",
  31529=>"111111001",
  31530=>"000000100",
  31531=>"111001111",
  31532=>"000001001",
  31533=>"111110000",
  31534=>"000111110",
  31535=>"000000000",
  31536=>"010000000",
  31537=>"001001000",
  31538=>"000000000",
  31539=>"000110010",
  31540=>"000010100",
  31541=>"000000000",
  31542=>"000000000",
  31543=>"101000000",
  31544=>"110110000",
  31545=>"100000000",
  31546=>"001000000",
  31547=>"111000000",
  31548=>"111111111",
  31549=>"011110000",
  31550=>"011111000",
  31551=>"001011000",
  31552=>"000000000",
  31553=>"000000000",
  31554=>"111111011",
  31555=>"000000000",
  31556=>"111000000",
  31557=>"101111111",
  31558=>"000000110",
  31559=>"000000000",
  31560=>"111100000",
  31561=>"010010000",
  31562=>"000100000",
  31563=>"000000111",
  31564=>"000100110",
  31565=>"111111000",
  31566=>"111111111",
  31567=>"000000000",
  31568=>"111111011",
  31569=>"011011000",
  31570=>"111111111",
  31571=>"011111111",
  31572=>"100000111",
  31573=>"011001001",
  31574=>"001100000",
  31575=>"000000111",
  31576=>"000001001",
  31577=>"000000000",
  31578=>"000000000",
  31579=>"111111111",
  31580=>"000000000",
  31581=>"110100110",
  31582=>"011111111",
  31583=>"111111111",
  31584=>"111000000",
  31585=>"000000000",
  31586=>"000000000",
  31587=>"111111111",
  31588=>"001110110",
  31589=>"000000000",
  31590=>"111100000",
  31591=>"111101111",
  31592=>"110010110",
  31593=>"000000111",
  31594=>"111111111",
  31595=>"111111111",
  31596=>"111110110",
  31597=>"000010001",
  31598=>"111111111",
  31599=>"001000000",
  31600=>"000000101",
  31601=>"111111111",
  31602=>"000000000",
  31603=>"111111001",
  31604=>"110000000",
  31605=>"000000000",
  31606=>"000000011",
  31607=>"010000000",
  31608=>"000010010",
  31609=>"011111100",
  31610=>"000000000",
  31611=>"111100000",
  31612=>"100000000",
  31613=>"100000011",
  31614=>"111111010",
  31615=>"111111111",
  31616=>"000000000",
  31617=>"000000000",
  31618=>"100111111",
  31619=>"000000000",
  31620=>"000100111",
  31621=>"011111111",
  31622=>"000100110",
  31623=>"111011011",
  31624=>"000000000",
  31625=>"001111111",
  31626=>"000011011",
  31627=>"000000001",
  31628=>"110011111",
  31629=>"100100100",
  31630=>"000000011",
  31631=>"000000000",
  31632=>"000000110",
  31633=>"111111111",
  31634=>"000110100",
  31635=>"111011001",
  31636=>"111011111",
  31637=>"011011000",
  31638=>"000011001",
  31639=>"000100111",
  31640=>"011010110",
  31641=>"000000000",
  31642=>"111011000",
  31643=>"111111001",
  31644=>"100000000",
  31645=>"000000101",
  31646=>"000000000",
  31647=>"110110000",
  31648=>"100000111",
  31649=>"000100100",
  31650=>"011011001",
  31651=>"111111000",
  31652=>"111110100",
  31653=>"111111001",
  31654=>"000000000",
  31655=>"000000000",
  31656=>"011011001",
  31657=>"111111111",
  31658=>"100001111",
  31659=>"111000000",
  31660=>"111111110",
  31661=>"000000011",
  31662=>"110000000",
  31663=>"110000001",
  31664=>"110101001",
  31665=>"000000000",
  31666=>"000000000",
  31667=>"000000000",
  31668=>"100000011",
  31669=>"011111011",
  31670=>"000000000",
  31671=>"001001111",
  31672=>"111110110",
  31673=>"101111111",
  31674=>"100110110",
  31675=>"101100111",
  31676=>"110100110",
  31677=>"011001001",
  31678=>"110111100",
  31679=>"001011000",
  31680=>"011011001",
  31681=>"000000000",
  31682=>"000111111",
  31683=>"110111111",
  31684=>"000000000",
  31685=>"001000000",
  31686=>"000000110",
  31687=>"000000111",
  31688=>"111001000",
  31689=>"111001000",
  31690=>"010100110",
  31691=>"111000000",
  31692=>"000000000",
  31693=>"000000010",
  31694=>"011010110",
  31695=>"101101110",
  31696=>"001011111",
  31697=>"111111011",
  31698=>"011000101",
  31699=>"001000100",
  31700=>"001001111",
  31701=>"000000111",
  31702=>"000000000",
  31703=>"111111111",
  31704=>"001000000",
  31705=>"010010011",
  31706=>"011000000",
  31707=>"000000000",
  31708=>"000000000",
  31709=>"111001000",
  31710=>"111011000",
  31711=>"110111111",
  31712=>"111111111",
  31713=>"000000000",
  31714=>"000000111",
  31715=>"011110110",
  31716=>"111111111",
  31717=>"111111000",
  31718=>"111111101",
  31719=>"110111010",
  31720=>"111100110",
  31721=>"000000000",
  31722=>"011010011",
  31723=>"111100000",
  31724=>"111000000",
  31725=>"000100000",
  31726=>"000000101",
  31727=>"111000001",
  31728=>"100100111",
  31729=>"000000000",
  31730=>"101000001",
  31731=>"000000000",
  31732=>"001001001",
  31733=>"100100000",
  31734=>"000101111",
  31735=>"000011111",
  31736=>"011011000",
  31737=>"111100000",
  31738=>"000100100",
  31739=>"111111111",
  31740=>"111011111",
  31741=>"111101101",
  31742=>"000101111",
  31743=>"111100110",
  31744=>"110110111",
  31745=>"111110110",
  31746=>"000000000",
  31747=>"111111000",
  31748=>"101111111",
  31749=>"000000000",
  31750=>"111111111",
  31751=>"111111111",
  31752=>"011000000",
  31753=>"110100011",
  31754=>"000000000",
  31755=>"100100000",
  31756=>"011110000",
  31757=>"000000000",
  31758=>"111111111",
  31759=>"001001001",
  31760=>"100100000",
  31761=>"111110011",
  31762=>"111111110",
  31763=>"101101101",
  31764=>"000000000",
  31765=>"011111000",
  31766=>"000000010",
  31767=>"001001001",
  31768=>"111111111",
  31769=>"001011111",
  31770=>"000000000",
  31771=>"110111111",
  31772=>"011001001",
  31773=>"000000000",
  31774=>"111111111",
  31775=>"001011111",
  31776=>"001001111",
  31777=>"000000100",
  31778=>"010010000",
  31779=>"110100110",
  31780=>"000000000",
  31781=>"011111111",
  31782=>"000000000",
  31783=>"000000000",
  31784=>"000000111",
  31785=>"000000000",
  31786=>"101101101",
  31787=>"000001111",
  31788=>"000000011",
  31789=>"000011011",
  31790=>"111001111",
  31791=>"000100100",
  31792=>"000000100",
  31793=>"011011001",
  31794=>"001000000",
  31795=>"100000100",
  31796=>"000010000",
  31797=>"111011011",
  31798=>"000010000",
  31799=>"111101001",
  31800=>"100111111",
  31801=>"000110110",
  31802=>"111111111",
  31803=>"111111111",
  31804=>"101000001",
  31805=>"000000001",
  31806=>"000000100",
  31807=>"000000000",
  31808=>"100000010",
  31809=>"111111111",
  31810=>"111111101",
  31811=>"111110111",
  31812=>"011111111",
  31813=>"001001111",
  31814=>"100100000",
  31815=>"100000000",
  31816=>"001001001",
  31817=>"111111110",
  31818=>"000000000",
  31819=>"101111111",
  31820=>"110111110",
  31821=>"010000000",
  31822=>"001000000",
  31823=>"000000111",
  31824=>"010111010",
  31825=>"110100100",
  31826=>"100000110",
  31827=>"100100000",
  31828=>"101111111",
  31829=>"111100000",
  31830=>"111111000",
  31831=>"001000000",
  31832=>"100000001",
  31833=>"100000100",
  31834=>"000000111",
  31835=>"010010000",
  31836=>"000100111",
  31837=>"001000000",
  31838=>"111111100",
  31839=>"010010000",
  31840=>"000000000",
  31841=>"000000001",
  31842=>"111110000",
  31843=>"011110011",
  31844=>"010000000",
  31845=>"110100100",
  31846=>"100100000",
  31847=>"100100000",
  31848=>"000100111",
  31849=>"001011111",
  31850=>"111111111",
  31851=>"111111110",
  31852=>"100111111",
  31853=>"111100100",
  31854=>"110100100",
  31855=>"000000000",
  31856=>"110111111",
  31857=>"001000100",
  31858=>"001000000",
  31859=>"110100100",
  31860=>"001000001",
  31861=>"000000001",
  31862=>"111011000",
  31863=>"111111111",
  31864=>"010000000",
  31865=>"001000111",
  31866=>"110100100",
  31867=>"000110110",
  31868=>"111111111",
  31869=>"000000000",
  31870=>"111111111",
  31871=>"000000000",
  31872=>"111111100",
  31873=>"111111111",
  31874=>"111111111",
  31875=>"000011001",
  31876=>"000000000",
  31877=>"111111111",
  31878=>"100111010",
  31879=>"000011011",
  31880=>"011000000",
  31881=>"000100100",
  31882=>"011001101",
  31883=>"001000000",
  31884=>"101000000",
  31885=>"110100110",
  31886=>"110111110",
  31887=>"011011011",
  31888=>"101111111",
  31889=>"000000001",
  31890=>"000000000",
  31891=>"011001000",
  31892=>"111111111",
  31893=>"111110111",
  31894=>"000001111",
  31895=>"001000000",
  31896=>"000000000",
  31897=>"000000111",
  31898=>"000010100",
  31899=>"011000001",
  31900=>"111111010",
  31901=>"101100100",
  31902=>"111111110",
  31903=>"110111101",
  31904=>"111111000",
  31905=>"110110111",
  31906=>"111101101",
  31907=>"000000000",
  31908=>"111100000",
  31909=>"000000001",
  31910=>"111101110",
  31911=>"000000000",
  31912=>"000000110",
  31913=>"000000000",
  31914=>"111111110",
  31915=>"000000000",
  31916=>"100000001",
  31917=>"111111011",
  31918=>"000000000",
  31919=>"011110110",
  31920=>"111111111",
  31921=>"111000000",
  31922=>"010111010",
  31923=>"000000000",
  31924=>"110110110",
  31925=>"101001000",
  31926=>"111000000",
  31927=>"101000111",
  31928=>"110111111",
  31929=>"011011000",
  31930=>"101100101",
  31931=>"010010000",
  31932=>"000000000",
  31933=>"011011011",
  31934=>"110111111",
  31935=>"000001101",
  31936=>"111100111",
  31937=>"111111111",
  31938=>"101001001",
  31939=>"111100000",
  31940=>"001001000",
  31941=>"000000000",
  31942=>"110100000",
  31943=>"111111110",
  31944=>"010010010",
  31945=>"111111111",
  31946=>"000000000",
  31947=>"111111111",
  31948=>"000000000",
  31949=>"111001001",
  31950=>"000001111",
  31951=>"111100110",
  31952=>"000010011",
  31953=>"001001111",
  31954=>"111111110",
  31955=>"000110100",
  31956=>"001001001",
  31957=>"111111111",
  31958=>"000000000",
  31959=>"001001001",
  31960=>"111111110",
  31961=>"001001111",
  31962=>"000111010",
  31963=>"011011011",
  31964=>"110100100",
  31965=>"000000100",
  31966=>"000000011",
  31967=>"111000111",
  31968=>"000100111",
  31969=>"010010110",
  31970=>"000000011",
  31971=>"011010010",
  31972=>"000000111",
  31973=>"110000000",
  31974=>"000111010",
  31975=>"101101000",
  31976=>"001111111",
  31977=>"000010111",
  31978=>"001011111",
  31979=>"001000110",
  31980=>"111111111",
  31981=>"000000000",
  31982=>"111000000",
  31983=>"000000000",
  31984=>"001000000",
  31985=>"111100111",
  31986=>"111111001",
  31987=>"001001111",
  31988=>"111111111",
  31989=>"000001001",
  31990=>"100100000",
  31991=>"000010111",
  31992=>"000101111",
  31993=>"111111111",
  31994=>"000000001",
  31995=>"011001101",
  31996=>"011000010",
  31997=>"111001100",
  31998=>"101000000",
  31999=>"111111111",
  32000=>"011011101",
  32001=>"000000000",
  32002=>"000001101",
  32003=>"000000001",
  32004=>"101101111",
  32005=>"000111111",
  32006=>"111111000",
  32007=>"110111100",
  32008=>"000001111",
  32009=>"111000111",
  32010=>"011011111",
  32011=>"111110010",
  32012=>"000000000",
  32013=>"111111111",
  32014=>"010010000",
  32015=>"011011011",
  32016=>"110110000",
  32017=>"010011010",
  32018=>"110000000",
  32019=>"011110110",
  32020=>"111111111",
  32021=>"110111001",
  32022=>"010110000",
  32023=>"000000001",
  32024=>"011001101",
  32025=>"111111111",
  32026=>"110110110",
  32027=>"001001000",
  32028=>"001011111",
  32029=>"111010011",
  32030=>"000000000",
  32031=>"001011011",
  32032=>"110110000",
  32033=>"000000111",
  32034=>"110110000",
  32035=>"111111000",
  32036=>"111111100",
  32037=>"010011111",
  32038=>"011010011",
  32039=>"111111111",
  32040=>"001000000",
  32041=>"001001101",
  32042=>"000010000",
  32043=>"010111111",
  32044=>"000010000",
  32045=>"100000011",
  32046=>"100111111",
  32047=>"000000000",
  32048=>"110110000",
  32049=>"011111000",
  32050=>"010000100",
  32051=>"111111010",
  32052=>"000000000",
  32053=>"000010000",
  32054=>"111111110",
  32055=>"000010011",
  32056=>"110110000",
  32057=>"100100100",
  32058=>"000000000",
  32059=>"111111110",
  32060=>"000001000",
  32061=>"000000000",
  32062=>"101101000",
  32063=>"001001000",
  32064=>"000000000",
  32065=>"000100000",
  32066=>"111111111",
  32067=>"010110100",
  32068=>"011011011",
  32069=>"000000000",
  32070=>"111111111",
  32071=>"111011000",
  32072=>"000000000",
  32073=>"100100100",
  32074=>"010110000",
  32075=>"110100100",
  32076=>"001000000",
  32077=>"111111111",
  32078=>"110100000",
  32079=>"000000001",
  32080=>"111001001",
  32081=>"001000110",
  32082=>"000000000",
  32083=>"000000000",
  32084=>"111111001",
  32085=>"011011011",
  32086=>"111111000",
  32087=>"000000101",
  32088=>"100100000",
  32089=>"000000000",
  32090=>"011001001",
  32091=>"100000111",
  32092=>"010110000",
  32093=>"001001001",
  32094=>"000000000",
  32095=>"111110110",
  32096=>"000100100",
  32097=>"111101101",
  32098=>"111111110",
  32099=>"111111010",
  32100=>"001001001",
  32101=>"101000101",
  32102=>"000000010",
  32103=>"000000000",
  32104=>"001111011",
  32105=>"111111110",
  32106=>"011011110",
  32107=>"010010000",
  32108=>"111111110",
  32109=>"100111001",
  32110=>"110010000",
  32111=>"001001011",
  32112=>"000000000",
  32113=>"111111111",
  32114=>"010000010",
  32115=>"001100100",
  32116=>"100000001",
  32117=>"000000001",
  32118=>"100000000",
  32119=>"000011000",
  32120=>"000000100",
  32121=>"000000111",
  32122=>"110100101",
  32123=>"000000001",
  32124=>"110110000",
  32125=>"010111000",
  32126=>"110110110",
  32127=>"111100000",
  32128=>"001111001",
  32129=>"100111110",
  32130=>"000000000",
  32131=>"100100100",
  32132=>"000000000",
  32133=>"111100100",
  32134=>"111111111",
  32135=>"110111110",
  32136=>"000000000",
  32137=>"000001111",
  32138=>"111110000",
  32139=>"100111111",
  32140=>"111111111",
  32141=>"000000000",
  32142=>"110010000",
  32143=>"000110100",
  32144=>"111111111",
  32145=>"111111000",
  32146=>"000000000",
  32147=>"110110110",
  32148=>"000000000",
  32149=>"000001000",
  32150=>"111111111",
  32151=>"011001000",
  32152=>"110111111",
  32153=>"111111101",
  32154=>"000000000",
  32155=>"001111110",
  32156=>"000000011",
  32157=>"000000001",
  32158=>"001001001",
  32159=>"000000011",
  32160=>"101100100",
  32161=>"001001000",
  32162=>"000000000",
  32163=>"100110110",
  32164=>"101101111",
  32165=>"111110111",
  32166=>"000000000",
  32167=>"010110110",
  32168=>"111111000",
  32169=>"011011011",
  32170=>"111111111",
  32171=>"001000011",
  32172=>"111111000",
  32173=>"000000000",
  32174=>"110010000",
  32175=>"111111111",
  32176=>"100100110",
  32177=>"011011000",
  32178=>"111111111",
  32179=>"000001001",
  32180=>"111101101",
  32181=>"100000000",
  32182=>"111111010",
  32183=>"000000000",
  32184=>"000000000",
  32185=>"000010010",
  32186=>"110100000",
  32187=>"001000000",
  32188=>"111010000",
  32189=>"000110000",
  32190=>"011000000",
  32191=>"000000000",
  32192=>"000000000",
  32193=>"110111111",
  32194=>"001001111",
  32195=>"000110111",
  32196=>"111110111",
  32197=>"101111111",
  32198=>"000000000",
  32199=>"000000111",
  32200=>"000001000",
  32201=>"000000110",
  32202=>"110110110",
  32203=>"000110111",
  32204=>"111110000",
  32205=>"000000011",
  32206=>"000001000",
  32207=>"101100000",
  32208=>"111111111",
  32209=>"100000011",
  32210=>"111111111",
  32211=>"001001011",
  32212=>"011111111",
  32213=>"001001111",
  32214=>"111110000",
  32215=>"011011001",
  32216=>"000001001",
  32217=>"000010111",
  32218=>"000000101",
  32219=>"111111000",
  32220=>"101011011",
  32221=>"001001001",
  32222=>"011111000",
  32223=>"000001000",
  32224=>"011011011",
  32225=>"000000000",
  32226=>"101111101",
  32227=>"111111111",
  32228=>"111111100",
  32229=>"000111111",
  32230=>"100100110",
  32231=>"110100000",
  32232=>"000111000",
  32233=>"001011000",
  32234=>"000000111",
  32235=>"111000111",
  32236=>"110111111",
  32237=>"000110111",
  32238=>"111101000",
  32239=>"110100111",
  32240=>"000000101",
  32241=>"000110011",
  32242=>"100000100",
  32243=>"000000000",
  32244=>"100101111",
  32245=>"011011111",
  32246=>"000000000",
  32247=>"111111000",
  32248=>"000000000",
  32249=>"001000001",
  32250=>"010000000",
  32251=>"000000000",
  32252=>"110111111",
  32253=>"000000001",
  32254=>"000000011",
  32255=>"111111011",
  32256=>"000000000",
  32257=>"111000000",
  32258=>"100110100",
  32259=>"001001000",
  32260=>"000000000",
  32261=>"110110011",
  32262=>"100100001",
  32263=>"111111111",
  32264=>"000000000",
  32265=>"000000100",
  32266=>"100100110",
  32267=>"111111111",
  32268=>"000000000",
  32269=>"100001001",
  32270=>"100001101",
  32271=>"111111101",
  32272=>"000000001",
  32273=>"100111111",
  32274=>"010000000",
  32275=>"111111111",
  32276=>"111110000",
  32277=>"001111111",
  32278=>"000000001",
  32279=>"111111111",
  32280=>"111111111",
  32281=>"000001001",
  32282=>"111100111",
  32283=>"000000001",
  32284=>"000000000",
  32285=>"000000000",
  32286=>"001011010",
  32287=>"111000010",
  32288=>"111111001",
  32289=>"000000000",
  32290=>"010011011",
  32291=>"000000000",
  32292=>"000000000",
  32293=>"111110100",
  32294=>"000000000",
  32295=>"111111111",
  32296=>"111011011",
  32297=>"000000000",
  32298=>"000000101",
  32299=>"111111111",
  32300=>"111111111",
  32301=>"000011111",
  32302=>"000000000",
  32303=>"011011011",
  32304=>"110000010",
  32305=>"111000000",
  32306=>"100100000",
  32307=>"111111000",
  32308=>"000111111",
  32309=>"000011111",
  32310=>"111100000",
  32311=>"000000000",
  32312=>"111111111",
  32313=>"001001001",
  32314=>"000000000",
  32315=>"011000000",
  32316=>"011001111",
  32317=>"000000001",
  32318=>"010010000",
  32319=>"000000000",
  32320=>"101101100",
  32321=>"100000000",
  32322=>"000000000",
  32323=>"111111111",
  32324=>"110000000",
  32325=>"000000100",
  32326=>"111111111",
  32327=>"011111111",
  32328=>"000110100",
  32329=>"000000000",
  32330=>"001011001",
  32331=>"111011011",
  32332=>"111011001",
  32333=>"111111111",
  32334=>"110111111",
  32335=>"001001001",
  32336=>"011001000",
  32337=>"001000111",
  32338=>"111111111",
  32339=>"000000000",
  32340=>"000000000",
  32341=>"111000000",
  32342=>"110111111",
  32343=>"000000000",
  32344=>"011000110",
  32345=>"111000000",
  32346=>"111011111",
  32347=>"000000000",
  32348=>"010010011",
  32349=>"111111111",
  32350=>"111111100",
  32351=>"000001111",
  32352=>"000000000",
  32353=>"111111111",
  32354=>"010110110",
  32355=>"101111100",
  32356=>"000111011",
  32357=>"100110110",
  32358=>"111111111",
  32359=>"000001001",
  32360=>"011011111",
  32361=>"000000000",
  32362=>"101000000",
  32363=>"000001111",
  32364=>"001000000",
  32365=>"111111111",
  32366=>"111111110",
  32367=>"000000000",
  32368=>"111111111",
  32369=>"000001111",
  32370=>"001001001",
  32371=>"111111011",
  32372=>"000000110",
  32373=>"100110111",
  32374=>"111000000",
  32375=>"111111111",
  32376=>"000000000",
  32377=>"111001000",
  32378=>"000000000",
  32379=>"100000000",
  32380=>"000111111",
  32381=>"111001001",
  32382=>"111111101",
  32383=>"000000110",
  32384=>"000000000",
  32385=>"000000111",
  32386=>"111111111",
  32387=>"000000000",
  32388=>"111111111",
  32389=>"001101111",
  32390=>"110100110",
  32391=>"000010111",
  32392=>"011000011",
  32393=>"110111111",
  32394=>"100111111",
  32395=>"000101111",
  32396=>"011000001",
  32397=>"111111111",
  32398=>"101111111",
  32399=>"111000110",
  32400=>"111001001",
  32401=>"011000000",
  32402=>"100000100",
  32403=>"010000000",
  32404=>"001000100",
  32405=>"110111111",
  32406=>"000000000",
  32407=>"111011000",
  32408=>"111111011",
  32409=>"100100111",
  32410=>"111001111",
  32411=>"111111000",
  32412=>"111101111",
  32413=>"110110111",
  32414=>"001001011",
  32415=>"111111111",
  32416=>"000110111",
  32417=>"111011111",
  32418=>"000000000",
  32419=>"110000000",
  32420=>"000011111",
  32421=>"000000111",
  32422=>"000000000",
  32423=>"001111111",
  32424=>"011000000",
  32425=>"001001000",
  32426=>"000000000",
  32427=>"000010111",
  32428=>"110101111",
  32429=>"111111000",
  32430=>"000000000",
  32431=>"001111111",
  32432=>"111111111",
  32433=>"000000011",
  32434=>"011111111",
  32435=>"111111000",
  32436=>"100101111",
  32437=>"000000000",
  32438=>"010000000",
  32439=>"100000000",
  32440=>"001000000",
  32441=>"000000111",
  32442=>"000101101",
  32443=>"000000001",
  32444=>"111111111",
  32445=>"100100000",
  32446=>"110100000",
  32447=>"000000000",
  32448=>"111111000",
  32449=>"110100111",
  32450=>"000000000",
  32451=>"111111111",
  32452=>"000000001",
  32453=>"101111111",
  32454=>"111111000",
  32455=>"111000000",
  32456=>"010001000",
  32457=>"100000100",
  32458=>"000100111",
  32459=>"111100100",
  32460=>"111111100",
  32461=>"111111111",
  32462=>"111000110",
  32463=>"100100111",
  32464=>"111111000",
  32465=>"000010011",
  32466=>"111100111",
  32467=>"000000000",
  32468=>"000000111",
  32469=>"000000000",
  32470=>"000110111",
  32471=>"000000000",
  32472=>"000000000",
  32473=>"111111110",
  32474=>"000000000",
  32475=>"111000000",
  32476=>"000000000",
  32477=>"111000000",
  32478=>"111111011",
  32479=>"111111011",
  32480=>"000000111",
  32481=>"000010000",
  32482=>"011111010",
  32483=>"111111011",
  32484=>"000011000",
  32485=>"111000000",
  32486=>"000000001",
  32487=>"001001000",
  32488=>"000000000",
  32489=>"111111111",
  32490=>"000111111",
  32491=>"111101000",
  32492=>"001011000",
  32493=>"000000000",
  32494=>"010010000",
  32495=>"111111000",
  32496=>"000000101",
  32497=>"110011000",
  32498=>"000000011",
  32499=>"001001111",
  32500=>"111100100",
  32501=>"001011000",
  32502=>"000111011",
  32503=>"111001000",
  32504=>"111111111",
  32505=>"011111011",
  32506=>"111111100",
  32507=>"111010000",
  32508=>"000000000",
  32509=>"001001001",
  32510=>"100000000",
  32511=>"011011010",
  32512=>"101001011",
  32513=>"000001001",
  32514=>"111111000",
  32515=>"111111111",
  32516=>"000000001",
  32517=>"111111111",
  32518=>"000001000",
  32519=>"000000000",
  32520=>"111101101",
  32521=>"000000000",
  32522=>"110111011",
  32523=>"100111111",
  32524=>"000000110",
  32525=>"110000010",
  32526=>"101001001",
  32527=>"111111111",
  32528=>"111111111",
  32529=>"000000101",
  32530=>"111110110",
  32531=>"000100110",
  32532=>"111111000",
  32533=>"000000000",
  32534=>"111111111",
  32535=>"111110000",
  32536=>"111111100",
  32537=>"000000000",
  32538=>"000000000",
  32539=>"000000000",
  32540=>"000011011",
  32541=>"000000000",
  32542=>"111111000",
  32543=>"111111111",
  32544=>"110100000",
  32545=>"000000000",
  32546=>"000000000",
  32547=>"000000000",
  32548=>"000000000",
  32549=>"111111111",
  32550=>"110100110",
  32551=>"111111000",
  32552=>"110111011",
  32553=>"000100100",
  32554=>"000100111",
  32555=>"000000000",
  32556=>"111111000",
  32557=>"111111000",
  32558=>"000100000",
  32559=>"000000000",
  32560=>"000100111",
  32561=>"000000000",
  32562=>"110000000",
  32563=>"100010011",
  32564=>"111100000",
  32565=>"000000000",
  32566=>"111000000",
  32567=>"000000000",
  32568=>"000000000",
  32569=>"111101111",
  32570=>"000100111",
  32571=>"000000000",
  32572=>"011001011",
  32573=>"000000100",
  32574=>"000001000",
  32575=>"111111001",
  32576=>"001000000",
  32577=>"100111111",
  32578=>"011011000",
  32579=>"000000000",
  32580=>"011000000",
  32581=>"000011010",
  32582=>"010000000",
  32583=>"011000001",
  32584=>"000000000",
  32585=>"110100000",
  32586=>"000000000",
  32587=>"111011011",
  32588=>"000000001",
  32589=>"100000000",
  32590=>"111000000",
  32591=>"100101111",
  32592=>"001000001",
  32593=>"111110000",
  32594=>"111111111",
  32595=>"110011001",
  32596=>"000000000",
  32597=>"011011011",
  32598=>"100100000",
  32599=>"000000000",
  32600=>"000000000",
  32601=>"000000100",
  32602=>"001011000",
  32603=>"000001001",
  32604=>"000000010",
  32605=>"011011111",
  32606=>"011001001",
  32607=>"001111111",
  32608=>"100100110",
  32609=>"100111000",
  32610=>"111101001",
  32611=>"001011011",
  32612=>"110010110",
  32613=>"000000001",
  32614=>"111111111",
  32615=>"001001001",
  32616=>"011011010",
  32617=>"111111011",
  32618=>"000000001",
  32619=>"000000111",
  32620=>"011111111",
  32621=>"101101011",
  32622=>"111100000",
  32623=>"000110110",
  32624=>"111001000",
  32625=>"000000000",
  32626=>"000111001",
  32627=>"000000000",
  32628=>"111111111",
  32629=>"111011000",
  32630=>"101101111",
  32631=>"110010000",
  32632=>"100000000",
  32633=>"000000000",
  32634=>"111111111",
  32635=>"110101111",
  32636=>"000000011",
  32637=>"111111011",
  32638=>"111111111",
  32639=>"000000111",
  32640=>"000000110",
  32641=>"011011111",
  32642=>"000000001",
  32643=>"111111111",
  32644=>"000000000",
  32645=>"010010000",
  32646=>"111111000",
  32647=>"000000111",
  32648=>"111111111",
  32649=>"000000000",
  32650=>"100100111",
  32651=>"111111111",
  32652=>"111101111",
  32653=>"000000000",
  32654=>"111111010",
  32655=>"111111010",
  32656=>"000000000",
  32657=>"000000000",
  32658=>"000000001",
  32659=>"110000111",
  32660=>"111111111",
  32661=>"000000000",
  32662=>"111110100",
  32663=>"001000111",
  32664=>"000000100",
  32665=>"110000011",
  32666=>"100110111",
  32667=>"000100111",
  32668=>"111111111",
  32669=>"111111011",
  32670=>"000000001",
  32671=>"000111011",
  32672=>"100100000",
  32673=>"111111011",
  32674=>"000001000",
  32675=>"110011111",
  32676=>"111100000",
  32677=>"111111111",
  32678=>"111000000",
  32679=>"000000000",
  32680=>"000000111",
  32681=>"011111110",
  32682=>"110111111",
  32683=>"000000111",
  32684=>"011011000",
  32685=>"111101101",
  32686=>"000100000",
  32687=>"000000000",
  32688=>"111111111",
  32689=>"110100000",
  32690=>"100111111",
  32691=>"000000000",
  32692=>"000110111",
  32693=>"000000000",
  32694=>"101111011",
  32695=>"101100000",
  32696=>"100111111",
  32697=>"111111111",
  32698=>"111111111",
  32699=>"011000101",
  32700=>"000000000",
  32701=>"000000100",
  32702=>"000000110",
  32703=>"011011001",
  32704=>"111111111",
  32705=>"000000000",
  32706=>"000000011",
  32707=>"111110000",
  32708=>"010000000",
  32709=>"000000111",
  32710=>"111100000",
  32711=>"011011001",
  32712=>"111101111",
  32713=>"100001011",
  32714=>"001111111",
  32715=>"011111000",
  32716=>"000000000",
  32717=>"111111110",
  32718=>"100100100",
  32719=>"111111111",
  32720=>"000000011",
  32721=>"011000110",
  32722=>"110000010",
  32723=>"111011011",
  32724=>"000000000",
  32725=>"111111111",
  32726=>"110000000",
  32727=>"000000001",
  32728=>"111000111",
  32729=>"011000000",
  32730=>"111111011",
  32731=>"111111001",
  32732=>"000000000",
  32733=>"000000101",
  32734=>"000000000",
  32735=>"000000001",
  32736=>"000000111",
  32737=>"000001001",
  32738=>"000000000",
  32739=>"000000000",
  32740=>"111111000",
  32741=>"000001001",
  32742=>"111000111",
  32743=>"111111111",
  32744=>"000000101",
  32745=>"111111111",
  32746=>"010000000",
  32747=>"111101111",
  32748=>"111111011",
  32749=>"111110001",
  32750=>"011011000",
  32751=>"100111111",
  32752=>"100000100",
  32753=>"000000000",
  32754=>"111110111",
  32755=>"101111111",
  32756=>"000000000",
  32757=>"110000000",
  32758=>"000000011",
  32759=>"111111111",
  32760=>"000000000",
  32761=>"111110000",
  32762=>"000000000",
  32763=>"111111111",
  32764=>"000000001",
  32765=>"111101000",
  32766=>"111111111",
  32767=>"000100110",
  32768=>"000000111",
  32769=>"111111000",
  32770=>"111111111",
  32771=>"000000111",
  32772=>"111111111",
  32773=>"111111111",
  32774=>"100000100",
  32775=>"000000000",
  32776=>"100111111",
  32777=>"000110111",
  32778=>"111111111",
  32779=>"000000000",
  32780=>"000011000",
  32781=>"000000010",
  32782=>"011111011",
  32783=>"001001000",
  32784=>"111111110",
  32785=>"000000000",
  32786=>"011111010",
  32787=>"000011011",
  32788=>"110111101",
  32789=>"001001001",
  32790=>"010000000",
  32791=>"000000001",
  32792=>"000000111",
  32793=>"000000000",
  32794=>"000000010",
  32795=>"000100100",
  32796=>"111111111",
  32797=>"111111110",
  32798=>"000000000",
  32799=>"000000100",
  32800=>"111111111",
  32801=>"000110111",
  32802=>"110010000",
  32803=>"000000110",
  32804=>"011000111",
  32805=>"111111111",
  32806=>"000010010",
  32807=>"001001111",
  32808=>"001111111",
  32809=>"000000000",
  32810=>"110000110",
  32811=>"000000000",
  32812=>"100000000",
  32813=>"001100100",
  32814=>"111111111",
  32815=>"111111111",
  32816=>"000011111",
  32817=>"111111111",
  32818=>"111110110",
  32819=>"111111111",
  32820=>"000000000",
  32821=>"100110000",
  32822=>"111111111",
  32823=>"000111111",
  32824=>"111111111",
  32825=>"000110111",
  32826=>"000000000",
  32827=>"000000000",
  32828=>"111111111",
  32829=>"000000000",
  32830=>"111111111",
  32831=>"111111111",
  32832=>"111111100",
  32833=>"110111111",
  32834=>"000000101",
  32835=>"000000001",
  32836=>"110000000",
  32837=>"111111110",
  32838=>"111111000",
  32839=>"000000000",
  32840=>"000000000",
  32841=>"000000000",
  32842=>"000000111",
  32843=>"000000011",
  32844=>"000111111",
  32845=>"011011100",
  32846=>"000000000",
  32847=>"100111111",
  32848=>"111111101",
  32849=>"111111111",
  32850=>"000000000",
  32851=>"010010000",
  32852=>"111111011",
  32853=>"001000000",
  32854=>"000000000",
  32855=>"011011011",
  32856=>"000000000",
  32857=>"100100111",
  32858=>"000000000",
  32859=>"000011111",
  32860=>"000000010",
  32861=>"000010011",
  32862=>"000000011",
  32863=>"100111100",
  32864=>"000000000",
  32865=>"011111111",
  32866=>"000000000",
  32867=>"001001000",
  32868=>"000000001",
  32869=>"101100111",
  32870=>"111111111",
  32871=>"010111111",
  32872=>"000111001",
  32873=>"000100111",
  32874=>"111110111",
  32875=>"000000000",
  32876=>"111000111",
  32877=>"110100111",
  32878=>"111111111",
  32879=>"001000100",
  32880=>"111111111",
  32881=>"100101111",
  32882=>"100100111",
  32883=>"011000111",
  32884=>"111110111",
  32885=>"111111110",
  32886=>"000000111",
  32887=>"111111111",
  32888=>"111111111",
  32889=>"000000000",
  32890=>"011011110",
  32891=>"000000000",
  32892=>"010110010",
  32893=>"111011111",
  32894=>"111111111",
  32895=>"111111111",
  32896=>"000001101",
  32897=>"111111011",
  32898=>"111111111",
  32899=>"011000000",
  32900=>"110100111",
  32901=>"111111111",
  32902=>"000000001",
  32903=>"000001111",
  32904=>"111111111",
  32905=>"111111111",
  32906=>"000100111",
  32907=>"111111111",
  32908=>"111111111",
  32909=>"110010000",
  32910=>"000000000",
  32911=>"111111110",
  32912=>"000000000",
  32913=>"101100111",
  32914=>"000000100",
  32915=>"111111111",
  32916=>"101111111",
  32917=>"111100000",
  32918=>"111111111",
  32919=>"110111000",
  32920=>"000000111",
  32921=>"111100111",
  32922=>"000000111",
  32923=>"111111111",
  32924=>"000001111",
  32925=>"011001100",
  32926=>"110000000",
  32927=>"111111111",
  32928=>"011000000",
  32929=>"111100000",
  32930=>"111101001",
  32931=>"111111111",
  32932=>"001011000",
  32933=>"111011001",
  32934=>"111101110",
  32935=>"011000000",
  32936=>"111111111",
  32937=>"011111000",
  32938=>"111111111",
  32939=>"101101001",
  32940=>"110000011",
  32941=>"000110111",
  32942=>"000000000",
  32943=>"001001000",
  32944=>"111111111",
  32945=>"100000000",
  32946=>"111111100",
  32947=>"111000000",
  32948=>"110110100",
  32949=>"111111111",
  32950=>"000000000",
  32951=>"001000000",
  32952=>"111111111",
  32953=>"001001011",
  32954=>"000000111",
  32955=>"011011000",
  32956=>"111111111",
  32957=>"000000000",
  32958=>"000000000",
  32959=>"101101111",
  32960=>"000110100",
  32961=>"101011111",
  32962=>"011000001",
  32963=>"000000000",
  32964=>"011011011",
  32965=>"000000000",
  32966=>"111111111",
  32967=>"000000111",
  32968=>"000000000",
  32969=>"111111111",
  32970=>"111111111",
  32971=>"000000000",
  32972=>"111111111",
  32973=>"111111101",
  32974=>"011000000",
  32975=>"000000000",
  32976=>"111000000",
  32977=>"001000000",
  32978=>"111101000",
  32979=>"111111111",
  32980=>"111111110",
  32981=>"000000000",
  32982=>"111111111",
  32983=>"000001000",
  32984=>"000000000",
  32985=>"011000000",
  32986=>"111111111",
  32987=>"111111011",
  32988=>"111000000",
  32989=>"111111111",
  32990=>"101111111",
  32991=>"110111111",
  32992=>"111111111",
  32993=>"111111111",
  32994=>"000000000",
  32995=>"011011111",
  32996=>"111011000",
  32997=>"110110110",
  32998=>"000000000",
  32999=>"001111000",
  33000=>"111000000",
  33001=>"111110110",
  33002=>"111100000",
  33003=>"111110111",
  33004=>"000111000",
  33005=>"111111111",
  33006=>"000000000",
  33007=>"011000000",
  33008=>"010010110",
  33009=>"000000000",
  33010=>"001001001",
  33011=>"001001000",
  33012=>"000000000",
  33013=>"110110110",
  33014=>"000110110",
  33015=>"001000001",
  33016=>"110111111",
  33017=>"000111111",
  33018=>"111000000",
  33019=>"000000000",
  33020=>"100100111",
  33021=>"001111111",
  33022=>"011111011",
  33023=>"111110111",
  33024=>"000000001",
  33025=>"011000011",
  33026=>"111111111",
  33027=>"011111111",
  33028=>"111111111",
  33029=>"101101111",
  33030=>"110000000",
  33031=>"000000010",
  33032=>"000000111",
  33033=>"000000000",
  33034=>"100111111",
  33035=>"111110111",
  33036=>"000000000",
  33037=>"000000000",
  33038=>"000000000",
  33039=>"111111111",
  33040=>"000000000",
  33041=>"000000001",
  33042=>"110100100",
  33043=>"111111111",
  33044=>"000111001",
  33045=>"000000000",
  33046=>"110110010",
  33047=>"001001111",
  33048=>"101101000",
  33049=>"111111111",
  33050=>"000000000",
  33051=>"100000000",
  33052=>"011011111",
  33053=>"000111111",
  33054=>"111111111",
  33055=>"000000000",
  33056=>"010111111",
  33057=>"000000000",
  33058=>"111111111",
  33059=>"000000000",
  33060=>"100110110",
  33061=>"101111101",
  33062=>"111111110",
  33063=>"111111111",
  33064=>"111111011",
  33065=>"111111111",
  33066=>"011101111",
  33067=>"110000111",
  33068=>"000001000",
  33069=>"000000011",
  33070=>"110100000",
  33071=>"000000000",
  33072=>"000000010",
  33073=>"110111111",
  33074=>"011000000",
  33075=>"011111111",
  33076=>"000010010",
  33077=>"011000000",
  33078=>"000000011",
  33079=>"000000000",
  33080=>"100000000",
  33081=>"000000000",
  33082=>"111111111",
  33083=>"010000000",
  33084=>"000000000",
  33085=>"001000000",
  33086=>"000000000",
  33087=>"000000000",
  33088=>"000000000",
  33089=>"001000000",
  33090=>"000111111",
  33091=>"000000011",
  33092=>"111111111",
  33093=>"000000000",
  33094=>"000000111",
  33095=>"111000000",
  33096=>"000000000",
  33097=>"000110100",
  33098=>"111000001",
  33099=>"001001000",
  33100=>"000001000",
  33101=>"000000000",
  33102=>"111111010",
  33103=>"000000110",
  33104=>"000000000",
  33105=>"001001001",
  33106=>"000100000",
  33107=>"000000000",
  33108=>"000000000",
  33109=>"011011011",
  33110=>"000000111",
  33111=>"111111001",
  33112=>"100000100",
  33113=>"000111111",
  33114=>"000110000",
  33115=>"111111111",
  33116=>"101111111",
  33117=>"000000000",
  33118=>"111111011",
  33119=>"110111010",
  33120=>"000000000",
  33121=>"000001000",
  33122=>"000000000",
  33123=>"000000000",
  33124=>"000000000",
  33125=>"000000111",
  33126=>"110111100",
  33127=>"011111111",
  33128=>"111000000",
  33129=>"110111111",
  33130=>"000010000",
  33131=>"111111111",
  33132=>"001001001",
  33133=>"111111000",
  33134=>"110100101",
  33135=>"000000000",
  33136=>"001101000",
  33137=>"111111111",
  33138=>"000000001",
  33139=>"001000000",
  33140=>"111111110",
  33141=>"101110110",
  33142=>"111011000",
  33143=>"000000000",
  33144=>"000000000",
  33145=>"000011000",
  33146=>"111001001",
  33147=>"100110111",
  33148=>"111111111",
  33149=>"111111111",
  33150=>"111111111",
  33151=>"101111111",
  33152=>"110110110",
  33153=>"011000000",
  33154=>"000011001",
  33155=>"111111111",
  33156=>"100100000",
  33157=>"000000000",
  33158=>"111000110",
  33159=>"000101111",
  33160=>"110111110",
  33161=>"111111111",
  33162=>"100010000",
  33163=>"000000000",
  33164=>"111111111",
  33165=>"011011110",
  33166=>"001011110",
  33167=>"111111111",
  33168=>"000001000",
  33169=>"111101111",
  33170=>"001100110",
  33171=>"000000000",
  33172=>"110111110",
  33173=>"000000110",
  33174=>"000000000",
  33175=>"000011111",
  33176=>"000000000",
  33177=>"111001100",
  33178=>"111111111",
  33179=>"000000000",
  33180=>"001011110",
  33181=>"000011000",
  33182=>"111001000",
  33183=>"011000001",
  33184=>"111111111",
  33185=>"011010000",
  33186=>"111111100",
  33187=>"111111000",
  33188=>"011111110",
  33189=>"000000000",
  33190=>"000000000",
  33191=>"000000000",
  33192=>"000011111",
  33193=>"000000000",
  33194=>"111111000",
  33195=>"001000011",
  33196=>"000000000",
  33197=>"000000001",
  33198=>"110111101",
  33199=>"000111011",
  33200=>"111111111",
  33201=>"111111111",
  33202=>"111101000",
  33203=>"000111111",
  33204=>"000000111",
  33205=>"100110110",
  33206=>"111111110",
  33207=>"001011111",
  33208=>"000111111",
  33209=>"111111101",
  33210=>"000000000",
  33211=>"000000000",
  33212=>"000000000",
  33213=>"001101111",
  33214=>"111110000",
  33215=>"010000000",
  33216=>"001000000",
  33217=>"111111000",
  33218=>"000000000",
  33219=>"111111111",
  33220=>"001100111",
  33221=>"110100100",
  33222=>"000011111",
  33223=>"001000000",
  33224=>"001011111",
  33225=>"110110110",
  33226=>"000000110",
  33227=>"000000000",
  33228=>"000000010",
  33229=>"111111000",
  33230=>"011100100",
  33231=>"111011010",
  33232=>"011001111",
  33233=>"000000001",
  33234=>"000000000",
  33235=>"111111111",
  33236=>"000000000",
  33237=>"111111111",
  33238=>"011011010",
  33239=>"101100110",
  33240=>"111011111",
  33241=>"111000000",
  33242=>"110111111",
  33243=>"000000000",
  33244=>"000000000",
  33245=>"111101100",
  33246=>"011011011",
  33247=>"111111110",
  33248=>"111111111",
  33249=>"111000000",
  33250=>"000000000",
  33251=>"111111000",
  33252=>"001001000",
  33253=>"111111111",
  33254=>"100000111",
  33255=>"111111111",
  33256=>"101101111",
  33257=>"000011100",
  33258=>"011001100",
  33259=>"000001011",
  33260=>"111100000",
  33261=>"001111111",
  33262=>"110110010",
  33263=>"111111111",
  33264=>"111101001",
  33265=>"111111111",
  33266=>"111111111",
  33267=>"111111000",
  33268=>"000000000",
  33269=>"110000010",
  33270=>"000000000",
  33271=>"111110000",
  33272=>"010010000",
  33273=>"000000010",
  33274=>"101000000",
  33275=>"000000000",
  33276=>"001111111",
  33277=>"111010110",
  33278=>"111111111",
  33279=>"111111111",
  33280=>"110111100",
  33281=>"111111111",
  33282=>"000111111",
  33283=>"100100111",
  33284=>"100100001",
  33285=>"000000000",
  33286=>"111111110",
  33287=>"000000000",
  33288=>"111110000",
  33289=>"000111001",
  33290=>"111111110",
  33291=>"111111111",
  33292=>"000110110",
  33293=>"111111001",
  33294=>"111111011",
  33295=>"000000000",
  33296=>"111111001",
  33297=>"111111111",
  33298=>"001100000",
  33299=>"000000111",
  33300=>"101011111",
  33301=>"111111000",
  33302=>"111111101",
  33303=>"000000111",
  33304=>"000100111",
  33305=>"100000000",
  33306=>"000000000",
  33307=>"110110100",
  33308=>"111111111",
  33309=>"111000111",
  33310=>"100100100",
  33311=>"000001000",
  33312=>"000000000",
  33313=>"000000000",
  33314=>"000000000",
  33315=>"011111000",
  33316=>"000000111",
  33317=>"111111110",
  33318=>"001111111",
  33319=>"111111111",
  33320=>"000000000",
  33321=>"000000000",
  33322=>"000000000",
  33323=>"111111111",
  33324=>"110011111",
  33325=>"000111111",
  33326=>"000001111",
  33327=>"000000000",
  33328=>"100011001",
  33329=>"010110000",
  33330=>"101111101",
  33331=>"101000000",
  33332=>"100110000",
  33333=>"000000000",
  33334=>"110111111",
  33335=>"110101101",
  33336=>"000000000",
  33337=>"101000100",
  33338=>"010011000",
  33339=>"111000001",
  33340=>"111111101",
  33341=>"001110111",
  33342=>"001000001",
  33343=>"000000001",
  33344=>"111011001",
  33345=>"111000000",
  33346=>"011011111",
  33347=>"000000000",
  33348=>"110100100",
  33349=>"000000000",
  33350=>"101111111",
  33351=>"001011111",
  33352=>"111111111",
  33353=>"111001000",
  33354=>"110110111",
  33355=>"101000000",
  33356=>"011111111",
  33357=>"000000000",
  33358=>"000000000",
  33359=>"010000000",
  33360=>"000000000",
  33361=>"101001001",
  33362=>"111001000",
  33363=>"111111110",
  33364=>"111111111",
  33365=>"000000000",
  33366=>"000000011",
  33367=>"111111111",
  33368=>"000000000",
  33369=>"101001111",
  33370=>"100111000",
  33371=>"000001001",
  33372=>"000111011",
  33373=>"111101111",
  33374=>"111111111",
  33375=>"110111111",
  33376=>"111111111",
  33377=>"100100100",
  33378=>"000001001",
  33379=>"000000000",
  33380=>"111111000",
  33381=>"101100000",
  33382=>"111111000",
  33383=>"100000111",
  33384=>"011011001",
  33385=>"000000000",
  33386=>"000000001",
  33387=>"111001000",
  33388=>"000100100",
  33389=>"000000000",
  33390=>"111101111",
  33391=>"000000000",
  33392=>"000000001",
  33393=>"000000101",
  33394=>"111001001",
  33395=>"000110101",
  33396=>"000000000",
  33397=>"011011111",
  33398=>"111000000",
  33399=>"000010111",
  33400=>"111111111",
  33401=>"000100100",
  33402=>"101111111",
  33403=>"101000001",
  33404=>"110110110",
  33405=>"000000000",
  33406=>"110100100",
  33407=>"000011111",
  33408=>"000000000",
  33409=>"000000000",
  33410=>"010110111",
  33411=>"000100011",
  33412=>"000000001",
  33413=>"011000000",
  33414=>"111111111",
  33415=>"010111111",
  33416=>"000000000",
  33417=>"100000100",
  33418=>"000000000",
  33419=>"111111111",
  33420=>"101101100",
  33421=>"100111111",
  33422=>"001000000",
  33423=>"111111111",
  33424=>"001000000",
  33425=>"000111111",
  33426=>"111111111",
  33427=>"110110110",
  33428=>"000000110",
  33429=>"000000110",
  33430=>"000000000",
  33431=>"000000000",
  33432=>"000000111",
  33433=>"110111000",
  33434=>"000000000",
  33435=>"111111111",
  33436=>"000010011",
  33437=>"110000000",
  33438=>"001111000",
  33439=>"000000100",
  33440=>"000000000",
  33441=>"111111110",
  33442=>"111111111",
  33443=>"000000000",
  33444=>"100111100",
  33445=>"111111111",
  33446=>"000000001",
  33447=>"100000011",
  33448=>"000000000",
  33449=>"111111111",
  33450=>"000000000",
  33451=>"111111111",
  33452=>"111111111",
  33453=>"000000000",
  33454=>"000000000",
  33455=>"010111111",
  33456=>"011111000",
  33457=>"011011011",
  33458=>"111111111",
  33459=>"000001111",
  33460=>"100110110",
  33461=>"110010000",
  33462=>"000010011",
  33463=>"111101000",
  33464=>"111111011",
  33465=>"111111111",
  33466=>"000000110",
  33467=>"001011111",
  33468=>"111001111",
  33469=>"000000000",
  33470=>"000000000",
  33471=>"111111111",
  33472=>"000000000",
  33473=>"111000000",
  33474=>"000000111",
  33475=>"000000000",
  33476=>"110110000",
  33477=>"111111111",
  33478=>"100100000",
  33479=>"010010000",
  33480=>"000000000",
  33481=>"111111111",
  33482=>"111111001",
  33483=>"100111100",
  33484=>"111111011",
  33485=>"110000000",
  33486=>"000110111",
  33487=>"000000111",
  33488=>"011001000",
  33489=>"000000000",
  33490=>"001000000",
  33491=>"000100111",
  33492=>"100100000",
  33493=>"000100000",
  33494=>"000000010",
  33495=>"000000001",
  33496=>"010110110",
  33497=>"111010000",
  33498=>"111111110",
  33499=>"111000010",
  33500=>"000000000",
  33501=>"101011111",
  33502=>"110110000",
  33503=>"000000000",
  33504=>"101101001",
  33505=>"000001111",
  33506=>"101011011",
  33507=>"111111010",
  33508=>"000000000",
  33509=>"000000000",
  33510=>"111111111",
  33511=>"111111101",
  33512=>"111111111",
  33513=>"010111111",
  33514=>"000000000",
  33515=>"100000100",
  33516=>"000000111",
  33517=>"000000111",
  33518=>"000000001",
  33519=>"110101101",
  33520=>"001101101",
  33521=>"000000000",
  33522=>"000000000",
  33523=>"000110000",
  33524=>"000000000",
  33525=>"111111111",
  33526=>"111111110",
  33527=>"111001111",
  33528=>"000000000",
  33529=>"000000111",
  33530=>"000000000",
  33531=>"000000000",
  33532=>"001000000",
  33533=>"001111011",
  33534=>"101100111",
  33535=>"000000000",
  33536=>"110110000",
  33537=>"101000101",
  33538=>"000001011",
  33539=>"000000000",
  33540=>"000000000",
  33541=>"000000000",
  33542=>"111110000",
  33543=>"111011001",
  33544=>"100000000",
  33545=>"000100111",
  33546=>"000000000",
  33547=>"111111001",
  33548=>"000000000",
  33549=>"000000000",
  33550=>"111000000",
  33551=>"001001011",
  33552=>"111101101",
  33553=>"000000000",
  33554=>"101000111",
  33555=>"111111111",
  33556=>"000000000",
  33557=>"001000100",
  33558=>"001000100",
  33559=>"000111111",
  33560=>"001011111",
  33561=>"000000001",
  33562=>"111111111",
  33563=>"001000000",
  33564=>"110111110",
  33565=>"110000000",
  33566=>"000000000",
  33567=>"111111111",
  33568=>"001011011",
  33569=>"111111111",
  33570=>"000000000",
  33571=>"111111110",
  33572=>"001000010",
  33573=>"000000000",
  33574=>"000000000",
  33575=>"110000101",
  33576=>"111111111",
  33577=>"111010011",
  33578=>"001111111",
  33579=>"111111101",
  33580=>"110110010",
  33581=>"111111111",
  33582=>"101111001",
  33583=>"100000111",
  33584=>"111111111",
  33585=>"110111100",
  33586=>"000000001",
  33587=>"000100111",
  33588=>"111001000",
  33589=>"010111111",
  33590=>"011000000",
  33591=>"011011011",
  33592=>"000010000",
  33593=>"000000000",
  33594=>"101001011",
  33595=>"110000010",
  33596=>"100110111",
  33597=>"111111010",
  33598=>"000001111",
  33599=>"111111111",
  33600=>"000011110",
  33601=>"000000000",
  33602=>"000000000",
  33603=>"000000001",
  33604=>"101011000",
  33605=>"000000000",
  33606=>"010111111",
  33607=>"110111111",
  33608=>"100000000",
  33609=>"011000000",
  33610=>"000000000",
  33611=>"011101111",
  33612=>"000111000",
  33613=>"000000001",
  33614=>"111110111",
  33615=>"011011011",
  33616=>"001001111",
  33617=>"001111111",
  33618=>"101111110",
  33619=>"110000000",
  33620=>"000100111",
  33621=>"001001011",
  33622=>"000000001",
  33623=>"001000000",
  33624=>"000000000",
  33625=>"101111111",
  33626=>"111111111",
  33627=>"000000000",
  33628=>"111111000",
  33629=>"001000000",
  33630=>"100111111",
  33631=>"110000000",
  33632=>"000000010",
  33633=>"111000000",
  33634=>"111011111",
  33635=>"111101111",
  33636=>"001011001",
  33637=>"000000100",
  33638=>"000000011",
  33639=>"111110110",
  33640=>"110101100",
  33641=>"000011011",
  33642=>"001000111",
  33643=>"000010000",
  33644=>"100000000",
  33645=>"000000000",
  33646=>"000000111",
  33647=>"100010000",
  33648=>"000000000",
  33649=>"000001011",
  33650=>"000011000",
  33651=>"111111011",
  33652=>"111111111",
  33653=>"000000000",
  33654=>"111111111",
  33655=>"000000000",
  33656=>"000000000",
  33657=>"100000000",
  33658=>"000000000",
  33659=>"011111111",
  33660=>"000001101",
  33661=>"000000000",
  33662=>"101101111",
  33663=>"000000000",
  33664=>"000001100",
  33665=>"000000000",
  33666=>"001000000",
  33667=>"101000000",
  33668=>"000000010",
  33669=>"001111000",
  33670=>"111100101",
  33671=>"011011111",
  33672=>"001101101",
  33673=>"101100111",
  33674=>"100100100",
  33675=>"000100111",
  33676=>"000000000",
  33677=>"100000000",
  33678=>"000001101",
  33679=>"000000101",
  33680=>"000000000",
  33681=>"111111111",
  33682=>"111111111",
  33683=>"011011001",
  33684=>"001001001",
  33685=>"000010010",
  33686=>"000000000",
  33687=>"000000100",
  33688=>"111111001",
  33689=>"100110111",
  33690=>"000010000",
  33691=>"111000011",
  33692=>"000000000",
  33693=>"111111111",
  33694=>"100000001",
  33695=>"000000111",
  33696=>"000100110",
  33697=>"111111111",
  33698=>"111111111",
  33699=>"000000011",
  33700=>"111111110",
  33701=>"000000000",
  33702=>"111111111",
  33703=>"111111111",
  33704=>"000000000",
  33705=>"011000000",
  33706=>"100100000",
  33707=>"111111000",
  33708=>"000000000",
  33709=>"110001000",
  33710=>"100001000",
  33711=>"000001111",
  33712=>"111100100",
  33713=>"000111111",
  33714=>"000000001",
  33715=>"000000000",
  33716=>"111011001",
  33717=>"000000000",
  33718=>"100100100",
  33719=>"000000101",
  33720=>"000000000",
  33721=>"000000000",
  33722=>"000010000",
  33723=>"111111111",
  33724=>"010001111",
  33725=>"111000100",
  33726=>"000000111",
  33727=>"101101110",
  33728=>"000000100",
  33729=>"000000100",
  33730=>"000000011",
  33731=>"111111111",
  33732=>"100010001",
  33733=>"111111000",
  33734=>"001000000",
  33735=>"111111111",
  33736=>"000000000",
  33737=>"000010111",
  33738=>"001000000",
  33739=>"000000000",
  33740=>"110111111",
  33741=>"100111111",
  33742=>"111111000",
  33743=>"000000000",
  33744=>"111000000",
  33745=>"000000000",
  33746=>"000000000",
  33747=>"110000011",
  33748=>"100110111",
  33749=>"000000000",
  33750=>"000111111",
  33751=>"000011011",
  33752=>"101100000",
  33753=>"011111000",
  33754=>"111111111",
  33755=>"000000110",
  33756=>"110110111",
  33757=>"000000000",
  33758=>"111110010",
  33759=>"100101011",
  33760=>"000111111",
  33761=>"001000100",
  33762=>"000000000",
  33763=>"100111111",
  33764=>"000001101",
  33765=>"101001000",
  33766=>"011000000",
  33767=>"110111111",
  33768=>"111111111",
  33769=>"000000000",
  33770=>"000000111",
  33771=>"000000000",
  33772=>"000000000",
  33773=>"000000000",
  33774=>"111111111",
  33775=>"001000000",
  33776=>"000001011",
  33777=>"000000101",
  33778=>"011001001",
  33779=>"001110110",
  33780=>"111111111",
  33781=>"000101000",
  33782=>"101101111",
  33783=>"111111000",
  33784=>"111111111",
  33785=>"001000001",
  33786=>"000000000",
  33787=>"011010000",
  33788=>"111101111",
  33789=>"101101111",
  33790=>"111111111",
  33791=>"111111111",
  33792=>"011011100",
  33793=>"000000000",
  33794=>"100101100",
  33795=>"100110100",
  33796=>"111111111",
  33797=>"011001001",
  33798=>"100000000",
  33799=>"000000000",
  33800=>"111111111",
  33801=>"000010110",
  33802=>"111111111",
  33803=>"000011111",
  33804=>"001000000",
  33805=>"001001001",
  33806=>"000000000",
  33807=>"111111001",
  33808=>"111101111",
  33809=>"111000000",
  33810=>"101000000",
  33811=>"011001001",
  33812=>"000000000",
  33813=>"111100000",
  33814=>"000111100",
  33815=>"111111011",
  33816=>"111101111",
  33817=>"111111110",
  33818=>"111000000",
  33819=>"000001001",
  33820=>"010111011",
  33821=>"011010111",
  33822=>"011011000",
  33823=>"101111111",
  33824=>"110100101",
  33825=>"111111111",
  33826=>"000000000",
  33827=>"000000011",
  33828=>"111111111",
  33829=>"111111000",
  33830=>"111111111",
  33831=>"000010000",
  33832=>"000000000",
  33833=>"000000000",
  33834=>"011011011",
  33835=>"000000111",
  33836=>"111111111",
  33837=>"001111111",
  33838=>"000000110",
  33839=>"000000000",
  33840=>"110100000",
  33841=>"000000000",
  33842=>"011011011",
  33843=>"010100100",
  33844=>"100100110",
  33845=>"001011011",
  33846=>"111111111",
  33847=>"011000000",
  33848=>"111111111",
  33849=>"010000000",
  33850=>"000000000",
  33851=>"000000011",
  33852=>"000000110",
  33853=>"111111111",
  33854=>"111100001",
  33855=>"000001001",
  33856=>"111011001",
  33857=>"000000000",
  33858=>"111001000",
  33859=>"000100100",
  33860=>"000000001",
  33861=>"100000000",
  33862=>"000110000",
  33863=>"100000000",
  33864=>"111011111",
  33865=>"000000000",
  33866=>"001000000",
  33867=>"111111111",
  33868=>"000111111",
  33869=>"111000100",
  33870=>"000000000",
  33871=>"000111111",
  33872=>"111010011",
  33873=>"010010000",
  33874=>"000000000",
  33875=>"011011001",
  33876=>"111111111",
  33877=>"111011010",
  33878=>"000000000",
  33879=>"011011011",
  33880=>"011010110",
  33881=>"000000000",
  33882=>"000000111",
  33883=>"111111011",
  33884=>"110111111",
  33885=>"101100000",
  33886=>"111001111",
  33887=>"111111110",
  33888=>"000000000",
  33889=>"000011111",
  33890=>"110110111",
  33891=>"000000000",
  33892=>"000011100",
  33893=>"001000000",
  33894=>"011001111",
  33895=>"000000000",
  33896=>"010111111",
  33897=>"100101101",
  33898=>"111110110",
  33899=>"110111111",
  33900=>"001000000",
  33901=>"000000000",
  33902=>"001000000",
  33903=>"000000000",
  33904=>"111111111",
  33905=>"000001110",
  33906=>"101001000",
  33907=>"111111111",
  33908=>"100100110",
  33909=>"111000100",
  33910=>"000000000",
  33911=>"000000000",
  33912=>"111111111",
  33913=>"000110111",
  33914=>"000000001",
  33915=>"111111111",
  33916=>"001000000",
  33917=>"000000111",
  33918=>"100000001",
  33919=>"000000001",
  33920=>"000000101",
  33921=>"111111000",
  33922=>"000000111",
  33923=>"111111111",
  33924=>"000000000",
  33925=>"111001000",
  33926=>"000000000",
  33927=>"101111001",
  33928=>"000000000",
  33929=>"110000110",
  33930=>"111111000",
  33931=>"011111011",
  33932=>"010000101",
  33933=>"000000100",
  33934=>"111000000",
  33935=>"000000100",
  33936=>"000000010",
  33937=>"111101111",
  33938=>"000111111",
  33939=>"100111111",
  33940=>"001000000",
  33941=>"111011000",
  33942=>"111111111",
  33943=>"000000000",
  33944=>"001001111",
  33945=>"111111111",
  33946=>"000000000",
  33947=>"000000000",
  33948=>"001000000",
  33949=>"101101100",
  33950=>"111100110",
  33951=>"000000001",
  33952=>"011011011",
  33953=>"000011111",
  33954=>"100000000",
  33955=>"111111111",
  33956=>"000000000",
  33957=>"111111110",
  33958=>"111111111",
  33959=>"100000010",
  33960=>"000111111",
  33961=>"000100001",
  33962=>"111111011",
  33963=>"001111111",
  33964=>"000100111",
  33965=>"011100001",
  33966=>"111011000",
  33967=>"011000000",
  33968=>"000111111",
  33969=>"111111111",
  33970=>"111111111",
  33971=>"000000000",
  33972=>"000000000",
  33973=>"111111100",
  33974=>"101001000",
  33975=>"110111111",
  33976=>"110111111",
  33977=>"000000000",
  33978=>"000000000",
  33979=>"001111111",
  33980=>"000000000",
  33981=>"111111110",
  33982=>"010111111",
  33983=>"100101001",
  33984=>"111111111",
  33985=>"111000001",
  33986=>"000000000",
  33987=>"000000111",
  33988=>"100111000",
  33989=>"010000000",
  33990=>"000001111",
  33991=>"111101111",
  33992=>"111100110",
  33993=>"011001000",
  33994=>"001001001",
  33995=>"001011011",
  33996=>"010110111",
  33997=>"000100001",
  33998=>"111111111",
  33999=>"110111111",
  34000=>"100100111",
  34001=>"000000000",
  34002=>"000000000",
  34003=>"000000000",
  34004=>"000000000",
  34005=>"111011001",
  34006=>"000000000",
  34007=>"000000000",
  34008=>"111111000",
  34009=>"111111111",
  34010=>"000000000",
  34011=>"111110010",
  34012=>"111101111",
  34013=>"000000000",
  34014=>"110111111",
  34015=>"001001000",
  34016=>"000000000",
  34017=>"000000000",
  34018=>"111111111",
  34019=>"111111111",
  34020=>"111111111",
  34021=>"111111110",
  34022=>"101000000",
  34023=>"000000000",
  34024=>"000000000",
  34025=>"000000000",
  34026=>"001000101",
  34027=>"111001000",
  34028=>"001001011",
  34029=>"011111111",
  34030=>"001111111",
  34031=>"111111111",
  34032=>"111111111",
  34033=>"011001000",
  34034=>"111111111",
  34035=>"000000111",
  34036=>"000110111",
  34037=>"111111011",
  34038=>"111110110",
  34039=>"110110000",
  34040=>"000000000",
  34041=>"111111111",
  34042=>"111111111",
  34043=>"000101111",
  34044=>"111111111",
  34045=>"010000110",
  34046=>"000000000",
  34047=>"111101101",
  34048=>"000010011",
  34049=>"000000001",
  34050=>"110100100",
  34051=>"000000000",
  34052=>"111111111",
  34053=>"011010000",
  34054=>"000000110",
  34055=>"001001001",
  34056=>"111111111",
  34057=>"000000000",
  34058=>"111111111",
  34059=>"100000111",
  34060=>"000000000",
  34061=>"100101101",
  34062=>"111111011",
  34063=>"011001111",
  34064=>"110111111",
  34065=>"000001100",
  34066=>"000000100",
  34067=>"000000101",
  34068=>"111111000",
  34069=>"111000000",
  34070=>"111111111",
  34071=>"111111111",
  34072=>"011111101",
  34073=>"011011110",
  34074=>"000000100",
  34075=>"111000111",
  34076=>"000000110",
  34077=>"000000000",
  34078=>"100000000",
  34079=>"111111111",
  34080=>"111101111",
  34081=>"000000110",
  34082=>"011111111",
  34083=>"100100001",
  34084=>"001001100",
  34085=>"000010000",
  34086=>"111111111",
  34087=>"000000000",
  34088=>"001000000",
  34089=>"011011111",
  34090=>"000111100",
  34091=>"000110110",
  34092=>"111011001",
  34093=>"100100110",
  34094=>"111111000",
  34095=>"000000000",
  34096=>"011011011",
  34097=>"111001000",
  34098=>"111111111",
  34099=>"100000111",
  34100=>"110001000",
  34101=>"000001111",
  34102=>"000000000",
  34103=>"000000000",
  34104=>"011000111",
  34105=>"000000000",
  34106=>"000001111",
  34107=>"011111000",
  34108=>"000000000",
  34109=>"010000000",
  34110=>"000000011",
  34111=>"000000001",
  34112=>"000000110",
  34113=>"000000001",
  34114=>"111111111",
  34115=>"000111111",
  34116=>"100111111",
  34117=>"000011000",
  34118=>"111111111",
  34119=>"111011000",
  34120=>"111111111",
  34121=>"000000000",
  34122=>"000000000",
  34123=>"111111111",
  34124=>"000000100",
  34125=>"100110111",
  34126=>"011000000",
  34127=>"001000000",
  34128=>"000010110",
  34129=>"000000111",
  34130=>"001000111",
  34131=>"000000000",
  34132=>"111011011",
  34133=>"000000001",
  34134=>"111111100",
  34135=>"001001001",
  34136=>"010000000",
  34137=>"111111011",
  34138=>"111001001",
  34139=>"011011100",
  34140=>"000100110",
  34141=>"111111101",
  34142=>"001000000",
  34143=>"111111111",
  34144=>"111111101",
  34145=>"111111111",
  34146=>"000100000",
  34147=>"000000001",
  34148=>"010110000",
  34149=>"000100111",
  34150=>"000000000",
  34151=>"000000111",
  34152=>"111111001",
  34153=>"110000000",
  34154=>"000000111",
  34155=>"000000111",
  34156=>"111011011",
  34157=>"000111111",
  34158=>"000111111",
  34159=>"001001000",
  34160=>"100111101",
  34161=>"110000100",
  34162=>"110111011",
  34163=>"001000000",
  34164=>"111111110",
  34165=>"000000000",
  34166=>"000000000",
  34167=>"000000000",
  34168=>"111111111",
  34169=>"000000000",
  34170=>"010011111",
  34171=>"000000000",
  34172=>"000000111",
  34173=>"000000000",
  34174=>"000000000",
  34175=>"000011011",
  34176=>"000000000",
  34177=>"100000111",
  34178=>"000000000",
  34179=>"111111011",
  34180=>"011000000",
  34181=>"000000111",
  34182=>"000000100",
  34183=>"111000000",
  34184=>"000111111",
  34185=>"000111111",
  34186=>"111001001",
  34187=>"111111000",
  34188=>"000001011",
  34189=>"000010000",
  34190=>"111110000",
  34191=>"011001011",
  34192=>"000100100",
  34193=>"100000110",
  34194=>"111111111",
  34195=>"000000000",
  34196=>"000001111",
  34197=>"100000000",
  34198=>"010000010",
  34199=>"001000111",
  34200=>"000000110",
  34201=>"100000101",
  34202=>"000100111",
  34203=>"110110000",
  34204=>"000000000",
  34205=>"111010111",
  34206=>"001011111",
  34207=>"000000000",
  34208=>"111111111",
  34209=>"001011011",
  34210=>"001111011",
  34211=>"000111101",
  34212=>"011011000",
  34213=>"100001001",
  34214=>"111111010",
  34215=>"011111111",
  34216=>"110000000",
  34217=>"010000000",
  34218=>"111111010",
  34219=>"000000000",
  34220=>"111111110",
  34221=>"001010111",
  34222=>"000100110",
  34223=>"010000001",
  34224=>"000000011",
  34225=>"000111111",
  34226=>"111100100",
  34227=>"000000000",
  34228=>"111111010",
  34229=>"100000000",
  34230=>"110000001",
  34231=>"011111001",
  34232=>"111010110",
  34233=>"111111111",
  34234=>"111101111",
  34235=>"001011101",
  34236=>"011111111",
  34237=>"111111111",
  34238=>"001001000",
  34239=>"000000000",
  34240=>"001000110",
  34241=>"110000011",
  34242=>"000000010",
  34243=>"111010000",
  34244=>"111001000",
  34245=>"000100110",
  34246=>"000000000",
  34247=>"000000000",
  34248=>"111011100",
  34249=>"111111000",
  34250=>"000000000",
  34251=>"000000100",
  34252=>"001101111",
  34253=>"000000110",
  34254=>"000100001",
  34255=>"100100100",
  34256=>"000000000",
  34257=>"000000111",
  34258=>"001101111",
  34259=>"111111111",
  34260=>"000000001",
  34261=>"111110111",
  34262=>"111100100",
  34263=>"110000000",
  34264=>"010111001",
  34265=>"111000111",
  34266=>"111000001",
  34267=>"011011111",
  34268=>"010011011",
  34269=>"011111011",
  34270=>"111111100",
  34271=>"000010000",
  34272=>"110110000",
  34273=>"111100111",
  34274=>"111111111",
  34275=>"000000111",
  34276=>"111101100",
  34277=>"000000100",
  34278=>"000100100",
  34279=>"000000000",
  34280=>"110100100",
  34281=>"111111111",
  34282=>"000011111",
  34283=>"000000000",
  34284=>"111011000",
  34285=>"111101111",
  34286=>"000111111",
  34287=>"101000100",
  34288=>"000000100",
  34289=>"001001111",
  34290=>"111001011",
  34291=>"000001011",
  34292=>"000011010",
  34293=>"111001000",
  34294=>"010000000",
  34295=>"000000110",
  34296=>"000000110",
  34297=>"010010000",
  34298=>"111000000",
  34299=>"111111111",
  34300=>"101111100",
  34301=>"111111111",
  34302=>"111111111",
  34303=>"000000000",
  34304=>"111111110",
  34305=>"011001000",
  34306=>"001001001",
  34307=>"000000000",
  34308=>"111111001",
  34309=>"000000000",
  34310=>"001011001",
  34311=>"111111111",
  34312=>"101101001",
  34313=>"000000110",
  34314=>"000000000",
  34315=>"000000000",
  34316=>"010111111",
  34317=>"100000100",
  34318=>"001001101",
  34319=>"001000000",
  34320=>"010110000",
  34321=>"000000000",
  34322=>"111011000",
  34323=>"000000000",
  34324=>"111111100",
  34325=>"010111111",
  34326=>"000000000",
  34327=>"000000100",
  34328=>"111100111",
  34329=>"111111000",
  34330=>"110000000",
  34331=>"001000100",
  34332=>"001000001",
  34333=>"010000000",
  34334=>"111111101",
  34335=>"001111111",
  34336=>"111101000",
  34337=>"111111111",
  34338=>"000100000",
  34339=>"000011011",
  34340=>"000000001",
  34341=>"000000000",
  34342=>"000000000",
  34343=>"110111111",
  34344=>"000111111",
  34345=>"000000000",
  34346=>"000100100",
  34347=>"100111111",
  34348=>"100101000",
  34349=>"001000000",
  34350=>"111011011",
  34351=>"100101111",
  34352=>"101000101",
  34353=>"111111111",
  34354=>"011111111",
  34355=>"000010111",
  34356=>"111010000",
  34357=>"111111110",
  34358=>"000000000",
  34359=>"011000000",
  34360=>"000000000",
  34361=>"110111000",
  34362=>"000110111",
  34363=>"111001000",
  34364=>"111110110",
  34365=>"111111000",
  34366=>"111111111",
  34367=>"100111111",
  34368=>"001000000",
  34369=>"010011011",
  34370=>"000000111",
  34371=>"110111100",
  34372=>"000100000",
  34373=>"001001111",
  34374=>"110010000",
  34375=>"000000000",
  34376=>"110111011",
  34377=>"111111111",
  34378=>"011111111",
  34379=>"111111100",
  34380=>"111001100",
  34381=>"101000100",
  34382=>"011000111",
  34383=>"100000100",
  34384=>"110111111",
  34385=>"000000010",
  34386=>"100100100",
  34387=>"110111110",
  34388=>"001001101",
  34389=>"000101101",
  34390=>"110111000",
  34391=>"101101111",
  34392=>"111111011",
  34393=>"100100100",
  34394=>"110100000",
  34395=>"111111101",
  34396=>"001000000",
  34397=>"111111011",
  34398=>"011111101",
  34399=>"111111111",
  34400=>"110000010",
  34401=>"000000100",
  34402=>"111001111",
  34403=>"100000000",
  34404=>"100000000",
  34405=>"111111101",
  34406=>"010010110",
  34407=>"111110110",
  34408=>"000000000",
  34409=>"000000000",
  34410=>"000011011",
  34411=>"000000011",
  34412=>"110000000",
  34413=>"010010000",
  34414=>"111111111",
  34415=>"000111111",
  34416=>"100000000",
  34417=>"101001111",
  34418=>"000000000",
  34419=>"011111110",
  34420=>"100000000",
  34421=>"011000110",
  34422=>"100000000",
  34423=>"101111011",
  34424=>"111111111",
  34425=>"100100011",
  34426=>"111111011",
  34427=>"100101100",
  34428=>"100000000",
  34429=>"000011011",
  34430=>"001000000",
  34431=>"100100100",
  34432=>"000000111",
  34433=>"111100111",
  34434=>"000000000",
  34435=>"111011111",
  34436=>"000000000",
  34437=>"111111011",
  34438=>"011111101",
  34439=>"000000100",
  34440=>"111111010",
  34441=>"000001001",
  34442=>"001111111",
  34443=>"000000000",
  34444=>"000011011",
  34445=>"110111111",
  34446=>"000001000",
  34447=>"110111111",
  34448=>"111111111",
  34449=>"111000000",
  34450=>"111100100",
  34451=>"111100110",
  34452=>"111011111",
  34453=>"111111111",
  34454=>"001011011",
  34455=>"100000000",
  34456=>"000000000",
  34457=>"111111001",
  34458=>"111111000",
  34459=>"001000001",
  34460=>"111000000",
  34461=>"000000000",
  34462=>"000000001",
  34463=>"000000000",
  34464=>"111111110",
  34465=>"110011000",
  34466=>"000010111",
  34467=>"000000000",
  34468=>"111111110",
  34469=>"011111111",
  34470=>"111111111",
  34471=>"111110111",
  34472=>"111111101",
  34473=>"110000110",
  34474=>"000111111",
  34475=>"111011111",
  34476=>"000100000",
  34477=>"000100101",
  34478=>"111101111",
  34479=>"111111100",
  34480=>"000000000",
  34481=>"101100110",
  34482=>"000000000",
  34483=>"010010111",
  34484=>"000110110",
  34485=>"010111100",
  34486=>"100100101",
  34487=>"111111111",
  34488=>"000000000",
  34489=>"110111111",
  34490=>"101001001",
  34491=>"111000100",
  34492=>"000101111",
  34493=>"111111111",
  34494=>"000000000",
  34495=>"011111111",
  34496=>"111000000",
  34497=>"000000010",
  34498=>"000110011",
  34499=>"000000000",
  34500=>"000000001",
  34501=>"000000000",
  34502=>"000000000",
  34503=>"100100100",
  34504=>"011011000",
  34505=>"000110101",
  34506=>"000000100",
  34507=>"111111111",
  34508=>"111101000",
  34509=>"001000000",
  34510=>"000000100",
  34511=>"111001011",
  34512=>"011000000",
  34513=>"001001000",
  34514=>"011000000",
  34515=>"100100100",
  34516=>"111111111",
  34517=>"001111110",
  34518=>"111001011",
  34519=>"111000100",
  34520=>"000000000",
  34521=>"000000000",
  34522=>"110111111",
  34523=>"111101001",
  34524=>"111111111",
  34525=>"111111111",
  34526=>"111111111",
  34527=>"111110000",
  34528=>"000000000",
  34529=>"000000001",
  34530=>"000100111",
  34531=>"111111001",
  34532=>"111111101",
  34533=>"000110110",
  34534=>"001101101",
  34535=>"110100000",
  34536=>"001011000",
  34537=>"000000000",
  34538=>"000010110",
  34539=>"000000000",
  34540=>"111111000",
  34541=>"111000000",
  34542=>"111111111",
  34543=>"111111111",
  34544=>"111111111",
  34545=>"111111111",
  34546=>"100111111",
  34547=>"000000000",
  34548=>"111111000",
  34549=>"000100111",
  34550=>"011000110",
  34551=>"011111000",
  34552=>"111000100",
  34553=>"100100100",
  34554=>"000111111",
  34555=>"011000001",
  34556=>"110110111",
  34557=>"100000101",
  34558=>"111111000",
  34559=>"110110000",
  34560=>"000111111",
  34561=>"100000100",
  34562=>"110111111",
  34563=>"111111111",
  34564=>"111111111",
  34565=>"000000000",
  34566=>"000001111",
  34567=>"111111110",
  34568=>"000000100",
  34569=>"000000001",
  34570=>"000000100",
  34571=>"111011011",
  34572=>"100000000",
  34573=>"101111000",
  34574=>"000000101",
  34575=>"000000110",
  34576=>"111111100",
  34577=>"000101111",
  34578=>"110110111",
  34579=>"000000011",
  34580=>"000000000",
  34581=>"000000000",
  34582=>"001001101",
  34583=>"000000000",
  34584=>"010010000",
  34585=>"111111111",
  34586=>"100000100",
  34587=>"000010110",
  34588=>"001001101",
  34589=>"101111111",
  34590=>"000000010",
  34591=>"011011111",
  34592=>"011111111",
  34593=>"111001101",
  34594=>"111100110",
  34595=>"110111011",
  34596=>"110000000",
  34597=>"001110110",
  34598=>"000000000",
  34599=>"100001011",
  34600=>"101101101",
  34601=>"111111111",
  34602=>"000010010",
  34603=>"000000111",
  34604=>"111111111",
  34605=>"100110110",
  34606=>"111111111",
  34607=>"111111000",
  34608=>"111111001",
  34609=>"100110111",
  34610=>"111100000",
  34611=>"000100111",
  34612=>"111000010",
  34613=>"111001010",
  34614=>"011000000",
  34615=>"111110110",
  34616=>"000000000",
  34617=>"010110000",
  34618=>"111111111",
  34619=>"011000000",
  34620=>"111111101",
  34621=>"110100000",
  34622=>"100101111",
  34623=>"000011111",
  34624=>"001010000",
  34625=>"000000000",
  34626=>"000000000",
  34627=>"101101111",
  34628=>"100100100",
  34629=>"111111111",
  34630=>"111101001",
  34631=>"000000000",
  34632=>"100000000",
  34633=>"000000011",
  34634=>"000010111",
  34635=>"110110110",
  34636=>"000110100",
  34637=>"011111111",
  34638=>"111110100",
  34639=>"100001001",
  34640=>"011111111",
  34641=>"100000000",
  34642=>"000000100",
  34643=>"111000000",
  34644=>"111100111",
  34645=>"001001011",
  34646=>"111101100",
  34647=>"011000100",
  34648=>"000111111",
  34649=>"000010000",
  34650=>"101111111",
  34651=>"111101100",
  34652=>"100110001",
  34653=>"000000100",
  34654=>"110000000",
  34655=>"000011111",
  34656=>"000000000",
  34657=>"001000000",
  34658=>"011011011",
  34659=>"100111000",
  34660=>"111111110",
  34661=>"010000000",
  34662=>"110000000",
  34663=>"000000000",
  34664=>"000000001",
  34665=>"000000100",
  34666=>"100000000",
  34667=>"100000000",
  34668=>"000000000",
  34669=>"000000111",
  34670=>"000000101",
  34671=>"110111111",
  34672=>"000000111",
  34673=>"001011000",
  34674=>"000000000",
  34675=>"111111111",
  34676=>"111111111",
  34677=>"011000000",
  34678=>"000000100",
  34679=>"100000000",
  34680=>"111111111",
  34681=>"111001000",
  34682=>"100001100",
  34683=>"000000100",
  34684=>"000010011",
  34685=>"111111111",
  34686=>"000111111",
  34687=>"000111111",
  34688=>"001111111",
  34689=>"000000000",
  34690=>"100100110",
  34691=>"100000110",
  34692=>"000101111",
  34693=>"000010011",
  34694=>"000000000",
  34695=>"111011000",
  34696=>"010000100",
  34697=>"111111110",
  34698=>"110110000",
  34699=>"111111111",
  34700=>"111111111",
  34701=>"111111111",
  34702=>"000011011",
  34703=>"000111111",
  34704=>"001000000",
  34705=>"100111111",
  34706=>"111011111",
  34707=>"111111101",
  34708=>"000000000",
  34709=>"000000000",
  34710=>"111101000",
  34711=>"110111000",
  34712=>"000100111",
  34713=>"001001000",
  34714=>"111101001",
  34715=>"111111111",
  34716=>"000100000",
  34717=>"000000100",
  34718=>"100100000",
  34719=>"001111111",
  34720=>"011000000",
  34721=>"101100101",
  34722=>"100111111",
  34723=>"000000000",
  34724=>"111111111",
  34725=>"111111110",
  34726=>"111111111",
  34727=>"000000000",
  34728=>"000000000",
  34729=>"000100100",
  34730=>"000111111",
  34731=>"000010100",
  34732=>"000000000",
  34733=>"000001111",
  34734=>"100100000",
  34735=>"101111111",
  34736=>"100110111",
  34737=>"110111111",
  34738=>"110110101",
  34739=>"010111110",
  34740=>"111111111",
  34741=>"010010110",
  34742=>"011011011",
  34743=>"111110111",
  34744=>"110100111",
  34745=>"001000100",
  34746=>"111111111",
  34747=>"111111111",
  34748=>"110000000",
  34749=>"111111001",
  34750=>"000011111",
  34751=>"101101101",
  34752=>"111110000",
  34753=>"000000000",
  34754=>"111111111",
  34755=>"011000000",
  34756=>"100000000",
  34757=>"000000101",
  34758=>"111011000",
  34759=>"001001000",
  34760=>"000000000",
  34761=>"001111111",
  34762=>"000000000",
  34763=>"000000000",
  34764=>"111111111",
  34765=>"101111001",
  34766=>"011001000",
  34767=>"001001000",
  34768=>"011001111",
  34769=>"100000100",
  34770=>"001001001",
  34771=>"000000000",
  34772=>"000110100",
  34773=>"110000000",
  34774=>"111111101",
  34775=>"111011001",
  34776=>"100100000",
  34777=>"111111100",
  34778=>"000000111",
  34779=>"111011000",
  34780=>"000000000",
  34781=>"000000000",
  34782=>"111100111",
  34783=>"111111111",
  34784=>"000000000",
  34785=>"000000111",
  34786=>"000111111",
  34787=>"000000000",
  34788=>"000010110",
  34789=>"110111111",
  34790=>"000010110",
  34791=>"000100000",
  34792=>"000000001",
  34793=>"101111111",
  34794=>"100000100",
  34795=>"111111111",
  34796=>"000000001",
  34797=>"001011101",
  34798=>"000000000",
  34799=>"111111011",
  34800=>"010010111",
  34801=>"001001100",
  34802=>"011001000",
  34803=>"010000010",
  34804=>"000110111",
  34805=>"001111111",
  34806=>"001111110",
  34807=>"001001001",
  34808=>"111001000",
  34809=>"000100001",
  34810=>"000000000",
  34811=>"010000000",
  34812=>"111111110",
  34813=>"000000000",
  34814=>"111001000",
  34815=>"111111111",
  34816=>"000100110",
  34817=>"001111000",
  34818=>"111111111",
  34819=>"110111111",
  34820=>"011011011",
  34821=>"100000100",
  34822=>"000000000",
  34823=>"111111111",
  34824=>"111111100",
  34825=>"111111111",
  34826=>"000000011",
  34827=>"110111111",
  34828=>"000100000",
  34829=>"011010010",
  34830=>"010110000",
  34831=>"111111111",
  34832=>"111001001",
  34833=>"000000000",
  34834=>"000000000",
  34835=>"111111111",
  34836=>"000000000",
  34837=>"001000100",
  34838=>"111111011",
  34839=>"001001001",
  34840=>"111111111",
  34841=>"111111111",
  34842=>"100000000",
  34843=>"110110110",
  34844=>"110111110",
  34845=>"000000000",
  34846=>"001000001",
  34847=>"101111000",
  34848=>"000010111",
  34849=>"110110111",
  34850=>"101100000",
  34851=>"000000000",
  34852=>"000000011",
  34853=>"111111111",
  34854=>"110000000",
  34855=>"111111000",
  34856=>"000000000",
  34857=>"001001001",
  34858=>"000110110",
  34859=>"011000000",
  34860=>"111111101",
  34861=>"111111111",
  34862=>"000111111",
  34863=>"110000000",
  34864=>"001000111",
  34865=>"001101101",
  34866=>"111110011",
  34867=>"110111110",
  34868=>"011011000",
  34869=>"111111111",
  34870=>"000000111",
  34871=>"000000000",
  34872=>"111111111",
  34873=>"111000000",
  34874=>"111100000",
  34875=>"111111010",
  34876=>"000000000",
  34877=>"111011111",
  34878=>"000000110",
  34879=>"111111111",
  34880=>"001001011",
  34881=>"111111111",
  34882=>"011111101",
  34883=>"110111010",
  34884=>"000000000",
  34885=>"100000000",
  34886=>"111111110",
  34887=>"000000000",
  34888=>"001011011",
  34889=>"000000000",
  34890=>"111111000",
  34891=>"110110111",
  34892=>"111111000",
  34893=>"000000010",
  34894=>"000010010",
  34895=>"111111111",
  34896=>"001000000",
  34897=>"000101111",
  34898=>"111111111",
  34899=>"110010010",
  34900=>"111001101",
  34901=>"110000000",
  34902=>"110001000",
  34903=>"110110000",
  34904=>"110111111",
  34905=>"000000000",
  34906=>"000000000",
  34907=>"100001001",
  34908=>"111111111",
  34909=>"111111111",
  34910=>"110111111",
  34911=>"111111111",
  34912=>"000000000",
  34913=>"101101100",
  34914=>"110100000",
  34915=>"000000000",
  34916=>"000110000",
  34917=>"000000111",
  34918=>"111111001",
  34919=>"100000100",
  34920=>"100111110",
  34921=>"000000111",
  34922=>"000000001",
  34923=>"101101111",
  34924=>"100000000",
  34925=>"110000100",
  34926=>"000111111",
  34927=>"000000000",
  34928=>"010110111",
  34929=>"111111110",
  34930=>"000000001",
  34931=>"111111111",
  34932=>"111111111",
  34933=>"000110111",
  34934=>"111111111",
  34935=>"000000000",
  34936=>"000100110",
  34937=>"000000000",
  34938=>"000000000",
  34939=>"000000001",
  34940=>"000000000",
  34941=>"000000000",
  34942=>"000000111",
  34943=>"000000000",
  34944=>"000000000",
  34945=>"000000000",
  34946=>"000000000",
  34947=>"000000000",
  34948=>"111110111",
  34949=>"111111111",
  34950=>"010111110",
  34951=>"000000010",
  34952=>"111111111",
  34953=>"001000000",
  34954=>"000110111",
  34955=>"111001011",
  34956=>"000100000",
  34957=>"111111111",
  34958=>"100000111",
  34959=>"000000000",
  34960=>"000011001",
  34961=>"011111111",
  34962=>"000000111",
  34963=>"010010010",
  34964=>"000100111",
  34965=>"000011111",
  34966=>"111111110",
  34967=>"000111111",
  34968=>"000000000",
  34969=>"000000000",
  34970=>"000000111",
  34971=>"100100100",
  34972=>"100110111",
  34973=>"000000000",
  34974=>"111111111",
  34975=>"111000000",
  34976=>"101111111",
  34977=>"000111010",
  34978=>"000000000",
  34979=>"111010111",
  34980=>"000110011",
  34981=>"110110000",
  34982=>"010000000",
  34983=>"001000000",
  34984=>"000010000",
  34985=>"011010000",
  34986=>"000000000",
  34987=>"100101111",
  34988=>"011000001",
  34989=>"100000001",
  34990=>"000001001",
  34991=>"000110000",
  34992=>"000000000",
  34993=>"111011001",
  34994=>"000001000",
  34995=>"000000000",
  34996=>"111111111",
  34997=>"110110000",
  34998=>"000001011",
  34999=>"000000011",
  35000=>"000011001",
  35001=>"110000110",
  35002=>"000000000",
  35003=>"100101001",
  35004=>"000000000",
  35005=>"100111111",
  35006=>"000000000",
  35007=>"000000111",
  35008=>"000101111",
  35009=>"001001111",
  35010=>"111111111",
  35011=>"011111111",
  35012=>"000000000",
  35013=>"111111110",
  35014=>"110110111",
  35015=>"110000111",
  35016=>"000000001",
  35017=>"111111111",
  35018=>"110110110",
  35019=>"000011011",
  35020=>"010111111",
  35021=>"111101111",
  35022=>"111111111",
  35023=>"000001011",
  35024=>"000000011",
  35025=>"000011001",
  35026=>"000000000",
  35027=>"100101101",
  35028=>"000110111",
  35029=>"001000100",
  35030=>"000010000",
  35031=>"000000000",
  35032=>"111100000",
  35033=>"011111111",
  35034=>"000000000",
  35035=>"000000010",
  35036=>"111111000",
  35037=>"010011000",
  35038=>"111111111",
  35039=>"111111101",
  35040=>"111110000",
  35041=>"101000111",
  35042=>"000000000",
  35043=>"100110000",
  35044=>"111111111",
  35045=>"111110110",
  35046=>"000100110",
  35047=>"000010111",
  35048=>"111111111",
  35049=>"000000000",
  35050=>"110110000",
  35051=>"111111111",
  35052=>"111111001",
  35053=>"000000000",
  35054=>"110100100",
  35055=>"010010000",
  35056=>"000000011",
  35057=>"000001101",
  35058=>"000001001",
  35059=>"010011001",
  35060=>"000010111",
  35061=>"111111101",
  35062=>"000000000",
  35063=>"111111111",
  35064=>"000000000",
  35065=>"111111110",
  35066=>"100111001",
  35067=>"100100000",
  35068=>"000000000",
  35069=>"110000000",
  35070=>"111111100",
  35071=>"000000010",
  35072=>"000011111",
  35073=>"110110110",
  35074=>"000000000",
  35075=>"110000011",
  35076=>"111111111",
  35077=>"111111000",
  35078=>"110111100",
  35079=>"111010000",
  35080=>"100101100",
  35081=>"001000000",
  35082=>"111111110",
  35083=>"111011000",
  35084=>"000000100",
  35085=>"110010001",
  35086=>"000111111",
  35087=>"111100010",
  35088=>"111110100",
  35089=>"000000000",
  35090=>"000000000",
  35091=>"110110011",
  35092=>"000000000",
  35093=>"110000111",
  35094=>"011111001",
  35095=>"000000001",
  35096=>"011011011",
  35097=>"000110000",
  35098=>"110111011",
  35099=>"000000000",
  35100=>"111011011",
  35101=>"101001001",
  35102=>"101000000",
  35103=>"011111111",
  35104=>"000000000",
  35105=>"110110000",
  35106=>"000000000",
  35107=>"111011000",
  35108=>"111111110",
  35109=>"000000000",
  35110=>"011111111",
  35111=>"011011110",
  35112=>"111111111",
  35113=>"110110110",
  35114=>"000001011",
  35115=>"000000111",
  35116=>"000011111",
  35117=>"000000100",
  35118=>"000000000",
  35119=>"000000000",
  35120=>"011001001",
  35121=>"111111111",
  35122=>"111111111",
  35123=>"111100100",
  35124=>"000000000",
  35125=>"000000000",
  35126=>"001000000",
  35127=>"000000000",
  35128=>"000000001",
  35129=>"111000110",
  35130=>"100001111",
  35131=>"101111111",
  35132=>"000000000",
  35133=>"111111000",
  35134=>"111111111",
  35135=>"000110000",
  35136=>"000000000",
  35137=>"000000000",
  35138=>"000100000",
  35139=>"000000000",
  35140=>"000000000",
  35141=>"101001000",
  35142=>"011110111",
  35143=>"110111111",
  35144=>"111111111",
  35145=>"000000000",
  35146=>"010111010",
  35147=>"011010110",
  35148=>"111111111",
  35149=>"110001111",
  35150=>"000111111",
  35151=>"011011001",
  35152=>"000000001",
  35153=>"000000000",
  35154=>"111111111",
  35155=>"000000111",
  35156=>"000000000",
  35157=>"000100100",
  35158=>"111001111",
  35159=>"111111111",
  35160=>"000100001",
  35161=>"000000000",
  35162=>"111100000",
  35163=>"110110111",
  35164=>"101101101",
  35165=>"101101000",
  35166=>"001001000",
  35167=>"000110001",
  35168=>"000000000",
  35169=>"111000000",
  35170=>"000010010",
  35171=>"000111111",
  35172=>"000000000",
  35173=>"111111111",
  35174=>"000000111",
  35175=>"100000000",
  35176=>"111001000",
  35177=>"000000000",
  35178=>"000000000",
  35179=>"111111000",
  35180=>"011111011",
  35181=>"000000001",
  35182=>"111111000",
  35183=>"010010000",
  35184=>"011011000",
  35185=>"111000000",
  35186=>"111000000",
  35187=>"000011000",
  35188=>"111111111",
  35189=>"111011011",
  35190=>"000000000",
  35191=>"111101101",
  35192=>"011011011",
  35193=>"000000111",
  35194=>"111111111",
  35195=>"110000001",
  35196=>"000111111",
  35197=>"010011111",
  35198=>"000000000",
  35199=>"000100000",
  35200=>"111111111",
  35201=>"100111111",
  35202=>"000010010",
  35203=>"111111111",
  35204=>"111000000",
  35205=>"000000000",
  35206=>"001000110",
  35207=>"001111001",
  35208=>"001111010",
  35209=>"111011111",
  35210=>"000100111",
  35211=>"001000000",
  35212=>"000000000",
  35213=>"101101000",
  35214=>"111111111",
  35215=>"000000000",
  35216=>"111111111",
  35217=>"111110110",
  35218=>"000100000",
  35219=>"000000000",
  35220=>"110111110",
  35221=>"000000111",
  35222=>"100100000",
  35223=>"111111111",
  35224=>"000111111",
  35225=>"111111111",
  35226=>"111111111",
  35227=>"000001101",
  35228=>"000000111",
  35229=>"100000010",
  35230=>"100000000",
  35231=>"000000000",
  35232=>"111111111",
  35233=>"100100100",
  35234=>"110110000",
  35235=>"000000000",
  35236=>"001111110",
  35237=>"111111100",
  35238=>"010010000",
  35239=>"111111001",
  35240=>"001000000",
  35241=>"010010011",
  35242=>"000000000",
  35243=>"000000000",
  35244=>"101000110",
  35245=>"101001000",
  35246=>"111011011",
  35247=>"000000001",
  35248=>"011000110",
  35249=>"000000000",
  35250=>"001011000",
  35251=>"000000000",
  35252=>"111111111",
  35253=>"011111111",
  35254=>"111111001",
  35255=>"000000000",
  35256=>"111010010",
  35257=>"111000000",
  35258=>"000100000",
  35259=>"100110100",
  35260=>"111111111",
  35261=>"011011111",
  35262=>"000000000",
  35263=>"010010010",
  35264=>"111111111",
  35265=>"111111011",
  35266=>"111111111",
  35267=>"000000000",
  35268=>"000011110",
  35269=>"001001000",
  35270=>"000000000",
  35271=>"101111111",
  35272=>"000000000",
  35273=>"000000111",
  35274=>"000000000",
  35275=>"000000000",
  35276=>"000000000",
  35277=>"010111111",
  35278=>"010000000",
  35279=>"111001001",
  35280=>"100110000",
  35281=>"000000000",
  35282=>"011001001",
  35283=>"111111111",
  35284=>"000110010",
  35285=>"000000000",
  35286=>"000100111",
  35287=>"000011111",
  35288=>"111111111",
  35289=>"111100100",
  35290=>"100110100",
  35291=>"000000111",
  35292=>"111111000",
  35293=>"000000000",
  35294=>"000100000",
  35295=>"010011010",
  35296=>"000000000",
  35297=>"000000111",
  35298=>"111111111",
  35299=>"111000000",
  35300=>"110110000",
  35301=>"111000000",
  35302=>"000011111",
  35303=>"001000101",
  35304=>"100000011",
  35305=>"111111111",
  35306=>"110000001",
  35307=>"011110000",
  35308=>"111111110",
  35309=>"000000100",
  35310=>"000100111",
  35311=>"111110000",
  35312=>"000000000",
  35313=>"111101101",
  35314=>"111000001",
  35315=>"111111111",
  35316=>"100111000",
  35317=>"000000000",
  35318=>"000000000",
  35319=>"001001001",
  35320=>"010000001",
  35321=>"000000100",
  35322=>"111111111",
  35323=>"000000111",
  35324=>"001001111",
  35325=>"000000100",
  35326=>"000000000",
  35327=>"000000000",
  35328=>"111111111",
  35329=>"100111111",
  35330=>"111110100",
  35331=>"000000000",
  35332=>"111111111",
  35333=>"110000111",
  35334=>"000000001",
  35335=>"000000111",
  35336=>"000000000",
  35337=>"101000000",
  35338=>"000000000",
  35339=>"100001011",
  35340=>"000000000",
  35341=>"111111111",
  35342=>"001111111",
  35343=>"001101111",
  35344=>"000000000",
  35345=>"000000000",
  35346=>"111111000",
  35347=>"000011111",
  35348=>"100111110",
  35349=>"000011000",
  35350=>"111111111",
  35351=>"011001001",
  35352=>"110000000",
  35353=>"001111111",
  35354=>"100111111",
  35355=>"000000000",
  35356=>"000000000",
  35357=>"111111000",
  35358=>"100110010",
  35359=>"011000111",
  35360=>"100111111",
  35361=>"000010010",
  35362=>"110110000",
  35363=>"111111111",
  35364=>"100100000",
  35365=>"000110110",
  35366=>"001001001",
  35367=>"111101101",
  35368=>"101001000",
  35369=>"000000000",
  35370=>"000000000",
  35371=>"000011111",
  35372=>"101001001",
  35373=>"111111101",
  35374=>"111111101",
  35375=>"000000011",
  35376=>"000000001",
  35377=>"111111000",
  35378=>"001100100",
  35379=>"000000101",
  35380=>"111101111",
  35381=>"000000000",
  35382=>"000000000",
  35383=>"100100111",
  35384=>"111101011",
  35385=>"000001001",
  35386=>"001001111",
  35387=>"111111101",
  35388=>"111110000",
  35389=>"000000101",
  35390=>"110100100",
  35391=>"111111111",
  35392=>"111011111",
  35393=>"000000100",
  35394=>"000000110",
  35395=>"000000101",
  35396=>"000110011",
  35397=>"001111111",
  35398=>"100000000",
  35399=>"111111111",
  35400=>"001001111",
  35401=>"000000100",
  35402=>"110111111",
  35403=>"111111100",
  35404=>"110000110",
  35405=>"010000101",
  35406=>"110111111",
  35407=>"000001111",
  35408=>"000000000",
  35409=>"101000000",
  35410=>"111111111",
  35411=>"000000000",
  35412=>"111111111",
  35413=>"000000010",
  35414=>"011111001",
  35415=>"111111110",
  35416=>"000000001",
  35417=>"111100000",
  35418=>"111111111",
  35419=>"000000000",
  35420=>"111111001",
  35421=>"010111111",
  35422=>"001000000",
  35423=>"111001000",
  35424=>"111111111",
  35425=>"000000000",
  35426=>"100111001",
  35427=>"000110010",
  35428=>"000000000",
  35429=>"000000000",
  35430=>"000000000",
  35431=>"000000000",
  35432=>"001000000",
  35433=>"101111111",
  35434=>"011000000",
  35435=>"001000111",
  35436=>"111111111",
  35437=>"110111000",
  35438=>"001000001",
  35439=>"111111111",
  35440=>"000000110",
  35441=>"000000000",
  35442=>"000000100",
  35443=>"111111111",
  35444=>"100111111",
  35445=>"111110000",
  35446=>"010011111",
  35447=>"101000101",
  35448=>"111111111",
  35449=>"111001111",
  35450=>"111000000",
  35451=>"001000000",
  35452=>"000100100",
  35453=>"000010010",
  35454=>"111111011",
  35455=>"000000101",
  35456=>"111111111",
  35457=>"001000000",
  35458=>"111111111",
  35459=>"000000000",
  35460=>"111111111",
  35461=>"001000000",
  35462=>"111011001",
  35463=>"111111111",
  35464=>"000000000",
  35465=>"111111111",
  35466=>"111111111",
  35467=>"111111111",
  35468=>"111100000",
  35469=>"000000000",
  35470=>"001000001",
  35471=>"111110100",
  35472=>"000000110",
  35473=>"000000000",
  35474=>"000000000",
  35475=>"000000000",
  35476=>"000001000",
  35477=>"111111111",
  35478=>"000101101",
  35479=>"001100111",
  35480=>"000000111",
  35481=>"111111000",
  35482=>"100101111",
  35483=>"000000000",
  35484=>"000000000",
  35485=>"000000000",
  35486=>"100101111",
  35487=>"000001011",
  35488=>"000000000",
  35489=>"011011100",
  35490=>"110111111",
  35491=>"111111111",
  35492=>"000000000",
  35493=>"000000000",
  35494=>"000000000",
  35495=>"011011011",
  35496=>"000000000",
  35497=>"000100100",
  35498=>"000000101",
  35499=>"000000111",
  35500=>"111010001",
  35501=>"111111110",
  35502=>"111111111",
  35503=>"011001000",
  35504=>"110000111",
  35505=>"001001001",
  35506=>"011111111",
  35507=>"000000110",
  35508=>"000000000",
  35509=>"111111001",
  35510=>"000111100",
  35511=>"111111111",
  35512=>"111111111",
  35513=>"101001000",
  35514=>"100100101",
  35515=>"000000001",
  35516=>"111111111",
  35517=>"000000110",
  35518=>"011011110",
  35519=>"000000111",
  35520=>"000000100",
  35521=>"000001001",
  35522=>"111111111",
  35523=>"001111000",
  35524=>"010011111",
  35525=>"001000000",
  35526=>"000000000",
  35527=>"111111111",
  35528=>"111111111",
  35529=>"111111101",
  35530=>"110000100",
  35531=>"111111111",
  35532=>"101001000",
  35533=>"000000101",
  35534=>"111101001",
  35535=>"111110110",
  35536=>"011000000",
  35537=>"000111111",
  35538=>"110111000",
  35539=>"100000111",
  35540=>"111011010",
  35541=>"111111000",
  35542=>"110110010",
  35543=>"000000000",
  35544=>"000000001",
  35545=>"000000111",
  35546=>"000000000",
  35547=>"011011111",
  35548=>"011001011",
  35549=>"111111111",
  35550=>"001000000",
  35551=>"000001001",
  35552=>"000000111",
  35553=>"000000000",
  35554=>"011001000",
  35555=>"001001001",
  35556=>"111010000",
  35557=>"000000000",
  35558=>"000000000",
  35559=>"111000000",
  35560=>"111111010",
  35561=>"000000000",
  35562=>"111001111",
  35563=>"000000101",
  35564=>"111111011",
  35565=>"000000001",
  35566=>"111111111",
  35567=>"000111111",
  35568=>"110000000",
  35569=>"111000001",
  35570=>"110111101",
  35571=>"000000000",
  35572=>"000000111",
  35573=>"111111000",
  35574=>"110111111",
  35575=>"111111111",
  35576=>"000000000",
  35577=>"111111100",
  35578=>"111111111",
  35579=>"110100000",
  35580=>"011011000",
  35581=>"110101111",
  35582=>"000000000",
  35583=>"111111111",
  35584=>"000000011",
  35585=>"000010010",
  35586=>"000000111",
  35587=>"001010111",
  35588=>"000100100",
  35589=>"111111111",
  35590=>"110111000",
  35591=>"000101111",
  35592=>"111111111",
  35593=>"000000000",
  35594=>"101000000",
  35595=>"000000000",
  35596=>"110100000",
  35597=>"111111000",
  35598=>"110100000",
  35599=>"111011000",
  35600=>"000000001",
  35601=>"111111100",
  35602=>"100000001",
  35603=>"111111111",
  35604=>"101111000",
  35605=>"111111011",
  35606=>"001111111",
  35607=>"111111111",
  35608=>"111101001",
  35609=>"000101100",
  35610=>"111010010",
  35611=>"100000000",
  35612=>"000000000",
  35613=>"111100101",
  35614=>"000000000",
  35615=>"001100110",
  35616=>"000000000",
  35617=>"111001011",
  35618=>"111100100",
  35619=>"111111111",
  35620=>"000110000",
  35621=>"100111111",
  35622=>"111001000",
  35623=>"011011111",
  35624=>"000000000",
  35625=>"000000000",
  35626=>"111000111",
  35627=>"000000000",
  35628=>"100111000",
  35629=>"110010000",
  35630=>"110000110",
  35631=>"011101001",
  35632=>"001001011",
  35633=>"100000000",
  35634=>"111111111",
  35635=>"111111111",
  35636=>"110101111",
  35637=>"111001001",
  35638=>"000111001",
  35639=>"000000000",
  35640=>"111111110",
  35641=>"111111111",
  35642=>"111111111",
  35643=>"000010110",
  35644=>"111111111",
  35645=>"000001100",
  35646=>"011001001",
  35647=>"111111000",
  35648=>"000001111",
  35649=>"101100100",
  35650=>"001000000",
  35651=>"100110111",
  35652=>"000000111",
  35653=>"000000111",
  35654=>"000000000",
  35655=>"111111111",
  35656=>"000011001",
  35657=>"111101101",
  35658=>"000000100",
  35659=>"000100100",
  35660=>"000000000",
  35661=>"111001001",
  35662=>"110111111",
  35663=>"110110110",
  35664=>"000001001",
  35665=>"111001000",
  35666=>"000100111",
  35667=>"111111111",
  35668=>"110000000",
  35669=>"011001001",
  35670=>"011100000",
  35671=>"111010010",
  35672=>"000000000",
  35673=>"110111111",
  35674=>"111111001",
  35675=>"111111011",
  35676=>"000011111",
  35677=>"000000111",
  35678=>"000000000",
  35679=>"111111111",
  35680=>"111111111",
  35681=>"111110000",
  35682=>"011111111",
  35683=>"000000000",
  35684=>"001000001",
  35685=>"000001001",
  35686=>"110111111",
  35687=>"101111111",
  35688=>"001001001",
  35689=>"000000111",
  35690=>"101111111",
  35691=>"010010000",
  35692=>"000011011",
  35693=>"101000000",
  35694=>"000000000",
  35695=>"000000000",
  35696=>"100000000",
  35697=>"111111111",
  35698=>"110100110",
  35699=>"111111001",
  35700=>"111111111",
  35701=>"100000000",
  35702=>"010000000",
  35703=>"000000111",
  35704=>"111111111",
  35705=>"110000000",
  35706=>"001000010",
  35707=>"000011111",
  35708=>"101001001",
  35709=>"000000111",
  35710=>"111101000",
  35711=>"111100000",
  35712=>"001101111",
  35713=>"111101011",
  35714=>"010111111",
  35715=>"000000000",
  35716=>"111111001",
  35717=>"111000000",
  35718=>"000011111",
  35719=>"110111111",
  35720=>"000000010",
  35721=>"001011011",
  35722=>"111111011",
  35723=>"110110111",
  35724=>"111111111",
  35725=>"111111110",
  35726=>"110010000",
  35727=>"000000000",
  35728=>"000000000",
  35729=>"001001001",
  35730=>"000000000",
  35731=>"111111111",
  35732=>"111111111",
  35733=>"000000000",
  35734=>"000000000",
  35735=>"000100101",
  35736=>"001011001",
  35737=>"100110000",
  35738=>"111111111",
  35739=>"100101111",
  35740=>"000000010",
  35741=>"110000000",
  35742=>"000000000",
  35743=>"000010010",
  35744=>"111000000",
  35745=>"111111111",
  35746=>"100000111",
  35747=>"111111111",
  35748=>"111101111",
  35749=>"001000000",
  35750=>"101101111",
  35751=>"100000111",
  35752=>"111111110",
  35753=>"000000000",
  35754=>"000000000",
  35755=>"011111100",
  35756=>"000111000",
  35757=>"000000001",
  35758=>"000011111",
  35759=>"000001001",
  35760=>"111111111",
  35761=>"111111110",
  35762=>"111111110",
  35763=>"111111111",
  35764=>"001100100",
  35765=>"011000100",
  35766=>"100111111",
  35767=>"111111111",
  35768=>"111111111",
  35769=>"000000000",
  35770=>"111111111",
  35771=>"100100100",
  35772=>"011111111",
  35773=>"000000000",
  35774=>"000000000",
  35775=>"000110010",
  35776=>"011000111",
  35777=>"000000000",
  35778=>"011001000",
  35779=>"000111111",
  35780=>"000000000",
  35781=>"001000110",
  35782=>"011001111",
  35783=>"000000000",
  35784=>"111011001",
  35785=>"111000000",
  35786=>"000001111",
  35787=>"000110000",
  35788=>"000000000",
  35789=>"000000001",
  35790=>"011001000",
  35791=>"000000000",
  35792=>"110000000",
  35793=>"011111101",
  35794=>"010000000",
  35795=>"111011011",
  35796=>"001000000",
  35797=>"001001111",
  35798=>"001000000",
  35799=>"000000000",
  35800=>"000000000",
  35801=>"100000000",
  35802=>"011001111",
  35803=>"111111101",
  35804=>"000000111",
  35805=>"000000000",
  35806=>"000000000",
  35807=>"000001000",
  35808=>"000000110",
  35809=>"111111111",
  35810=>"111111110",
  35811=>"111111111",
  35812=>"111111011",
  35813=>"000001111",
  35814=>"001000100",
  35815=>"111111111",
  35816=>"001101100",
  35817=>"000011111",
  35818=>"000000000",
  35819=>"011111111",
  35820=>"111111111",
  35821=>"011011111",
  35822=>"111111111",
  35823=>"111111100",
  35824=>"000000000",
  35825=>"001111111",
  35826=>"000000000",
  35827=>"000000000",
  35828=>"111111000",
  35829=>"000110111",
  35830=>"111111000",
  35831=>"111111110",
  35832=>"111111111",
  35833=>"001000001",
  35834=>"000000000",
  35835=>"011011011",
  35836=>"111110111",
  35837=>"000000000",
  35838=>"111011011",
  35839=>"001000000",
  35840=>"000000000",
  35841=>"000000000",
  35842=>"111111111",
  35843=>"101111101",
  35844=>"011111111",
  35845=>"111111101",
  35846=>"000000000",
  35847=>"000111111",
  35848=>"111110000",
  35849=>"111111111",
  35850=>"000010000",
  35851=>"000000111",
  35852=>"000110110",
  35853=>"111111111",
  35854=>"111111011",
  35855=>"000010000",
  35856=>"100000110",
  35857=>"000000001",
  35858=>"011111110",
  35859=>"100000000",
  35860=>"110010111",
  35861=>"000000000",
  35862=>"000000000",
  35863=>"001001011",
  35864=>"110110110",
  35865=>"011111111",
  35866=>"000000000",
  35867=>"000100100",
  35868=>"000000000",
  35869=>"111111111",
  35870=>"000001000",
  35871=>"011111111",
  35872=>"111111110",
  35873=>"000000000",
  35874=>"000000000",
  35875=>"000000000",
  35876=>"111111111",
  35877=>"111000100",
  35878=>"000000011",
  35879=>"111010110",
  35880=>"000000000",
  35881=>"000000000",
  35882=>"111100111",
  35883=>"101111111",
  35884=>"000000011",
  35885=>"001001001",
  35886=>"000000101",
  35887=>"001000000",
  35888=>"111111001",
  35889=>"000010000",
  35890=>"111001000",
  35891=>"000000000",
  35892=>"001100000",
  35893=>"100000000",
  35894=>"110000111",
  35895=>"110000000",
  35896=>"110110111",
  35897=>"000000111",
  35898=>"000100110",
  35899=>"000000111",
  35900=>"111111111",
  35901=>"000011111",
  35902=>"101111111",
  35903=>"011001101",
  35904=>"001000000",
  35905=>"110111111",
  35906=>"000001111",
  35907=>"000000000",
  35908=>"000110110",
  35909=>"111111011",
  35910=>"010110110",
  35911=>"011011000",
  35912=>"111111111",
  35913=>"111111111",
  35914=>"100000001",
  35915=>"000000111",
  35916=>"101001000",
  35917=>"000000111",
  35918=>"000010000",
  35919=>"101111111",
  35920=>"001001000",
  35921=>"111000000",
  35922=>"111111111",
  35923=>"101101100",
  35924=>"111111001",
  35925=>"000000001",
  35926=>"000010110",
  35927=>"111101101",
  35928=>"000010010",
  35929=>"000000000",
  35930=>"101001000",
  35931=>"000100100",
  35932=>"000000000",
  35933=>"111111100",
  35934=>"000001000",
  35935=>"110110110",
  35936=>"000000000",
  35937=>"000000000",
  35938=>"000010000",
  35939=>"000000111",
  35940=>"010111000",
  35941=>"111011000",
  35942=>"100100100",
  35943=>"001000010",
  35944=>"000111111",
  35945=>"111111110",
  35946=>"000000001",
  35947=>"000000000",
  35948=>"011111111",
  35949=>"111111111",
  35950=>"111111111",
  35951=>"111111110",
  35952=>"111101101",
  35953=>"000000000",
  35954=>"011011001",
  35955=>"000000000",
  35956=>"111111000",
  35957=>"000010000",
  35958=>"110000000",
  35959=>"000000000",
  35960=>"111111111",
  35961=>"111111111",
  35962=>"000110111",
  35963=>"100100100",
  35964=>"110110110",
  35965=>"000000000",
  35966=>"000000000",
  35967=>"000000000",
  35968=>"000000110",
  35969=>"111111111",
  35970=>"111000000",
  35971=>"000000000",
  35972=>"111111110",
  35973=>"111011111",
  35974=>"111110110",
  35975=>"000010010",
  35976=>"111111111",
  35977=>"100111000",
  35978=>"000000010",
  35979=>"100111111",
  35980=>"000100111",
  35981=>"000000000",
  35982=>"000001011",
  35983=>"000000000",
  35984=>"111111111",
  35985=>"111111101",
  35986=>"111110110",
  35987=>"000001001",
  35988=>"000011111",
  35989=>"000000011",
  35990=>"111111000",
  35991=>"110110111",
  35992=>"111110010",
  35993=>"001100110",
  35994=>"111111111",
  35995=>"010111111",
  35996=>"100000111",
  35997=>"000010110",
  35998=>"111001011",
  35999=>"001111111",
  36000=>"000000001",
  36001=>"001000000",
  36002=>"000000000",
  36003=>"011001000",
  36004=>"000000000",
  36005=>"000000110",
  36006=>"000000000",
  36007=>"011001001",
  36008=>"001001000",
  36009=>"000000000",
  36010=>"111111111",
  36011=>"111111110",
  36012=>"110110110",
  36013=>"111111110",
  36014=>"000000000",
  36015=>"111101000",
  36016=>"000000000",
  36017=>"111110101",
  36018=>"010011111",
  36019=>"111111000",
  36020=>"001001111",
  36021=>"000000000",
  36022=>"000100111",
  36023=>"000000000",
  36024=>"100000100",
  36025=>"000000000",
  36026=>"000000111",
  36027=>"111011111",
  36028=>"101100100",
  36029=>"000000000",
  36030=>"111111000",
  36031=>"000000000",
  36032=>"011100111",
  36033=>"111111011",
  36034=>"000010011",
  36035=>"001000000",
  36036=>"111111111",
  36037=>"000101111",
  36038=>"000000000",
  36039=>"001001111",
  36040=>"011000000",
  36041=>"000001111",
  36042=>"000001001",
  36043=>"000001100",
  36044=>"111111111",
  36045=>"001001101",
  36046=>"111001111",
  36047=>"100000000",
  36048=>"000111011",
  36049=>"000000101",
  36050=>"111111111",
  36051=>"111111111",
  36052=>"000000000",
  36053=>"100100000",
  36054=>"001001011",
  36055=>"000000101",
  36056=>"111110111",
  36057=>"000110110",
  36058=>"000000000",
  36059=>"111111111",
  36060=>"100111111",
  36061=>"111111111",
  36062=>"111111111",
  36063=>"111000000",
  36064=>"100000010",
  36065=>"000100000",
  36066=>"111111100",
  36067=>"000000000",
  36068=>"000101111",
  36069=>"000001111",
  36070=>"111111111",
  36071=>"000000110",
  36072=>"110110000",
  36073=>"000110001",
  36074=>"000111111",
  36075=>"001001111",
  36076=>"111111111",
  36077=>"111000000",
  36078=>"111100111",
  36079=>"111111111",
  36080=>"001000101",
  36081=>"000011001",
  36082=>"111111111",
  36083=>"111111111",
  36084=>"000000111",
  36085=>"111001001",
  36086=>"111111011",
  36087=>"111111110",
  36088=>"000000000",
  36089=>"000000000",
  36090=>"000011001",
  36091=>"000010010",
  36092=>"000000000",
  36093=>"100000000",
  36094=>"111001000",
  36095=>"111100100",
  36096=>"110111111",
  36097=>"111111100",
  36098=>"111000000",
  36099=>"111111000",
  36100=>"111111000",
  36101=>"110000000",
  36102=>"111111111",
  36103=>"111111111",
  36104=>"000000000",
  36105=>"111011011",
  36106=>"000001101",
  36107=>"100110111",
  36108=>"110000000",
  36109=>"111000000",
  36110=>"000000000",
  36111=>"000111111",
  36112=>"111100000",
  36113=>"000000101",
  36114=>"011111111",
  36115=>"101111110",
  36116=>"000000000",
  36117=>"000000000",
  36118=>"100110100",
  36119=>"111111111",
  36120=>"000001000",
  36121=>"111110110",
  36122=>"000000000",
  36123=>"000000001",
  36124=>"000111111",
  36125=>"111111011",
  36126=>"111010000",
  36127=>"111111111",
  36128=>"101011000",
  36129=>"000000100",
  36130=>"111111000",
  36131=>"100111000",
  36132=>"111000000",
  36133=>"111001101",
  36134=>"000000111",
  36135=>"011010000",
  36136=>"000000000",
  36137=>"000111011",
  36138=>"000010010",
  36139=>"111111111",
  36140=>"110110110",
  36141=>"101111111",
  36142=>"000000000",
  36143=>"000000000",
  36144=>"000011010",
  36145=>"111111111",
  36146=>"000000000",
  36147=>"000000111",
  36148=>"111111110",
  36149=>"111111111",
  36150=>"000000000",
  36151=>"111111110",
  36152=>"001011000",
  36153=>"000000000",
  36154=>"000110110",
  36155=>"111111000",
  36156=>"100100111",
  36157=>"000010000",
  36158=>"100101100",
  36159=>"111111111",
  36160=>"000000000",
  36161=>"000000000",
  36162=>"000110000",
  36163=>"111000000",
  36164=>"111000000",
  36165=>"000111111",
  36166=>"000111111",
  36167=>"111000001",
  36168=>"111111101",
  36169=>"110111111",
  36170=>"010010000",
  36171=>"001000000",
  36172=>"001000000",
  36173=>"000000010",
  36174=>"000000001",
  36175=>"111111000",
  36176=>"000110110",
  36177=>"000000000",
  36178=>"011000000",
  36179=>"111000010",
  36180=>"000000000",
  36181=>"001000001",
  36182=>"100100100",
  36183=>"101001111",
  36184=>"000000011",
  36185=>"000000000",
  36186=>"000000000",
  36187=>"000000000",
  36188=>"010000000",
  36189=>"100111100",
  36190=>"100110000",
  36191=>"111111111",
  36192=>"001000001",
  36193=>"111111000",
  36194=>"100000001",
  36195=>"111111111",
  36196=>"111111111",
  36197=>"100000111",
  36198=>"111111101",
  36199=>"110110110",
  36200=>"101000000",
  36201=>"000000000",
  36202=>"011111111",
  36203=>"000001000",
  36204=>"000100100",
  36205=>"011000000",
  36206=>"000000001",
  36207=>"100000000",
  36208=>"000000000",
  36209=>"111010000",
  36210=>"111000000",
  36211=>"000000001",
  36212=>"111110000",
  36213=>"111111111",
  36214=>"111111111",
  36215=>"111111110",
  36216=>"111011111",
  36217=>"111111111",
  36218=>"000000000",
  36219=>"010111000",
  36220=>"000000000",
  36221=>"101000000",
  36222=>"111111000",
  36223=>"001101111",
  36224=>"110111111",
  36225=>"101000000",
  36226=>"111011011",
  36227=>"111111110",
  36228=>"111010111",
  36229=>"111111000",
  36230=>"000000100",
  36231=>"100111010",
  36232=>"110010000",
  36233=>"000000111",
  36234=>"111111101",
  36235=>"111111110",
  36236=>"111111111",
  36237=>"101001001",
  36238=>"000111111",
  36239=>"000000000",
  36240=>"111111000",
  36241=>"111111111",
  36242=>"111111110",
  36243=>"001001111",
  36244=>"111111111",
  36245=>"000010010",
  36246=>"000000000",
  36247=>"001001000",
  36248=>"000000100",
  36249=>"111111110",
  36250=>"100110110",
  36251=>"110110000",
  36252=>"001001000",
  36253=>"111111011",
  36254=>"011001111",
  36255=>"000000000",
  36256=>"000000000",
  36257=>"111011001",
  36258=>"100110111",
  36259=>"111111001",
  36260=>"000000000",
  36261=>"000000000",
  36262=>"111000000",
  36263=>"001000100",
  36264=>"111111000",
  36265=>"111101111",
  36266=>"000111110",
  36267=>"111000111",
  36268=>"000000010",
  36269=>"000000000",
  36270=>"111111111",
  36271=>"000111111",
  36272=>"000100100",
  36273=>"000010010",
  36274=>"111000100",
  36275=>"100000000",
  36276=>"111011111",
  36277=>"000000001",
  36278=>"001111111",
  36279=>"110111000",
  36280=>"010010010",
  36281=>"000100000",
  36282=>"001001000",
  36283=>"111100000",
  36284=>"000101111",
  36285=>"111111111",
  36286=>"101011111",
  36287=>"111101001",
  36288=>"001001000",
  36289=>"000011111",
  36290=>"111111111",
  36291=>"110000000",
  36292=>"001000000",
  36293=>"011001000",
  36294=>"100000011",
  36295=>"000000010",
  36296=>"001001011",
  36297=>"000111000",
  36298=>"001000001",
  36299=>"111111111",
  36300=>"000011000",
  36301=>"101111110",
  36302=>"111111111",
  36303=>"000001111",
  36304=>"011011011",
  36305=>"000000000",
  36306=>"111011011",
  36307=>"111111111",
  36308=>"111101111",
  36309=>"111100100",
  36310=>"011001001",
  36311=>"000011111",
  36312=>"001111001",
  36313=>"111001001",
  36314=>"111111110",
  36315=>"111111111",
  36316=>"000000001",
  36317=>"111111101",
  36318=>"111111111",
  36319=>"001001001",
  36320=>"000000011",
  36321=>"110111111",
  36322=>"000000111",
  36323=>"111111111",
  36324=>"111111100",
  36325=>"111111110",
  36326=>"111100100",
  36327=>"000000000",
  36328=>"011011111",
  36329=>"000111111",
  36330=>"001001001",
  36331=>"000000101",
  36332=>"110111111",
  36333=>"111111001",
  36334=>"000000111",
  36335=>"111011111",
  36336=>"000000000",
  36337=>"000000000",
  36338=>"000011000",
  36339=>"000101111",
  36340=>"000001111",
  36341=>"111111111",
  36342=>"000000000",
  36343=>"111101000",
  36344=>"001001011",
  36345=>"101001001",
  36346=>"110110111",
  36347=>"010010010",
  36348=>"011010111",
  36349=>"010000000",
  36350=>"101000000",
  36351=>"111111111",
  36352=>"000100110",
  36353=>"111001100",
  36354=>"100000000",
  36355=>"111111000",
  36356=>"110111111",
  36357=>"111111111",
  36358=>"001000000",
  36359=>"111111111",
  36360=>"011011111",
  36361=>"100100000",
  36362=>"000010111",
  36363=>"000010110",
  36364=>"111011101",
  36365=>"111101110",
  36366=>"010000110",
  36367=>"111111111",
  36368=>"111011001",
  36369=>"001011010",
  36370=>"000111111",
  36371=>"111111111",
  36372=>"100111111",
  36373=>"001000100",
  36374=>"111110000",
  36375=>"101000000",
  36376=>"001000000",
  36377=>"100101100",
  36378=>"000100110",
  36379=>"001111111",
  36380=>"111111000",
  36381=>"000111011",
  36382=>"011000000",
  36383=>"111000000",
  36384=>"000000100",
  36385=>"000011011",
  36386=>"000000101",
  36387=>"000011001",
  36388=>"010110111",
  36389=>"100110111",
  36390=>"000010000",
  36391=>"111110111",
  36392=>"001111111",
  36393=>"110110010",
  36394=>"111000011",
  36395=>"011001001",
  36396=>"111011000",
  36397=>"101000101",
  36398=>"000000000",
  36399=>"111111111",
  36400=>"001000010",
  36401=>"111111111",
  36402=>"111111101",
  36403=>"111000000",
  36404=>"110110000",
  36405=>"101101000",
  36406=>"111000000",
  36407=>"101110010",
  36408=>"110111111",
  36409=>"111111011",
  36410=>"100000000",
  36411=>"000000100",
  36412=>"000000000",
  36413=>"000000011",
  36414=>"010011011",
  36415=>"000000000",
  36416=>"001000000",
  36417=>"000000000",
  36418=>"111111000",
  36419=>"101100100",
  36420=>"111011011",
  36421=>"011100100",
  36422=>"111010010",
  36423=>"000000000",
  36424=>"100011000",
  36425=>"001000111",
  36426=>"000111000",
  36427=>"000000000",
  36428=>"111110110",
  36429=>"101101111",
  36430=>"111100111",
  36431=>"111000001",
  36432=>"000111111",
  36433=>"111111111",
  36434=>"111111100",
  36435=>"101100110",
  36436=>"111001111",
  36437=>"000000100",
  36438=>"011001000",
  36439=>"001001001",
  36440=>"000000110",
  36441=>"101100000",
  36442=>"000000000",
  36443=>"011111111",
  36444=>"100100100",
  36445=>"000000000",
  36446=>"011010100",
  36447=>"000000000",
  36448=>"000000000",
  36449=>"001011001",
  36450=>"011010000",
  36451=>"001111100",
  36452=>"111111111",
  36453=>"000011010",
  36454=>"000000000",
  36455=>"110000111",
  36456=>"001000000",
  36457=>"100110110",
  36458=>"111111011",
  36459=>"111000000",
  36460=>"000001000",
  36461=>"111101001",
  36462=>"111010010",
  36463=>"000000100",
  36464=>"001010000",
  36465=>"110100100",
  36466=>"011011011",
  36467=>"011011000",
  36468=>"111111111",
  36469=>"110000011",
  36470=>"111111111",
  36471=>"000010000",
  36472=>"011111110",
  36473=>"000000010",
  36474=>"111011000",
  36475=>"000010111",
  36476=>"100000000",
  36477=>"011011011",
  36478=>"000000000",
  36479=>"000011111",
  36480=>"100001001",
  36481=>"111111010",
  36482=>"111001111",
  36483=>"110110110",
  36484=>"110100100",
  36485=>"000111111",
  36486=>"001000000",
  36487=>"111111000",
  36488=>"111011001",
  36489=>"001110110",
  36490=>"000000111",
  36491=>"100100100",
  36492=>"100000100",
  36493=>"110001000",
  36494=>"000000000",
  36495=>"000100101",
  36496=>"011001001",
  36497=>"111110110",
  36498=>"111000001",
  36499=>"001100111",
  36500=>"110111110",
  36501=>"000000100",
  36502=>"000100111",
  36503=>"000000000",
  36504=>"110010010",
  36505=>"011000100",
  36506=>"111111111",
  36507=>"000000000",
  36508=>"000000100",
  36509=>"001110110",
  36510=>"000111111",
  36511=>"111110011",
  36512=>"000000000",
  36513=>"111011000",
  36514=>"001001111",
  36515=>"011111111",
  36516=>"111100011",
  36517=>"100101100",
  36518=>"101101101",
  36519=>"000001001",
  36520=>"000001000",
  36521=>"001011111",
  36522=>"110111111",
  36523=>"000100000",
  36524=>"000000000",
  36525=>"001001000",
  36526=>"000000000",
  36527=>"000000111",
  36528=>"111111101",
  36529=>"000111001",
  36530=>"101101101",
  36531=>"111101111",
  36532=>"111111111",
  36533=>"100111111",
  36534=>"000000000",
  36535=>"100000000",
  36536=>"010011111",
  36537=>"000000000",
  36538=>"011011010",
  36539=>"100000000",
  36540=>"000000000",
  36541=>"101000000",
  36542=>"111111111",
  36543=>"001000000",
  36544=>"110111011",
  36545=>"110111111",
  36546=>"111111011",
  36547=>"011011010",
  36548=>"000000000",
  36549=>"111111011",
  36550=>"111111111",
  36551=>"000000010",
  36552=>"000000000",
  36553=>"000000000",
  36554=>"111111111",
  36555=>"000000000",
  36556=>"111111000",
  36557=>"111111101",
  36558=>"111111111",
  36559=>"001000000",
  36560=>"011101100",
  36561=>"110100100",
  36562=>"001000111",
  36563=>"000000101",
  36564=>"111101000",
  36565=>"111111110",
  36566=>"000101111",
  36567=>"000011111",
  36568=>"011000111",
  36569=>"110010000",
  36570=>"111101111",
  36571=>"000000000",
  36572=>"001000000",
  36573=>"010110111",
  36574=>"111111110",
  36575=>"000000000",
  36576=>"000000000",
  36577=>"001001111",
  36578=>"111111111",
  36579=>"100100110",
  36580=>"110111111",
  36581=>"011001100",
  36582=>"010000000",
  36583=>"011001011",
  36584=>"001001011",
  36585=>"111101111",
  36586=>"101101100",
  36587=>"000000011",
  36588=>"111111111",
  36589=>"000000100",
  36590=>"111111111",
  36591=>"111111111",
  36592=>"011000000",
  36593=>"111111111",
  36594=>"100111100",
  36595=>"100100100",
  36596=>"110100110",
  36597=>"000100100",
  36598=>"011001011",
  36599=>"111111111",
  36600=>"111111100",
  36601=>"001001100",
  36602=>"111111111",
  36603=>"111111001",
  36604=>"000110111",
  36605=>"001001010",
  36606=>"001011010",
  36607=>"000000001",
  36608=>"111000000",
  36609=>"001011011",
  36610=>"000110000",
  36611=>"101110011",
  36612=>"011111011",
  36613=>"011001001",
  36614=>"111000000",
  36615=>"100111100",
  36616=>"111111011",
  36617=>"000000011",
  36618=>"000000000",
  36619=>"111111000",
  36620=>"100100000",
  36621=>"000000000",
  36622=>"111001000",
  36623=>"011010000",
  36624=>"001011001",
  36625=>"111100111",
  36626=>"100111110",
  36627=>"100100000",
  36628=>"000100111",
  36629=>"010000000",
  36630=>"011001001",
  36631=>"000000111",
  36632=>"111000000",
  36633=>"000100111",
  36634=>"010011110",
  36635=>"011000011",
  36636=>"011111001",
  36637=>"111111001",
  36638=>"110111111",
  36639=>"111100000",
  36640=>"111011111",
  36641=>"111000000",
  36642=>"100100000",
  36643=>"111011111",
  36644=>"111111111",
  36645=>"000000001",
  36646=>"110110110",
  36647=>"111111111",
  36648=>"011011111",
  36649=>"101001001",
  36650=>"011000000",
  36651=>"000010011",
  36652=>"001011001",
  36653=>"110110111",
  36654=>"000001111",
  36655=>"100000100",
  36656=>"011000000",
  36657=>"011011011",
  36658=>"000000011",
  36659=>"101000000",
  36660=>"110100000",
  36661=>"001011011",
  36662=>"001111111",
  36663=>"000000000",
  36664=>"101011111",
  36665=>"000000000",
  36666=>"101101101",
  36667=>"100000100",
  36668=>"001001000",
  36669=>"111111111",
  36670=>"111111111",
  36671=>"111111111",
  36672=>"000000000",
  36673=>"000000110",
  36674=>"001101111",
  36675=>"001011011",
  36676=>"000000000",
  36677=>"111001001",
  36678=>"001001101",
  36679=>"000000000",
  36680=>"111111000",
  36681=>"010111111",
  36682=>"111100111",
  36683=>"000100000",
  36684=>"000000111",
  36685=>"000000110",
  36686=>"111111111",
  36687=>"100000000",
  36688=>"001111001",
  36689=>"111100100",
  36690=>"000101000",
  36691=>"000110111",
  36692=>"000010000",
  36693=>"111111111",
  36694=>"000000001",
  36695=>"111111110",
  36696=>"111111001",
  36697=>"000000001",
  36698=>"011111000",
  36699=>"011000000",
  36700=>"101000100",
  36701=>"111100101",
  36702=>"001000100",
  36703=>"110000001",
  36704=>"111111111",
  36705=>"011011011",
  36706=>"001001000",
  36707=>"000001001",
  36708=>"010110110",
  36709=>"000000000",
  36710=>"111111000",
  36711=>"000000110",
  36712=>"001001011",
  36713=>"000010000",
  36714=>"001111011",
  36715=>"011001111",
  36716=>"110111111",
  36717=>"111010000",
  36718=>"000000000",
  36719=>"101111111",
  36720=>"000000111",
  36721=>"111111001",
  36722=>"111011100",
  36723=>"100000100",
  36724=>"001101111",
  36725=>"000000000",
  36726=>"101000000",
  36727=>"101111111",
  36728=>"111000000",
  36729=>"111111111",
  36730=>"111111111",
  36731=>"111100100",
  36732=>"000001101",
  36733=>"000000111",
  36734=>"110000000",
  36735=>"111001111",
  36736=>"100110000",
  36737=>"000011000",
  36738=>"111111111",
  36739=>"111111111",
  36740=>"000000111",
  36741=>"111111111",
  36742=>"011001011",
  36743=>"001100111",
  36744=>"011001000",
  36745=>"110010000",
  36746=>"000001011",
  36747=>"000111111",
  36748=>"000000000",
  36749=>"011000000",
  36750=>"000000000",
  36751=>"001011111",
  36752=>"001001001",
  36753=>"111001111",
  36754=>"010000000",
  36755=>"110110110",
  36756=>"000000000",
  36757=>"000111111",
  36758=>"111111000",
  36759=>"101111111",
  36760=>"000000000",
  36761=>"001001000",
  36762=>"111000000",
  36763=>"000011111",
  36764=>"001000111",
  36765=>"111111111",
  36766=>"011011001",
  36767=>"000000000",
  36768=>"000000000",
  36769=>"000011010",
  36770=>"110000000",
  36771=>"100000111",
  36772=>"110110000",
  36773=>"000000000",
  36774=>"011111111",
  36775=>"011011111",
  36776=>"110110000",
  36777=>"011011011",
  36778=>"101001111",
  36779=>"111110110",
  36780=>"000100100",
  36781=>"111011111",
  36782=>"101101001",
  36783=>"110111111",
  36784=>"111111000",
  36785=>"000010011",
  36786=>"111101100",
  36787=>"111111110",
  36788=>"011111111",
  36789=>"001111000",
  36790=>"000011011",
  36791=>"110100000",
  36792=>"100000000",
  36793=>"111111111",
  36794=>"000000100",
  36795=>"001010010",
  36796=>"111111111",
  36797=>"011011010",
  36798=>"111010000",
  36799=>"011011011",
  36800=>"000010111",
  36801=>"111000111",
  36802=>"011000000",
  36803=>"111000000",
  36804=>"000000000",
  36805=>"110110000",
  36806=>"000000000",
  36807=>"011011111",
  36808=>"111001010",
  36809=>"111110111",
  36810=>"000000010",
  36811=>"111111111",
  36812=>"100000000",
  36813=>"000000000",
  36814=>"011000000",
  36815=>"101111111",
  36816=>"111001111",
  36817=>"111000111",
  36818=>"000111111",
  36819=>"111111111",
  36820=>"001111110",
  36821=>"000000010",
  36822=>"010011000",
  36823=>"000000000",
  36824=>"111111110",
  36825=>"000011111",
  36826=>"100100111",
  36827=>"111111100",
  36828=>"000000001",
  36829=>"111100001",
  36830=>"000001000",
  36831=>"011001001",
  36832=>"011000000",
  36833=>"001000000",
  36834=>"000111000",
  36835=>"011011111",
  36836=>"000000111",
  36837=>"110000000",
  36838=>"000010110",
  36839=>"111111111",
  36840=>"001111111",
  36841=>"000001111",
  36842=>"111110100",
  36843=>"000000000",
  36844=>"111111111",
  36845=>"101111010",
  36846=>"000000111",
  36847=>"110000011",
  36848=>"111111100",
  36849=>"000000000",
  36850=>"000110010",
  36851=>"011000000",
  36852=>"111111111",
  36853=>"100000101",
  36854=>"000111110",
  36855=>"000010111",
  36856=>"010011000",
  36857=>"101100000",
  36858=>"001111111",
  36859=>"000000000",
  36860=>"010010000",
  36861=>"000111111",
  36862=>"011111110",
  36863=>"000001101",
  36864=>"111111100",
  36865=>"010111010",
  36866=>"101100101",
  36867=>"001000000",
  36868=>"001001111",
  36869=>"000001011",
  36870=>"000111111",
  36871=>"000000000",
  36872=>"000000111",
  36873=>"011011111",
  36874=>"111111011",
  36875=>"000110000",
  36876=>"110110000",
  36877=>"000000001",
  36878=>"011111111",
  36879=>"111000000",
  36880=>"000110110",
  36881=>"010011001",
  36882=>"000000011",
  36883=>"111111111",
  36884=>"100000000",
  36885=>"011010110",
  36886=>"001100100",
  36887=>"011111111",
  36888=>"111111101",
  36889=>"000011111",
  36890=>"000000000",
  36891=>"000000000",
  36892=>"000000001",
  36893=>"000000001",
  36894=>"111101100",
  36895=>"111111111",
  36896=>"101011110",
  36897=>"100111111",
  36898=>"110111111",
  36899=>"000000000",
  36900=>"000000000",
  36901=>"010110000",
  36902=>"101111111",
  36903=>"111000000",
  36904=>"111101111",
  36905=>"111111111",
  36906=>"000000000",
  36907=>"001001011",
  36908=>"000110111",
  36909=>"010110000",
  36910=>"000111111",
  36911=>"111101111",
  36912=>"011000000",
  36913=>"001101111",
  36914=>"001000000",
  36915=>"010010010",
  36916=>"111101100",
  36917=>"111100110",
  36918=>"111011011",
  36919=>"000000111",
  36920=>"001000000",
  36921=>"110111000",
  36922=>"110111110",
  36923=>"000000000",
  36924=>"000000000",
  36925=>"101000000",
  36926=>"000001000",
  36927=>"000000001",
  36928=>"111001000",
  36929=>"000000000",
  36930=>"110110111",
  36931=>"111111111",
  36932=>"000000000",
  36933=>"000001001",
  36934=>"111011000",
  36935=>"111111111",
  36936=>"011011001",
  36937=>"000011011",
  36938=>"111000000",
  36939=>"000000001",
  36940=>"000000100",
  36941=>"100100111",
  36942=>"011010000",
  36943=>"000010000",
  36944=>"110100110",
  36945=>"110011001",
  36946=>"011000000",
  36947=>"000000000",
  36948=>"001001000",
  36949=>"000000101",
  36950=>"000000000",
  36951=>"001001001",
  36952=>"111111001",
  36953=>"001000000",
  36954=>"000101111",
  36955=>"001011111",
  36956=>"000000000",
  36957=>"000000000",
  36958=>"000100110",
  36959=>"000000000",
  36960=>"111111111",
  36961=>"000000000",
  36962=>"010000000",
  36963=>"111111111",
  36964=>"110010111",
  36965=>"001000000",
  36966=>"110011001",
  36967=>"111111000",
  36968=>"000111111",
  36969=>"111001001",
  36970=>"100111000",
  36971=>"000000000",
  36972=>"111110010",
  36973=>"100101111",
  36974=>"110101111",
  36975=>"111111110",
  36976=>"000000000",
  36977=>"111000000",
  36978=>"011011011",
  36979=>"011001111",
  36980=>"001111111",
  36981=>"111001011",
  36982=>"000100111",
  36983=>"111111111",
  36984=>"001001000",
  36985=>"101100000",
  36986=>"000000000",
  36987=>"000000000",
  36988=>"001001000",
  36989=>"010111010",
  36990=>"101000000",
  36991=>"111111110",
  36992=>"111100000",
  36993=>"010000000",
  36994=>"111111111",
  36995=>"000000000",
  36996=>"100111111",
  36997=>"011001101",
  36998=>"100110111",
  36999=>"001001111",
  37000=>"000010010",
  37001=>"011001001",
  37002=>"001111111",
  37003=>"111111010",
  37004=>"110111001",
  37005=>"000000001",
  37006=>"111101000",
  37007=>"000000000",
  37008=>"000000000",
  37009=>"011111111",
  37010=>"000000000",
  37011=>"100000100",
  37012=>"000001111",
  37013=>"000000000",
  37014=>"010111110",
  37015=>"000000000",
  37016=>"101001111",
  37017=>"100000000",
  37018=>"000110000",
  37019=>"000000101",
  37020=>"111011001",
  37021=>"001000000",
  37022=>"111111000",
  37023=>"011111111",
  37024=>"111111111",
  37025=>"111100000",
  37026=>"000001111",
  37027=>"001100000",
  37028=>"001000000",
  37029=>"111111111",
  37030=>"000000000",
  37031=>"000011001",
  37032=>"000000000",
  37033=>"000001001",
  37034=>"000000000",
  37035=>"000001001",
  37036=>"000000010",
  37037=>"001001001",
  37038=>"011001000",
  37039=>"001001100",
  37040=>"000011111",
  37041=>"111111111",
  37042=>"011111111",
  37043=>"101000000",
  37044=>"000000100",
  37045=>"101000000",
  37046=>"000000000",
  37047=>"110111111",
  37048=>"001101111",
  37049=>"000010010",
  37050=>"001001000",
  37051=>"000000000",
  37052=>"001101000",
  37053=>"111111011",
  37054=>"111010001",
  37055=>"000111111",
  37056=>"011011111",
  37057=>"111001111",
  37058=>"110111111",
  37059=>"111000000",
  37060=>"110110000",
  37061=>"000000000",
  37062=>"000010111",
  37063=>"010011111",
  37064=>"000000000",
  37065=>"101101011",
  37066=>"000000000",
  37067=>"011111111",
  37068=>"000000000",
  37069=>"111000000",
  37070=>"111001000",
  37071=>"111111110",
  37072=>"001001011",
  37073=>"000000000",
  37074=>"000000000",
  37075=>"000010000",
  37076=>"111011001",
  37077=>"000000110",
  37078=>"111101111",
  37079=>"111111001",
  37080=>"111111111",
  37081=>"111010000",
  37082=>"010010011",
  37083=>"000011110",
  37084=>"110100000",
  37085=>"111000110",
  37086=>"000000000",
  37087=>"111111111",
  37088=>"111111111",
  37089=>"110011010",
  37090=>"111000000",
  37091=>"111111111",
  37092=>"111111100",
  37093=>"100100100",
  37094=>"110111111",
  37095=>"000000000",
  37096=>"100000000",
  37097=>"111111110",
  37098=>"001101011",
  37099=>"011001000",
  37100=>"000000000",
  37101=>"100000111",
  37102=>"011001000",
  37103=>"011111111",
  37104=>"101111111",
  37105=>"000001111",
  37106=>"000111111",
  37107=>"000000011",
  37108=>"111111111",
  37109=>"011000000",
  37110=>"100101111",
  37111=>"111001000",
  37112=>"000000000",
  37113=>"001001010",
  37114=>"000000001",
  37115=>"111111111",
  37116=>"001100100",
  37117=>"111111111",
  37118=>"101000000",
  37119=>"111111111",
  37120=>"111111110",
  37121=>"000000000",
  37122=>"111111111",
  37123=>"001011001",
  37124=>"101101001",
  37125=>"000000000",
  37126=>"000000000",
  37127=>"000000001",
  37128=>"111111111",
  37129=>"111000000",
  37130=>"000110110",
  37131=>"111111110",
  37132=>"110100100",
  37133=>"101100101",
  37134=>"000101111",
  37135=>"111001000",
  37136=>"000110000",
  37137=>"000000000",
  37138=>"000000000",
  37139=>"001110100",
  37140=>"000000000",
  37141=>"011011100",
  37142=>"111110010",
  37143=>"111111111",
  37144=>"000000000",
  37145=>"000001101",
  37146=>"000001111",
  37147=>"001000000",
  37148=>"110110000",
  37149=>"000111111",
  37150=>"111111010",
  37151=>"000000011",
  37152=>"000000000",
  37153=>"111111000",
  37154=>"111111110",
  37155=>"001001111",
  37156=>"111001011",
  37157=>"001011000",
  37158=>"011111111",
  37159=>"111110111",
  37160=>"010001111",
  37161=>"001000111",
  37162=>"011000001",
  37163=>"000000000",
  37164=>"111000000",
  37165=>"000100111",
  37166=>"000000000",
  37167=>"001000001",
  37168=>"100100000",
  37169=>"001000000",
  37170=>"001000000",
  37171=>"011001001",
  37172=>"111000000",
  37173=>"011111111",
  37174=>"000110111",
  37175=>"011111011",
  37176=>"111011011",
  37177=>"001000001",
  37178=>"101000000",
  37179=>"000000000",
  37180=>"111111011",
  37181=>"000111111",
  37182=>"011111111",
  37183=>"111111011",
  37184=>"111111111",
  37185=>"000001011",
  37186=>"111111111",
  37187=>"000010010",
  37188=>"111111001",
  37189=>"111111111",
  37190=>"000000000",
  37191=>"001111111",
  37192=>"111001011",
  37193=>"001011000",
  37194=>"010000000",
  37195=>"000000000",
  37196=>"000000000",
  37197=>"000000000",
  37198=>"111110100",
  37199=>"111111001",
  37200=>"111100110",
  37201=>"001000000",
  37202=>"111111011",
  37203=>"000001001",
  37204=>"111111111",
  37205=>"001011001",
  37206=>"011111111",
  37207=>"111000001",
  37208=>"101100111",
  37209=>"111000000",
  37210=>"001000000",
  37211=>"100100111",
  37212=>"000001111",
  37213=>"000000111",
  37214=>"110110000",
  37215=>"110000000",
  37216=>"111111111",
  37217=>"111111111",
  37218=>"101001001",
  37219=>"000000000",
  37220=>"111111111",
  37221=>"000000000",
  37222=>"110111111",
  37223=>"011011111",
  37224=>"000000000",
  37225=>"001111000",
  37226=>"001001001",
  37227=>"111111110",
  37228=>"101111111",
  37229=>"111111011",
  37230=>"000100000",
  37231=>"111011111",
  37232=>"111111111",
  37233=>"111001001",
  37234=>"000010011",
  37235=>"100000000",
  37236=>"111111111",
  37237=>"101111111",
  37238=>"100000001",
  37239=>"100000100",
  37240=>"000000000",
  37241=>"000000111",
  37242=>"001011111",
  37243=>"001000001",
  37244=>"000000100",
  37245=>"111111111",
  37246=>"000000000",
  37247=>"000000000",
  37248=>"001001001",
  37249=>"000000000",
  37250=>"110100110",
  37251=>"000110110",
  37252=>"111100100",
  37253=>"110111111",
  37254=>"011001001",
  37255=>"001000000",
  37256=>"000000000",
  37257=>"111111111",
  37258=>"110110000",
  37259=>"101111000",
  37260=>"000000001",
  37261=>"000000000",
  37262=>"111010000",
  37263=>"000000000",
  37264=>"111101100",
  37265=>"001000000",
  37266=>"111111111",
  37267=>"111111011",
  37268=>"110111111",
  37269=>"000000011",
  37270=>"000000000",
  37271=>"110100100",
  37272=>"111100111",
  37273=>"000000000",
  37274=>"111111111",
  37275=>"111011000",
  37276=>"111111110",
  37277=>"000000000",
  37278=>"001001000",
  37279=>"111111110",
  37280=>"101000101",
  37281=>"001001001",
  37282=>"100100100",
  37283=>"110001111",
  37284=>"000000001",
  37285=>"011111111",
  37286=>"001001001",
  37287=>"111000011",
  37288=>"000000111",
  37289=>"000000101",
  37290=>"000000100",
  37291=>"000000111",
  37292=>"111111010",
  37293=>"000000111",
  37294=>"000000001",
  37295=>"000000000",
  37296=>"110000000",
  37297=>"001001111",
  37298=>"000000000",
  37299=>"000100000",
  37300=>"001100000",
  37301=>"110110111",
  37302=>"000000000",
  37303=>"111110110",
  37304=>"111111001",
  37305=>"011011001",
  37306=>"001000000",
  37307=>"111111111",
  37308=>"000000000",
  37309=>"110000000",
  37310=>"000000110",
  37311=>"011011000",
  37312=>"000000001",
  37313=>"101001111",
  37314=>"010000000",
  37315=>"011000000",
  37316=>"000111111",
  37317=>"101100100",
  37318=>"110000000",
  37319=>"111111111",
  37320=>"001000001",
  37321=>"111111111",
  37322=>"000000101",
  37323=>"000000000",
  37324=>"111111111",
  37325=>"000000111",
  37326=>"111001001",
  37327=>"000111111",
  37328=>"000100000",
  37329=>"001101111",
  37330=>"111110100",
  37331=>"000011111",
  37332=>"000000001",
  37333=>"000000110",
  37334=>"110000000",
  37335=>"011011000",
  37336=>"000011010",
  37337=>"000000000",
  37338=>"000000000",
  37339=>"111111111",
  37340=>"000000000",
  37341=>"110100001",
  37342=>"101000000",
  37343=>"011111110",
  37344=>"000000000",
  37345=>"111101000",
  37346=>"000000001",
  37347=>"010110111",
  37348=>"101100000",
  37349=>"000000000",
  37350=>"010010010",
  37351=>"111101111",
  37352=>"000000000",
  37353=>"111000000",
  37354=>"001011111",
  37355=>"011000001",
  37356=>"110111111",
  37357=>"101111111",
  37358=>"000000010",
  37359=>"111111111",
  37360=>"001100111",
  37361=>"111111111",
  37362=>"011111011",
  37363=>"110111111",
  37364=>"000001000",
  37365=>"111111111",
  37366=>"001000000",
  37367=>"011011001",
  37368=>"111100000",
  37369=>"001001110",
  37370=>"001001101",
  37371=>"110100111",
  37372=>"111111111",
  37373=>"111111111",
  37374=>"111110000",
  37375=>"101101011",
  37376=>"001001111",
  37377=>"111001001",
  37378=>"010110000",
  37379=>"101101111",
  37380=>"010010000",
  37381=>"111111111",
  37382=>"001001000",
  37383=>"000000000",
  37384=>"111111010",
  37385=>"111111111",
  37386=>"100111111",
  37387=>"111111000",
  37388=>"001011011",
  37389=>"110111011",
  37390=>"000000111",
  37391=>"001000000",
  37392=>"000000000",
  37393=>"111111111",
  37394=>"000000000",
  37395=>"011111111",
  37396=>"111010110",
  37397=>"000111111",
  37398=>"000000000",
  37399=>"111100110",
  37400=>"011000000",
  37401=>"001011111",
  37402=>"000010000",
  37403=>"110000001",
  37404=>"100111111",
  37405=>"100111111",
  37406=>"100100000",
  37407=>"100000001",
  37408=>"110110110",
  37409=>"000110100",
  37410=>"000100001",
  37411=>"000110011",
  37412=>"000000000",
  37413=>"111111111",
  37414=>"000000111",
  37415=>"011000000",
  37416=>"000000000",
  37417=>"111011011",
  37418=>"111111111",
  37419=>"000000100",
  37420=>"111110000",
  37421=>"001001000",
  37422=>"010111111",
  37423=>"111111111",
  37424=>"110000000",
  37425=>"000000000",
  37426=>"000000100",
  37427=>"011011011",
  37428=>"011111111",
  37429=>"011011111",
  37430=>"111111111",
  37431=>"110010000",
  37432=>"110111110",
  37433=>"110111111",
  37434=>"001111110",
  37435=>"111011101",
  37436=>"000000111",
  37437=>"011111111",
  37438=>"111111111",
  37439=>"111111111",
  37440=>"010000001",
  37441=>"001101100",
  37442=>"100000000",
  37443=>"000010001",
  37444=>"111111111",
  37445=>"000100100",
  37446=>"111111111",
  37447=>"000011111",
  37448=>"100110110",
  37449=>"001001000",
  37450=>"111111111",
  37451=>"010110110",
  37452=>"000000000",
  37453=>"000010101",
  37454=>"111100100",
  37455=>"000001000",
  37456=>"111111111",
  37457=>"111011011",
  37458=>"001000000",
  37459=>"100100110",
  37460=>"011000000",
  37461=>"110100100",
  37462=>"000010011",
  37463=>"000000000",
  37464=>"111111111",
  37465=>"000000111",
  37466=>"011010010",
  37467=>"000001001",
  37468=>"111111111",
  37469=>"000000000",
  37470=>"000000001",
  37471=>"000000000",
  37472=>"000110110",
  37473=>"001000000",
  37474=>"000001000",
  37475=>"001000000",
  37476=>"001100100",
  37477=>"110110000",
  37478=>"000100110",
  37479=>"100100000",
  37480=>"111111000",
  37481=>"000000000",
  37482=>"110111111",
  37483=>"101010111",
  37484=>"110111111",
  37485=>"000000000",
  37486=>"111101001",
  37487=>"110111111",
  37488=>"000001001",
  37489=>"000001010",
  37490=>"101101001",
  37491=>"000011011",
  37492=>"011011110",
  37493=>"111100100",
  37494=>"111111111",
  37495=>"011000000",
  37496=>"111111111",
  37497=>"000000000",
  37498=>"100111111",
  37499=>"111111001",
  37500=>"001011011",
  37501=>"111111110",
  37502=>"000000000",
  37503=>"011111111",
  37504=>"111111111",
  37505=>"111110110",
  37506=>"111111111",
  37507=>"011000000",
  37508=>"111111011",
  37509=>"000000000",
  37510=>"111111111",
  37511=>"100100111",
  37512=>"001000000",
  37513=>"111111111",
  37514=>"010101000",
  37515=>"000100110",
  37516=>"111111111",
  37517=>"111111011",
  37518=>"111111111",
  37519=>"111000000",
  37520=>"000000000",
  37521=>"111111111",
  37522=>"011011001",
  37523=>"000000000",
  37524=>"110110000",
  37525=>"011000000",
  37526=>"000101000",
  37527=>"000000000",
  37528=>"111001011",
  37529=>"011011011",
  37530=>"110010010",
  37531=>"111101111",
  37532=>"010110111",
  37533=>"011011001",
  37534=>"000111110",
  37535=>"111010110",
  37536=>"110010111",
  37537=>"001111001",
  37538=>"010100000",
  37539=>"111111100",
  37540=>"001101111",
  37541=>"000000000",
  37542=>"001001001",
  37543=>"111111011",
  37544=>"111111000",
  37545=>"001011000",
  37546=>"111111111",
  37547=>"011010110",
  37548=>"111111111",
  37549=>"111111111",
  37550=>"000011011",
  37551=>"010000001",
  37552=>"001111101",
  37553=>"000000111",
  37554=>"001001000",
  37555=>"111111000",
  37556=>"110010000",
  37557=>"111100000",
  37558=>"111110111",
  37559=>"111111111",
  37560=>"000010111",
  37561=>"101001111",
  37562=>"110100111",
  37563=>"000010110",
  37564=>"111111011",
  37565=>"110110011",
  37566=>"001111111",
  37567=>"111111011",
  37568=>"111110111",
  37569=>"000000100",
  37570=>"011001011",
  37571=>"000010111",
  37572=>"111111111",
  37573=>"000000000",
  37574=>"111000001",
  37575=>"110111111",
  37576=>"111000011",
  37577=>"000000000",
  37578=>"111111011",
  37579=>"001001111",
  37580=>"000111111",
  37581=>"111111111",
  37582=>"000110111",
  37583=>"000111100",
  37584=>"111110101",
  37585=>"000001011",
  37586=>"000000011",
  37587=>"111000000",
  37588=>"111010011",
  37589=>"000000001",
  37590=>"111111111",
  37591=>"010111010",
  37592=>"111111111",
  37593=>"000000000",
  37594=>"111111100",
  37595=>"011111111",
  37596=>"000000000",
  37597=>"000000000",
  37598=>"000100110",
  37599=>"010110110",
  37600=>"001011110",
  37601=>"101101101",
  37602=>"111000000",
  37603=>"000000000",
  37604=>"111111111",
  37605=>"001001011",
  37606=>"111111111",
  37607=>"000000011",
  37608=>"000000000",
  37609=>"111111111",
  37610=>"000000000",
  37611=>"000111111",
  37612=>"111111111",
  37613=>"111111000",
  37614=>"000111000",
  37615=>"111111010",
  37616=>"110100111",
  37617=>"100000100",
  37618=>"110111111",
  37619=>"110111111",
  37620=>"000000000",
  37621=>"111100000",
  37622=>"011011000",
  37623=>"010000000",
  37624=>"111111111",
  37625=>"111111111",
  37626=>"000100111",
  37627=>"111111111",
  37628=>"111111110",
  37629=>"010011111",
  37630=>"001011011",
  37631=>"111110100",
  37632=>"111111111",
  37633=>"111111011",
  37634=>"001000000",
  37635=>"110111111",
  37636=>"000000000",
  37637=>"000110111",
  37638=>"000010000",
  37639=>"010100100",
  37640=>"000000000",
  37641=>"101111111",
  37642=>"111111111",
  37643=>"001011011",
  37644=>"010000000",
  37645=>"111111111",
  37646=>"111111011",
  37647=>"111111111",
  37648=>"110110110",
  37649=>"100111111",
  37650=>"000110000",
  37651=>"000000000",
  37652=>"000000011",
  37653=>"110100000",
  37654=>"111111100",
  37655=>"111111111",
  37656=>"111111111",
  37657=>"110001001",
  37658=>"111111001",
  37659=>"100101111",
  37660=>"000011000",
  37661=>"110010110",
  37662=>"010011011",
  37663=>"011000000",
  37664=>"100101111",
  37665=>"111111111",
  37666=>"000111010",
  37667=>"000000000",
  37668=>"000000000",
  37669=>"111110111",
  37670=>"101010010",
  37671=>"011111111",
  37672=>"111110111",
  37673=>"011111111",
  37674=>"000000011",
  37675=>"001100100",
  37676=>"100000000",
  37677=>"011001101",
  37678=>"101111000",
  37679=>"111000000",
  37680=>"000000100",
  37681=>"000000000",
  37682=>"000110111",
  37683=>"101111111",
  37684=>"111001000",
  37685=>"111111101",
  37686=>"100111111",
  37687=>"111111111",
  37688=>"111111010",
  37689=>"000000000",
  37690=>"110100000",
  37691=>"111111111",
  37692=>"010010010",
  37693=>"000100110",
  37694=>"100110101",
  37695=>"010000000",
  37696=>"000000001",
  37697=>"000000111",
  37698=>"111111000",
  37699=>"100111111",
  37700=>"110111111",
  37701=>"010010010",
  37702=>"111111111",
  37703=>"001001011",
  37704=>"000000000",
  37705=>"111111101",
  37706=>"011001001",
  37707=>"010010000",
  37708=>"111111111",
  37709=>"000000000",
  37710=>"111110111",
  37711=>"111111000",
  37712=>"001000100",
  37713=>"010011110",
  37714=>"111001111",
  37715=>"111111111",
  37716=>"000111110",
  37717=>"100100111",
  37718=>"010110100",
  37719=>"000000000",
  37720=>"000000000",
  37721=>"111111110",
  37722=>"000000011",
  37723=>"010011010",
  37724=>"111111001",
  37725=>"111111111",
  37726=>"011011001",
  37727=>"110110000",
  37728=>"110100000",
  37729=>"000000000",
  37730=>"010010010",
  37731=>"111111111",
  37732=>"000000111",
  37733=>"000000000",
  37734=>"111111011",
  37735=>"000110000",
  37736=>"011011011",
  37737=>"001100000",
  37738=>"000001000",
  37739=>"111001011",
  37740=>"100100100",
  37741=>"000000011",
  37742=>"111111111",
  37743=>"000000111",
  37744=>"100000000",
  37745=>"001000000",
  37746=>"111011011",
  37747=>"000000100",
  37748=>"000001100",
  37749=>"000000000",
  37750=>"110111000",
  37751=>"001001111",
  37752=>"000000000",
  37753=>"000000000",
  37754=>"110111110",
  37755=>"111111111",
  37756=>"111100000",
  37757=>"111111111",
  37758=>"111111111",
  37759=>"111111111",
  37760=>"111100100",
  37761=>"110110000",
  37762=>"011011011",
  37763=>"000000000",
  37764=>"111011000",
  37765=>"111111111",
  37766=>"101111111",
  37767=>"000000001",
  37768=>"111111111",
  37769=>"111111101",
  37770=>"111111111",
  37771=>"000000000",
  37772=>"001000001",
  37773=>"111111111",
  37774=>"010100000",
  37775=>"111111000",
  37776=>"010111010",
  37777=>"110110000",
  37778=>"000000000",
  37779=>"000001011",
  37780=>"111111111",
  37781=>"111111111",
  37782=>"000000000",
  37783=>"111001011",
  37784=>"110110001",
  37785=>"110110111",
  37786=>"010010000",
  37787=>"000000000",
  37788=>"100101111",
  37789=>"000011000",
  37790=>"111110111",
  37791=>"000000000",
  37792=>"110110100",
  37793=>"111111110",
  37794=>"010000000",
  37795=>"000111010",
  37796=>"110110011",
  37797=>"101111111",
  37798=>"111000000",
  37799=>"111111111",
  37800=>"111111111",
  37801=>"110110111",
  37802=>"000000000",
  37803=>"111000001",
  37804=>"111111110",
  37805=>"111110111",
  37806=>"111111110",
  37807=>"111111111",
  37808=>"111111100",
  37809=>"000000010",
  37810=>"011011111",
  37811=>"010010000",
  37812=>"100000111",
  37813=>"011011111",
  37814=>"011010000",
  37815=>"000000000",
  37816=>"000100100",
  37817=>"000000000",
  37818=>"111110000",
  37819=>"000000000",
  37820=>"000011000",
  37821=>"000000000",
  37822=>"011011001",
  37823=>"111111111",
  37824=>"101111111",
  37825=>"000001111",
  37826=>"111111111",
  37827=>"000000000",
  37828=>"000111111",
  37829=>"011111000",
  37830=>"111111111",
  37831=>"111010000",
  37832=>"000111111",
  37833=>"000100000",
  37834=>"000000000",
  37835=>"000010000",
  37836=>"100111111",
  37837=>"011111011",
  37838=>"110110111",
  37839=>"111110000",
  37840=>"001000000",
  37841=>"011011111",
  37842=>"111110111",
  37843=>"000011111",
  37844=>"111111111",
  37845=>"110110000",
  37846=>"011001111",
  37847=>"100110110",
  37848=>"100000001",
  37849=>"110110110",
  37850=>"100100000",
  37851=>"000001100",
  37852=>"000000110",
  37853=>"000000111",
  37854=>"111100000",
  37855=>"100101001",
  37856=>"010000000",
  37857=>"100000000",
  37858=>"000000100",
  37859=>"111111111",
  37860=>"000000000",
  37861=>"000000100",
  37862=>"111111111",
  37863=>"111111111",
  37864=>"000100001",
  37865=>"111111111",
  37866=>"111111111",
  37867=>"000000000",
  37868=>"000000001",
  37869=>"111111111",
  37870=>"111111111",
  37871=>"111111111",
  37872=>"110100111",
  37873=>"111110111",
  37874=>"011011000",
  37875=>"111111001",
  37876=>"110111111",
  37877=>"100100001",
  37878=>"000000000",
  37879=>"101101101",
  37880=>"101111111",
  37881=>"001000000",
  37882=>"011010000",
  37883=>"000000000",
  37884=>"011011000",
  37885=>"111111111",
  37886=>"011111111",
  37887=>"000000000",
  37888=>"111111111",
  37889=>"111111111",
  37890=>"101001111",
  37891=>"000000000",
  37892=>"000000000",
  37893=>"000000010",
  37894=>"000000000",
  37895=>"000000000",
  37896=>"011000000",
  37897=>"111011001",
  37898=>"010000111",
  37899=>"100000000",
  37900=>"000000000",
  37901=>"111111111",
  37902=>"000100110",
  37903=>"111111111",
  37904=>"111111111",
  37905=>"010001101",
  37906=>"111111111",
  37907=>"000111111",
  37908=>"001000000",
  37909=>"000000000",
  37910=>"000100100",
  37911=>"100100111",
  37912=>"001001101",
  37913=>"011110111",
  37914=>"001111111",
  37915=>"000000100",
  37916=>"000011111",
  37917=>"101111111",
  37918=>"111011011",
  37919=>"010001011",
  37920=>"111111110",
  37921=>"110100000",
  37922=>"000000100",
  37923=>"111111111",
  37924=>"000000100",
  37925=>"001111111",
  37926=>"110111111",
  37927=>"100110000",
  37928=>"000000000",
  37929=>"101101000",
  37930=>"111111111",
  37931=>"101000000",
  37932=>"001000000",
  37933=>"010110110",
  37934=>"100100100",
  37935=>"111100111",
  37936=>"111000101",
  37937=>"001111111",
  37938=>"111110000",
  37939=>"100100100",
  37940=>"101101100",
  37941=>"111111000",
  37942=>"100111111",
  37943=>"101111000",
  37944=>"001000000",
  37945=>"001000111",
  37946=>"111111111",
  37947=>"000000111",
  37948=>"000000000",
  37949=>"001001000",
  37950=>"000000000",
  37951=>"111111111",
  37952=>"111111111",
  37953=>"010110110",
  37954=>"000000000",
  37955=>"000000101",
  37956=>"000000100",
  37957=>"011011000",
  37958=>"010000000",
  37959=>"111111111",
  37960=>"011011011",
  37961=>"111001001",
  37962=>"111111111",
  37963=>"111011011",
  37964=>"011111111",
  37965=>"111011000",
  37966=>"001110111",
  37967=>"000111111",
  37968=>"000001011",
  37969=>"111111100",
  37970=>"111111000",
  37971=>"111111111",
  37972=>"000000000",
  37973=>"001000000",
  37974=>"000000000",
  37975=>"101111100",
  37976=>"100001000",
  37977=>"111000100",
  37978=>"111111111",
  37979=>"000000000",
  37980=>"000000000",
  37981=>"000111111",
  37982=>"000100110",
  37983=>"110110100",
  37984=>"000000110",
  37985=>"000100100",
  37986=>"000000000",
  37987=>"000000000",
  37988=>"000000111",
  37989=>"011011001",
  37990=>"111111111",
  37991=>"111000000",
  37992=>"000000000",
  37993=>"100000000",
  37994=>"000010010",
  37995=>"111111111",
  37996=>"000000000",
  37997=>"001001000",
  37998=>"001001111",
  37999=>"000000000",
  38000=>"000000000",
  38001=>"011010110",
  38002=>"111011011",
  38003=>"111000000",
  38004=>"000000000",
  38005=>"000000000",
  38006=>"000000000",
  38007=>"000000000",
  38008=>"110000000",
  38009=>"111111110",
  38010=>"000000000",
  38011=>"011111111",
  38012=>"100100100",
  38013=>"000000000",
  38014=>"111111111",
  38015=>"111101111",
  38016=>"000000000",
  38017=>"111101000",
  38018=>"110110111",
  38019=>"111111111",
  38020=>"111101111",
  38021=>"111111111",
  38022=>"000000111",
  38023=>"111011001",
  38024=>"111111111",
  38025=>"000000001",
  38026=>"001000000",
  38027=>"111111000",
  38028=>"100100100",
  38029=>"111111111",
  38030=>"000000000",
  38031=>"000010000",
  38032=>"111111111",
  38033=>"000000000",
  38034=>"000000000",
  38035=>"000001111",
  38036=>"000000110",
  38037=>"110000100",
  38038=>"100000011",
  38039=>"111110111",
  38040=>"000000000",
  38041=>"111111100",
  38042=>"111101111",
  38043=>"111110110",
  38044=>"100111110",
  38045=>"000000000",
  38046=>"111111111",
  38047=>"000000000",
  38048=>"111111111",
  38049=>"001101111",
  38050=>"001001111",
  38051=>"111111111",
  38052=>"100000000",
  38053=>"000001011",
  38054=>"000000000",
  38055=>"011011000",
  38056=>"100100000",
  38057=>"000000100",
  38058=>"111111111",
  38059=>"000110111",
  38060=>"011000000",
  38061=>"001001111",
  38062=>"111111111",
  38063=>"000000110",
  38064=>"000000000",
  38065=>"100000111",
  38066=>"101101111",
  38067=>"000000000",
  38068=>"111111111",
  38069=>"111000110",
  38070=>"001101101",
  38071=>"000000000",
  38072=>"111111110",
  38073=>"000000000",
  38074=>"100000000",
  38075=>"001111001",
  38076=>"000000101",
  38077=>"000000000",
  38078=>"111111111",
  38079=>"101011111",
  38080=>"000000000",
  38081=>"000000011",
  38082=>"111111111",
  38083=>"000000000",
  38084=>"001101001",
  38085=>"000000111",
  38086=>"100100000",
  38087=>"001100000",
  38088=>"100000000",
  38089=>"001000001",
  38090=>"111111111",
  38091=>"000001001",
  38092=>"111111111",
  38093=>"111011000",
  38094=>"000110110",
  38095=>"000110110",
  38096=>"101101111",
  38097=>"111110001",
  38098=>"111111001",
  38099=>"111111111",
  38100=>"111000000",
  38101=>"011110110",
  38102=>"110000100",
  38103=>"000101111",
  38104=>"001000000",
  38105=>"111110110",
  38106=>"000000111",
  38107=>"000000011",
  38108=>"000000000",
  38109=>"111000001",
  38110=>"111111111",
  38111=>"110100000",
  38112=>"111000000",
  38113=>"000000011",
  38114=>"010111100",
  38115=>"111000001",
  38116=>"110110110",
  38117=>"000100000",
  38118=>"101101000",
  38119=>"000000000",
  38120=>"110110000",
  38121=>"111110100",
  38122=>"111000000",
  38123=>"111110110",
  38124=>"000000001",
  38125=>"111111111",
  38126=>"000000111",
  38127=>"100100000",
  38128=>"110111111",
  38129=>"100000000",
  38130=>"111111111",
  38131=>"111000000",
  38132=>"100110000",
  38133=>"011001000",
  38134=>"100100000",
  38135=>"001000000",
  38136=>"111111111",
  38137=>"111111111",
  38138=>"001000000",
  38139=>"000000000",
  38140=>"000000110",
  38141=>"101101000",
  38142=>"000000000",
  38143=>"010000000",
  38144=>"000000000",
  38145=>"111011001",
  38146=>"110111000",
  38147=>"000000000",
  38148=>"000000000",
  38149=>"101000000",
  38150=>"000000000",
  38151=>"111110110",
  38152=>"000000000",
  38153=>"000000000",
  38154=>"111111111",
  38155=>"111111000",
  38156=>"000000000",
  38157=>"111000000",
  38158=>"000000000",
  38159=>"010110100",
  38160=>"111011010",
  38161=>"001000011",
  38162=>"111111111",
  38163=>"000001001",
  38164=>"111111111",
  38165=>"111111111",
  38166=>"100100110",
  38167=>"101111101",
  38168=>"111111101",
  38169=>"000000000",
  38170=>"000001000",
  38171=>"000000000",
  38172=>"110100110",
  38173=>"111101101",
  38174=>"111001001",
  38175=>"111001000",
  38176=>"111111001",
  38177=>"000000100",
  38178=>"111111111",
  38179=>"000111111",
  38180=>"000000000",
  38181=>"000110010",
  38182=>"101111111",
  38183=>"010110011",
  38184=>"111101001",
  38185=>"111111000",
  38186=>"101101001",
  38187=>"111111111",
  38188=>"000100010",
  38189=>"001111111",
  38190=>"111111000",
  38191=>"111111000",
  38192=>"000000101",
  38193=>"110111110",
  38194=>"111111111",
  38195=>"000000000",
  38196=>"000000000",
  38197=>"000110100",
  38198=>"101101101",
  38199=>"000000000",
  38200=>"011000000",
  38201=>"111101111",
  38202=>"111111011",
  38203=>"000111111",
  38204=>"100001111",
  38205=>"000000110",
  38206=>"000100110",
  38207=>"000010111",
  38208=>"000000000",
  38209=>"000000000",
  38210=>"000000000",
  38211=>"000010010",
  38212=>"111111100",
  38213=>"010000000",
  38214=>"000000000",
  38215=>"111101001",
  38216=>"001001111",
  38217=>"000000011",
  38218=>"111111111",
  38219=>"110100100",
  38220=>"101111111",
  38221=>"110111111",
  38222=>"001000000",
  38223=>"111111111",
  38224=>"000000100",
  38225=>"111011000",
  38226=>"100110111",
  38227=>"000000000",
  38228=>"111001101",
  38229=>"011010011",
  38230=>"000000010",
  38231=>"111111111",
  38232=>"111111111",
  38233=>"000000000",
  38234=>"000000000",
  38235=>"000000000",
  38236=>"001000000",
  38237=>"001000011",
  38238=>"111111111",
  38239=>"111110110",
  38240=>"111111111",
  38241=>"000000000",
  38242=>"110100110",
  38243=>"111111111",
  38244=>"000000000",
  38245=>"111100000",
  38246=>"111111111",
  38247=>"001101011",
  38248=>"111111111",
  38249=>"011111000",
  38250=>"000011111",
  38251=>"111111000",
  38252=>"011011111",
  38253=>"111111111",
  38254=>"000000000",
  38255=>"111010000",
  38256=>"000000010",
  38257=>"000000000",
  38258=>"000001000",
  38259=>"000000000",
  38260=>"111111111",
  38261=>"110000100",
  38262=>"111000000",
  38263=>"000000000",
  38264=>"111001001",
  38265=>"000000100",
  38266=>"001001011",
  38267=>"000011011",
  38268=>"011000000",
  38269=>"001000010",
  38270=>"100110010",
  38271=>"000000000",
  38272=>"000010011",
  38273=>"001000111",
  38274=>"100000000",
  38275=>"111111111",
  38276=>"011111111",
  38277=>"001101011",
  38278=>"000000000",
  38279=>"000000000",
  38280=>"111111111",
  38281=>"111111111",
  38282=>"100100000",
  38283=>"000000100",
  38284=>"101111111",
  38285=>"011111111",
  38286=>"000000110",
  38287=>"000000000",
  38288=>"000000000",
  38289=>"100000000",
  38290=>"011000000",
  38291=>"111001101",
  38292=>"110111000",
  38293=>"000011000",
  38294=>"100001101",
  38295=>"000000000",
  38296=>"000000110",
  38297=>"111111111",
  38298=>"111000000",
  38299=>"101100111",
  38300=>"110111100",
  38301=>"111111111",
  38302=>"000110011",
  38303=>"000000110",
  38304=>"011000000",
  38305=>"100001001",
  38306=>"111111101",
  38307=>"101101101",
  38308=>"111111111",
  38309=>"000000110",
  38310=>"000000111",
  38311=>"111111111",
  38312=>"000000000",
  38313=>"111111111",
  38314=>"111000110",
  38315=>"100000100",
  38316=>"011000001",
  38317=>"000000000",
  38318=>"001111111",
  38319=>"000000000",
  38320=>"110111111",
  38321=>"000001000",
  38322=>"011111111",
  38323=>"111001001",
  38324=>"000000000",
  38325=>"011011011",
  38326=>"100111111",
  38327=>"001011111",
  38328=>"111111000",
  38329=>"101001111",
  38330=>"000001000",
  38331=>"110110101",
  38332=>"111111000",
  38333=>"010111010",
  38334=>"101000000",
  38335=>"000000000",
  38336=>"000000000",
  38337=>"000111111",
  38338=>"111111000",
  38339=>"000000000",
  38340=>"000000100",
  38341=>"011111110",
  38342=>"111001000",
  38343=>"111000000",
  38344=>"100100000",
  38345=>"110110010",
  38346=>"000000000",
  38347=>"110111111",
  38348=>"000000000",
  38349=>"011000000",
  38350=>"001001101",
  38351=>"111100111",
  38352=>"000100111",
  38353=>"000001001",
  38354=>"000001001",
  38355=>"111111111",
  38356=>"001000000",
  38357=>"111111111",
  38358=>"000000000",
  38359=>"000000010",
  38360=>"111111111",
  38361=>"111111110",
  38362=>"111001001",
  38363=>"000010000",
  38364=>"000101111",
  38365=>"111101100",
  38366=>"100001000",
  38367=>"001001011",
  38368=>"100110000",
  38369=>"000000000",
  38370=>"111111111",
  38371=>"000000000",
  38372=>"111111111",
  38373=>"000001000",
  38374=>"000000011",
  38375=>"011000001",
  38376=>"000000000",
  38377=>"000000000",
  38378=>"111111000",
  38379=>"000010011",
  38380=>"000110111",
  38381=>"000000000",
  38382=>"000001000",
  38383=>"000000100",
  38384=>"000000000",
  38385=>"000000000",
  38386=>"100100111",
  38387=>"001000000",
  38388=>"000000000",
  38389=>"000000000",
  38390=>"000000111",
  38391=>"001001111",
  38392=>"000000001",
  38393=>"001001000",
  38394=>"100000111",
  38395=>"111111111",
  38396=>"010000011",
  38397=>"000000000",
  38398=>"000000000",
  38399=>"110110110",
  38400=>"110111100",
  38401=>"101000100",
  38402=>"111111001",
  38403=>"100000101",
  38404=>"100001111",
  38405=>"111111111",
  38406=>"111111000",
  38407=>"111100110",
  38408=>"011111111",
  38409=>"111111000",
  38410=>"011000111",
  38411=>"111011011",
  38412=>"000000000",
  38413=>"100100001",
  38414=>"000000001",
  38415=>"001000100",
  38416=>"111101111",
  38417=>"010110111",
  38418=>"001000111",
  38419=>"000111111",
  38420=>"000000000",
  38421=>"111111000",
  38422=>"000000111",
  38423=>"000000000",
  38424=>"111111111",
  38425=>"111111111",
  38426=>"111111011",
  38427=>"000000110",
  38428=>"010000000",
  38429=>"001111111",
  38430=>"000000000",
  38431=>"000000000",
  38432=>"000000101",
  38433=>"110111111",
  38434=>"000000110",
  38435=>"111001111",
  38436=>"111111111",
  38437=>"000000000",
  38438=>"001111111",
  38439=>"111000000",
  38440=>"001000000",
  38441=>"111000000",
  38442=>"000000000",
  38443=>"111111111",
  38444=>"111101111",
  38445=>"111000000",
  38446=>"110111111",
  38447=>"011000001",
  38448=>"000000001",
  38449=>"111001000",
  38450=>"110000000",
  38451=>"011011101",
  38452=>"011101100",
  38453=>"110000000",
  38454=>"111111000",
  38455=>"100000001",
  38456=>"010111000",
  38457=>"000000011",
  38458=>"000000001",
  38459=>"111000111",
  38460=>"111000000",
  38461=>"000000000",
  38462=>"111000000",
  38463=>"111011111",
  38464=>"000000000",
  38465=>"110111111",
  38466=>"100111111",
  38467=>"000110111",
  38468=>"011001111",
  38469=>"111000000",
  38470=>"111000111",
  38471=>"111111111",
  38472=>"011000001",
  38473=>"011001001",
  38474=>"111111111",
  38475=>"010111000",
  38476=>"111000000",
  38477=>"000000000",
  38478=>"000111111",
  38479=>"000000000",
  38480=>"000000000",
  38481=>"111000000",
  38482=>"100100100",
  38483=>"111111111",
  38484=>"000011111",
  38485=>"011000000",
  38486=>"001001111",
  38487=>"110010010",
  38488=>"010010010",
  38489=>"111001000",
  38490=>"111011001",
  38491=>"100111111",
  38492=>"000000000",
  38493=>"000000001",
  38494=>"111101111",
  38495=>"111111111",
  38496=>"111111000",
  38497=>"101111111",
  38498=>"111000111",
  38499=>"001000011",
  38500=>"000000000",
  38501=>"111000000",
  38502=>"111111110",
  38503=>"000000100",
  38504=>"000111010",
  38505=>"111111010",
  38506=>"000101001",
  38507=>"001111111",
  38508=>"101011000",
  38509=>"101000000",
  38510=>"000100111",
  38511=>"111101000",
  38512=>"000000011",
  38513=>"111111110",
  38514=>"111111001",
  38515=>"001111111",
  38516=>"111111110",
  38517=>"000111110",
  38518=>"000000000",
  38519=>"100100000",
  38520=>"111111111",
  38521=>"111001000",
  38522=>"000000111",
  38523=>"000000000",
  38524=>"101000000",
  38525=>"111111011",
  38526=>"111111111",
  38527=>"111000000",
  38528=>"000000000",
  38529=>"000011111",
  38530=>"111111111",
  38531=>"001111111",
  38532=>"111000000",
  38533=>"111001111",
  38534=>"111111000",
  38535=>"001000010",
  38536=>"101111100",
  38537=>"100111111",
  38538=>"000000000",
  38539=>"111111111",
  38540=>"011000000",
  38541=>"101000000",
  38542=>"101000000",
  38543=>"111000001",
  38544=>"111000000",
  38545=>"111111111",
  38546=>"000111111",
  38547=>"000000000",
  38548=>"000000111",
  38549=>"111111111",
  38550=>"111111111",
  38551=>"111111000",
  38552=>"001001001",
  38553=>"111000000",
  38554=>"001000000",
  38555=>"010000000",
  38556=>"001001000",
  38557=>"100110000",
  38558=>"000000101",
  38559=>"000000111",
  38560=>"000000000",
  38561=>"111000001",
  38562=>"111011000",
  38563=>"000000000",
  38564=>"000000000",
  38565=>"000000000",
  38566=>"111111110",
  38567=>"111110000",
  38568=>"111101000",
  38569=>"000000000",
  38570=>"101100111",
  38571=>"000000000",
  38572=>"000000110",
  38573=>"111111111",
  38574=>"000011011",
  38575=>"000000000",
  38576=>"111111111",
  38577=>"111100000",
  38578=>"111111111",
  38579=>"111111111",
  38580=>"000000110",
  38581=>"111111110",
  38582=>"001001000",
  38583=>"100000111",
  38584=>"111000000",
  38585=>"111111111",
  38586=>"111001000",
  38587=>"001001111",
  38588=>"101000100",
  38589=>"000000000",
  38590=>"001001111",
  38591=>"100100111",
  38592=>"001001101",
  38593=>"000000000",
  38594=>"111111000",
  38595=>"111000000",
  38596=>"111111111",
  38597=>"000111111",
  38598=>"000101111",
  38599=>"111111001",
  38600=>"111111111",
  38601=>"000001111",
  38602=>"000111111",
  38603=>"000000001",
  38604=>"101100111",
  38605=>"000000101",
  38606=>"000000000",
  38607=>"000000000",
  38608=>"000000011",
  38609=>"111000111",
  38610=>"111001111",
  38611=>"000000101",
  38612=>"111001001",
  38613=>"000001111",
  38614=>"111111111",
  38615=>"010000010",
  38616=>"000000000",
  38617=>"011111110",
  38618=>"111000000",
  38619=>"111111111",
  38620=>"101111100",
  38621=>"111000000",
  38622=>"000111111",
  38623=>"000000000",
  38624=>"010000000",
  38625=>"000011011",
  38626=>"111111100",
  38627=>"111000000",
  38628=>"111111101",
  38629=>"011111111",
  38630=>"000111111",
  38631=>"111101000",
  38632=>"101111111",
  38633=>"111000000",
  38634=>"000111111",
  38635=>"100001000",
  38636=>"000000111",
  38637=>"001111111",
  38638=>"100000111",
  38639=>"111111111",
  38640=>"000000011",
  38641=>"001001011",
  38642=>"111111000",
  38643=>"000000000",
  38644=>"111111000",
  38645=>"111111111",
  38646=>"010110000",
  38647=>"000010110",
  38648=>"111101101",
  38649=>"111111111",
  38650=>"000000000",
  38651=>"000010010",
  38652=>"000111001",
  38653=>"100100111",
  38654=>"111000000",
  38655=>"111000111",
  38656=>"111011111",
  38657=>"011011011",
  38658=>"111111001",
  38659=>"000000000",
  38660=>"001011011",
  38661=>"000000000",
  38662=>"111100100",
  38663=>"000000111",
  38664=>"000000000",
  38665=>"001000000",
  38666=>"111101100",
  38667=>"000111111",
  38668=>"000000110",
  38669=>"011000000",
  38670=>"000100000",
  38671=>"111111000",
  38672=>"000000111",
  38673=>"000000011",
  38674=>"111000001",
  38675=>"011100100",
  38676=>"111111001",
  38677=>"111111000",
  38678=>"001001001",
  38679=>"110111101",
  38680=>"110110000",
  38681=>"111111001",
  38682=>"100011000",
  38683=>"000000000",
  38684=>"000000000",
  38685=>"011111111",
  38686=>"000000011",
  38687=>"111111100",
  38688=>"111111000",
  38689=>"110110111",
  38690=>"111011000",
  38691=>"111111111",
  38692=>"100000000",
  38693=>"000000000",
  38694=>"111000000",
  38695=>"111111100",
  38696=>"111111111",
  38697=>"111000101",
  38698=>"001111111",
  38699=>"001111000",
  38700=>"111000000",
  38701=>"111111100",
  38702=>"111000101",
  38703=>"000111000",
  38704=>"000001011",
  38705=>"000000001",
  38706=>"111000000",
  38707=>"010000000",
  38708=>"111101011",
  38709=>"111111000",
  38710=>"000011011",
  38711=>"100110111",
  38712=>"011111000",
  38713=>"111000000",
  38714=>"001001000",
  38715=>"000001111",
  38716=>"111000000",
  38717=>"111111111",
  38718=>"000010110",
  38719=>"111111111",
  38720=>"000000000",
  38721=>"111111111",
  38722=>"000000000",
  38723=>"000000011",
  38724=>"000111111",
  38725=>"000111111",
  38726=>"000000000",
  38727=>"001001001",
  38728=>"100110111",
  38729=>"111111111",
  38730=>"111111111",
  38731=>"111111100",
  38732=>"111111111",
  38733=>"000001011",
  38734=>"000000000",
  38735=>"000111111",
  38736=>"000000000",
  38737=>"111101100",
  38738=>"011111000",
  38739=>"111111111",
  38740=>"000000000",
  38741=>"011010010",
  38742=>"000000000",
  38743=>"000000111",
  38744=>"111111001",
  38745=>"000000000",
  38746=>"111000000",
  38747=>"100000000",
  38748=>"110001111",
  38749=>"000000111",
  38750=>"101111111",
  38751=>"100110111",
  38752=>"000110111",
  38753=>"111111011",
  38754=>"010010000",
  38755=>"100000111",
  38756=>"110110100",
  38757=>"011111111",
  38758=>"000111111",
  38759=>"000000111",
  38760=>"100000011",
  38761=>"011111111",
  38762=>"000000111",
  38763=>"111000000",
  38764=>"100111111",
  38765=>"000000000",
  38766=>"000000010",
  38767=>"000000001",
  38768=>"000001111",
  38769=>"100000000",
  38770=>"111101101",
  38771=>"000000000",
  38772=>"111111000",
  38773=>"111011111",
  38774=>"000000111",
  38775=>"000001001",
  38776=>"111111111",
  38777=>"111110110",
  38778=>"111111111",
  38779=>"111111110",
  38780=>"111111010",
  38781=>"111110110",
  38782=>"100100000",
  38783=>"111111001",
  38784=>"111111111",
  38785=>"011100000",
  38786=>"101001000",
  38787=>"010011111",
  38788=>"000000111",
  38789=>"011111000",
  38790=>"000000000",
  38791=>"111011000",
  38792=>"001111111",
  38793=>"000000000",
  38794=>"000111111",
  38795=>"000101000",
  38796=>"111111111",
  38797=>"000011000",
  38798=>"000000000",
  38799=>"000000000",
  38800=>"000100111",
  38801=>"111111111",
  38802=>"100110111",
  38803=>"111000000",
  38804=>"101101111",
  38805=>"011101000",
  38806=>"111011011",
  38807=>"110110111",
  38808=>"110111111",
  38809=>"000111100",
  38810=>"111110111",
  38811=>"111111011",
  38812=>"100111111",
  38813=>"100000000",
  38814=>"111101001",
  38815=>"111001000",
  38816=>"000110111",
  38817=>"100111011",
  38818=>"111111111",
  38819=>"110111111",
  38820=>"111000111",
  38821=>"111111000",
  38822=>"100111111",
  38823=>"000111111",
  38824=>"001000000",
  38825=>"000000001",
  38826=>"101000000",
  38827=>"100011101",
  38828=>"111111100",
  38829=>"111111001",
  38830=>"000000000",
  38831=>"000000000",
  38832=>"001000000",
  38833=>"010010111",
  38834=>"001000000",
  38835=>"111111111",
  38836=>"111001000",
  38837=>"111100101",
  38838=>"111111111",
  38839=>"111111000",
  38840=>"010111010",
  38841=>"011111110",
  38842=>"100101111",
  38843=>"111111101",
  38844=>"111000000",
  38845=>"111111111",
  38846=>"111110010",
  38847=>"000000000",
  38848=>"100000000",
  38849=>"000111001",
  38850=>"111111101",
  38851=>"101100111",
  38852=>"111000100",
  38853=>"000000000",
  38854=>"110011001",
  38855=>"011110110",
  38856=>"001001101",
  38857=>"111000000",
  38858=>"100100001",
  38859=>"111101000",
  38860=>"110111000",
  38861=>"111000000",
  38862=>"000111111",
  38863=>"011000000",
  38864=>"000000000",
  38865=>"000000000",
  38866=>"000001111",
  38867=>"000101111",
  38868=>"111111111",
  38869=>"111000111",
  38870=>"100111100",
  38871=>"000000011",
  38872=>"111110001",
  38873=>"000100100",
  38874=>"111111000",
  38875=>"000001111",
  38876=>"000111001",
  38877=>"000111111",
  38878=>"111000000",
  38879=>"000000101",
  38880=>"001000111",
  38881=>"000000000",
  38882=>"111111010",
  38883=>"000111111",
  38884=>"000000000",
  38885=>"111111111",
  38886=>"111010100",
  38887=>"000111111",
  38888=>"110110011",
  38889=>"000000000",
  38890=>"010000000",
  38891=>"000000000",
  38892=>"111110111",
  38893=>"011111111",
  38894=>"000000000",
  38895=>"000000000",
  38896=>"111000000",
  38897=>"111111111",
  38898=>"111000110",
  38899=>"110110110",
  38900=>"000000100",
  38901=>"011001011",
  38902=>"000011111",
  38903=>"001000100",
  38904=>"110111000",
  38905=>"100000000",
  38906=>"000000110",
  38907=>"011111011",
  38908=>"000000111",
  38909=>"111101000",
  38910=>"000000000",
  38911=>"100111111",
  38912=>"111111111",
  38913=>"100000011",
  38914=>"111111111",
  38915=>"000000001",
  38916=>"011001001",
  38917=>"100110000",
  38918=>"000100100",
  38919=>"000000000",
  38920=>"000000000",
  38921=>"111111111",
  38922=>"110000000",
  38923=>"001111111",
  38924=>"000100000",
  38925=>"111111101",
  38926=>"001001000",
  38927=>"000000110",
  38928=>"010000100",
  38929=>"000000000",
  38930=>"011011111",
  38931=>"111111111",
  38932=>"111000100",
  38933=>"111111111",
  38934=>"000000001",
  38935=>"111110110",
  38936=>"111110110",
  38937=>"000000010",
  38938=>"111111111",
  38939=>"001101001",
  38940=>"000000000",
  38941=>"011000000",
  38942=>"001001001",
  38943=>"011000100",
  38944=>"000110100",
  38945=>"111111111",
  38946=>"111111110",
  38947=>"011000100",
  38948=>"111111100",
  38949=>"000000000",
  38950=>"000000011",
  38951=>"100000000",
  38952=>"111111011",
  38953=>"000000000",
  38954=>"010111111",
  38955=>"011011000",
  38956=>"000101111",
  38957=>"111111111",
  38958=>"111111000",
  38959=>"000000000",
  38960=>"111111111",
  38961=>"000000000",
  38962=>"001111111",
  38963=>"100100011",
  38964=>"000000000",
  38965=>"000011000",
  38966=>"111001111",
  38967=>"111001111",
  38968=>"110100110",
  38969=>"000000001",
  38970=>"111111111",
  38971=>"000000000",
  38972=>"111101000",
  38973=>"001000000",
  38974=>"011010011",
  38975=>"000000000",
  38976=>"000000000",
  38977=>"000000110",
  38978=>"111011011",
  38979=>"111111111",
  38980=>"110100100",
  38981=>"011011011",
  38982=>"000000001",
  38983=>"011111111",
  38984=>"000100000",
  38985=>"000000001",
  38986=>"111111111",
  38987=>"111011111",
  38988=>"000000000",
  38989=>"000000000",
  38990=>"110110100",
  38991=>"111111111",
  38992=>"000000001",
  38993=>"000000000",
  38994=>"011001111",
  38995=>"011000000",
  38996=>"000000000",
  38997=>"111001001",
  38998=>"111111111",
  38999=>"111111111",
  39000=>"011111100",
  39001=>"000000000",
  39002=>"011011111",
  39003=>"000000000",
  39004=>"000000000",
  39005=>"001111111",
  39006=>"011011111",
  39007=>"110100000",
  39008=>"000000000",
  39009=>"000000000",
  39010=>"111110000",
  39011=>"111111111",
  39012=>"011111110",
  39013=>"111111111",
  39014=>"000000000",
  39015=>"011001100",
  39016=>"000000000",
  39017=>"000000000",
  39018=>"111111111",
  39019=>"011011011",
  39020=>"001000101",
  39021=>"000000000",
  39022=>"010000000",
  39023=>"000000111",
  39024=>"010110110",
  39025=>"011010000",
  39026=>"000000000",
  39027=>"000000000",
  39028=>"000000000",
  39029=>"001000111",
  39030=>"000000000",
  39031=>"101111111",
  39032=>"001011111",
  39033=>"001000000",
  39034=>"000000000",
  39035=>"000000000",
  39036=>"110110110",
  39037=>"000000011",
  39038=>"111000000",
  39039=>"111111111",
  39040=>"001000101",
  39041=>"000001111",
  39042=>"111111111",
  39043=>"000000000",
  39044=>"111111111",
  39045=>"111111111",
  39046=>"000000000",
  39047=>"000000110",
  39048=>"100111001",
  39049=>"010111110",
  39050=>"111110100",
  39051=>"100001000",
  39052=>"000000000",
  39053=>"111101111",
  39054=>"000011111",
  39055=>"000001111",
  39056=>"000000000",
  39057=>"000000000",
  39058=>"111110111",
  39059=>"100000000",
  39060=>"111110011",
  39061=>"110000000",
  39062=>"111111111",
  39063=>"101000110",
  39064=>"010000000",
  39065=>"000000000",
  39066=>"111001000",
  39067=>"000110000",
  39068=>"110100111",
  39069=>"011000000",
  39070=>"111111111",
  39071=>"000000000",
  39072=>"000000000",
  39073=>"111111111",
  39074=>"111111111",
  39075=>"011000100",
  39076=>"000000000",
  39077=>"111111111",
  39078=>"000000110",
  39079=>"110111111",
  39080=>"111111101",
  39081=>"001001011",
  39082=>"010000000",
  39083=>"111111111",
  39084=>"000101111",
  39085=>"111111111",
  39086=>"011001001",
  39087=>"001001000",
  39088=>"000000000",
  39089=>"000000000",
  39090=>"000000000",
  39091=>"111101111",
  39092=>"000000001",
  39093=>"000000000",
  39094=>"000000000",
  39095=>"111111111",
  39096=>"111011111",
  39097=>"000000111",
  39098=>"111001101",
  39099=>"001001111",
  39100=>"111011000",
  39101=>"100000011",
  39102=>"000000000",
  39103=>"111111111",
  39104=>"110000000",
  39105=>"110000000",
  39106=>"000000000",
  39107=>"001001001",
  39108=>"111111111",
  39109=>"000001001",
  39110=>"111101101",
  39111=>"000000000",
  39112=>"000000000",
  39113=>"111000000",
  39114=>"111000000",
  39115=>"111111111",
  39116=>"100111111",
  39117=>"100111101",
  39118=>"000000001",
  39119=>"100101000",
  39120=>"111110110",
  39121=>"111111111",
  39122=>"111111001",
  39123=>"000000000",
  39124=>"000000111",
  39125=>"000000000",
  39126=>"111111111",
  39127=>"110110110",
  39128=>"001000000",
  39129=>"001000100",
  39130=>"111001101",
  39131=>"111110000",
  39132=>"000111111",
  39133=>"101111111",
  39134=>"000000000",
  39135=>"000000000",
  39136=>"000110110",
  39137=>"000000000",
  39138=>"111110100",
  39139=>"111101111",
  39140=>"000111110",
  39141=>"000000000",
  39142=>"111111001",
  39143=>"010000000",
  39144=>"000000000",
  39145=>"111111000",
  39146=>"111111111",
  39147=>"111111111",
  39148=>"011111111",
  39149=>"000010111",
  39150=>"000000000",
  39151=>"000000000",
  39152=>"001011111",
  39153=>"111111111",
  39154=>"111111001",
  39155=>"111100000",
  39156=>"111111111",
  39157=>"011001001",
  39158=>"000110110",
  39159=>"111111011",
  39160=>"000000000",
  39161=>"111011011",
  39162=>"001000000",
  39163=>"000000111",
  39164=>"000001001",
  39165=>"001001101",
  39166=>"110111111",
  39167=>"111111100",
  39168=>"111011001",
  39169=>"111111111",
  39170=>"000000000",
  39171=>"111110110",
  39172=>"101000000",
  39173=>"000000000",
  39174=>"001000000",
  39175=>"011011111",
  39176=>"000000000",
  39177=>"110000000",
  39178=>"001001001",
  39179=>"110110110",
  39180=>"111111111",
  39181=>"110111001",
  39182=>"000000000",
  39183=>"000000000",
  39184=>"111001000",
  39185=>"100000111",
  39186=>"001001111",
  39187=>"111111111",
  39188=>"111111111",
  39189=>"000000110",
  39190=>"111001001",
  39191=>"011011000",
  39192=>"000100100",
  39193=>"100100100",
  39194=>"000000111",
  39195=>"000001011",
  39196=>"000000000",
  39197=>"111111111",
  39198=>"000111111",
  39199=>"000110000",
  39200=>"111111111",
  39201=>"000110000",
  39202=>"111111111",
  39203=>"000000000",
  39204=>"011001000",
  39205=>"111111111",
  39206=>"110110111",
  39207=>"011010000",
  39208=>"000000000",
  39209=>"000000000",
  39210=>"000001111",
  39211=>"000000000",
  39212=>"110000111",
  39213=>"101111101",
  39214=>"111111111",
  39215=>"000000000",
  39216=>"001001101",
  39217=>"000000000",
  39218=>"000000000",
  39219=>"011110110",
  39220=>"010111011",
  39221=>"000000001",
  39222=>"000010001",
  39223=>"111111001",
  39224=>"000000000",
  39225=>"000000000",
  39226=>"001001000",
  39227=>"000000000",
  39228=>"000000000",
  39229=>"001011111",
  39230=>"010000000",
  39231=>"111111111",
  39232=>"000000000",
  39233=>"000000000",
  39234=>"111101111",
  39235=>"111111111",
  39236=>"111111100",
  39237=>"111111110",
  39238=>"010000000",
  39239=>"111110000",
  39240=>"000100100",
  39241=>"000000000",
  39242=>"111111011",
  39243=>"100000000",
  39244=>"000000100",
  39245=>"111000000",
  39246=>"111111111",
  39247=>"000000000",
  39248=>"000000110",
  39249=>"111111111",
  39250=>"000000000",
  39251=>"000000100",
  39252=>"011000111",
  39253=>"011011000",
  39254=>"000111111",
  39255=>"111111000",
  39256=>"111111111",
  39257=>"111000000",
  39258=>"000011111",
  39259=>"111000001",
  39260=>"101001001",
  39261=>"111111111",
  39262=>"000000000",
  39263=>"010011111",
  39264=>"100100000",
  39265=>"111111111",
  39266=>"001100110",
  39267=>"111111100",
  39268=>"110110000",
  39269=>"111111011",
  39270=>"000110100",
  39271=>"000000000",
  39272=>"100000001",
  39273=>"000000000",
  39274=>"000000000",
  39275=>"111111111",
  39276=>"111110100",
  39277=>"111001101",
  39278=>"100100100",
  39279=>"000100111",
  39280=>"000000111",
  39281=>"000000001",
  39282=>"100000110",
  39283=>"010000000",
  39284=>"111110000",
  39285=>"111111111",
  39286=>"001000100",
  39287=>"000000111",
  39288=>"111000000",
  39289=>"110110000",
  39290=>"000000000",
  39291=>"000000000",
  39292=>"001000100",
  39293=>"000111111",
  39294=>"000100100",
  39295=>"000000111",
  39296=>"110110000",
  39297=>"111111111",
  39298=>"110110000",
  39299=>"111111111",
  39300=>"111111111",
  39301=>"001111001",
  39302=>"000000000",
  39303=>"111110111",
  39304=>"000000110",
  39305=>"000100111",
  39306=>"111111000",
  39307=>"000011111",
  39308=>"000000000",
  39309=>"000111011",
  39310=>"000100111",
  39311=>"000000000",
  39312=>"111111111",
  39313=>"000000000",
  39314=>"001011000",
  39315=>"111010000",
  39316=>"010000000",
  39317=>"010000000",
  39318=>"111111101",
  39319=>"111000000",
  39320=>"000000011",
  39321=>"010111100",
  39322=>"100001000",
  39323=>"111111111",
  39324=>"011000000",
  39325=>"000010010",
  39326=>"001001001",
  39327=>"110111000",
  39328=>"001111111",
  39329=>"001000000",
  39330=>"100000001",
  39331=>"111011011",
  39332=>"001001001",
  39333=>"000111111",
  39334=>"000000111",
  39335=>"000001001",
  39336=>"000100011",
  39337=>"111011000",
  39338=>"111000000",
  39339=>"100000011",
  39340=>"000000000",
  39341=>"000100100",
  39342=>"101111111",
  39343=>"000000000",
  39344=>"111111111",
  39345=>"000000000",
  39346=>"111111111",
  39347=>"111000000",
  39348=>"000000001",
  39349=>"100110111",
  39350=>"111001101",
  39351=>"000000000",
  39352=>"111111111",
  39353=>"000000000",
  39354=>"000000100",
  39355=>"111000100",
  39356=>"000000011",
  39357=>"111111111",
  39358=>"100100100",
  39359=>"001001001",
  39360=>"100111111",
  39361=>"000001011",
  39362=>"111111111",
  39363=>"000100111",
  39364=>"111111111",
  39365=>"001101111",
  39366=>"111011000",
  39367=>"011000111",
  39368=>"000000000",
  39369=>"111111111",
  39370=>"000000000",
  39371=>"000000000",
  39372=>"111111111",
  39373=>"000000000",
  39374=>"000011000",
  39375=>"100100111",
  39376=>"000110010",
  39377=>"000000111",
  39378=>"000000000",
  39379=>"111111111",
  39380=>"001001000",
  39381=>"111100001",
  39382=>"111000001",
  39383=>"000100100",
  39384=>"001000110",
  39385=>"111001111",
  39386=>"111111111",
  39387=>"011111111",
  39388=>"000000000",
  39389=>"111000100",
  39390=>"111000001",
  39391=>"111111000",
  39392=>"110000000",
  39393=>"000100000",
  39394=>"000011001",
  39395=>"001000000",
  39396=>"000000100",
  39397=>"011011111",
  39398=>"000001011",
  39399=>"000000100",
  39400=>"000011111",
  39401=>"011000000",
  39402=>"011010110",
  39403=>"000000000",
  39404=>"001000000",
  39405=>"011001111",
  39406=>"000000000",
  39407=>"000000000",
  39408=>"111001000",
  39409=>"000000111",
  39410=>"000000000",
  39411=>"101000000",
  39412=>"100000000",
  39413=>"000000000",
  39414=>"111111111",
  39415=>"100000000",
  39416=>"000000000",
  39417=>"001001101",
  39418=>"110100000",
  39419=>"101111111",
  39420=>"000000111",
  39421=>"111111100",
  39422=>"000000000",
  39423=>"110000000",
  39424=>"111100101",
  39425=>"011000000",
  39426=>"111000111",
  39427=>"111001000",
  39428=>"111111111",
  39429=>"101100000",
  39430=>"011111011",
  39431=>"000000110",
  39432=>"111111010",
  39433=>"000000111",
  39434=>"111101000",
  39435=>"000000111",
  39436=>"000110111",
  39437=>"110110110",
  39438=>"001101011",
  39439=>"111011001",
  39440=>"100001000",
  39441=>"000011111",
  39442=>"000101111",
  39443=>"111100000",
  39444=>"101000000",
  39445=>"111111100",
  39446=>"101001000",
  39447=>"100111101",
  39448=>"000001111",
  39449=>"111001111",
  39450=>"000100111",
  39451=>"000000010",
  39452=>"010000001",
  39453=>"000100111",
  39454=>"100110100",
  39455=>"111111110",
  39456=>"100101111",
  39457=>"111111101",
  39458=>"000000110",
  39459=>"111111111",
  39460=>"000000000",
  39461=>"110000001",
  39462=>"001000000",
  39463=>"000001000",
  39464=>"000000000",
  39465=>"000010110",
  39466=>"000000000",
  39467=>"000000000",
  39468=>"111000000",
  39469=>"000110001",
  39470=>"000000000",
  39471=>"111111111",
  39472=>"000100110",
  39473=>"000000000",
  39474=>"000000000",
  39475=>"000001111",
  39476=>"000000100",
  39477=>"011011000",
  39478=>"111101011",
  39479=>"000100001",
  39480=>"101111000",
  39481=>"000000101",
  39482=>"000000110",
  39483=>"110111111",
  39484=>"000000000",
  39485=>"101000100",
  39486=>"111111100",
  39487=>"111000111",
  39488=>"111100111",
  39489=>"000100000",
  39490=>"100000001",
  39491=>"111001001",
  39492=>"000000111",
  39493=>"011111001",
  39494=>"111111000",
  39495=>"011000000",
  39496=>"000111111",
  39497=>"111100111",
  39498=>"111001000",
  39499=>"000000000",
  39500=>"011111110",
  39501=>"111111000",
  39502=>"001000000",
  39503=>"111001000",
  39504=>"101000000",
  39505=>"111110000",
  39506=>"000000000",
  39507=>"111111000",
  39508=>"011011010",
  39509=>"000000011",
  39510=>"111111111",
  39511=>"101000000",
  39512=>"000000000",
  39513=>"111000000",
  39514=>"000000000",
  39515=>"000001000",
  39516=>"000011111",
  39517=>"111000000",
  39518=>"000000000",
  39519=>"000011111",
  39520=>"110111111",
  39521=>"000110111",
  39522=>"111111111",
  39523=>"100111000",
  39524=>"111111111",
  39525=>"000111111",
  39526=>"110011111",
  39527=>"000000111",
  39528=>"111110100",
  39529=>"110000111",
  39530=>"000000001",
  39531=>"111000000",
  39532=>"111111010",
  39533=>"011000000",
  39534=>"000000000",
  39535=>"111111110",
  39536=>"001001001",
  39537=>"101000000",
  39538=>"010000000",
  39539=>"111111000",
  39540=>"000000000",
  39541=>"000110111",
  39542=>"100000100",
  39543=>"000001001",
  39544=>"100111111",
  39545=>"000000000",
  39546=>"111001000",
  39547=>"111111111",
  39548=>"111110110",
  39549=>"101011001",
  39550=>"001000000",
  39551=>"111100000",
  39552=>"111111111",
  39553=>"001000000",
  39554=>"111111000",
  39555=>"001001100",
  39556=>"000000000",
  39557=>"111111111",
  39558=>"111101100",
  39559=>"101000000",
  39560=>"000000000",
  39561=>"000001000",
  39562=>"111111011",
  39563=>"000001011",
  39564=>"100111111",
  39565=>"000000001",
  39566=>"101111100",
  39567=>"000000111",
  39568=>"001000000",
  39569=>"000000101",
  39570=>"000000010",
  39571=>"000011111",
  39572=>"111110000",
  39573=>"000000111",
  39574=>"000110111",
  39575=>"011000000",
  39576=>"011000000",
  39577=>"111111111",
  39578=>"111000000",
  39579=>"000110110",
  39580=>"100100111",
  39581=>"001001000",
  39582=>"111111001",
  39583=>"000101111",
  39584=>"000001000",
  39585=>"000100111",
  39586=>"111111111",
  39587=>"110111111",
  39588=>"111111011",
  39589=>"101000011",
  39590=>"111111111",
  39591=>"110010000",
  39592=>"100111001",
  39593=>"000010110",
  39594=>"101000000",
  39595=>"111011001",
  39596=>"000000101",
  39597=>"100101100",
  39598=>"001001001",
  39599=>"000101111",
  39600=>"111110000",
  39601=>"100101111",
  39602=>"111111111",
  39603=>"000000000",
  39604=>"000001000",
  39605=>"100000000",
  39606=>"010111111",
  39607=>"110111111",
  39608=>"000000000",
  39609=>"000100111",
  39610=>"111111011",
  39611=>"110111111",
  39612=>"111111111",
  39613=>"000000111",
  39614=>"000110111",
  39615=>"000000000",
  39616=>"111110000",
  39617=>"111111111",
  39618=>"011010111",
  39619=>"000000000",
  39620=>"111011111",
  39621=>"000000111",
  39622=>"000101000",
  39623=>"000000001",
  39624=>"110000000",
  39625=>"111001011",
  39626=>"000000000",
  39627=>"011001000",
  39628=>"101000100",
  39629=>"000000000",
  39630=>"100110111",
  39631=>"001000000",
  39632=>"111000000",
  39633=>"111111111",
  39634=>"000000000",
  39635=>"000111111",
  39636=>"001011011",
  39637=>"001111110",
  39638=>"011000000",
  39639=>"000000000",
  39640=>"000000000",
  39641=>"001111110",
  39642=>"000110111",
  39643=>"111011011",
  39644=>"101100111",
  39645=>"111001001",
  39646=>"000000000",
  39647=>"000000000",
  39648=>"111000000",
  39649=>"110111111",
  39650=>"111111000",
  39651=>"000000000",
  39652=>"000000010",
  39653=>"000001001",
  39654=>"111011000",
  39655=>"010111111",
  39656=>"111111011",
  39657=>"000000000",
  39658=>"101000000",
  39659=>"000000000",
  39660=>"011001111",
  39661=>"111000111",
  39662=>"011111111",
  39663=>"111100000",
  39664=>"011011001",
  39665=>"100110100",
  39666=>"111111011",
  39667=>"110000001",
  39668=>"000111111",
  39669=>"110110111",
  39670=>"001001001",
  39671=>"111111000",
  39672=>"001001000",
  39673=>"011000000",
  39674=>"111000000",
  39675=>"111111111",
  39676=>"000001000",
  39677=>"111111000",
  39678=>"001000000",
  39679=>"111001000",
  39680=>"000000111",
  39681=>"001101000",
  39682=>"000111111",
  39683=>"110000000",
  39684=>"000101111",
  39685=>"111100110",
  39686=>"000000000",
  39687=>"111111111",
  39688=>"000000111",
  39689=>"111000001",
  39690=>"101111111",
  39691=>"000001111",
  39692=>"111111000",
  39693=>"110110111",
  39694=>"000000001",
  39695=>"110111000",
  39696=>"000011000",
  39697=>"000100111",
  39698=>"000001111",
  39699=>"010000000",
  39700=>"000000010",
  39701=>"011111111",
  39702=>"000111111",
  39703=>"000000111",
  39704=>"000101111",
  39705=>"111111000",
  39706=>"101111011",
  39707=>"000111111",
  39708=>"000001001",
  39709=>"111101000",
  39710=>"000000000",
  39711=>"000001111",
  39712=>"100110000",
  39713=>"111111101",
  39714=>"111001000",
  39715=>"111101000",
  39716=>"100000000",
  39717=>"111000000",
  39718=>"111111111",
  39719=>"001101000",
  39720=>"111111111",
  39721=>"000111000",
  39722=>"000101111",
  39723=>"111100100",
  39724=>"111111000",
  39725=>"111111111",
  39726=>"000000000",
  39727=>"000000000",
  39728=>"000110011",
  39729=>"111000000",
  39730=>"100000000",
  39731=>"000111111",
  39732=>"000100111",
  39733=>"011000000",
  39734=>"000000000",
  39735=>"000110111",
  39736=>"111111001",
  39737=>"000000000",
  39738=>"111000000",
  39739=>"111010000",
  39740=>"000000000",
  39741=>"100111001",
  39742=>"111111111",
  39743=>"001111111",
  39744=>"110111000",
  39745=>"111111000",
  39746=>"010111111",
  39747=>"111111000",
  39748=>"111111000",
  39749=>"100100100",
  39750=>"000000111",
  39751=>"111111000",
  39752=>"000000000",
  39753=>"000111111",
  39754=>"001000111",
  39755=>"100100000",
  39756=>"000111111",
  39757=>"000011010",
  39758=>"111011011",
  39759=>"110001000",
  39760=>"001111011",
  39761=>"000011111",
  39762=>"100111000",
  39763=>"000000001",
  39764=>"111000111",
  39765=>"011011001",
  39766=>"111111111",
  39767=>"101000000",
  39768=>"000111111",
  39769=>"111111000",
  39770=>"000000000",
  39771=>"111000000",
  39772=>"001100100",
  39773=>"000111111",
  39774=>"000000001",
  39775=>"000011011",
  39776=>"000000000",
  39777=>"111100000",
  39778=>"001010000",
  39779=>"111111111",
  39780=>"110111110",
  39781=>"001001000",
  39782=>"001000111",
  39783=>"100000000",
  39784=>"001111101",
  39785=>"111111111",
  39786=>"000000000",
  39787=>"111100100",
  39788=>"011001000",
  39789=>"111111001",
  39790=>"000000000",
  39791=>"111111111",
  39792=>"000000000",
  39793=>"111111000",
  39794=>"111111101",
  39795=>"011111111",
  39796=>"001111111",
  39797=>"100111000",
  39798=>"000000110",
  39799=>"000000001",
  39800=>"111101010",
  39801=>"000111110",
  39802=>"111111111",
  39803=>"111011000",
  39804=>"110000000",
  39805=>"000000111",
  39806=>"000011010",
  39807=>"111111011",
  39808=>"000000001",
  39809=>"000111111",
  39810=>"110011001",
  39811=>"000000000",
  39812=>"000000000",
  39813=>"111111110",
  39814=>"111110100",
  39815=>"001000000",
  39816=>"000000000",
  39817=>"110111010",
  39818=>"000000100",
  39819=>"010110111",
  39820=>"000000000",
  39821=>"001111111",
  39822=>"100100110",
  39823=>"000111111",
  39824=>"000000011",
  39825=>"111111111",
  39826=>"000100000",
  39827=>"000000000",
  39828=>"111000000",
  39829=>"000011010",
  39830=>"110000000",
  39831=>"011011011",
  39832=>"000000000",
  39833=>"000100110",
  39834=>"110110010",
  39835=>"111001001",
  39836=>"111000000",
  39837=>"000000111",
  39838=>"101000000",
  39839=>"000000000",
  39840=>"011111111",
  39841=>"111110110",
  39842=>"111000000",
  39843=>"111111000",
  39844=>"101000000",
  39845=>"000111111",
  39846=>"000000000",
  39847=>"000000000",
  39848=>"111111111",
  39849=>"101000000",
  39850=>"111001011",
  39851=>"111111100",
  39852=>"001000000",
  39853=>"111111110",
  39854=>"111111000",
  39855=>"000000000",
  39856=>"111111001",
  39857=>"111010000",
  39858=>"110100100",
  39859=>"111111000",
  39860=>"110000000",
  39861=>"111111011",
  39862=>"000000100",
  39863=>"000000000",
  39864=>"000000001",
  39865=>"111111010",
  39866=>"110000000",
  39867=>"111111000",
  39868=>"111111000",
  39869=>"000011111",
  39870=>"111001000",
  39871=>"111111111",
  39872=>"000000000",
  39873=>"100000000",
  39874=>"111111111",
  39875=>"000000111",
  39876=>"100111111",
  39877=>"000000110",
  39878=>"000000001",
  39879=>"111111001",
  39880=>"101001000",
  39881=>"011100010",
  39882=>"011000010",
  39883=>"000000000",
  39884=>"000001000",
  39885=>"011000001",
  39886=>"111000001",
  39887=>"000000110",
  39888=>"000011010",
  39889=>"111111111",
  39890=>"000000001",
  39891=>"111100100",
  39892=>"000000111",
  39893=>"111111000",
  39894=>"001111111",
  39895=>"010111111",
  39896=>"111111111",
  39897=>"111111000",
  39898=>"000100111",
  39899=>"000100110",
  39900=>"000000111",
  39901=>"111101101",
  39902=>"001000000",
  39903=>"101111000",
  39904=>"100111111",
  39905=>"100100000",
  39906=>"000000000",
  39907=>"000000000",
  39908=>"110011001",
  39909=>"111010000",
  39910=>"001000000",
  39911=>"111000000",
  39912=>"000000100",
  39913=>"110111111",
  39914=>"011001000",
  39915=>"111011000",
  39916=>"111111111",
  39917=>"011001001",
  39918=>"101000000",
  39919=>"111101000",
  39920=>"111010001",
  39921=>"000111111",
  39922=>"000011111",
  39923=>"100100100",
  39924=>"011111111",
  39925=>"111111011",
  39926=>"000111111",
  39927=>"011011001",
  39928=>"000000000",
  39929=>"000001111",
  39930=>"111000000",
  39931=>"101100100",
  39932=>"001000100",
  39933=>"100111111",
  39934=>"111111110",
  39935=>"110110010",
  39936=>"111110110",
  39937=>"000000101",
  39938=>"101000000",
  39939=>"000010111",
  39940=>"000110100",
  39941=>"000001001",
  39942=>"111111111",
  39943=>"111111111",
  39944=>"100100111",
  39945=>"000000000",
  39946=>"011111111",
  39947=>"010100000",
  39948=>"011011111",
  39949=>"110111111",
  39950=>"000000000",
  39951=>"101111111",
  39952=>"000000000",
  39953=>"000000000",
  39954=>"111111111",
  39955=>"000000000",
  39956=>"000000000",
  39957=>"111100000",
  39958=>"111111000",
  39959=>"001000001",
  39960=>"111111111",
  39961=>"001001001",
  39962=>"000000000",
  39963=>"100100100",
  39964=>"001111111",
  39965=>"000000000",
  39966=>"100100000",
  39967=>"000000000",
  39968=>"000000000",
  39969=>"111111111",
  39970=>"111001001",
  39971=>"000000010",
  39972=>"111111111",
  39973=>"000000111",
  39974=>"011011000",
  39975=>"001000000",
  39976=>"111111001",
  39977=>"000110110",
  39978=>"001001000",
  39979=>"111111111",
  39980=>"000011011",
  39981=>"111111100",
  39982=>"000010011",
  39983=>"100100000",
  39984=>"000000000",
  39985=>"000101111",
  39986=>"001011111",
  39987=>"000000000",
  39988=>"111111000",
  39989=>"010110110",
  39990=>"010000000",
  39991=>"110110111",
  39992=>"011000000",
  39993=>"111110100",
  39994=>"001001111",
  39995=>"000011111",
  39996=>"111111011",
  39997=>"000111111",
  39998=>"111111110",
  39999=>"000001000",
  40000=>"000000001",
  40001=>"110110001",
  40002=>"110111111",
  40003=>"101111111",
  40004=>"000000100",
  40005=>"001001000",
  40006=>"111111111",
  40007=>"111111111",
  40008=>"001011011",
  40009=>"111111111",
  40010=>"111111111",
  40011=>"111111111",
  40012=>"000000100",
  40013=>"011011011",
  40014=>"000000000",
  40015=>"001111000",
  40016=>"000000000",
  40017=>"000000100",
  40018=>"011000001",
  40019=>"111111110",
  40020=>"001011000",
  40021=>"000000011",
  40022=>"001100000",
  40023=>"000000000",
  40024=>"111010100",
  40025=>"001000100",
  40026=>"110111111",
  40027=>"010111001",
  40028=>"000000000",
  40029=>"000000000",
  40030=>"001001000",
  40031=>"000000000",
  40032=>"000000100",
  40033=>"111111000",
  40034=>"101000100",
  40035=>"111011001",
  40036=>"110110111",
  40037=>"000000001",
  40038=>"000000000",
  40039=>"111111000",
  40040=>"111111111",
  40041=>"000000000",
  40042=>"111111111",
  40043=>"111111111",
  40044=>"111100000",
  40045=>"000000000",
  40046=>"000111111",
  40047=>"110110000",
  40048=>"000000111",
  40049=>"000000000",
  40050=>"000000000",
  40051=>"000000000",
  40052=>"111111111",
  40053=>"000000000",
  40054=>"000000000",
  40055=>"111111111",
  40056=>"101111111",
  40057=>"110110101",
  40058=>"111111000",
  40059=>"011010000",
  40060=>"000000001",
  40061=>"010010000",
  40062=>"111111111",
  40063=>"011001000",
  40064=>"110111111",
  40065=>"111111010",
  40066=>"110100100",
  40067=>"000111111",
  40068=>"111111111",
  40069=>"111111111",
  40070=>"111000111",
  40071=>"111111111",
  40072=>"011000111",
  40073=>"000000000",
  40074=>"111111111",
  40075=>"111111111",
  40076=>"010010110",
  40077=>"000110000",
  40078=>"000000100",
  40079=>"001011111",
  40080=>"111111111",
  40081=>"000011111",
  40082=>"000111111",
  40083=>"000000111",
  40084=>"111111111",
  40085=>"111111111",
  40086=>"000000111",
  40087=>"000000000",
  40088=>"000111111",
  40089=>"011011111",
  40090=>"100000110",
  40091=>"000000111",
  40092=>"000000000",
  40093=>"111001001",
  40094=>"000000000",
  40095=>"000000000",
  40096=>"101001100",
  40097=>"000000000",
  40098=>"000001111",
  40099=>"111110111",
  40100=>"111001011",
  40101=>"011111111",
  40102=>"000000000",
  40103=>"010011011",
  40104=>"010111000",
  40105=>"011001111",
  40106=>"111000000",
  40107=>"001001000",
  40108=>"111111000",
  40109=>"110000000",
  40110=>"011110111",
  40111=>"111011111",
  40112=>"000111111",
  40113=>"000100110",
  40114=>"111101111",
  40115=>"111111111",
  40116=>"110111111",
  40117=>"111111111",
  40118=>"000000110",
  40119=>"000000000",
  40120=>"111111111",
  40121=>"000000000",
  40122=>"111000011",
  40123=>"101001000",
  40124=>"111111111",
  40125=>"000000000",
  40126=>"111000000",
  40127=>"111111111",
  40128=>"111111100",
  40129=>"000001001",
  40130=>"111110111",
  40131=>"111111111",
  40132=>"000001000",
  40133=>"111111111",
  40134=>"100000010",
  40135=>"001100100",
  40136=>"000111000",
  40137=>"111011000",
  40138=>"111001001",
  40139=>"111100000",
  40140=>"001111111",
  40141=>"110110000",
  40142=>"111111111",
  40143=>"111110000",
  40144=>"000010111",
  40145=>"000000100",
  40146=>"111111111",
  40147=>"100110000",
  40148=>"000000000",
  40149=>"000000010",
  40150=>"000000000",
  40151=>"111110000",
  40152=>"111110110",
  40153=>"000000111",
  40154=>"010111110",
  40155=>"000000111",
  40156=>"000000000",
  40157=>"111111111",
  40158=>"111111111",
  40159=>"111111011",
  40160=>"111111111",
  40161=>"110111010",
  40162=>"000011000",
  40163=>"011001001",
  40164=>"111111111",
  40165=>"100100100",
  40166=>"000000000",
  40167=>"011111111",
  40168=>"000000000",
  40169=>"011000000",
  40170=>"000000000",
  40171=>"111111100",
  40172=>"111111110",
  40173=>"000000000",
  40174=>"111111111",
  40175=>"111001111",
  40176=>"111000101",
  40177=>"000000100",
  40178=>"010110110",
  40179=>"000000010",
  40180=>"111001111",
  40181=>"000000010",
  40182=>"111001001",
  40183=>"111001000",
  40184=>"111111111",
  40185=>"000000111",
  40186=>"001011001",
  40187=>"000000000",
  40188=>"111111111",
  40189=>"011011001",
  40190=>"101100000",
  40191=>"111111111",
  40192=>"001001000",
  40193=>"110110111",
  40194=>"111111000",
  40195=>"000000000",
  40196=>"101110100",
  40197=>"111000000",
  40198=>"110110000",
  40199=>"111001111",
  40200=>"001011000",
  40201=>"100100100",
  40202=>"101111011",
  40203=>"001010000",
  40204=>"000000101",
  40205=>"000000111",
  40206=>"101011110",
  40207=>"000000000",
  40208=>"111111111",
  40209=>"000110111",
  40210=>"111011001",
  40211=>"000000000",
  40212=>"000000111",
  40213=>"100000000",
  40214=>"011010010",
  40215=>"001101111",
  40216=>"000100100",
  40217=>"010111000",
  40218=>"111011000",
  40219=>"111111001",
  40220=>"000000000",
  40221=>"000000000",
  40222=>"000000011",
  40223=>"000111111",
  40224=>"000110011",
  40225=>"010011111",
  40226=>"100000000",
  40227=>"001011011",
  40228=>"000100111",
  40229=>"111100011",
  40230=>"000100111",
  40231=>"011000000",
  40232=>"111111111",
  40233=>"000000000",
  40234=>"000000000",
  40235=>"000111110",
  40236=>"101100000",
  40237=>"000100100",
  40238=>"111111111",
  40239=>"111111101",
  40240=>"001000000",
  40241=>"111111111",
  40242=>"000000001",
  40243=>"000000000",
  40244=>"000000000",
  40245=>"000100100",
  40246=>"000000000",
  40247=>"000000000",
  40248=>"000000000",
  40249=>"010110111",
  40250=>"100100000",
  40251=>"000000000",
  40252=>"011001000",
  40253=>"111111111",
  40254=>"111111101",
  40255=>"001001111",
  40256=>"000110111",
  40257=>"000000000",
  40258=>"000111111",
  40259=>"000000000",
  40260=>"000000110",
  40261=>"010111111",
  40262=>"000001000",
  40263=>"100101111",
  40264=>"000000000",
  40265=>"100110111",
  40266=>"011101111",
  40267=>"000100101",
  40268=>"011111011",
  40269=>"111011001",
  40270=>"000011111",
  40271=>"000001001",
  40272=>"001001001",
  40273=>"011011111",
  40274=>"110110110",
  40275=>"101101111",
  40276=>"111111001",
  40277=>"111111011",
  40278=>"111111111",
  40279=>"100000000",
  40280=>"000001001",
  40281=>"111011111",
  40282=>"000000001",
  40283=>"000011111",
  40284=>"010010000",
  40285=>"111111111",
  40286=>"010000111",
  40287=>"111111111",
  40288=>"011000000",
  40289=>"001000000",
  40290=>"000000000",
  40291=>"000000000",
  40292=>"111111111",
  40293=>"111101000",
  40294=>"000000001",
  40295=>"000101111",
  40296=>"000000110",
  40297=>"000000000",
  40298=>"101000000",
  40299=>"000001011",
  40300=>"010110000",
  40301=>"001000011",
  40302=>"100100110",
  40303=>"000000101",
  40304=>"001101001",
  40305=>"000000000",
  40306=>"111111111",
  40307=>"100100100",
  40308=>"111111111",
  40309=>"000000110",
  40310=>"110010000",
  40311=>"111111111",
  40312=>"010000000",
  40313=>"111100111",
  40314=>"111111111",
  40315=>"001101111",
  40316=>"111111111",
  40317=>"111111111",
  40318=>"110110110",
  40319=>"100111111",
  40320=>"001011011",
  40321=>"111001000",
  40322=>"000000000",
  40323=>"000001000",
  40324=>"000000000",
  40325=>"000000000",
  40326=>"011111001",
  40327=>"000000000",
  40328=>"000000000",
  40329=>"000000000",
  40330=>"001001001",
  40331=>"000000010",
  40332=>"111111111",
  40333=>"110110110",
  40334=>"000010000",
  40335=>"000000000",
  40336=>"000000000",
  40337=>"111111111",
  40338=>"011000000",
  40339=>"000110100",
  40340=>"001101111",
  40341=>"000010000",
  40342=>"111111111",
  40343=>"000001000",
  40344=>"000000000",
  40345=>"001000001",
  40346=>"000001000",
  40347=>"111101100",
  40348=>"000000000",
  40349=>"000000000",
  40350=>"000101000",
  40351=>"111111111",
  40352=>"111111100",
  40353=>"011011011",
  40354=>"000011011",
  40355=>"011000110",
  40356=>"000000110",
  40357=>"111111111",
  40358=>"011111101",
  40359=>"000000000",
  40360=>"000010000",
  40361=>"000111110",
  40362=>"000001111",
  40363=>"011111111",
  40364=>"000011111",
  40365=>"111111111",
  40366=>"000000111",
  40367=>"111111111",
  40368=>"010000000",
  40369=>"111111101",
  40370=>"111111111",
  40371=>"001000000",
  40372=>"000111001",
  40373=>"000000000",
  40374=>"000000000",
  40375=>"111111111",
  40376=>"000000111",
  40377=>"010011111",
  40378=>"011111111",
  40379=>"100100001",
  40380=>"000000000",
  40381=>"011111001",
  40382=>"111111000",
  40383=>"000000000",
  40384=>"111111000",
  40385=>"111111111",
  40386=>"000000111",
  40387=>"111111111",
  40388=>"001001000",
  40389=>"111110111",
  40390=>"111111111",
  40391=>"000110100",
  40392=>"000100111",
  40393=>"111111111",
  40394=>"000000000",
  40395=>"000000000",
  40396=>"100000000",
  40397=>"001001111",
  40398=>"100111110",
  40399=>"000111111",
  40400=>"110100111",
  40401=>"000111111",
  40402=>"100110111",
  40403=>"111111111",
  40404=>"010010110",
  40405=>"001011111",
  40406=>"111111111",
  40407=>"001111111",
  40408=>"000111011",
  40409=>"001001000",
  40410=>"010111111",
  40411=>"000000000",
  40412=>"000000011",
  40413=>"011001111",
  40414=>"001001111",
  40415=>"110110100",
  40416=>"000000000",
  40417=>"100110111",
  40418=>"000001111",
  40419=>"000000000",
  40420=>"000000001",
  40421=>"110000000",
  40422=>"000000110",
  40423=>"000000000",
  40424=>"111111000",
  40425=>"000000000",
  40426=>"000000000",
  40427=>"000000111",
  40428=>"111111101",
  40429=>"001001000",
  40430=>"000000000",
  40431=>"111110110",
  40432=>"100101111",
  40433=>"000110000",
  40434=>"111111111",
  40435=>"000000000",
  40436=>"111011111",
  40437=>"110111111",
  40438=>"000000100",
  40439=>"111110110",
  40440=>"000000000",
  40441=>"101001001",
  40442=>"000000000",
  40443=>"111000000",
  40444=>"111101100",
  40445=>"000000000",
  40446=>"000000000",
  40447=>"001011111",
  40448=>"000000110",
  40449=>"111111111",
  40450=>"111111111",
  40451=>"011111111",
  40452=>"111110111",
  40453=>"010000000",
  40454=>"000000000",
  40455=>"111111111",
  40456=>"011111111",
  40457=>"000000110",
  40458=>"000000000",
  40459=>"000000000",
  40460=>"000000000",
  40461=>"000001100",
  40462=>"000000110",
  40463=>"111111111",
  40464=>"111011000",
  40465=>"011111111",
  40466=>"111111111",
  40467=>"111010000",
  40468=>"111111111",
  40469=>"010010000",
  40470=>"001001001",
  40471=>"000001001",
  40472=>"110110111",
  40473=>"000010110",
  40474=>"111111111",
  40475=>"111110000",
  40476=>"111111111",
  40477=>"000000000",
  40478=>"111111111",
  40479=>"000000000",
  40480=>"000000110",
  40481=>"000000000",
  40482=>"111111000",
  40483=>"000000000",
  40484=>"111111111",
  40485=>"111110000",
  40486=>"111110111",
  40487=>"111111111",
  40488=>"001111100",
  40489=>"100111111",
  40490=>"000000100",
  40491=>"111000000",
  40492=>"111111010",
  40493=>"000000001",
  40494=>"111111111",
  40495=>"111111111",
  40496=>"000000100",
  40497=>"000101001",
  40498=>"011001000",
  40499=>"111100000",
  40500=>"000010000",
  40501=>"000000000",
  40502=>"000000000",
  40503=>"111111101",
  40504=>"111111111",
  40505=>"111111111",
  40506=>"000000000",
  40507=>"000000000",
  40508=>"111101101",
  40509=>"111111100",
  40510=>"000001101",
  40511=>"111111111",
  40512=>"000000000",
  40513=>"100101011",
  40514=>"110100100",
  40515=>"000100000",
  40516=>"100111111",
  40517=>"100000001",
  40518=>"000000000",
  40519=>"111000000",
  40520=>"000000000",
  40521=>"000000110",
  40522=>"110111110",
  40523=>"000110100",
  40524=>"111100100",
  40525=>"011111111",
  40526=>"000000000",
  40527=>"000101111",
  40528=>"000000000",
  40529=>"000000110",
  40530=>"000000000",
  40531=>"100100110",
  40532=>"000000000",
  40533=>"111111000",
  40534=>"100110110",
  40535=>"000000000",
  40536=>"111011000",
  40537=>"000000000",
  40538=>"001000110",
  40539=>"000000001",
  40540=>"010011011",
  40541=>"111111111",
  40542=>"000000000",
  40543=>"000000000",
  40544=>"100000010",
  40545=>"000000000",
  40546=>"100000111",
  40547=>"111111111",
  40548=>"111101100",
  40549=>"000000111",
  40550=>"110000000",
  40551=>"111111111",
  40552=>"100110111",
  40553=>"000000110",
  40554=>"000000111",
  40555=>"100000010",
  40556=>"100001001",
  40557=>"000000000",
  40558=>"000000000",
  40559=>"111110110",
  40560=>"111111111",
  40561=>"000000000",
  40562=>"000010000",
  40563=>"000000101",
  40564=>"111111111",
  40565=>"111000000",
  40566=>"000000100",
  40567=>"111011110",
  40568=>"000000000",
  40569=>"000101111",
  40570=>"001001000",
  40571=>"111010000",
  40572=>"100110000",
  40573=>"000101111",
  40574=>"000000000",
  40575=>"111111111",
  40576=>"000000000",
  40577=>"111110000",
  40578=>"000010111",
  40579=>"111111111",
  40580=>"110011000",
  40581=>"111111000",
  40582=>"111110000",
  40583=>"011000000",
  40584=>"111011000",
  40585=>"001001111",
  40586=>"001000001",
  40587=>"111111111",
  40588=>"110110111",
  40589=>"010111110",
  40590=>"000000000",
  40591=>"000100110",
  40592=>"111111111",
  40593=>"000000000",
  40594=>"111111000",
  40595=>"111111111",
  40596=>"000100110",
  40597=>"010110010",
  40598=>"100111111",
  40599=>"111111011",
  40600=>"111101100",
  40601=>"110111111",
  40602=>"111111111",
  40603=>"000000000",
  40604=>"111111100",
  40605=>"000000000",
  40606=>"111110000",
  40607=>"111111111",
  40608=>"000000000",
  40609=>"111000000",
  40610=>"011011111",
  40611=>"000000000",
  40612=>"000000000",
  40613=>"001001011",
  40614=>"110111111",
  40615=>"000011001",
  40616=>"111111010",
  40617=>"111111111",
  40618=>"000000000",
  40619=>"111001011",
  40620=>"111110111",
  40621=>"000000000",
  40622=>"111111111",
  40623=>"000111110",
  40624=>"100111111",
  40625=>"100000000",
  40626=>"111111110",
  40627=>"000111010",
  40628=>"000000001",
  40629=>"001110000",
  40630=>"010110110",
  40631=>"000000000",
  40632=>"000000000",
  40633=>"111101000",
  40634=>"000000000",
  40635=>"001000100",
  40636=>"000000000",
  40637=>"000000110",
  40638=>"111111111",
  40639=>"000010110",
  40640=>"000000000",
  40641=>"010101110",
  40642=>"111111111",
  40643=>"000110111",
  40644=>"000000000",
  40645=>"111000000",
  40646=>"000000000",
  40647=>"011000111",
  40648=>"000001111",
  40649=>"011011111",
  40650=>"000000000",
  40651=>"000000000",
  40652=>"000000000",
  40653=>"010000000",
  40654=>"111111111",
  40655=>"000000000",
  40656=>"011000000",
  40657=>"000000000",
  40658=>"011111111",
  40659=>"111111111",
  40660=>"000000000",
  40661=>"100100000",
  40662=>"001011000",
  40663=>"000100000",
  40664=>"100110110",
  40665=>"000000100",
  40666=>"111111000",
  40667=>"001111111",
  40668=>"000100000",
  40669=>"011001011",
  40670=>"111110111",
  40671=>"000000000",
  40672=>"000000000",
  40673=>"000000110",
  40674=>"000010000",
  40675=>"101000001",
  40676=>"000000010",
  40677=>"000000000",
  40678=>"100001111",
  40679=>"000000101",
  40680=>"111111100",
  40681=>"000000000",
  40682=>"111101111",
  40683=>"111111011",
  40684=>"111111111",
  40685=>"000111010",
  40686=>"111111011",
  40687=>"000010110",
  40688=>"110111111",
  40689=>"001000101",
  40690=>"111111111",
  40691=>"000000000",
  40692=>"000111111",
  40693=>"000000000",
  40694=>"011011011",
  40695=>"111111000",
  40696=>"111011111",
  40697=>"000000011",
  40698=>"001011111",
  40699=>"000000000",
  40700=>"111111111",
  40701=>"000000000",
  40702=>"000000000",
  40703=>"100000001",
  40704=>"000000000",
  40705=>"110100100",
  40706=>"100000000",
  40707=>"111111111",
  40708=>"000000001",
  40709=>"011001111",
  40710=>"111101000",
  40711=>"110111111",
  40712=>"111100111",
  40713=>"000010111",
  40714=>"100100100",
  40715=>"000000000",
  40716=>"111111111",
  40717=>"000011010",
  40718=>"000110010",
  40719=>"000000000",
  40720=>"000000000",
  40721=>"110000000",
  40722=>"011010000",
  40723=>"110000000",
  40724=>"000000000",
  40725=>"000000000",
  40726=>"110100000",
  40727=>"011111011",
  40728=>"111111111",
  40729=>"111110111",
  40730=>"111010000",
  40731=>"000000000",
  40732=>"010111111",
  40733=>"010010010",
  40734=>"111111111",
  40735=>"011010010",
  40736=>"000000000",
  40737=>"110010111",
  40738=>"000000000",
  40739=>"110111111",
  40740=>"110111100",
  40741=>"111001001",
  40742=>"000000001",
  40743=>"010000100",
  40744=>"110000000",
  40745=>"100111111",
  40746=>"111100111",
  40747=>"111100000",
  40748=>"000000000",
  40749=>"110110110",
  40750=>"111111111",
  40751=>"000100111",
  40752=>"000000000",
  40753=>"000000111",
  40754=>"010111000",
  40755=>"001000100",
  40756=>"111110110",
  40757=>"001011011",
  40758=>"000000000",
  40759=>"000000000",
  40760=>"000000000",
  40761=>"011000100",
  40762=>"000000000",
  40763=>"001000000",
  40764=>"111111111",
  40765=>"001010111",
  40766=>"100100100",
  40767=>"000000111",
  40768=>"111000100",
  40769=>"111111111",
  40770=>"111111111",
  40771=>"111100100",
  40772=>"110111111",
  40773=>"111110110",
  40774=>"000000011",
  40775=>"100000000",
  40776=>"111111010",
  40777=>"000000000",
  40778=>"110000001",
  40779=>"011111111",
  40780=>"000000011",
  40781=>"000100100",
  40782=>"000100111",
  40783=>"000000000",
  40784=>"000110110",
  40785=>"000000000",
  40786=>"010111010",
  40787=>"000001000",
  40788=>"000000000",
  40789=>"001001001",
  40790=>"101111010",
  40791=>"100000000",
  40792=>"001000001",
  40793=>"111011011",
  40794=>"000010001",
  40795=>"000000000",
  40796=>"000000000",
  40797=>"011011000",
  40798=>"100000000",
  40799=>"100100111",
  40800=>"110000000",
  40801=>"111111111",
  40802=>"111111110",
  40803=>"000111111",
  40804=>"000100101",
  40805=>"000000000",
  40806=>"111111111",
  40807=>"111111111",
  40808=>"111111111",
  40809=>"100000110",
  40810=>"111111111",
  40811=>"010011000",
  40812=>"110000001",
  40813=>"000011011",
  40814=>"111111111",
  40815=>"100000100",
  40816=>"111110000",
  40817=>"000000000",
  40818=>"010111111",
  40819=>"111111111",
  40820=>"111111111",
  40821=>"111111111",
  40822=>"000000000",
  40823=>"111101000",
  40824=>"011010110",
  40825=>"000110110",
  40826=>"010010010",
  40827=>"111110111",
  40828=>"011111111",
  40829=>"010000000",
  40830=>"010110111",
  40831=>"111111111",
  40832=>"011001111",
  40833=>"111011000",
  40834=>"001001001",
  40835=>"111111111",
  40836=>"010010000",
  40837=>"000000001",
  40838=>"010010100",
  40839=>"111111111",
  40840=>"000000000",
  40841=>"000000000",
  40842=>"000000000",
  40843=>"111111111",
  40844=>"000000111",
  40845=>"001000110",
  40846=>"000000110",
  40847=>"000000010",
  40848=>"000000000",
  40849=>"000000011",
  40850=>"011011111",
  40851=>"111111111",
  40852=>"000000000",
  40853=>"000000000",
  40854=>"111011001",
  40855=>"110110111",
  40856=>"010000000",
  40857=>"000000000",
  40858=>"111111111",
  40859=>"111111000",
  40860=>"111000001",
  40861=>"111111111",
  40862=>"000000000",
  40863=>"111110110",
  40864=>"001000000",
  40865=>"010110110",
  40866=>"111111111",
  40867=>"000111011",
  40868=>"111111110",
  40869=>"111011000",
  40870=>"011111111",
  40871=>"000000110",
  40872=>"000000001",
  40873=>"000111111",
  40874=>"100000000",
  40875=>"011000001",
  40876=>"000000000",
  40877=>"000000000",
  40878=>"000100100",
  40879=>"011111111",
  40880=>"111011011",
  40881=>"011111111",
  40882=>"000000000",
  40883=>"000000000",
  40884=>"000000000",
  40885=>"111111110",
  40886=>"110010111",
  40887=>"111011010",
  40888=>"111111111",
  40889=>"011011011",
  40890=>"000000000",
  40891=>"001101111",
  40892=>"111011011",
  40893=>"111111111",
  40894=>"000000000",
  40895=>"111111111",
  40896=>"111111111",
  40897=>"000000111",
  40898=>"111111111",
  40899=>"111111111",
  40900=>"111111100",
  40901=>"101001011",
  40902=>"111111111",
  40903=>"110110110",
  40904=>"000101111",
  40905=>"111111111",
  40906=>"000000000",
  40907=>"010011011",
  40908=>"110000000",
  40909=>"000111111",
  40910=>"111111111",
  40911=>"011011011",
  40912=>"111111111",
  40913=>"111111111",
  40914=>"111111000",
  40915=>"111111111",
  40916=>"000000000",
  40917=>"101111100",
  40918=>"001000000",
  40919=>"000000000",
  40920=>"111111111",
  40921=>"010011111",
  40922=>"011000000",
  40923=>"111111111",
  40924=>"000000000",
  40925=>"111111110",
  40926=>"000000000",
  40927=>"111111111",
  40928=>"111111111",
  40929=>"010110110",
  40930=>"110111111",
  40931=>"110100000",
  40932=>"111111100",
  40933=>"001111001",
  40934=>"000000110",
  40935=>"000001000",
  40936=>"111111111",
  40937=>"111111111",
  40938=>"011000000",
  40939=>"111111111",
  40940=>"000000100",
  40941=>"001000000",
  40942=>"111111111",
  40943=>"111111111",
  40944=>"000000000",
  40945=>"000011001",
  40946=>"001000000",
  40947=>"000000000",
  40948=>"100100000",
  40949=>"100000000",
  40950=>"111100100",
  40951=>"011111100",
  40952=>"000000000",
  40953=>"001001001",
  40954=>"110110000",
  40955=>"010011000",
  40956=>"000100111",
  40957=>"011000000",
  40958=>"111111111",
  40959=>"000000000",
  40960=>"111111111",
  40961=>"000000111",
  40962=>"110100111",
  40963=>"000100110",
  40964=>"000110111",
  40965=>"001001011",
  40966=>"001000000",
  40967=>"111111111",
  40968=>"000000110",
  40969=>"011010011",
  40970=>"000000000",
  40971=>"111000111",
  40972=>"001001001",
  40973=>"000001111",
  40974=>"000001000",
  40975=>"000000000",
  40976=>"110100110",
  40977=>"000110111",
  40978=>"111110110",
  40979=>"111110000",
  40980=>"010111111",
  40981=>"111010111",
  40982=>"000000111",
  40983=>"111111111",
  40984=>"100111111",
  40985=>"001000000",
  40986=>"101000011",
  40987=>"111100101",
  40988=>"101000111",
  40989=>"111111110",
  40990=>"111110000",
  40991=>"001001000",
  40992=>"111011001",
  40993=>"100100110",
  40994=>"111111110",
  40995=>"111111101",
  40996=>"001111001",
  40997=>"101000101",
  40998=>"100000000",
  40999=>"000000001",
  41000=>"111011101",
  41001=>"010000010",
  41002=>"110111111",
  41003=>"111111111",
  41004=>"000011111",
  41005=>"000111111",
  41006=>"111110110",
  41007=>"000000000",
  41008=>"111111111",
  41009=>"100111111",
  41010=>"001111111",
  41011=>"011111111",
  41012=>"011010000",
  41013=>"000000001",
  41014=>"000110110",
  41015=>"000000110",
  41016=>"111111111",
  41017=>"011000110",
  41018=>"000110000",
  41019=>"000110100",
  41020=>"111100000",
  41021=>"000001000",
  41022=>"000011111",
  41023=>"000000000",
  41024=>"111000000",
  41025=>"001011111",
  41026=>"001111111",
  41027=>"001011110",
  41028=>"000100000",
  41029=>"011011000",
  41030=>"000011111",
  41031=>"010000100",
  41032=>"011011000",
  41033=>"000000000",
  41034=>"111011011",
  41035=>"010000000",
  41036=>"000111111",
  41037=>"000000000",
  41038=>"111000000",
  41039=>"111001000",
  41040=>"000000000",
  41041=>"111111111",
  41042=>"000000000",
  41043=>"000000000",
  41044=>"111010100",
  41045=>"111110100",
  41046=>"111001111",
  41047=>"110111111",
  41048=>"100100100",
  41049=>"000111111",
  41050=>"110000000",
  41051=>"001000000",
  41052=>"110111111",
  41053=>"111111111",
  41054=>"000110000",
  41055=>"000100111",
  41056=>"100000000",
  41057=>"000000111",
  41058=>"000111111",
  41059=>"000010110",
  41060=>"111110100",
  41061=>"000100110",
  41062=>"111110000",
  41063=>"100000000",
  41064=>"000100000",
  41065=>"000001111",
  41066=>"110100111",
  41067=>"000110000",
  41068=>"010111111",
  41069=>"001111111",
  41070=>"000100111",
  41071=>"111110000",
  41072=>"011111111",
  41073=>"100000000",
  41074=>"101000000",
  41075=>"001000000",
  41076=>"100111000",
  41077=>"110111001",
  41078=>"000000000",
  41079=>"111111111",
  41080=>"000000000",
  41081=>"000000000",
  41082=>"001100000",
  41083=>"000000000",
  41084=>"111111110",
  41085=>"011011000",
  41086=>"000000101",
  41087=>"011111111",
  41088=>"000000000",
  41089=>"100110110",
  41090=>"111111111",
  41091=>"000001111",
  41092=>"000000000",
  41093=>"001101001",
  41094=>"111111111",
  41095=>"000000000",
  41096=>"111111000",
  41097=>"111111111",
  41098=>"111001111",
  41099=>"111111011",
  41100=>"110000000",
  41101=>"000000110",
  41102=>"111000000",
  41103=>"100110110",
  41104=>"000000010",
  41105=>"001111111",
  41106=>"000000000",
  41107=>"110111111",
  41108=>"111111111",
  41109=>"000000011",
  41110=>"111110110",
  41111=>"000111111",
  41112=>"000111111",
  41113=>"111001111",
  41114=>"111111111",
  41115=>"110000000",
  41116=>"000000000",
  41117=>"111000000",
  41118=>"111111111",
  41119=>"111111111",
  41120=>"000000000",
  41121=>"000000000",
  41122=>"111110100",
  41123=>"010000000",
  41124=>"001001001",
  41125=>"000100111",
  41126=>"000111111",
  41127=>"110000011",
  41128=>"111111111",
  41129=>"000000000",
  41130=>"010000000",
  41131=>"111100110",
  41132=>"010000100",
  41133=>"111011010",
  41134=>"001001111",
  41135=>"000000100",
  41136=>"000010111",
  41137=>"000000110",
  41138=>"111110110",
  41139=>"011000000",
  41140=>"011011111",
  41141=>"000000100",
  41142=>"100100110",
  41143=>"111110000",
  41144=>"000000000",
  41145=>"000001101",
  41146=>"001000000",
  41147=>"000000111",
  41148=>"000000111",
  41149=>"000000111",
  41150=>"111000000",
  41151=>"000000000",
  41152=>"001001111",
  41153=>"100000111",
  41154=>"011000000",
  41155=>"011111111",
  41156=>"000010110",
  41157=>"110111111",
  41158=>"011011000",
  41159=>"011001111",
  41160=>"110000000",
  41161=>"111100100",
  41162=>"111100110",
  41163=>"000001101",
  41164=>"001111111",
  41165=>"000000100",
  41166=>"000000100",
  41167=>"000000000",
  41168=>"000100000",
  41169=>"111000000",
  41170=>"000110000",
  41171=>"000000000",
  41172=>"110000111",
  41173=>"000000000",
  41174=>"110010110",
  41175=>"000000001",
  41176=>"101000000",
  41177=>"001001100",
  41178=>"000000000",
  41179=>"000000111",
  41180=>"000000000",
  41181=>"000000000",
  41182=>"011111111",
  41183=>"110110111",
  41184=>"110111000",
  41185=>"100000100",
  41186=>"101111011",
  41187=>"111111111",
  41188=>"111111000",
  41189=>"100000011",
  41190=>"101000001",
  41191=>"111111111",
  41192=>"000000000",
  41193=>"111111111",
  41194=>"111111111",
  41195=>"101001000",
  41196=>"111000000",
  41197=>"110111111",
  41198=>"011000000",
  41199=>"100000000",
  41200=>"000011000",
  41201=>"111000000",
  41202=>"111111110",
  41203=>"000000000",
  41204=>"000000000",
  41205=>"000000110",
  41206=>"101111111",
  41207=>"111000000",
  41208=>"111110000",
  41209=>"000000000",
  41210=>"000000110",
  41211=>"001101000",
  41212=>"000000111",
  41213=>"100100000",
  41214=>"110011111",
  41215=>"000000000",
  41216=>"000000000",
  41217=>"111111111",
  41218=>"000000000",
  41219=>"110000000",
  41220=>"101000000",
  41221=>"111000000",
  41222=>"001000110",
  41223=>"000110111",
  41224=>"111001111",
  41225=>"111000000",
  41226=>"111111111",
  41227=>"110111100",
  41228=>"111110110",
  41229=>"000000000",
  41230=>"000000110",
  41231=>"000000001",
  41232=>"000000001",
  41233=>"111111110",
  41234=>"111000000",
  41235=>"000000000",
  41236=>"000000000",
  41237=>"111111111",
  41238=>"111111101",
  41239=>"000100000",
  41240=>"111111111",
  41241=>"111111000",
  41242=>"000111110",
  41243=>"111111111",
  41244=>"000000000",
  41245=>"101000000",
  41246=>"111101101",
  41247=>"000000000",
  41248=>"000000000",
  41249=>"000000111",
  41250=>"111111011",
  41251=>"111001000",
  41252=>"111110100",
  41253=>"000001000",
  41254=>"111111000",
  41255=>"111111111",
  41256=>"111111110",
  41257=>"000111111",
  41258=>"100110110",
  41259=>"010111111",
  41260=>"000000000",
  41261=>"111111110",
  41262=>"101010111",
  41263=>"000000000",
  41264=>"100100000",
  41265=>"111000001",
  41266=>"000010011",
  41267=>"000000000",
  41268=>"111111000",
  41269=>"000111110",
  41270=>"000000000",
  41271=>"111111111",
  41272=>"000000000",
  41273=>"111000000",
  41274=>"000000000",
  41275=>"111000000",
  41276=>"111111111",
  41277=>"100110110",
  41278=>"001000000",
  41279=>"000000001",
  41280=>"111100000",
  41281=>"111111111",
  41282=>"111111110",
  41283=>"000111111",
  41284=>"110110000",
  41285=>"110000000",
  41286=>"110000000",
  41287=>"000111111",
  41288=>"000000000",
  41289=>"110000000",
  41290=>"111101000",
  41291=>"111110000",
  41292=>"111101111",
  41293=>"001110110",
  41294=>"100000110",
  41295=>"111011001",
  41296=>"000000000",
  41297=>"111111000",
  41298=>"110100000",
  41299=>"000000000",
  41300=>"111000001",
  41301=>"000000000",
  41302=>"111100111",
  41303=>"111110000",
  41304=>"111101001",
  41305=>"000100000",
  41306=>"100000000",
  41307=>"000000000",
  41308=>"010110000",
  41309=>"010010000",
  41310=>"000000000",
  41311=>"100011000",
  41312=>"000000000",
  41313=>"011111000",
  41314=>"100001011",
  41315=>"111101000",
  41316=>"111111111",
  41317=>"000111111",
  41318=>"000100110",
  41319=>"000000000",
  41320=>"111000000",
  41321=>"111111111",
  41322=>"001010111",
  41323=>"000000110",
  41324=>"000000000",
  41325=>"001001010",
  41326=>"000000000",
  41327=>"110110110",
  41328=>"110000100",
  41329=>"011111111",
  41330=>"000111110",
  41331=>"100100111",
  41332=>"111110111",
  41333=>"000001111",
  41334=>"000000000",
  41335=>"111111110",
  41336=>"111000000",
  41337=>"011010010",
  41338=>"111011000",
  41339=>"111111111",
  41340=>"100110110",
  41341=>"110011011",
  41342=>"110011111",
  41343=>"111000000",
  41344=>"001111111",
  41345=>"010110111",
  41346=>"110110011",
  41347=>"000000111",
  41348=>"111111111",
  41349=>"101001111",
  41350=>"000000000",
  41351=>"111111111",
  41352=>"000000000",
  41353=>"100100111",
  41354=>"111110000",
  41355=>"111111011",
  41356=>"111110100",
  41357=>"111111111",
  41358=>"110010111",
  41359=>"000111111",
  41360=>"000011111",
  41361=>"111111000",
  41362=>"111101010",
  41363=>"111001000",
  41364=>"001000001",
  41365=>"000001001",
  41366=>"111111101",
  41367=>"000000010",
  41368=>"111111111",
  41369=>"000000000",
  41370=>"100000000",
  41371=>"111111110",
  41372=>"000000000",
  41373=>"111111110",
  41374=>"000000100",
  41375=>"000111111",
  41376=>"111001000",
  41377=>"110111101",
  41378=>"110000110",
  41379=>"100110100",
  41380=>"000100100",
  41381=>"101001000",
  41382=>"111101111",
  41383=>"000111111",
  41384=>"000000000",
  41385=>"000111000",
  41386=>"111110000",
  41387=>"100110110",
  41388=>"010111110",
  41389=>"111000000",
  41390=>"111001101",
  41391=>"111000000",
  41392=>"011000000",
  41393=>"000000010",
  41394=>"111111111",
  41395=>"111000000",
  41396=>"000000011",
  41397=>"000000000",
  41398=>"010111101",
  41399=>"011000110",
  41400=>"100000110",
  41401=>"100111111",
  41402=>"000000000",
  41403=>"000001000",
  41404=>"100000001",
  41405=>"111101000",
  41406=>"001000000",
  41407=>"111111111",
  41408=>"000000111",
  41409=>"000011111",
  41410=>"000111111",
  41411=>"000001111",
  41412=>"011110111",
  41413=>"111000111",
  41414=>"011000111",
  41415=>"001100100",
  41416=>"000001111",
  41417=>"001101111",
  41418=>"000010110",
  41419=>"000000000",
  41420=>"111111000",
  41421=>"110110000",
  41422=>"101000000",
  41423=>"000000000",
  41424=>"111111001",
  41425=>"111111111",
  41426=>"111011111",
  41427=>"111111111",
  41428=>"100110000",
  41429=>"111110111",
  41430=>"000000000",
  41431=>"000000001",
  41432=>"111000000",
  41433=>"011000000",
  41434=>"110100111",
  41435=>"111111111",
  41436=>"100100110",
  41437=>"000010111",
  41438=>"000000000",
  41439=>"100000000",
  41440=>"110111111",
  41441=>"111111111",
  41442=>"111111111",
  41443=>"000000000",
  41444=>"110000000",
  41445=>"000000000",
  41446=>"001000000",
  41447=>"110110110",
  41448=>"000001111",
  41449=>"111000000",
  41450=>"111111000",
  41451=>"011101111",
  41452=>"000111111",
  41453=>"011110111",
  41454=>"000011111",
  41455=>"111111000",
  41456=>"100100111",
  41457=>"000011111",
  41458=>"111111111",
  41459=>"000000000",
  41460=>"101111111",
  41461=>"111011000",
  41462=>"111111111",
  41463=>"010011111",
  41464=>"000000000",
  41465=>"111101001",
  41466=>"000000111",
  41467=>"000000000",
  41468=>"000000000",
  41469=>"111011000",
  41470=>"001011000",
  41471=>"101001000",
  41472=>"101111001",
  41473=>"101100000",
  41474=>"111000000",
  41475=>"111111111",
  41476=>"000000111",
  41477=>"000000100",
  41478=>"111101000",
  41479=>"111111111",
  41480=>"111111001",
  41481=>"111111010",
  41482=>"111111001",
  41483=>"110111111",
  41484=>"101101100",
  41485=>"001000001",
  41486=>"111111011",
  41487=>"000000000",
  41488=>"110110110",
  41489=>"111111111",
  41490=>"000000011",
  41491=>"000001001",
  41492=>"010000000",
  41493=>"111001001",
  41494=>"000010011",
  41495=>"111111011",
  41496=>"110110100",
  41497=>"000001000",
  41498=>"000000000",
  41499=>"110000000",
  41500=>"101111111",
  41501=>"000001111",
  41502=>"110100000",
  41503=>"110110110",
  41504=>"100111001",
  41505=>"110000000",
  41506=>"110110110",
  41507=>"001000001",
  41508=>"000000001",
  41509=>"011011111",
  41510=>"100000100",
  41511=>"010000111",
  41512=>"111000001",
  41513=>"111111111",
  41514=>"000000000",
  41515=>"111111110",
  41516=>"110110110",
  41517=>"000000001",
  41518=>"000000001",
  41519=>"101111011",
  41520=>"001000110",
  41521=>"110111110",
  41522=>"000010010",
  41523=>"010010000",
  41524=>"001101001",
  41525=>"000000110",
  41526=>"110110000",
  41527=>"011111000",
  41528=>"111111111",
  41529=>"001001111",
  41530=>"101101000",
  41531=>"001101111",
  41532=>"000000001",
  41533=>"111111000",
  41534=>"000000000",
  41535=>"000000110",
  41536=>"111111001",
  41537=>"111000000",
  41538=>"101111111",
  41539=>"111111111",
  41540=>"110110100",
  41541=>"000000111",
  41542=>"001001001",
  41543=>"000000101",
  41544=>"000000000",
  41545=>"111001011",
  41546=>"000000000",
  41547=>"001001000",
  41548=>"001001000",
  41549=>"110110000",
  41550=>"000000000",
  41551=>"000000000",
  41552=>"000000000",
  41553=>"011001111",
  41554=>"000000000",
  41555=>"110110000",
  41556=>"000000000",
  41557=>"011111110",
  41558=>"111111101",
  41559=>"000101111",
  41560=>"000000000",
  41561=>"110110110",
  41562=>"001001011",
  41563=>"010010011",
  41564=>"111111111",
  41565=>"100100000",
  41566=>"000000110",
  41567=>"010000000",
  41568=>"000011110",
  41569=>"110110110",
  41570=>"111111110",
  41571=>"000100111",
  41572=>"111111011",
  41573=>"110110011",
  41574=>"000110111",
  41575=>"111111111",
  41576=>"010111010",
  41577=>"111100000",
  41578=>"001000110",
  41579=>"001001111",
  41580=>"100000100",
  41581=>"101101000",
  41582=>"001000000",
  41583=>"111111111",
  41584=>"110110010",
  41585=>"000001111",
  41586=>"100000000",
  41587=>"110110000",
  41588=>"000101111",
  41589=>"100000100",
  41590=>"001101111",
  41591=>"110110011",
  41592=>"101111111",
  41593=>"000010000",
  41594=>"001000000",
  41595=>"111000000",
  41596=>"100100100",
  41597=>"111111011",
  41598=>"010000000",
  41599=>"110111010",
  41600=>"001001001",
  41601=>"101000111",
  41602=>"010000000",
  41603=>"111111111",
  41604=>"001001001",
  41605=>"111111011",
  41606=>"011111111",
  41607=>"001001001",
  41608=>"000111111",
  41609=>"110000110",
  41610=>"011111000",
  41611=>"111111111",
  41612=>"110110110",
  41613=>"000000000",
  41614=>"111111101",
  41615=>"111101000",
  41616=>"100001111",
  41617=>"110111000",
  41618=>"000110111",
  41619=>"110110110",
  41620=>"000000000",
  41621=>"110010000",
  41622=>"001001101",
  41623=>"111100000",
  41624=>"000000000",
  41625=>"000000000",
  41626=>"110110000",
  41627=>"011111111",
  41628=>"111111101",
  41629=>"111111011",
  41630=>"100100110",
  41631=>"000001111",
  41632=>"100100000",
  41633=>"000000001",
  41634=>"000000111",
  41635=>"000110110",
  41636=>"101000000",
  41637=>"000000100",
  41638=>"111111001",
  41639=>"000000000",
  41640=>"111111011",
  41641=>"000000000",
  41642=>"100101000",
  41643=>"000110000",
  41644=>"111011110",
  41645=>"000100100",
  41646=>"100111111",
  41647=>"000101011",
  41648=>"111110111",
  41649=>"011010010",
  41650=>"111111111",
  41651=>"111001000",
  41652=>"100110110",
  41653=>"101101111",
  41654=>"100000000",
  41655=>"000000000",
  41656=>"001001001",
  41657=>"000111111",
  41658=>"111001000",
  41659=>"010010001",
  41660=>"000001111",
  41661=>"001001000",
  41662=>"010000000",
  41663=>"001001001",
  41664=>"100000000",
  41665=>"100000101",
  41666=>"111111111",
  41667=>"111111111",
  41668=>"000000001",
  41669=>"111101000",
  41670=>"010111110",
  41671=>"000000111",
  41672=>"111101101",
  41673=>"010000000",
  41674=>"111000000",
  41675=>"001000100",
  41676=>"111111111",
  41677=>"010000000",
  41678=>"001000000",
  41679=>"000000111",
  41680=>"000000000",
  41681=>"000000000",
  41682=>"111111111",
  41683=>"111110110",
  41684=>"000000111",
  41685=>"100000000",
  41686=>"000000000",
  41687=>"111111011",
  41688=>"000110111",
  41689=>"100001101",
  41690=>"000000100",
  41691=>"001001111",
  41692=>"110110110",
  41693=>"000000000",
  41694=>"000001001",
  41695=>"100001001",
  41696=>"011101111",
  41697=>"011000111",
  41698=>"010110000",
  41699=>"111011010",
  41700=>"000101101",
  41701=>"010000100",
  41702=>"000000000",
  41703=>"100000000",
  41704=>"111000000",
  41705=>"100100010",
  41706=>"000010010",
  41707=>"111111100",
  41708=>"000000011",
  41709=>"111111001",
  41710=>"000000001",
  41711=>"000111111",
  41712=>"101000000",
  41713=>"000001011",
  41714=>"100011011",
  41715=>"101001111",
  41716=>"011111111",
  41717=>"000000000",
  41718=>"100110100",
  41719=>"000000000",
  41720=>"000001101",
  41721=>"101111110",
  41722=>"000000001",
  41723=>"000001101",
  41724=>"111011011",
  41725=>"011011011",
  41726=>"111111001",
  41727=>"101100101",
  41728=>"110000000",
  41729=>"100101101",
  41730=>"001001111",
  41731=>"010000000",
  41732=>"000111111",
  41733=>"011010000",
  41734=>"000000100",
  41735=>"100110111",
  41736=>"110000000",
  41737=>"000000111",
  41738=>"110111111",
  41739=>"100000001",
  41740=>"001001000",
  41741=>"000000000",
  41742=>"110110010",
  41743=>"000001111",
  41744=>"010000000",
  41745=>"101000001",
  41746=>"001001101",
  41747=>"110110110",
  41748=>"111111111",
  41749=>"110010010",
  41750=>"100100111",
  41751=>"000111101",
  41752=>"011110000",
  41753=>"101000001",
  41754=>"000000000",
  41755=>"011001000",
  41756=>"101101101",
  41757=>"000011111",
  41758=>"100000000",
  41759=>"110111001",
  41760=>"011111111",
  41761=>"001011011",
  41762=>"111011001",
  41763=>"000000101",
  41764=>"011010110",
  41765=>"101001101",
  41766=>"011101111",
  41767=>"100111011",
  41768=>"110110010",
  41769=>"000000000",
  41770=>"110011001",
  41771=>"101101111",
  41772=>"000000010",
  41773=>"100110111",
  41774=>"111111000",
  41775=>"000110110",
  41776=>"000001000",
  41777=>"001000000",
  41778=>"111110111",
  41779=>"011011000",
  41780=>"000000001",
  41781=>"100100000",
  41782=>"011001000",
  41783=>"111000000",
  41784=>"001001011",
  41785=>"001000111",
  41786=>"111111111",
  41787=>"111111111",
  41788=>"000000000",
  41789=>"010110110",
  41790=>"000001000",
  41791=>"011111111",
  41792=>"111111001",
  41793=>"110000000",
  41794=>"001001001",
  41795=>"001000001",
  41796=>"000000000",
  41797=>"001000000",
  41798=>"000000000",
  41799=>"001001000",
  41800=>"111100111",
  41801=>"111010000",
  41802=>"000000000",
  41803=>"001001011",
  41804=>"110010110",
  41805=>"000000000",
  41806=>"110110110",
  41807=>"010010110",
  41808=>"111111010",
  41809=>"000000011",
  41810=>"111100110",
  41811=>"000000101",
  41812=>"100101100",
  41813=>"011011011",
  41814=>"001001001",
  41815=>"001011011",
  41816=>"101111101",
  41817=>"111010000",
  41818=>"000000000",
  41819=>"000000000",
  41820=>"101101101",
  41821=>"100000001",
  41822=>"111111111",
  41823=>"110110011",
  41824=>"111111111",
  41825=>"001001001",
  41826=>"100011011",
  41827=>"000000111",
  41828=>"111111111",
  41829=>"100000111",
  41830=>"001101101",
  41831=>"000000111",
  41832=>"111100100",
  41833=>"000000000",
  41834=>"100111111",
  41835=>"000011011",
  41836=>"001100110",
  41837=>"111000000",
  41838=>"001001000",
  41839=>"000000000",
  41840=>"110110110",
  41841=>"110110110",
  41842=>"000011110",
  41843=>"011111111",
  41844=>"000000001",
  41845=>"000000000",
  41846=>"000000001",
  41847=>"011101000",
  41848=>"010111110",
  41849=>"001000111",
  41850=>"000011110",
  41851=>"100000000",
  41852=>"010010110",
  41853=>"110110110",
  41854=>"111100111",
  41855=>"111000011",
  41856=>"001001000",
  41857=>"000000110",
  41858=>"000000000",
  41859=>"111001000",
  41860=>"111111111",
  41861=>"010001000",
  41862=>"111100100",
  41863=>"000001001",
  41864=>"100000001",
  41865=>"000000001",
  41866=>"100100110",
  41867=>"000010010",
  41868=>"000000001",
  41869=>"000000101",
  41870=>"000110111",
  41871=>"000111111",
  41872=>"000010010",
  41873=>"010110110",
  41874=>"000000000",
  41875=>"101100000",
  41876=>"000010010",
  41877=>"000000000",
  41878=>"000000000",
  41879=>"000000110",
  41880=>"000100001",
  41881=>"010110110",
  41882=>"001000000",
  41883=>"111111111",
  41884=>"110111110",
  41885=>"111111000",
  41886=>"001001101",
  41887=>"110010000",
  41888=>"000000000",
  41889=>"001101000",
  41890=>"100000001",
  41891=>"000001001",
  41892=>"111110000",
  41893=>"111111101",
  41894=>"010010000",
  41895=>"111110100",
  41896=>"100100000",
  41897=>"000110110",
  41898=>"110110111",
  41899=>"000000000",
  41900=>"101001111",
  41901=>"101001101",
  41902=>"000111111",
  41903=>"100000001",
  41904=>"111100000",
  41905=>"000000110",
  41906=>"111111111",
  41907=>"000000100",
  41908=>"001001110",
  41909=>"111111111",
  41910=>"111111111",
  41911=>"100111111",
  41912=>"011111011",
  41913=>"000111111",
  41914=>"000000000",
  41915=>"111100111",
  41916=>"111111000",
  41917=>"001001111",
  41918=>"100001001",
  41919=>"000000000",
  41920=>"000000000",
  41921=>"111111111",
  41922=>"000000010",
  41923=>"111111110",
  41924=>"001001001",
  41925=>"001011111",
  41926=>"001111111",
  41927=>"101100100",
  41928=>"111001001",
  41929=>"100100100",
  41930=>"101001001",
  41931=>"111111111",
  41932=>"110110111",
  41933=>"000000000",
  41934=>"001110111",
  41935=>"000000000",
  41936=>"000000001",
  41937=>"010000000",
  41938=>"111111010",
  41939=>"111100100",
  41940=>"000000000",
  41941=>"111000100",
  41942=>"000000000",
  41943=>"111111111",
  41944=>"001000111",
  41945=>"100101101",
  41946=>"111111000",
  41947=>"000001101",
  41948=>"000000000",
  41949=>"000000000",
  41950=>"101100000",
  41951=>"100000001",
  41952=>"001101100",
  41953=>"101000000",
  41954=>"111111000",
  41955=>"001000001",
  41956=>"000000001",
  41957=>"001111111",
  41958=>"111001000",
  41959=>"000000011",
  41960=>"101111111",
  41961=>"001001011",
  41962=>"111101001",
  41963=>"111111111",
  41964=>"000001101",
  41965=>"000001011",
  41966=>"001001101",
  41967=>"110110110",
  41968=>"000000110",
  41969=>"000000000",
  41970=>"010000011",
  41971=>"111111000",
  41972=>"000000010",
  41973=>"000001101",
  41974=>"100000000",
  41975=>"000111111",
  41976=>"111011000",
  41977=>"001011011",
  41978=>"000001101",
  41979=>"111111011",
  41980=>"011000000",
  41981=>"100000000",
  41982=>"001111111",
  41983=>"000000000",
  41984=>"110110011",
  41985=>"111011001",
  41986=>"101000000",
  41987=>"111000000",
  41988=>"000000000",
  41989=>"101001011",
  41990=>"100111000",
  41991=>"101101101",
  41992=>"000000110",
  41993=>"000000100",
  41994=>"011010000",
  41995=>"111111111",
  41996=>"011111111",
  41997=>"000000000",
  41998=>"000000000",
  41999=>"010000000",
  42000=>"110111111",
  42001=>"010111111",
  42002=>"000000000",
  42003=>"111111111",
  42004=>"001000000",
  42005=>"001101111",
  42006=>"000000001",
  42007=>"110110111",
  42008=>"000000000",
  42009=>"000000000",
  42010=>"000000000",
  42011=>"111111111",
  42012=>"001000000",
  42013=>"001001111",
  42014=>"000000000",
  42015=>"000101111",
  42016=>"110101111",
  42017=>"111111111",
  42018=>"000110111",
  42019=>"000000001",
  42020=>"100100000",
  42021=>"111111101",
  42022=>"101000000",
  42023=>"000111110",
  42024=>"000111111",
  42025=>"011011111",
  42026=>"000000000",
  42027=>"011111111",
  42028=>"111111111",
  42029=>"100110110",
  42030=>"111111111",
  42031=>"111111111",
  42032=>"101101111",
  42033=>"010000000",
  42034=>"010010000",
  42035=>"111111111",
  42036=>"000100000",
  42037=>"111111010",
  42038=>"100100000",
  42039=>"000100110",
  42040=>"000000000",
  42041=>"011100110",
  42042=>"111110111",
  42043=>"111111100",
  42044=>"000000000",
  42045=>"011111011",
  42046=>"111111111",
  42047=>"000000000",
  42048=>"000001111",
  42049=>"000000000",
  42050=>"000000000",
  42051=>"001100111",
  42052=>"011111011",
  42053=>"001001001",
  42054=>"000000000",
  42055=>"111111111",
  42056=>"011011111",
  42057=>"101111111",
  42058=>"111111111",
  42059=>"000000000",
  42060=>"111111111",
  42061=>"111111111",
  42062=>"111111011",
  42063=>"000001111",
  42064=>"000001111",
  42065=>"000100000",
  42066=>"000000000",
  42067=>"000000000",
  42068=>"111111111",
  42069=>"111101000",
  42070=>"001001100",
  42071=>"000000110",
  42072=>"101111110",
  42073=>"111101001",
  42074=>"111111000",
  42075=>"000000000",
  42076=>"111111111",
  42077=>"000011111",
  42078=>"001011110",
  42079=>"001000000",
  42080=>"111111010",
  42081=>"011111010",
  42082=>"111111111",
  42083=>"111001000",
  42084=>"000111000",
  42085=>"000000000",
  42086=>"000111111",
  42087=>"000010111",
  42088=>"111111001",
  42089=>"100100000",
  42090=>"111000000",
  42091=>"111111111",
  42092=>"111111111",
  42093=>"111111111",
  42094=>"001001111",
  42095=>"111111001",
  42096=>"111111111",
  42097=>"111111111",
  42098=>"100100110",
  42099=>"000000000",
  42100=>"011011001",
  42101=>"111111010",
  42102=>"111111111",
  42103=>"000000000",
  42104=>"000000100",
  42105=>"111101111",
  42106=>"000000000",
  42107=>"000000000",
  42108=>"010010000",
  42109=>"011011000",
  42110=>"111111111",
  42111=>"001100111",
  42112=>"000011000",
  42113=>"111111111",
  42114=>"100100100",
  42115=>"000000100",
  42116=>"000000000",
  42117=>"111000000",
  42118=>"111111111",
  42119=>"110111111",
  42120=>"000010011",
  42121=>"110111111",
  42122=>"011011001",
  42123=>"111111111",
  42124=>"101111111",
  42125=>"111111111",
  42126=>"111111111",
  42127=>"111111111",
  42128=>"000001001",
  42129=>"000000100",
  42130=>"000001000",
  42131=>"001001011",
  42132=>"011000000",
  42133=>"000011011",
  42134=>"000000000",
  42135=>"000000000",
  42136=>"000000000",
  42137=>"111111111",
  42138=>"111100100",
  42139=>"000000000",
  42140=>"000000000",
  42141=>"100111001",
  42142=>"111111111",
  42143=>"011111011",
  42144=>"111111111",
  42145=>"001101001",
  42146=>"000000000",
  42147=>"000000010",
  42148=>"000000100",
  42149=>"000000000",
  42150=>"001000000",
  42151=>"000010000",
  42152=>"000101001",
  42153=>"111111111",
  42154=>"100000100",
  42155=>"000000000",
  42156=>"000000000",
  42157=>"110111111",
  42158=>"111111111",
  42159=>"000000000",
  42160=>"111011000",
  42161=>"000110010",
  42162=>"110111010",
  42163=>"111000000",
  42164=>"110010000",
  42165=>"000000000",
  42166=>"000000000",
  42167=>"100111111",
  42168=>"000000000",
  42169=>"111111111",
  42170=>"001000000",
  42171=>"111111100",
  42172=>"000011111",
  42173=>"100101101",
  42174=>"100111111",
  42175=>"111111111",
  42176=>"110110010",
  42177=>"111111100",
  42178=>"000000000",
  42179=>"000110110",
  42180=>"111000000",
  42181=>"000100111",
  42182=>"111111111",
  42183=>"111111111",
  42184=>"000001000",
  42185=>"000000010",
  42186=>"111000000",
  42187=>"111111111",
  42188=>"001000111",
  42189=>"000001001",
  42190=>"000000000",
  42191=>"000001001",
  42192=>"011001000",
  42193=>"111111111",
  42194=>"011111111",
  42195=>"100100001",
  42196=>"000000000",
  42197=>"111111111",
  42198=>"010111000",
  42199=>"000000110",
  42200=>"000000000",
  42201=>"110111111",
  42202=>"111000000",
  42203=>"000000000",
  42204=>"000000001",
  42205=>"000000011",
  42206=>"000000000",
  42207=>"000000000",
  42208=>"000000000",
  42209=>"010000110",
  42210=>"000000000",
  42211=>"000000000",
  42212=>"111011000",
  42213=>"001001011",
  42214=>"111111110",
  42215=>"000100100",
  42216=>"111111111",
  42217=>"000111110",
  42218=>"111101000",
  42219=>"101100111",
  42220=>"111111111",
  42221=>"000111110",
  42222=>"111110110",
  42223=>"111111111",
  42224=>"101111111",
  42225=>"011000000",
  42226=>"111111111",
  42227=>"101100101",
  42228=>"111111111",
  42229=>"000000000",
  42230=>"100100110",
  42231=>"000000111",
  42232=>"111111001",
  42233=>"011001111",
  42234=>"011111010",
  42235=>"110110000",
  42236=>"001001001",
  42237=>"111111110",
  42238=>"000100111",
  42239=>"110010000",
  42240=>"111011001",
  42241=>"011001001",
  42242=>"000000000",
  42243=>"010010110",
  42244=>"000000111",
  42245=>"100000000",
  42246=>"100101111",
  42247=>"111111000",
  42248=>"000000000",
  42249=>"000000000",
  42250=>"111000000",
  42251=>"111111111",
  42252=>"000000000",
  42253=>"011111111",
  42254=>"001001000",
  42255=>"000011111",
  42256=>"000111111",
  42257=>"000000000",
  42258=>"000000000",
  42259=>"010000000",
  42260=>"111100111",
  42261=>"011011011",
  42262=>"100100100",
  42263=>"000000000",
  42264=>"111111111",
  42265=>"111111111",
  42266=>"111111010",
  42267=>"000111001",
  42268=>"000000100",
  42269=>"000111111",
  42270=>"000000000",
  42271=>"000001011",
  42272=>"000000000",
  42273=>"000000011",
  42274=>"111111111",
  42275=>"001001111",
  42276=>"000000000",
  42277=>"111000000",
  42278=>"000000000",
  42279=>"000101111",
  42280=>"111111000",
  42281=>"001000101",
  42282=>"000000000",
  42283=>"000000000",
  42284=>"000001010",
  42285=>"111111111",
  42286=>"011011000",
  42287=>"000000000",
  42288=>"111111111",
  42289=>"000000000",
  42290=>"001011011",
  42291=>"110111111",
  42292=>"001000000",
  42293=>"100111011",
  42294=>"100100101",
  42295=>"100000000",
  42296=>"011010000",
  42297=>"001000000",
  42298=>"000110010",
  42299=>"000000000",
  42300=>"000000100",
  42301=>"000000010",
  42302=>"110000000",
  42303=>"000000000",
  42304=>"111111111",
  42305=>"000000100",
  42306=>"000000000",
  42307=>"111111111",
  42308=>"100100101",
  42309=>"001000111",
  42310=>"000011000",
  42311=>"000000000",
  42312=>"000000000",
  42313=>"111011000",
  42314=>"000000000",
  42315=>"100000000",
  42316=>"111110000",
  42317=>"111110000",
  42318=>"111101111",
  42319=>"000000000",
  42320=>"000111100",
  42321=>"101111100",
  42322=>"000000000",
  42323=>"000000000",
  42324=>"000000000",
  42325=>"011011011",
  42326=>"100111111",
  42327=>"000000000",
  42328=>"111111111",
  42329=>"000001111",
  42330=>"011111111",
  42331=>"111111111",
  42332=>"111111111",
  42333=>"000000001",
  42334=>"001111111",
  42335=>"101000000",
  42336=>"110111111",
  42337=>"001011111",
  42338=>"000000001",
  42339=>"111001111",
  42340=>"011010000",
  42341=>"001001001",
  42342=>"011011011",
  42343=>"000000000",
  42344=>"001000000",
  42345=>"111011000",
  42346=>"001111111",
  42347=>"000000000",
  42348=>"111111000",
  42349=>"001100110",
  42350=>"000000000",
  42351=>"000000000",
  42352=>"110100100",
  42353=>"110010000",
  42354=>"111111111",
  42355=>"111111111",
  42356=>"000000001",
  42357=>"000000000",
  42358=>"000000110",
  42359=>"000000101",
  42360=>"111111000",
  42361=>"000110111",
  42362=>"000000000",
  42363=>"111111111",
  42364=>"111111111",
  42365=>"111111111",
  42366=>"000000000",
  42367=>"111111010",
  42368=>"111111011",
  42369=>"111111111",
  42370=>"000000000",
  42371=>"111100000",
  42372=>"000000000",
  42373=>"111111111",
  42374=>"000000000",
  42375=>"000110111",
  42376=>"111111000",
  42377=>"011001000",
  42378=>"111000000",
  42379=>"100000000",
  42380=>"111111111",
  42381=>"001101111",
  42382=>"111111110",
  42383=>"000000000",
  42384=>"000000000",
  42385=>"000110111",
  42386=>"000000001",
  42387=>"000000000",
  42388=>"000000010",
  42389=>"000010000",
  42390=>"111111110",
  42391=>"110011010",
  42392=>"100111111",
  42393=>"111001001",
  42394=>"000000000",
  42395=>"001111110",
  42396=>"000000000",
  42397=>"111111000",
  42398=>"000000000",
  42399=>"011000000",
  42400=>"111111111",
  42401=>"101001000",
  42402=>"001000001",
  42403=>"111111111",
  42404=>"111111111",
  42405=>"111111111",
  42406=>"111111001",
  42407=>"000000001",
  42408=>"111011111",
  42409=>"001000001",
  42410=>"000000101",
  42411=>"011111001",
  42412=>"101000100",
  42413=>"111111111",
  42414=>"100101111",
  42415=>"000000000",
  42416=>"111111111",
  42417=>"000000000",
  42418=>"000000000",
  42419=>"111111111",
  42420=>"000000000",
  42421=>"000000011",
  42422=>"111111111",
  42423=>"100101100",
  42424=>"111111000",
  42425=>"111000000",
  42426=>"000011000",
  42427=>"111111000",
  42428=>"111111000",
  42429=>"000000000",
  42430=>"000000000",
  42431=>"001000110",
  42432=>"000000000",
  42433=>"110110111",
  42434=>"111011111",
  42435=>"000000000",
  42436=>"000100111",
  42437=>"000000010",
  42438=>"100111111",
  42439=>"101111111",
  42440=>"000000100",
  42441=>"000000000",
  42442=>"001001001",
  42443=>"001000000",
  42444=>"000000000",
  42445=>"111111111",
  42446=>"111111111",
  42447=>"111111111",
  42448=>"110110000",
  42449=>"001101000",
  42450=>"111011011",
  42451=>"001000111",
  42452=>"100100111",
  42453=>"111000000",
  42454=>"101111111",
  42455=>"110110110",
  42456=>"100000000",
  42457=>"000111111",
  42458=>"000000000",
  42459=>"000000001",
  42460=>"100000000",
  42461=>"101101001",
  42462=>"100110000",
  42463=>"100100110",
  42464=>"000000000",
  42465=>"000000000",
  42466=>"111111111",
  42467=>"111111111",
  42468=>"010100111",
  42469=>"000010111",
  42470=>"000000100",
  42471=>"000000000",
  42472=>"011001011",
  42473=>"100000111",
  42474=>"100111110",
  42475=>"000011011",
  42476=>"111011000",
  42477=>"011111111",
  42478=>"111111111",
  42479=>"111111110",
  42480=>"000000000",
  42481=>"000110000",
  42482=>"000011011",
  42483=>"000000000",
  42484=>"101111111",
  42485=>"000000000",
  42486=>"111111111",
  42487=>"001011000",
  42488=>"000111111",
  42489=>"110011011",
  42490=>"000100110",
  42491=>"101000000",
  42492=>"000100000",
  42493=>"001001001",
  42494=>"011001111",
  42495=>"000110011",
  42496=>"011011111",
  42497=>"000000000",
  42498=>"001000000",
  42499=>"110111111",
  42500=>"111111000",
  42501=>"000000000",
  42502=>"110000001",
  42503=>"001001111",
  42504=>"000001111",
  42505=>"111010000",
  42506=>"110100000",
  42507=>"001000000",
  42508=>"100000111",
  42509=>"000001111",
  42510=>"100101111",
  42511=>"111111111",
  42512=>"111111111",
  42513=>"010111110",
  42514=>"110111110",
  42515=>"110100111",
  42516=>"000000000",
  42517=>"001101111",
  42518=>"111111111",
  42519=>"110000001",
  42520=>"100000111",
  42521=>"000011100",
  42522=>"011001001",
  42523=>"001000001",
  42524=>"111111111",
  42525=>"111111111",
  42526=>"111000000",
  42527=>"101011000",
  42528=>"000011011",
  42529=>"110111111",
  42530=>"111111000",
  42531=>"000000000",
  42532=>"000000000",
  42533=>"000110111",
  42534=>"111011000",
  42535=>"101000101",
  42536=>"111001101",
  42537=>"010111111",
  42538=>"101101000",
  42539=>"000000011",
  42540=>"000000001",
  42541=>"111111110",
  42542=>"111111100",
  42543=>"110100100",
  42544=>"011011000",
  42545=>"001111111",
  42546=>"111111011",
  42547=>"111111111",
  42548=>"011011011",
  42549=>"101111111",
  42550=>"110111010",
  42551=>"000000111",
  42552=>"000110000",
  42553=>"001001000",
  42554=>"111000001",
  42555=>"111100101",
  42556=>"000000000",
  42557=>"111100110",
  42558=>"111011000",
  42559=>"000100111",
  42560=>"000111100",
  42561=>"011010000",
  42562=>"111111111",
  42563=>"111111001",
  42564=>"110111100",
  42565=>"000110111",
  42566=>"000000000",
  42567=>"111110100",
  42568=>"011011111",
  42569=>"001000000",
  42570=>"011011110",
  42571=>"101101111",
  42572=>"001001001",
  42573=>"111111111",
  42574=>"000111000",
  42575=>"001001000",
  42576=>"111111100",
  42577=>"110111111",
  42578=>"110111110",
  42579=>"001001001",
  42580=>"000000000",
  42581=>"100101000",
  42582=>"101000000",
  42583=>"101111111",
  42584=>"001001111",
  42585=>"101001001",
  42586=>"000000000",
  42587=>"100000000",
  42588=>"010000000",
  42589=>"000000000",
  42590=>"000000000",
  42591=>"111111000",
  42592=>"011000000",
  42593=>"000100100",
  42594=>"110110000",
  42595=>"000010000",
  42596=>"000010001",
  42597=>"001000000",
  42598=>"111111000",
  42599=>"000000010",
  42600=>"111110000",
  42601=>"111111111",
  42602=>"100000010",
  42603=>"000000000",
  42604=>"001001000",
  42605=>"000111111",
  42606=>"000000000",
  42607=>"001111111",
  42608=>"110110000",
  42609=>"001001000",
  42610=>"011000000",
  42611=>"111110000",
  42612=>"000110111",
  42613=>"110110110",
  42614=>"011111111",
  42615=>"100000000",
  42616=>"100000011",
  42617=>"000000001",
  42618=>"111000000",
  42619=>"000000000",
  42620=>"100000000",
  42621=>"000110111",
  42622=>"111111000",
  42623=>"000000000",
  42624=>"000000000",
  42625=>"111101001",
  42626=>"111111111",
  42627=>"000000111",
  42628=>"001000000",
  42629=>"001001101",
  42630=>"101000100",
  42631=>"111001011",
  42632=>"101111111",
  42633=>"110111111",
  42634=>"110100000",
  42635=>"101111111",
  42636=>"000000000",
  42637=>"111000000",
  42638=>"111111001",
  42639=>"000000000",
  42640=>"000000000",
  42641=>"110010010",
  42642=>"111111110",
  42643=>"000010011",
  42644=>"000100111",
  42645=>"100100100",
  42646=>"000000000",
  42647=>"001001001",
  42648=>"011001111",
  42649=>"111111010",
  42650=>"111111111",
  42651=>"000000000",
  42652=>"001001101",
  42653=>"100000011",
  42654=>"100001111",
  42655=>"111111100",
  42656=>"111111111",
  42657=>"000000111",
  42658=>"111111000",
  42659=>"011111011",
  42660=>"110001111",
  42661=>"000100111",
  42662=>"011111000",
  42663=>"110111110",
  42664=>"101101011",
  42665=>"000000000",
  42666=>"000000101",
  42667=>"110111110",
  42668=>"111111111",
  42669=>"111111000",
  42670=>"000000001",
  42671=>"111111010",
  42672=>"111000110",
  42673=>"100110100",
  42674=>"111111110",
  42675=>"000101000",
  42676=>"001111111",
  42677=>"000000000",
  42678=>"000000001",
  42679=>"000000001",
  42680=>"111111110",
  42681=>"110000111",
  42682=>"001001000",
  42683=>"111001001",
  42684=>"000000000",
  42685=>"000000111",
  42686=>"111111111",
  42687=>"000000001",
  42688=>"000000100",
  42689=>"001000000",
  42690=>"111000001",
  42691=>"000000000",
  42692=>"000000000",
  42693=>"000000000",
  42694=>"000001111",
  42695=>"000000111",
  42696=>"111111111",
  42697=>"100101111",
  42698=>"000010000",
  42699=>"000001111",
  42700=>"100000000",
  42701=>"000011011",
  42702=>"001000000",
  42703=>"100111010",
  42704=>"110000010",
  42705=>"000000000",
  42706=>"000000010",
  42707=>"000000000",
  42708=>"100101101",
  42709=>"000110100",
  42710=>"000111010",
  42711=>"001000101",
  42712=>"000000000",
  42713=>"111110111",
  42714=>"101111111",
  42715=>"110111110",
  42716=>"000000111",
  42717=>"001101111",
  42718=>"100000101",
  42719=>"111001001",
  42720=>"000000000",
  42721=>"000000111",
  42722=>"000010000",
  42723=>"111011000",
  42724=>"000000000",
  42725=>"111111001",
  42726=>"111111111",
  42727=>"111101110",
  42728=>"111000000",
  42729=>"000000000",
  42730=>"101101110",
  42731=>"111111111",
  42732=>"111111111",
  42733=>"000000000",
  42734=>"010001000",
  42735=>"000000000",
  42736=>"111000000",
  42737=>"111111111",
  42738=>"010010000",
  42739=>"111001111",
  42740=>"001101111",
  42741=>"101101111",
  42742=>"100000000",
  42743=>"111100000",
  42744=>"111111111",
  42745=>"111111001",
  42746=>"111110000",
  42747=>"111111111",
  42748=>"000110110",
  42749=>"110100101",
  42750=>"100000000",
  42751=>"111101010",
  42752=>"110100000",
  42753=>"100110100",
  42754=>"111111111",
  42755=>"000000001",
  42756=>"000000000",
  42757=>"110010100",
  42758=>"001001111",
  42759=>"011001111",
  42760=>"111000000",
  42761=>"000000000",
  42762=>"000000000",
  42763=>"001000101",
  42764=>"101101111",
  42765=>"110110000",
  42766=>"100111111",
  42767=>"010000000",
  42768=>"100000000",
  42769=>"101000000",
  42770=>"000001111",
  42771=>"110110010",
  42772=>"010111111",
  42773=>"100000000",
  42774=>"111110111",
  42775=>"111000101",
  42776=>"100110110",
  42777=>"111111111",
  42778=>"111111000",
  42779=>"110010011",
  42780=>"000000000",
  42781=>"111111000",
  42782=>"000000000",
  42783=>"111000000",
  42784=>"101001001",
  42785=>"011011000",
  42786=>"111110000",
  42787=>"111111000",
  42788=>"011111111",
  42789=>"110000000",
  42790=>"001001000",
  42791=>"111001111",
  42792=>"000100000",
  42793=>"111111010",
  42794=>"111111000",
  42795=>"111101111",
  42796=>"111000000",
  42797=>"111110000",
  42798=>"000000000",
  42799=>"101000000",
  42800=>"000000000",
  42801=>"111111110",
  42802=>"000101111",
  42803=>"000000111",
  42804=>"010101011",
  42805=>"000000001",
  42806=>"101111111",
  42807=>"111111111",
  42808=>"011011011",
  42809=>"001000011",
  42810=>"000001111",
  42811=>"111111010",
  42812=>"100000001",
  42813=>"001111000",
  42814=>"001011001",
  42815=>"111000000",
  42816=>"000100000",
  42817=>"001001000",
  42818=>"000000000",
  42819=>"001000000",
  42820=>"000000011",
  42821=>"111000001",
  42822=>"000001111",
  42823=>"101110110",
  42824=>"111001111",
  42825=>"000000000",
  42826=>"111000000",
  42827=>"100100011",
  42828=>"000110111",
  42829=>"111111101",
  42830=>"111110000",
  42831=>"111111111",
  42832=>"101001001",
  42833=>"111000000",
  42834=>"111001001",
  42835=>"111111111",
  42836=>"000000000",
  42837=>"001011010",
  42838=>"000111111",
  42839=>"011001111",
  42840=>"111111111",
  42841=>"011011110",
  42842=>"111000001",
  42843=>"101001101",
  42844=>"111010000",
  42845=>"000000101",
  42846=>"011010000",
  42847=>"111110110",
  42848=>"011001000",
  42849=>"000000001",
  42850=>"100000000",
  42851=>"111101111",
  42852=>"000000111",
  42853=>"111111111",
  42854=>"111111100",
  42855=>"111111111",
  42856=>"000001101",
  42857=>"111101101",
  42858=>"111111111",
  42859=>"111111111",
  42860=>"110110000",
  42861=>"111001000",
  42862=>"110111111",
  42863=>"111000100",
  42864=>"001001110",
  42865=>"000000100",
  42866=>"010111111",
  42867=>"000100110",
  42868=>"000000000",
  42869=>"110101000",
  42870=>"111001000",
  42871=>"000101111",
  42872=>"001001111",
  42873=>"111000111",
  42874=>"000111110",
  42875=>"111111100",
  42876=>"000000000",
  42877=>"110111010",
  42878=>"111000000",
  42879=>"000000000",
  42880=>"100111111",
  42881=>"111101000",
  42882=>"100111111",
  42883=>"010010000",
  42884=>"100000000",
  42885=>"011111111",
  42886=>"000000000",
  42887=>"100000000",
  42888=>"000000000",
  42889=>"101101001",
  42890=>"000111110",
  42891=>"111111011",
  42892=>"101101111",
  42893=>"110100100",
  42894=>"111100000",
  42895=>"001000011",
  42896=>"000000000",
  42897=>"111000000",
  42898=>"000000000",
  42899=>"111001001",
  42900=>"000110111",
  42901=>"000000000",
  42902=>"111111010",
  42903=>"101111111",
  42904=>"111111111",
  42905=>"000001111",
  42906=>"000001101",
  42907=>"001001111",
  42908=>"101101001",
  42909=>"000000001",
  42910=>"111111010",
  42911=>"110100000",
  42912=>"111111000",
  42913=>"011011000",
  42914=>"111010111",
  42915=>"111000111",
  42916=>"101001000",
  42917=>"010000011",
  42918=>"000000000",
  42919=>"010000100",
  42920=>"011011000",
  42921=>"001000000",
  42922=>"111111011",
  42923=>"000000000",
  42924=>"000000011",
  42925=>"111111111",
  42926=>"111000000",
  42927=>"111100000",
  42928=>"001001001",
  42929=>"110100001",
  42930=>"111111111",
  42931=>"111110000",
  42932=>"000000000",
  42933=>"110111111",
  42934=>"111100000",
  42935=>"000000000",
  42936=>"111000100",
  42937=>"001111000",
  42938=>"000000000",
  42939=>"000111111",
  42940=>"011010011",
  42941=>"000000000",
  42942=>"000000101",
  42943=>"111101100",
  42944=>"000010001",
  42945=>"111111111",
  42946=>"111111000",
  42947=>"011000000",
  42948=>"111011111",
  42949=>"101111111",
  42950=>"011011111",
  42951=>"011000000",
  42952=>"101000111",
  42953=>"100100000",
  42954=>"111111000",
  42955=>"110111000",
  42956=>"110000111",
  42957=>"011011000",
  42958=>"011011000",
  42959=>"011000100",
  42960=>"000000000",
  42961=>"000110110",
  42962=>"111111001",
  42963=>"011001111",
  42964=>"111111000",
  42965=>"111110000",
  42966=>"111000100",
  42967=>"111011011",
  42968=>"110000000",
  42969=>"111101010",
  42970=>"111111010",
  42971=>"010010111",
  42972=>"101111111",
  42973=>"001001000",
  42974=>"111011000",
  42975=>"000001111",
  42976=>"000000001",
  42977=>"001111111",
  42978=>"100100111",
  42979=>"001000111",
  42980=>"100000100",
  42981=>"011011011",
  42982=>"000000111",
  42983=>"111111110",
  42984=>"101001111",
  42985=>"111111110",
  42986=>"000001001",
  42987=>"110110000",
  42988=>"001000000",
  42989=>"111111010",
  42990=>"000001011",
  42991=>"001000000",
  42992=>"111111111",
  42993=>"110000000",
  42994=>"110000000",
  42995=>"000000000",
  42996=>"111110111",
  42997=>"111111111",
  42998=>"000100010",
  42999=>"000100111",
  43000=>"011111011",
  43001=>"111101001",
  43002=>"110110110",
  43003=>"111111111",
  43004=>"010010000",
  43005=>"111111111",
  43006=>"000000000",
  43007=>"000000111",
  43008=>"000000000",
  43009=>"011000000",
  43010=>"111111111",
  43011=>"000000000",
  43012=>"111000000",
  43013=>"000111110",
  43014=>"111111111",
  43015=>"111000000",
  43016=>"111001111",
  43017=>"100000000",
  43018=>"011111111",
  43019=>"101001001",
  43020=>"000000100",
  43021=>"101111111",
  43022=>"111000000",
  43023=>"111000000",
  43024=>"111111100",
  43025=>"111001001",
  43026=>"010000000",
  43027=>"111111101",
  43028=>"111111100",
  43029=>"000000111",
  43030=>"100111011",
  43031=>"011000111",
  43032=>"100001111",
  43033=>"000101111",
  43034=>"111101111",
  43035=>"110000000",
  43036=>"001111111",
  43037=>"111111111",
  43038=>"000110100",
  43039=>"111000000",
  43040=>"111111111",
  43041=>"111111111",
  43042=>"000111111",
  43043=>"001000001",
  43044=>"000000001",
  43045=>"111011111",
  43046=>"111111000",
  43047=>"101011000",
  43048=>"101000000",
  43049=>"000000111",
  43050=>"011011111",
  43051=>"111110111",
  43052=>"110000110",
  43053=>"110110000",
  43054=>"000000110",
  43055=>"100000111",
  43056=>"111111111",
  43057=>"111111000",
  43058=>"001011000",
  43059=>"111111000",
  43060=>"001000110",
  43061=>"011011011",
  43062=>"111000000",
  43063=>"111110000",
  43064=>"001000111",
  43065=>"111100111",
  43066=>"111111111",
  43067=>"001111111",
  43068=>"111111000",
  43069=>"000000000",
  43070=>"100000000",
  43071=>"000010011",
  43072=>"100110111",
  43073=>"110111000",
  43074=>"000101111",
  43075=>"111000011",
  43076=>"110100000",
  43077=>"001000001",
  43078=>"111111000",
  43079=>"111111111",
  43080=>"001011111",
  43081=>"101001111",
  43082=>"011110110",
  43083=>"111111011",
  43084=>"001111111",
  43085=>"100000000",
  43086=>"100000000",
  43087=>"001000000",
  43088=>"000000000",
  43089=>"001001010",
  43090=>"111011000",
  43091=>"111111000",
  43092=>"000000000",
  43093=>"000000001",
  43094=>"111101100",
  43095=>"000111111",
  43096=>"111000000",
  43097=>"111111000",
  43098=>"000100110",
  43099=>"100110110",
  43100=>"000111000",
  43101=>"000110111",
  43102=>"000011111",
  43103=>"111110100",
  43104=>"010000000",
  43105=>"011001011",
  43106=>"000011000",
  43107=>"111001000",
  43108=>"111111111",
  43109=>"111111001",
  43110=>"001000000",
  43111=>"000000000",
  43112=>"001111001",
  43113=>"011111110",
  43114=>"000000111",
  43115=>"111111000",
  43116=>"000000000",
  43117=>"110110000",
  43118=>"110010111",
  43119=>"111111111",
  43120=>"000110000",
  43121=>"111000001",
  43122=>"001011000",
  43123=>"111110111",
  43124=>"100000000",
  43125=>"000111111",
  43126=>"001111010",
  43127=>"000111111",
  43128=>"000000000",
  43129=>"011000110",
  43130=>"111100000",
  43131=>"111000000",
  43132=>"100000100",
  43133=>"000100111",
  43134=>"100110111",
  43135=>"010000000",
  43136=>"000000000",
  43137=>"111000111",
  43138=>"001000000",
  43139=>"111011000",
  43140=>"100000011",
  43141=>"000000000",
  43142=>"111000001",
  43143=>"110110111",
  43144=>"111100111",
  43145=>"111111111",
  43146=>"001011011",
  43147=>"000000000",
  43148=>"000000000",
  43149=>"000111111",
  43150=>"111011111",
  43151=>"111110000",
  43152=>"000111111",
  43153=>"000000000",
  43154=>"100000111",
  43155=>"000001000",
  43156=>"000000001",
  43157=>"111100111",
  43158=>"111110100",
  43159=>"111000110",
  43160=>"000100110",
  43161=>"111011010",
  43162=>"111111110",
  43163=>"111110010",
  43164=>"000000000",
  43165=>"111111100",
  43166=>"000000111",
  43167=>"000000000",
  43168=>"000100000",
  43169=>"111111111",
  43170=>"011111111",
  43171=>"000110110",
  43172=>"111001000",
  43173=>"100100011",
  43174=>"110100000",
  43175=>"100110111",
  43176=>"111100000",
  43177=>"111111000",
  43178=>"111111111",
  43179=>"000000111",
  43180=>"100100111",
  43181=>"001110110",
  43182=>"000000000",
  43183=>"100110111",
  43184=>"111101000",
  43185=>"110000000",
  43186=>"111111011",
  43187=>"000000000",
  43188=>"111111111",
  43189=>"100000000",
  43190=>"000111111",
  43191=>"000011000",
  43192=>"000000000",
  43193=>"011000000",
  43194=>"111101000",
  43195=>"100100111",
  43196=>"000000000",
  43197=>"010010111",
  43198=>"111100111",
  43199=>"000000001",
  43200=>"100111001",
  43201=>"000000111",
  43202=>"111111000",
  43203=>"110000100",
  43204=>"111111111",
  43205=>"111000000",
  43206=>"101000100",
  43207=>"000110000",
  43208=>"011111111",
  43209=>"111111011",
  43210=>"111000000",
  43211=>"000010011",
  43212=>"000111111",
  43213=>"110100100",
  43214=>"111110000",
  43215=>"111111111",
  43216=>"100100000",
  43217=>"011010000",
  43218=>"110100100",
  43219=>"100000100",
  43220=>"111111111",
  43221=>"011001111",
  43222=>"000000000",
  43223=>"111111101",
  43224=>"000111111",
  43225=>"111111111",
  43226=>"001011000",
  43227=>"000000111",
  43228=>"000000000",
  43229=>"111111111",
  43230=>"001001111",
  43231=>"110011111",
  43232=>"111111000",
  43233=>"000000010",
  43234=>"010000100",
  43235=>"000000000",
  43236=>"011010111",
  43237=>"010000000",
  43238=>"111111000",
  43239=>"111110111",
  43240=>"111111111",
  43241=>"110100000",
  43242=>"110000000",
  43243=>"100000000",
  43244=>"000100111",
  43245=>"111000000",
  43246=>"111111001",
  43247=>"101000000",
  43248=>"110000000",
  43249=>"111000000",
  43250=>"111111011",
  43251=>"110000000",
  43252=>"000000000",
  43253=>"010111001",
  43254=>"001001011",
  43255=>"000000111",
  43256=>"111111000",
  43257=>"100000000",
  43258=>"111111111",
  43259=>"011001000",
  43260=>"000000100",
  43261=>"001011111",
  43262=>"111111111",
  43263=>"111100111",
  43264=>"100000000",
  43265=>"001001000",
  43266=>"000000000",
  43267=>"100101111",
  43268=>"011110111",
  43269=>"000000000",
  43270=>"001110111",
  43271=>"110000010",
  43272=>"101100000",
  43273=>"000000000",
  43274=>"100000001",
  43275=>"111111011",
  43276=>"111000000",
  43277=>"000110111",
  43278=>"000000000",
  43279=>"001111111",
  43280=>"110000000",
  43281=>"111110111",
  43282=>"001001111",
  43283=>"000000011",
  43284=>"101011001",
  43285=>"000000000",
  43286=>"001001001",
  43287=>"111111111",
  43288=>"000000000",
  43289=>"110100100",
  43290=>"111111111",
  43291=>"000000000",
  43292=>"100111111",
  43293=>"000000000",
  43294=>"011111111",
  43295=>"000110000",
  43296=>"111111111",
  43297=>"011000000",
  43298=>"000011111",
  43299=>"000000000",
  43300=>"011001000",
  43301=>"101000000",
  43302=>"000111001",
  43303=>"111110110",
  43304=>"010110100",
  43305=>"010010110",
  43306=>"111111111",
  43307=>"111000000",
  43308=>"111111000",
  43309=>"110111111",
  43310=>"000101000",
  43311=>"111001000",
  43312=>"000000110",
  43313=>"000100110",
  43314=>"111111011",
  43315=>"000010011",
  43316=>"100110100",
  43317=>"100000111",
  43318=>"000111111",
  43319=>"001000000",
  43320=>"111000000",
  43321=>"111000000",
  43322=>"000100111",
  43323=>"110111111",
  43324=>"000000000",
  43325=>"100000000",
  43326=>"001000000",
  43327=>"110111111",
  43328=>"111000100",
  43329=>"000000110",
  43330=>"111011111",
  43331=>"000001011",
  43332=>"101001000",
  43333=>"000101111",
  43334=>"111101000",
  43335=>"100000000",
  43336=>"000000000",
  43337=>"110111111",
  43338=>"001000000",
  43339=>"110110000",
  43340=>"000100110",
  43341=>"011011000",
  43342=>"100111100",
  43343=>"001001001",
  43344=>"111111111",
  43345=>"110010111",
  43346=>"000000000",
  43347=>"111111000",
  43348=>"111111000",
  43349=>"001001011",
  43350=>"110110111",
  43351=>"100000011",
  43352=>"110010011",
  43353=>"111111000",
  43354=>"011000000",
  43355=>"111111011",
  43356=>"000000111",
  43357=>"000000000",
  43358=>"111111000",
  43359=>"000000000",
  43360=>"000000100",
  43361=>"111111001",
  43362=>"000001001",
  43363=>"111111000",
  43364=>"010000000",
  43365=>"000000000",
  43366=>"111000000",
  43367=>"111111000",
  43368=>"001110111",
  43369=>"010000000",
  43370=>"000011111",
  43371=>"111111000",
  43372=>"100110110",
  43373=>"100000100",
  43374=>"000000000",
  43375=>"111001000",
  43376=>"110110010",
  43377=>"000010001",
  43378=>"111111100",
  43379=>"100100000",
  43380=>"111000011",
  43381=>"111111111",
  43382=>"001000111",
  43383=>"001000000",
  43384=>"111111000",
  43385=>"111111111",
  43386=>"000000000",
  43387=>"000000000",
  43388=>"111111111",
  43389=>"111000000",
  43390=>"111111111",
  43391=>"001000111",
  43392=>"111111011",
  43393=>"000000111",
  43394=>"100110111",
  43395=>"111001001",
  43396=>"111111000",
  43397=>"110010110",
  43398=>"101111000",
  43399=>"111111111",
  43400=>"000011111",
  43401=>"100001101",
  43402=>"111111010",
  43403=>"000110000",
  43404=>"001000111",
  43405=>"000000000",
  43406=>"010001011",
  43407=>"111000000",
  43408=>"110110000",
  43409=>"111111111",
  43410=>"111111110",
  43411=>"100100111",
  43412=>"111111000",
  43413=>"010010000",
  43414=>"111111111",
  43415=>"001001001",
  43416=>"000011111",
  43417=>"011001011",
  43418=>"111111111",
  43419=>"001000001",
  43420=>"111111111",
  43421=>"000100110",
  43422=>"000000000",
  43423=>"111111111",
  43424=>"110110111",
  43425=>"011011011",
  43426=>"111001001",
  43427=>"000000010",
  43428=>"111001011",
  43429=>"011011010",
  43430=>"111000000",
  43431=>"101111111",
  43432=>"000011010",
  43433=>"000010110",
  43434=>"111111000",
  43435=>"111111000",
  43436=>"111110000",
  43437=>"000000000",
  43438=>"000100111",
  43439=>"001111011",
  43440=>"000000000",
  43441=>"010110111",
  43442=>"001001000",
  43443=>"111111000",
  43444=>"100000000",
  43445=>"011011111",
  43446=>"000000011",
  43447=>"110110110",
  43448=>"000000111",
  43449=>"100000000",
  43450=>"111111110",
  43451=>"111111111",
  43452=>"000101001",
  43453=>"111101011",
  43454=>"000111111",
  43455=>"000111000",
  43456=>"111111111",
  43457=>"001101111",
  43458=>"111000000",
  43459=>"111111000",
  43460=>"101001000",
  43461=>"101001111",
  43462=>"100000000",
  43463=>"111111110",
  43464=>"100000000",
  43465=>"111101110",
  43466=>"100000000",
  43467=>"011000000",
  43468=>"111010000",
  43469=>"011000000",
  43470=>"000000010",
  43471=>"111010011",
  43472=>"000010111",
  43473=>"000001001",
  43474=>"100000010",
  43475=>"010011111",
  43476=>"111001000",
  43477=>"001111000",
  43478=>"000000000",
  43479=>"011011001",
  43480=>"000000000",
  43481=>"000001111",
  43482=>"000000000",
  43483=>"011111111",
  43484=>"000000111",
  43485=>"111100111",
  43486=>"011011011",
  43487=>"100100111",
  43488=>"011011111",
  43489=>"111111111",
  43490=>"111111110",
  43491=>"000110111",
  43492=>"000111111",
  43493=>"111011001",
  43494=>"111100110",
  43495=>"111111111",
  43496=>"001010000",
  43497=>"110100000",
  43498=>"000011000",
  43499=>"000000111",
  43500=>"011001101",
  43501=>"100000000",
  43502=>"001011111",
  43503=>"111111000",
  43504=>"111111100",
  43505=>"000000011",
  43506=>"111011011",
  43507=>"101110111",
  43508=>"111000111",
  43509=>"110111100",
  43510=>"000000000",
  43511=>"110100110",
  43512=>"111111111",
  43513=>"111101101",
  43514=>"111000000",
  43515=>"110000111",
  43516=>"111111111",
  43517=>"111110000",
  43518=>"101000000",
  43519=>"001001001",
  43520=>"111111111",
  43521=>"000000000",
  43522=>"111000000",
  43523=>"000000000",
  43524=>"000000011",
  43525=>"100000000",
  43526=>"110010000",
  43527=>"000001101",
  43528=>"000000000",
  43529=>"011000100",
  43530=>"100100000",
  43531=>"000001011",
  43532=>"100010010",
  43533=>"000011111",
  43534=>"000001001",
  43535=>"111111111",
  43536=>"100100000",
  43537=>"000000100",
  43538=>"110001000",
  43539=>"111111111",
  43540=>"000110111",
  43541=>"010000000",
  43542=>"111111111",
  43543=>"111111111",
  43544=>"111111111",
  43545=>"100000000",
  43546=>"000011111",
  43547=>"101100000",
  43548=>"000001111",
  43549=>"011001111",
  43550=>"111111011",
  43551=>"000000000",
  43552=>"111111111",
  43553=>"100000000",
  43554=>"011001000",
  43555=>"010110111",
  43556=>"000100110",
  43557=>"010111100",
  43558=>"111111111",
  43559=>"110111111",
  43560=>"000101011",
  43561=>"000000000",
  43562=>"110111101",
  43563=>"000110000",
  43564=>"111111111",
  43565=>"000111111",
  43566=>"000010000",
  43567=>"111110010",
  43568=>"111010111",
  43569=>"110010010",
  43570=>"111111111",
  43571=>"000000011",
  43572=>"111011111",
  43573=>"111111111",
  43574=>"000001011",
  43575=>"000000111",
  43576=>"000000000",
  43577=>"011000101",
  43578=>"110010000",
  43579=>"011011010",
  43580=>"111111111",
  43581=>"111111011",
  43582=>"111111101",
  43583=>"000000000",
  43584=>"000000000",
  43585=>"111111111",
  43586=>"000000000",
  43587=>"000000000",
  43588=>"110110110",
  43589=>"111111111",
  43590=>"000010011",
  43591=>"110010111",
  43592=>"110011011",
  43593=>"001001000",
  43594=>"100111111",
  43595=>"000000001",
  43596=>"111111111",
  43597=>"000000000",
  43598=>"000000000",
  43599=>"000001111",
  43600=>"111111111",
  43601=>"110110101",
  43602=>"000000000",
  43603=>"000110110",
  43604=>"000000010",
  43605=>"000000000",
  43606=>"000000011",
  43607=>"001000111",
  43608=>"000000000",
  43609=>"100101101",
  43610=>"000000000",
  43611=>"100110110",
  43612=>"000000000",
  43613=>"110000111",
  43614=>"000100111",
  43615=>"000000000",
  43616=>"000000010",
  43617=>"110000110",
  43618=>"001011000",
  43619=>"000110000",
  43620=>"000000000",
  43621=>"101000000",
  43622=>"000000110",
  43623=>"000000000",
  43624=>"111011001",
  43625=>"111000000",
  43626=>"000000111",
  43627=>"000000000",
  43628=>"000000111",
  43629=>"000000000",
  43630=>"111111100",
  43631=>"010010000",
  43632=>"000000000",
  43633=>"000110111",
  43634=>"111111011",
  43635=>"111011000",
  43636=>"100000101",
  43637=>"000000000",
  43638=>"000000001",
  43639=>"100111111",
  43640=>"111000011",
  43641=>"100010010",
  43642=>"000000000",
  43643=>"000010111",
  43644=>"110110110",
  43645=>"110110111",
  43646=>"000000000",
  43647=>"000000011",
  43648=>"111111011",
  43649=>"000000110",
  43650=>"000000000",
  43651=>"000011011",
  43652=>"001111111",
  43653=>"001011111",
  43654=>"111110100",
  43655=>"111111011",
  43656=>"000100000",
  43657=>"100000110",
  43658=>"000000000",
  43659=>"000000011",
  43660=>"111111001",
  43661=>"110011011",
  43662=>"000000111",
  43663=>"110111111",
  43664=>"000000000",
  43665=>"011001111",
  43666=>"100100111",
  43667=>"111001011",
  43668=>"110000000",
  43669=>"110111000",
  43670=>"000011111",
  43671=>"111111111",
  43672=>"000001000",
  43673=>"000011111",
  43674=>"110000011",
  43675=>"000000000",
  43676=>"000000111",
  43677=>"000000000",
  43678=>"100001111",
  43679=>"111111110",
  43680=>"111000111",
  43681=>"110000000",
  43682=>"110110110",
  43683=>"011111111",
  43684=>"011011000",
  43685=>"000000000",
  43686=>"111010010",
  43687=>"111011011",
  43688=>"011111111",
  43689=>"011001000",
  43690=>"111111111",
  43691=>"001001111",
  43692=>"001111111",
  43693=>"000001100",
  43694=>"111111111",
  43695=>"111111000",
  43696=>"000000000",
  43697=>"111011011",
  43698=>"111111011",
  43699=>"000000111",
  43700=>"111110110",
  43701=>"100000000",
  43702=>"010000110",
  43703=>"000000000",
  43704=>"000000001",
  43705=>"111111111",
  43706=>"010000000",
  43707=>"000000000",
  43708=>"000000000",
  43709=>"000000000",
  43710=>"000101100",
  43711=>"100110111",
  43712=>"000100111",
  43713=>"000000011",
  43714=>"111111100",
  43715=>"000000000",
  43716=>"111111111",
  43717=>"111111001",
  43718=>"111111111",
  43719=>"001101111",
  43720=>"000111101",
  43721=>"100101111",
  43722=>"001111011",
  43723=>"111110100",
  43724=>"101100011",
  43725=>"000111111",
  43726=>"010010010",
  43727=>"111101001",
  43728=>"000000000",
  43729=>"000000000",
  43730=>"000000000",
  43731=>"000000000",
  43732=>"111000011",
  43733=>"111001111",
  43734=>"000000000",
  43735=>"100111111",
  43736=>"000000000",
  43737=>"111111111",
  43738=>"000000010",
  43739=>"111110000",
  43740=>"000000010",
  43741=>"000000010",
  43742=>"111000101",
  43743=>"111111101",
  43744=>"000000000",
  43745=>"000000111",
  43746=>"111111111",
  43747=>"111111100",
  43748=>"101111000",
  43749=>"001111111",
  43750=>"000000000",
  43751=>"111111001",
  43752=>"001000111",
  43753=>"110011001",
  43754=>"001111000",
  43755=>"101111111",
  43756=>"111111010",
  43757=>"000000000",
  43758=>"111111100",
  43759=>"000010000",
  43760=>"000000111",
  43761=>"011111001",
  43762=>"000000110",
  43763=>"000000100",
  43764=>"111110111",
  43765=>"000000000",
  43766=>"111111011",
  43767=>"000000000",
  43768=>"000000000",
  43769=>"111111100",
  43770=>"000000010",
  43771=>"111111111",
  43772=>"011011111",
  43773=>"111100100",
  43774=>"010000011",
  43775=>"000000000",
  43776=>"110100011",
  43777=>"111011011",
  43778=>"000000000",
  43779=>"000000000",
  43780=>"001000000",
  43781=>"110100000",
  43782=>"111111111",
  43783=>"100100110",
  43784=>"000000111",
  43785=>"000000000",
  43786=>"111111100",
  43787=>"000000001",
  43788=>"001001001",
  43789=>"111001001",
  43790=>"000001011",
  43791=>"111111111",
  43792=>"000000000",
  43793=>"111111111",
  43794=>"011011010",
  43795=>"111111101",
  43796=>"111011000",
  43797=>"010000011",
  43798=>"111001001",
  43799=>"000000000",
  43800=>"110110111",
  43801=>"111111110",
  43802=>"000000001",
  43803=>"111110000",
  43804=>"000000110",
  43805=>"111110000",
  43806=>"111111111",
  43807=>"000000000",
  43808=>"110011000",
  43809=>"000000000",
  43810=>"000010100",
  43811=>"000110010",
  43812=>"111111111",
  43813=>"111000001",
  43814=>"111011011",
  43815=>"000000000",
  43816=>"111101000",
  43817=>"001001111",
  43818=>"110000000",
  43819=>"100111001",
  43820=>"000000111",
  43821=>"001001111",
  43822=>"000000000",
  43823=>"111111011",
  43824=>"111111111",
  43825=>"000000000",
  43826=>"111111010",
  43827=>"110000000",
  43828=>"010000110",
  43829=>"100000101",
  43830=>"001001001",
  43831=>"000000001",
  43832=>"111111101",
  43833=>"000000000",
  43834=>"000000000",
  43835=>"000111110",
  43836=>"111111011",
  43837=>"101001000",
  43838=>"111111000",
  43839=>"111111111",
  43840=>"111000000",
  43841=>"010000100",
  43842=>"000000000",
  43843=>"111111111",
  43844=>"111111011",
  43845=>"000000000",
  43846=>"000000001",
  43847=>"100000000",
  43848=>"111111111",
  43849=>"000000000",
  43850=>"000000000",
  43851=>"001001001",
  43852=>"111111000",
  43853=>"011000011",
  43854=>"000111111",
  43855=>"001001001",
  43856=>"100000000",
  43857=>"110110100",
  43858=>"110011011",
  43859=>"111111111",
  43860=>"111000000",
  43861=>"011011111",
  43862=>"111000000",
  43863=>"011000000",
  43864=>"000000001",
  43865=>"111111000",
  43866=>"111011000",
  43867=>"000000000",
  43868=>"111111100",
  43869=>"000000110",
  43870=>"000000000",
  43871=>"110111001",
  43872=>"000000000",
  43873=>"011110011",
  43874=>"111111110",
  43875=>"110010111",
  43876=>"010000110",
  43877=>"111111101",
  43878=>"100100110",
  43879=>"111111111",
  43880=>"110010000",
  43881=>"000000000",
  43882=>"000000100",
  43883=>"111101011",
  43884=>"110001001",
  43885=>"000000111",
  43886=>"111111101",
  43887=>"011111111",
  43888=>"110110000",
  43889=>"000000000",
  43890=>"011011100",
  43891=>"011011011",
  43892=>"000000111",
  43893=>"111111111",
  43894=>"010111010",
  43895=>"000000000",
  43896=>"000000111",
  43897=>"100000011",
  43898=>"000000000",
  43899=>"111111100",
  43900=>"000001000",
  43901=>"000001111",
  43902=>"111011000",
  43903=>"111111100",
  43904=>"110010011",
  43905=>"010110111",
  43906=>"110011011",
  43907=>"000000000",
  43908=>"000000000",
  43909=>"000000000",
  43910=>"100111111",
  43911=>"100000000",
  43912=>"110010000",
  43913=>"000100000",
  43914=>"110111111",
  43915=>"100000000",
  43916=>"000000000",
  43917=>"100000011",
  43918=>"000101111",
  43919=>"111111111",
  43920=>"111110111",
  43921=>"000100110",
  43922=>"110110100",
  43923=>"111111000",
  43924=>"111111110",
  43925=>"000000111",
  43926=>"011001011",
  43927=>"111001100",
  43928=>"000000000",
  43929=>"110110111",
  43930=>"000000000",
  43931=>"000011011",
  43932=>"000000001",
  43933=>"111111111",
  43934=>"010000000",
  43935=>"100100100",
  43936=>"011000000",
  43937=>"110000000",
  43938=>"000010111",
  43939=>"010011111",
  43940=>"000001000",
  43941=>"000010111",
  43942=>"010000000",
  43943=>"000000000",
  43944=>"111100010",
  43945=>"000000000",
  43946=>"000000000",
  43947=>"000001000",
  43948=>"000000000",
  43949=>"111111000",
  43950=>"000100111",
  43951=>"000000000",
  43952=>"000000000",
  43953=>"000000000",
  43954=>"011001001",
  43955=>"110100110",
  43956=>"001000000",
  43957=>"000000000",
  43958=>"111101111",
  43959=>"100101111",
  43960=>"000100000",
  43961=>"000000000",
  43962=>"111000000",
  43963=>"000101111",
  43964=>"000000111",
  43965=>"100111111",
  43966=>"111000000",
  43967=>"111000000",
  43968=>"110010010",
  43969=>"000001001",
  43970=>"111011111",
  43971=>"111111100",
  43972=>"100111100",
  43973=>"001001100",
  43974=>"111111111",
  43975=>"000000000",
  43976=>"000000000",
  43977=>"000000111",
  43978=>"000000110",
  43979=>"001111111",
  43980=>"000000000",
  43981=>"001000000",
  43982=>"111000000",
  43983=>"111111000",
  43984=>"000000000",
  43985=>"011111111",
  43986=>"111111001",
  43987=>"001011111",
  43988=>"001011011",
  43989=>"100000001",
  43990=>"111011111",
  43991=>"011001001",
  43992=>"000110110",
  43993=>"111000111",
  43994=>"001111000",
  43995=>"110000000",
  43996=>"111011011",
  43997=>"000101111",
  43998=>"111011001",
  43999=>"011011111",
  44000=>"111100100",
  44001=>"000000001",
  44002=>"000000000",
  44003=>"111111111",
  44004=>"111010000",
  44005=>"000000000",
  44006=>"111000000",
  44007=>"000000000",
  44008=>"111000001",
  44009=>"110011001",
  44010=>"000000011",
  44011=>"000000011",
  44012=>"000000000",
  44013=>"001000001",
  44014=>"111111111",
  44015=>"011001001",
  44016=>"000000000",
  44017=>"111000111",
  44018=>"111110000",
  44019=>"000000000",
  44020=>"000110011",
  44021=>"000000100",
  44022=>"111111111",
  44023=>"111000000",
  44024=>"000000111",
  44025=>"111101101",
  44026=>"111101001",
  44027=>"111111111",
  44028=>"100111110",
  44029=>"110111111",
  44030=>"111111110",
  44031=>"111111000",
  44032=>"111111111",
  44033=>"001000000",
  44034=>"111111111",
  44035=>"000000000",
  44036=>"000000000",
  44037=>"111111111",
  44038=>"000000000",
  44039=>"111111111",
  44040=>"111111111",
  44041=>"000000000",
  44042=>"000000000",
  44043=>"011110010",
  44044=>"110000000",
  44045=>"101111111",
  44046=>"000111111",
  44047=>"001001001",
  44048=>"111111111",
  44049=>"000001111",
  44050=>"011001101",
  44051=>"100000000",
  44052=>"111111111",
  44053=>"100000100",
  44054=>"111110000",
  44055=>"011011001",
  44056=>"010000001",
  44057=>"000000000",
  44058=>"000000000",
  44059=>"000001011",
  44060=>"000000111",
  44061=>"000000000",
  44062=>"001010010",
  44063=>"000000011",
  44064=>"000001001",
  44065=>"000000010",
  44066=>"000101111",
  44067=>"000101111",
  44068=>"111000000",
  44069=>"001111011",
  44070=>"111111111",
  44071=>"000000001",
  44072=>"111111111",
  44073=>"110010110",
  44074=>"000011011",
  44075=>"110100000",
  44076=>"110111000",
  44077=>"000000000",
  44078=>"111111111",
  44079=>"000000000",
  44080=>"110111110",
  44081=>"000000000",
  44082=>"001000000",
  44083=>"000000000",
  44084=>"111101100",
  44085=>"000000000",
  44086=>"111111110",
  44087=>"000000000",
  44088=>"111111111",
  44089=>"000000000",
  44090=>"100100110",
  44091=>"110100000",
  44092=>"111111000",
  44093=>"111111110",
  44094=>"011000100",
  44095=>"011000000",
  44096=>"110001001",
  44097=>"000110110",
  44098=>"000111011",
  44099=>"000011000",
  44100=>"001001000",
  44101=>"001011001",
  44102=>"110000100",
  44103=>"100000000",
  44104=>"001001000",
  44105=>"111111010",
  44106=>"000000000",
  44107=>"111111111",
  44108=>"111110010",
  44109=>"000001111",
  44110=>"111111111",
  44111=>"111010000",
  44112=>"000100111",
  44113=>"000000100",
  44114=>"011111000",
  44115=>"011111111",
  44116=>"001000110",
  44117=>"110110110",
  44118=>"000100000",
  44119=>"000000000",
  44120=>"101100101",
  44121=>"111000000",
  44122=>"110110111",
  44123=>"011111111",
  44124=>"111111111",
  44125=>"000000000",
  44126=>"001001001",
  44127=>"111111100",
  44128=>"111111111",
  44129=>"111110010",
  44130=>"110111100",
  44131=>"111111000",
  44132=>"111111110",
  44133=>"111101001",
  44134=>"000000000",
  44135=>"000100111",
  44136=>"000111111",
  44137=>"111111111",
  44138=>"110111111",
  44139=>"011000000",
  44140=>"110111001",
  44141=>"111011111",
  44142=>"111111111",
  44143=>"111111111",
  44144=>"000000000",
  44145=>"000001011",
  44146=>"111100111",
  44147=>"111111111",
  44148=>"000000100",
  44149=>"111111001",
  44150=>"100000000",
  44151=>"000000011",
  44152=>"000000000",
  44153=>"001000000",
  44154=>"000000111",
  44155=>"010000000",
  44156=>"000000000",
  44157=>"111111111",
  44158=>"000000000",
  44159=>"111111111",
  44160=>"111111000",
  44161=>"111010000",
  44162=>"111000000",
  44163=>"111111111",
  44164=>"100100111",
  44165=>"000110111",
  44166=>"000000000",
  44167=>"100000010",
  44168=>"111111111",
  44169=>"010000000",
  44170=>"111111111",
  44171=>"000000000",
  44172=>"111111111",
  44173=>"000100111",
  44174=>"111111000",
  44175=>"001010111",
  44176=>"100100111",
  44177=>"111101111",
  44178=>"101101111",
  44179=>"110110111",
  44180=>"000000000",
  44181=>"111111111",
  44182=>"101100100",
  44183=>"111111111",
  44184=>"000000000",
  44185=>"000001000",
  44186=>"010000000",
  44187=>"000100111",
  44188=>"010110111",
  44189=>"011111111",
  44190=>"011000111",
  44191=>"000000000",
  44192=>"000100000",
  44193=>"011111111",
  44194=>"111111111",
  44195=>"111111111",
  44196=>"000111000",
  44197=>"111111011",
  44198=>"000000100",
  44199=>"010010010",
  44200=>"110010000",
  44201=>"001011011",
  44202=>"001001000",
  44203=>"111000000",
  44204=>"110111111",
  44205=>"010000000",
  44206=>"001111111",
  44207=>"101100111",
  44208=>"111111111",
  44209=>"011111111",
  44210=>"111111111",
  44211=>"110100000",
  44212=>"011111111",
  44213=>"111111111",
  44214=>"101101100",
  44215=>"110111111",
  44216=>"111000000",
  44217=>"000000000",
  44218=>"111101000",
  44219=>"000000111",
  44220=>"000000001",
  44221=>"101000100",
  44222=>"110111110",
  44223=>"011111000",
  44224=>"001000001",
  44225=>"111000001",
  44226=>"011011000",
  44227=>"000000000",
  44228=>"111111111",
  44229=>"000000111",
  44230=>"001100111",
  44231=>"000110111",
  44232=>"100100111",
  44233=>"000000000",
  44234=>"111011001",
  44235=>"111111111",
  44236=>"000111111",
  44237=>"000000011",
  44238=>"100011000",
  44239=>"111111111",
  44240=>"111001011",
  44241=>"111001011",
  44242=>"110111111",
  44243=>"000010111",
  44244=>"111001101",
  44245=>"000111111",
  44246=>"000000110",
  44247=>"111111111",
  44248=>"000011111",
  44249=>"000100110",
  44250=>"111111111",
  44251=>"111111111",
  44252=>"000000100",
  44253=>"111110000",
  44254=>"111100111",
  44255=>"000000000",
  44256=>"010011111",
  44257=>"000011011",
  44258=>"000000110",
  44259=>"111111111",
  44260=>"011010011",
  44261=>"100100110",
  44262=>"000000001",
  44263=>"111111111",
  44264=>"111111001",
  44265=>"000000000",
  44266=>"000100111",
  44267=>"001111111",
  44268=>"111111111",
  44269=>"111110000",
  44270=>"000111111",
  44271=>"000000000",
  44272=>"100100000",
  44273=>"100000000",
  44274=>"111000111",
  44275=>"000000011",
  44276=>"000000110",
  44277=>"110100000",
  44278=>"011010111",
  44279=>"000000100",
  44280=>"000000000",
  44281=>"111111111",
  44282=>"000000000",
  44283=>"111111111",
  44284=>"111111111",
  44285=>"000000000",
  44286=>"000000111",
  44287=>"001000000",
  44288=>"001111111",
  44289=>"111000000",
  44290=>"010001001",
  44291=>"111111111",
  44292=>"001111011",
  44293=>"101000111",
  44294=>"000000000",
  44295=>"111111111",
  44296=>"100111110",
  44297=>"010000110",
  44298=>"000111111",
  44299=>"000000000",
  44300=>"110000000",
  44301=>"111111111",
  44302=>"000000111",
  44303=>"000000011",
  44304=>"000000000",
  44305=>"001000000",
  44306=>"111000000",
  44307=>"001000000",
  44308=>"111011011",
  44309=>"111001000",
  44310=>"000000000",
  44311=>"001111011",
  44312=>"011000001",
  44313=>"111111111",
  44314=>"111111011",
  44315=>"111111111",
  44316=>"110111110",
  44317=>"000000000",
  44318=>"000000000",
  44319=>"111001111",
  44320=>"000101011",
  44321=>"011001000",
  44322=>"000111111",
  44323=>"000011011",
  44324=>"111111000",
  44325=>"000000000",
  44326=>"000000111",
  44327=>"111111111",
  44328=>"100000111",
  44329=>"000111111",
  44330=>"111101111",
  44331=>"100111000",
  44332=>"110111111",
  44333=>"000000000",
  44334=>"000111111",
  44335=>"111110000",
  44336=>"011111111",
  44337=>"011111111",
  44338=>"111110111",
  44339=>"000000010",
  44340=>"111100110",
  44341=>"100100100",
  44342=>"001011000",
  44343=>"100100100",
  44344=>"000000000",
  44345=>"000000100",
  44346=>"000000011",
  44347=>"000111111",
  44348=>"000000000",
  44349=>"000000000",
  44350=>"011101001",
  44351=>"000011111",
  44352=>"111111111",
  44353=>"111111111",
  44354=>"001000000",
  44355=>"111000000",
  44356=>"000000000",
  44357=>"110111110",
  44358=>"000000000",
  44359=>"100111111",
  44360=>"000000000",
  44361=>"111111100",
  44362=>"011011001",
  44363=>"110100100",
  44364=>"111111111",
  44365=>"100110111",
  44366=>"001111111",
  44367=>"111111111",
  44368=>"110001011",
  44369=>"000000000",
  44370=>"000000100",
  44371=>"000001000",
  44372=>"000101111",
  44373=>"011011011",
  44374=>"000000000",
  44375=>"101100000",
  44376=>"000000000",
  44377=>"000000000",
  44378=>"111000000",
  44379=>"001111111",
  44380=>"111111111",
  44381=>"101101000",
  44382=>"011001001",
  44383=>"000001000",
  44384=>"001001000",
  44385=>"001000000",
  44386=>"000111111",
  44387=>"111001111",
  44388=>"011000000",
  44389=>"000000000",
  44390=>"011001111",
  44391=>"000000100",
  44392=>"010011011",
  44393=>"111011000",
  44394=>"000000111",
  44395=>"111111000",
  44396=>"010001101",
  44397=>"101000000",
  44398=>"000000000",
  44399=>"100100000",
  44400=>"100100100",
  44401=>"000000000",
  44402=>"111111011",
  44403=>"000000001",
  44404=>"000010011",
  44405=>"000100101",
  44406=>"000001000",
  44407=>"000000000",
  44408=>"111011111",
  44409=>"000000000",
  44410=>"000000011",
  44411=>"000000111",
  44412=>"111111001",
  44413=>"111111111",
  44414=>"111111111",
  44415=>"111111111",
  44416=>"011111111",
  44417=>"000001001",
  44418=>"110110110",
  44419=>"000000100",
  44420=>"010011001",
  44421=>"111111000",
  44422=>"110110111",
  44423=>"000000000",
  44424=>"111111111",
  44425=>"011111111",
  44426=>"011011011",
  44427=>"111000100",
  44428=>"111111000",
  44429=>"100000000",
  44430=>"000000011",
  44431=>"100111000",
  44432=>"111011011",
  44433=>"111111111",
  44434=>"111100111",
  44435=>"000000000",
  44436=>"000011111",
  44437=>"010011000",
  44438=>"111110000",
  44439=>"011111000",
  44440=>"011111111",
  44441=>"111001000",
  44442=>"000000000",
  44443=>"011111111",
  44444=>"000000000",
  44445=>"111111111",
  44446=>"100000110",
  44447=>"000000000",
  44448=>"001000000",
  44449=>"111110111",
  44450=>"111111110",
  44451=>"000000000",
  44452=>"111111000",
  44453=>"110111111",
  44454=>"000000111",
  44455=>"101001001",
  44456=>"000000100",
  44457=>"111011111",
  44458=>"001000000",
  44459=>"001000100",
  44460=>"000000000",
  44461=>"000000110",
  44462=>"100111011",
  44463=>"111000000",
  44464=>"000100100",
  44465=>"110110011",
  44466=>"111000000",
  44467=>"110000011",
  44468=>"000000000",
  44469=>"110000000",
  44470=>"000000000",
  44471=>"110100000",
  44472=>"000000111",
  44473=>"000011111",
  44474=>"001100000",
  44475=>"111111111",
  44476=>"100100000",
  44477=>"001100010",
  44478=>"000000100",
  44479=>"000010000",
  44480=>"000000000",
  44481=>"111111000",
  44482=>"001000000",
  44483=>"000000000",
  44484=>"000000100",
  44485=>"000000001",
  44486=>"000001111",
  44487=>"100110000",
  44488=>"000100000",
  44489=>"111111001",
  44490=>"000000000",
  44491=>"000000000",
  44492=>"000101111",
  44493=>"001001011",
  44494=>"111001111",
  44495=>"000000011",
  44496=>"111000110",
  44497=>"000000101",
  44498=>"101001001",
  44499=>"000000000",
  44500=>"011011011",
  44501=>"000000101",
  44502=>"011011111",
  44503=>"111111001",
  44504=>"001111000",
  44505=>"011000000",
  44506=>"000000000",
  44507=>"110000000",
  44508=>"001000000",
  44509=>"001101111",
  44510=>"100100110",
  44511=>"000011011",
  44512=>"111100000",
  44513=>"000000111",
  44514=>"001111111",
  44515=>"000000000",
  44516=>"100000111",
  44517=>"011001000",
  44518=>"000110110",
  44519=>"111011111",
  44520=>"000000011",
  44521=>"000000000",
  44522=>"100100000",
  44523=>"111111100",
  44524=>"110011011",
  44525=>"000000000",
  44526=>"110000000",
  44527=>"010110111",
  44528=>"111111010",
  44529=>"110111101",
  44530=>"000000000",
  44531=>"000110111",
  44532=>"001000000",
  44533=>"111111000",
  44534=>"010000000",
  44535=>"111111010",
  44536=>"111111000",
  44537=>"110000000",
  44538=>"010000000",
  44539=>"111111111",
  44540=>"111111111",
  44541=>"000100111",
  44542=>"001111101",
  44543=>"000000000",
  44544=>"111111001",
  44545=>"111011000",
  44546=>"111000000",
  44547=>"111111110",
  44548=>"000000101",
  44549=>"001001000",
  44550=>"000000000",
  44551=>"111111111",
  44552=>"001011001",
  44553=>"000100111",
  44554=>"001000000",
  44555=>"111111111",
  44556=>"001011111",
  44557=>"000000111",
  44558=>"100110000",
  44559=>"111111111",
  44560=>"100110000",
  44561=>"000101101",
  44562=>"111111111",
  44563=>"000000000",
  44564=>"000000111",
  44565=>"000000001",
  44566=>"111110100",
  44567=>"100111111",
  44568=>"110111000",
  44569=>"011011111",
  44570=>"111110100",
  44571=>"111111111",
  44572=>"111000110",
  44573=>"111100100",
  44574=>"011111110",
  44575=>"100101101",
  44576=>"001000111",
  44577=>"000000000",
  44578=>"011111111",
  44579=>"100100100",
  44580=>"000000010",
  44581=>"100101111",
  44582=>"011010110",
  44583=>"000010111",
  44584=>"111100110",
  44585=>"011111010",
  44586=>"000000111",
  44587=>"100000100",
  44588=>"011011001",
  44589=>"110111111",
  44590=>"000000000",
  44591=>"111111100",
  44592=>"000000101",
  44593=>"000000000",
  44594=>"000111001",
  44595=>"111111111",
  44596=>"000011111",
  44597=>"111111011",
  44598=>"001111111",
  44599=>"000010001",
  44600=>"000000010",
  44601=>"100111111",
  44602=>"111111111",
  44603=>"001000000",
  44604=>"110000101",
  44605=>"000100111",
  44606=>"111111111",
  44607=>"110000000",
  44608=>"100100111",
  44609=>"000010000",
  44610=>"000010010",
  44611=>"100110111",
  44612=>"110111110",
  44613=>"011110110",
  44614=>"000000000",
  44615=>"011000011",
  44616=>"000000011",
  44617=>"111001111",
  44618=>"111111111",
  44619=>"100011001",
  44620=>"100000100",
  44621=>"110100111",
  44622=>"111001000",
  44623=>"100100111",
  44624=>"100111100",
  44625=>"001000001",
  44626=>"000000000",
  44627=>"001001011",
  44628=>"101101111",
  44629=>"000000000",
  44630=>"100111110",
  44631=>"000000110",
  44632=>"000010010",
  44633=>"000000000",
  44634=>"111111000",
  44635=>"000101001",
  44636=>"000111000",
  44637=>"000000111",
  44638=>"101111000",
  44639=>"111111100",
  44640=>"100000000",
  44641=>"001000011",
  44642=>"011011111",
  44643=>"000000000",
  44644=>"000000000",
  44645=>"101000001",
  44646=>"101111011",
  44647=>"000000100",
  44648=>"111001111",
  44649=>"000000001",
  44650=>"000000111",
  44651=>"000111111",
  44652=>"011011010",
  44653=>"000000100",
  44654=>"000000000",
  44655=>"000010001",
  44656=>"001001001",
  44657=>"111110110",
  44658=>"001010111",
  44659=>"000000000",
  44660=>"111111111",
  44661=>"000101111",
  44662=>"000000111",
  44663=>"000000000",
  44664=>"111111111",
  44665=>"111000000",
  44666=>"000101101",
  44667=>"110000000",
  44668=>"010010010",
  44669=>"000000000",
  44670=>"000000000",
  44671=>"001000111",
  44672=>"000000100",
  44673=>"000000111",
  44674=>"001000000",
  44675=>"100111111",
  44676=>"101100000",
  44677=>"111111111",
  44678=>"000100110",
  44679=>"001111111",
  44680=>"111000000",
  44681=>"111111010",
  44682=>"000111111",
  44683=>"111111111",
  44684=>"111111101",
  44685=>"111101000",
  44686=>"111000010",
  44687=>"000000001",
  44688=>"000000111",
  44689=>"010100111",
  44690=>"111111001",
  44691=>"000011011",
  44692=>"100100000",
  44693=>"111111111",
  44694=>"000000000",
  44695=>"000000000",
  44696=>"000000000",
  44697=>"111110111",
  44698=>"111111111",
  44699=>"111111000",
  44700=>"110110110",
  44701=>"111001001",
  44702=>"100100110",
  44703=>"000000000",
  44704=>"111111111",
  44705=>"111011011",
  44706=>"000000000",
  44707=>"000011000",
  44708=>"001001001",
  44709=>"111111000",
  44710=>"111011000",
  44711=>"011101001",
  44712=>"000000001",
  44713=>"000000011",
  44714=>"111111111",
  44715=>"111110110",
  44716=>"110111111",
  44717=>"111011000",
  44718=>"111100111",
  44719=>"111010001",
  44720=>"111000000",
  44721=>"110111111",
  44722=>"011111001",
  44723=>"111000000",
  44724=>"010010000",
  44725=>"100111110",
  44726=>"111100100",
  44727=>"110110111",
  44728=>"011010111",
  44729=>"111111110",
  44730=>"110100111",
  44731=>"000001001",
  44732=>"111111110",
  44733=>"111111010",
  44734=>"010000010",
  44735=>"000000000",
  44736=>"000000011",
  44737=>"111111110",
  44738=>"000000000",
  44739=>"010111111",
  44740=>"011011111",
  44741=>"000000101",
  44742=>"101111001",
  44743=>"111111000",
  44744=>"011111111",
  44745=>"000000111",
  44746=>"111111110",
  44747=>"110000000",
  44748=>"011000000",
  44749=>"011011001",
  44750=>"000000000",
  44751=>"111101100",
  44752=>"111011001",
  44753=>"111110000",
  44754=>"111001001",
  44755=>"000000111",
  44756=>"111111001",
  44757=>"100000111",
  44758=>"000000000",
  44759=>"111110110",
  44760=>"111111001",
  44761=>"100100000",
  44762=>"000000000",
  44763=>"101100000",
  44764=>"000000000",
  44765=>"111111111",
  44766=>"001000101",
  44767=>"000101111",
  44768=>"011011001",
  44769=>"000000000",
  44770=>"100000001",
  44771=>"100111111",
  44772=>"000000000",
  44773=>"110110110",
  44774=>"111111000",
  44775=>"000000111",
  44776=>"111111110",
  44777=>"001011111",
  44778=>"000100111",
  44779=>"111111011",
  44780=>"001000000",
  44781=>"001000000",
  44782=>"111111111",
  44783=>"000000000",
  44784=>"100001111",
  44785=>"111111011",
  44786=>"110010011",
  44787=>"001001111",
  44788=>"000100000",
  44789=>"011111111",
  44790=>"001000000",
  44791=>"010010001",
  44792=>"000111111",
  44793=>"110111100",
  44794=>"000000010",
  44795=>"000000011",
  44796=>"110111110",
  44797=>"000000000",
  44798=>"000001101",
  44799=>"000000111",
  44800=>"001111111",
  44801=>"101111111",
  44802=>"000000100",
  44803=>"111111111",
  44804=>"000100111",
  44805=>"011111111",
  44806=>"000000010",
  44807=>"101111000",
  44808=>"000000001",
  44809=>"000000010",
  44810=>"000000000",
  44811=>"111111111",
  44812=>"000001001",
  44813=>"111111001",
  44814=>"000000111",
  44815=>"111110110",
  44816=>"000000001",
  44817=>"011011111",
  44818=>"000000111",
  44819=>"000001000",
  44820=>"011011011",
  44821=>"101001000",
  44822=>"101100100",
  44823=>"100101101",
  44824=>"000100111",
  44825=>"111011000",
  44826=>"011111010",
  44827=>"111111011",
  44828=>"100000111",
  44829=>"111111011",
  44830=>"111111111",
  44831=>"000000011",
  44832=>"000000001",
  44833=>"011000001",
  44834=>"111111111",
  44835=>"000000111",
  44836=>"011111000",
  44837=>"011011111",
  44838=>"111111111",
  44839=>"011111000",
  44840=>"111000000",
  44841=>"000111111",
  44842=>"101000011",
  44843=>"000000000",
  44844=>"000000011",
  44845=>"101101100",
  44846=>"111000000",
  44847=>"100100100",
  44848=>"011111111",
  44849=>"000000000",
  44850=>"000000001",
  44851=>"111111111",
  44852=>"001000000",
  44853=>"000100000",
  44854=>"000101111",
  44855=>"000011111",
  44856=>"100110000",
  44857=>"000000000",
  44858=>"000000000",
  44859=>"100010111",
  44860=>"000100000",
  44861=>"111111011",
  44862=>"100000000",
  44863=>"110111111",
  44864=>"111111001",
  44865=>"100000000",
  44866=>"101111111",
  44867=>"000000000",
  44868=>"111101001",
  44869=>"000111111",
  44870=>"011000111",
  44871=>"111111111",
  44872=>"001001111",
  44873=>"100000000",
  44874=>"111010000",
  44875=>"000000001",
  44876=>"111001000",
  44877=>"010000111",
  44878=>"001000100",
  44879=>"000000111",
  44880=>"001111100",
  44881=>"111110000",
  44882=>"000001111",
  44883=>"101001000",
  44884=>"000101111",
  44885=>"011011001",
  44886=>"000000001",
  44887=>"000000011",
  44888=>"110000000",
  44889=>"011011111",
  44890=>"111111000",
  44891=>"101101101",
  44892=>"111000110",
  44893=>"011111111",
  44894=>"001000011",
  44895=>"110111111",
  44896=>"100000110",
  44897=>"111110000",
  44898=>"110110110",
  44899=>"000000111",
  44900=>"011011111",
  44901=>"001000101",
  44902=>"000000000",
  44903=>"101001001",
  44904=>"011100100",
  44905=>"000000000",
  44906=>"000000001",
  44907=>"100111111",
  44908=>"011001000",
  44909=>"000000111",
  44910=>"000000000",
  44911=>"111100000",
  44912=>"111011001",
  44913=>"111111111",
  44914=>"001111100",
  44915=>"111111111",
  44916=>"000000000",
  44917=>"000000000",
  44918=>"111111000",
  44919=>"001001111",
  44920=>"111000100",
  44921=>"000000100",
  44922=>"000000001",
  44923=>"111111101",
  44924=>"111111111",
  44925=>"000000000",
  44926=>"000000000",
  44927=>"000000100",
  44928=>"110111110",
  44929=>"000000001",
  44930=>"100111111",
  44931=>"000000110",
  44932=>"010111110",
  44933=>"111100000",
  44934=>"100101111",
  44935=>"101000000",
  44936=>"000000000",
  44937=>"111100000",
  44938=>"111001000",
  44939=>"011000000",
  44940=>"001000111",
  44941=>"000100100",
  44942=>"011010111",
  44943=>"011011111",
  44944=>"110111000",
  44945=>"100100000",
  44946=>"111111111",
  44947=>"000001000",
  44948=>"000000000",
  44949=>"010001000",
  44950=>"000000000",
  44951=>"101001001",
  44952=>"000001001",
  44953=>"110001000",
  44954=>"100111111",
  44955=>"000000001",
  44956=>"001011000",
  44957=>"000000100",
  44958=>"111111101",
  44959=>"001011111",
  44960=>"000000000",
  44961=>"111111111",
  44962=>"100100110",
  44963=>"000111011",
  44964=>"111110111",
  44965=>"011001000",
  44966=>"011000000",
  44967=>"111111111",
  44968=>"101000000",
  44969=>"111100111",
  44970=>"000000010",
  44971=>"111100000",
  44972=>"000111000",
  44973=>"100000000",
  44974=>"000111111",
  44975=>"111111110",
  44976=>"101101000",
  44977=>"000000000",
  44978=>"000111011",
  44979=>"000110111",
  44980=>"000010111",
  44981=>"001001111",
  44982=>"000000000",
  44983=>"110111111",
  44984=>"111011000",
  44985=>"111101011",
  44986=>"000100110",
  44987=>"111110110",
  44988=>"101001100",
  44989=>"110010100",
  44990=>"000000000",
  44991=>"100100111",
  44992=>"100111000",
  44993=>"111011111",
  44994=>"000000000",
  44995=>"101000000",
  44996=>"101010011",
  44997=>"010100100",
  44998=>"100000000",
  44999=>"001011000",
  45000=>"110111101",
  45001=>"111111001",
  45002=>"000011111",
  45003=>"111111111",
  45004=>"111000000",
  45005=>"000000001",
  45006=>"011000011",
  45007=>"000000000",
  45008=>"000000000",
  45009=>"111111011",
  45010=>"010011000",
  45011=>"100111111",
  45012=>"111011111",
  45013=>"111111111",
  45014=>"111111111",
  45015=>"100111111",
  45016=>"100111011",
  45017=>"111111111",
  45018=>"111010000",
  45019=>"000001001",
  45020=>"011111111",
  45021=>"101001011",
  45022=>"100000111",
  45023=>"111111111",
  45024=>"001111101",
  45025=>"000111111",
  45026=>"111111111",
  45027=>"111111011",
  45028=>"111011000",
  45029=>"000000100",
  45030=>"010000000",
  45031=>"011111111",
  45032=>"111000000",
  45033=>"000000110",
  45034=>"111111000",
  45035=>"001000100",
  45036=>"010001000",
  45037=>"101111111",
  45038=>"111111111",
  45039=>"100011110",
  45040=>"000100110",
  45041=>"111111101",
  45042=>"110010111",
  45043=>"000000000",
  45044=>"100000000",
  45045=>"000000000",
  45046=>"010010100",
  45047=>"111001000",
  45048=>"000110111",
  45049=>"011001010",
  45050=>"000000111",
  45051=>"111011001",
  45052=>"111110111",
  45053=>"001001001",
  45054=>"111111000",
  45055=>"111111000",
  45056=>"100001011",
  45057=>"111000000",
  45058=>"101000000",
  45059=>"111100101",
  45060=>"000000111",
  45061=>"110000011",
  45062=>"100000000",
  45063=>"000111111",
  45064=>"001011001",
  45065=>"111111100",
  45066=>"010011011",
  45067=>"111111101",
  45068=>"000000010",
  45069=>"000100111",
  45070=>"110111101",
  45071=>"100100110",
  45072=>"000000000",
  45073=>"000000010",
  45074=>"000000000",
  45075=>"000000000",
  45076=>"111111001",
  45077=>"100100000",
  45078=>"001001100",
  45079=>"000101111",
  45080=>"111111111",
  45081=>"001000000",
  45082=>"000000110",
  45083=>"000000111",
  45084=>"111111110",
  45085=>"111111111",
  45086=>"000000111",
  45087=>"010000000",
  45088=>"111111111",
  45089=>"100110111",
  45090=>"000001111",
  45091=>"000111111",
  45092=>"000000111",
  45093=>"000000101",
  45094=>"000000000",
  45095=>"101000101",
  45096=>"111111111",
  45097=>"011001101",
  45098=>"011111111",
  45099=>"001000000",
  45100=>"000001000",
  45101=>"111111000",
  45102=>"111010000",
  45103=>"000000000",
  45104=>"000110010",
  45105=>"111111111",
  45106=>"000000101",
  45107=>"000000000",
  45108=>"110110110",
  45109=>"000001001",
  45110=>"000110100",
  45111=>"001111111",
  45112=>"111111001",
  45113=>"011000110",
  45114=>"111100000",
  45115=>"010111111",
  45116=>"000000111",
  45117=>"010110100",
  45118=>"111000000",
  45119=>"111111000",
  45120=>"001001101",
  45121=>"011000000",
  45122=>"000000001",
  45123=>"001100100",
  45124=>"000001111",
  45125=>"000000110",
  45126=>"000111111",
  45127=>"000000000",
  45128=>"100111101",
  45129=>"000111110",
  45130=>"000111111",
  45131=>"111111001",
  45132=>"011011111",
  45133=>"111110111",
  45134=>"000000000",
  45135=>"111111111",
  45136=>"110110000",
  45137=>"010010110",
  45138=>"111111111",
  45139=>"111111110",
  45140=>"000101000",
  45141=>"110111111",
  45142=>"000000000",
  45143=>"000000000",
  45144=>"111110110",
  45145=>"111101111",
  45146=>"011111111",
  45147=>"000000110",
  45148=>"111111011",
  45149=>"000000000",
  45150=>"001000000",
  45151=>"111111110",
  45152=>"010000000",
  45153=>"000000000",
  45154=>"001001000",
  45155=>"111110110",
  45156=>"000001101",
  45157=>"111100000",
  45158=>"000001110",
  45159=>"011001000",
  45160=>"000001000",
  45161=>"111111111",
  45162=>"001011000",
  45163=>"111001001",
  45164=>"000000000",
  45165=>"000000000",
  45166=>"000000000",
  45167=>"000000000",
  45168=>"000000011",
  45169=>"111111000",
  45170=>"010000000",
  45171=>"000000111",
  45172=>"100111111",
  45173=>"000010000",
  45174=>"000000000",
  45175=>"110111000",
  45176=>"111110010",
  45177=>"000110111",
  45178=>"111111011",
  45179=>"111111000",
  45180=>"111111100",
  45181=>"000000100",
  45182=>"001001001",
  45183=>"000000111",
  45184=>"000000111",
  45185=>"111111111",
  45186=>"000000000",
  45187=>"000000011",
  45188=>"000000000",
  45189=>"111111100",
  45190=>"100000000",
  45191=>"111111111",
  45192=>"000000000",
  45193=>"111111111",
  45194=>"111000000",
  45195=>"001000000",
  45196=>"011111111",
  45197=>"000111111",
  45198=>"111101000",
  45199=>"000000000",
  45200=>"110111110",
  45201=>"111010000",
  45202=>"000000000",
  45203=>"111111110",
  45204=>"011010110",
  45205=>"001001111",
  45206=>"111101101",
  45207=>"111001000",
  45208=>"111111000",
  45209=>"000000111",
  45210=>"111111000",
  45211=>"111110111",
  45212=>"001000100",
  45213=>"111111111",
  45214=>"000101111",
  45215=>"010111110",
  45216=>"000000000",
  45217=>"111010000",
  45218=>"000000111",
  45219=>"111111100",
  45220=>"101001011",
  45221=>"000000100",
  45222=>"000000011",
  45223=>"001111011",
  45224=>"000101111",
  45225=>"110000001",
  45226=>"111001011",
  45227=>"010010111",
  45228=>"000111111",
  45229=>"000000100",
  45230=>"111111000",
  45231=>"111111111",
  45232=>"000000000",
  45233=>"100111110",
  45234=>"010010111",
  45235=>"111000000",
  45236=>"111000000",
  45237=>"000000100",
  45238=>"111111111",
  45239=>"111111000",
  45240=>"000000000",
  45241=>"111111110",
  45242=>"111111111",
  45243=>"001111111",
  45244=>"111111111",
  45245=>"111111111",
  45246=>"110111111",
  45247=>"100111111",
  45248=>"111000111",
  45249=>"000111111",
  45250=>"000000100",
  45251=>"000000111",
  45252=>"111111110",
  45253=>"101101101",
  45254=>"111111001",
  45255=>"000100000",
  45256=>"001001111",
  45257=>"000001111",
  45258=>"011001011",
  45259=>"111110100",
  45260=>"111111111",
  45261=>"100100000",
  45262=>"000110110",
  45263=>"000000000",
  45264=>"111000000",
  45265=>"000000000",
  45266=>"101111111",
  45267=>"000100000",
  45268=>"000000000",
  45269=>"000011010",
  45270=>"010000000",
  45271=>"111111110",
  45272=>"000001111",
  45273=>"000101111",
  45274=>"000100100",
  45275=>"000000111",
  45276=>"111001111",
  45277=>"111111111",
  45278=>"111101111",
  45279=>"000001101",
  45280=>"111011000",
  45281=>"111111000",
  45282=>"000000000",
  45283=>"111111001",
  45284=>"000000111",
  45285=>"100111111",
  45286=>"011000111",
  45287=>"111111111",
  45288=>"101111000",
  45289=>"111111011",
  45290=>"000100110",
  45291=>"100000111",
  45292=>"111000000",
  45293=>"000000000",
  45294=>"000010011",
  45295=>"111111111",
  45296=>"100111001",
  45297=>"000000001",
  45298=>"001000000",
  45299=>"111111000",
  45300=>"101001001",
  45301=>"001011111",
  45302=>"000000000",
  45303=>"111111000",
  45304=>"101111000",
  45305=>"001000000",
  45306=>"001001011",
  45307=>"011111000",
  45308=>"000000101",
  45309=>"011001100",
  45310=>"000000000",
  45311=>"101001001",
  45312=>"101111101",
  45313=>"000001111",
  45314=>"111111000",
  45315=>"111111000",
  45316=>"111111111",
  45317=>"111010000",
  45318=>"101000000",
  45319=>"111111111",
  45320=>"000100111",
  45321=>"111100000",
  45322=>"001001100",
  45323=>"001001111",
  45324=>"110100100",
  45325=>"111111000",
  45326=>"100101111",
  45327=>"000111111",
  45328=>"000000001",
  45329=>"000100100",
  45330=>"111111000",
  45331=>"111001111",
  45332=>"001000000",
  45333=>"001001111",
  45334=>"000000100",
  45335=>"101100000",
  45336=>"111111000",
  45337=>"111000000",
  45338=>"000000111",
  45339=>"111100101",
  45340=>"000000111",
  45341=>"111110101",
  45342=>"011111111",
  45343=>"011000111",
  45344=>"111111000",
  45345=>"111111111",
  45346=>"111111000",
  45347=>"011001001",
  45348=>"000000100",
  45349=>"000010010",
  45350=>"100100101",
  45351=>"111111001",
  45352=>"000000000",
  45353=>"111111000",
  45354=>"111101111",
  45355=>"111111011",
  45356=>"000011111",
  45357=>"110110100",
  45358=>"111111111",
  45359=>"111101100",
  45360=>"001001111",
  45361=>"011101001",
  45362=>"000000000",
  45363=>"000000000",
  45364=>"111111000",
  45365=>"100111000",
  45366=>"001001001",
  45367=>"111110110",
  45368=>"111111000",
  45369=>"111111111",
  45370=>"011011001",
  45371=>"001001000",
  45372=>"000000000",
  45373=>"100110110",
  45374=>"001000000",
  45375=>"000000111",
  45376=>"111111100",
  45377=>"011111111",
  45378=>"110111111",
  45379=>"111111111",
  45380=>"100000100",
  45381=>"011111111",
  45382=>"101111111",
  45383=>"000000000",
  45384=>"000000000",
  45385=>"111111000",
  45386=>"000001111",
  45387=>"111001101",
  45388=>"000000100",
  45389=>"000001001",
  45390=>"001100111",
  45391=>"001000001",
  45392=>"000000101",
  45393=>"001000001",
  45394=>"111111111",
  45395=>"111111111",
  45396=>"111111111",
  45397=>"011011001",
  45398=>"110000000",
  45399=>"111111111",
  45400=>"000000000",
  45401=>"111110111",
  45402=>"111111111",
  45403=>"101111111",
  45404=>"110110000",
  45405=>"111111111",
  45406=>"111111110",
  45407=>"100000001",
  45408=>"000000000",
  45409=>"000000100",
  45410=>"111111111",
  45411=>"000111111",
  45412=>"000000001",
  45413=>"111101000",
  45414=>"111111111",
  45415=>"011111000",
  45416=>"000000100",
  45417=>"111111110",
  45418=>"100000111",
  45419=>"000000011",
  45420=>"000000000",
  45421=>"111111011",
  45422=>"110111111",
  45423=>"000000101",
  45424=>"110001001",
  45425=>"111111000",
  45426=>"111111011",
  45427=>"100000110",
  45428=>"011011001",
  45429=>"111111111",
  45430=>"000000000",
  45431=>"111000000",
  45432=>"111111111",
  45433=>"111001100",
  45434=>"000000001",
  45435=>"001000111",
  45436=>"000011011",
  45437=>"111000001",
  45438=>"000111111",
  45439=>"111000000",
  45440=>"000110111",
  45441=>"101111111",
  45442=>"000110111",
  45443=>"000000111",
  45444=>"111111001",
  45445=>"010110000",
  45446=>"000001111",
  45447=>"110111111",
  45448=>"000000000",
  45449=>"100000100",
  45450=>"001000000",
  45451=>"111111000",
  45452=>"111101111",
  45453=>"000110110",
  45454=>"000111111",
  45455=>"001010100",
  45456=>"000111111",
  45457=>"001001111",
  45458=>"111000000",
  45459=>"001000001",
  45460=>"111111100",
  45461=>"000010000",
  45462=>"111111011",
  45463=>"000100000",
  45464=>"100100000",
  45465=>"111011000",
  45466=>"111000000",
  45467=>"101000000",
  45468=>"111111111",
  45469=>"100000101",
  45470=>"000110101",
  45471=>"000000000",
  45472=>"001001001",
  45473=>"111011000",
  45474=>"001001011",
  45475=>"011000000",
  45476=>"111111111",
  45477=>"101111101",
  45478=>"000000000",
  45479=>"000011110",
  45480=>"110110000",
  45481=>"000000000",
  45482=>"011111001",
  45483=>"000000111",
  45484=>"011000000",
  45485=>"011000000",
  45486=>"001011111",
  45487=>"011100111",
  45488=>"111100110",
  45489=>"001111111",
  45490=>"111000000",
  45491=>"000000001",
  45492=>"110110000",
  45493=>"000001111",
  45494=>"001111111",
  45495=>"000000000",
  45496=>"001000000",
  45497=>"000000000",
  45498=>"011111110",
  45499=>"100000000",
  45500=>"010000100",
  45501=>"000100111",
  45502=>"000001000",
  45503=>"000010110",
  45504=>"010000000",
  45505=>"000111111",
  45506=>"000000111",
  45507=>"111110000",
  45508=>"000000011",
  45509=>"111111100",
  45510=>"010000000",
  45511=>"011011001",
  45512=>"000111101",
  45513=>"111111111",
  45514=>"000000001",
  45515=>"110110111",
  45516=>"000110111",
  45517=>"001110111",
  45518=>"000001011",
  45519=>"000000000",
  45520=>"000000000",
  45521=>"100111110",
  45522=>"010011111",
  45523=>"011111111",
  45524=>"011011000",
  45525=>"000111111",
  45526=>"000000111",
  45527=>"000000100",
  45528=>"000000000",
  45529=>"111111111",
  45530=>"111111111",
  45531=>"111111001",
  45532=>"111111001",
  45533=>"111101111",
  45534=>"101100111",
  45535=>"000011010",
  45536=>"000000111",
  45537=>"000000000",
  45538=>"100100000",
  45539=>"000000100",
  45540=>"000000011",
  45541=>"000001100",
  45542=>"111000000",
  45543=>"000000000",
  45544=>"101101100",
  45545=>"000100111",
  45546=>"111111111",
  45547=>"000000101",
  45548=>"111111111",
  45549=>"000000001",
  45550=>"111110111",
  45551=>"111111101",
  45552=>"100100111",
  45553=>"000000000",
  45554=>"111100111",
  45555=>"100000000",
  45556=>"000001011",
  45557=>"000111111",
  45558=>"000000000",
  45559=>"100100000",
  45560=>"000100000",
  45561=>"000100111",
  45562=>"011000000",
  45563=>"000000110",
  45564=>"011000000",
  45565=>"000110110",
  45566=>"000000110",
  45567=>"111111101",
  45568=>"000000000",
  45569=>"001001011",
  45570=>"000000111",
  45571=>"001000000",
  45572=>"111111111",
  45573=>"100000000",
  45574=>"010110110",
  45575=>"000000000",
  45576=>"000001000",
  45577=>"000000111",
  45578=>"111111000",
  45579=>"000000000",
  45580=>"111111011",
  45581=>"110000111",
  45582=>"111011111",
  45583=>"110100000",
  45584=>"000000000",
  45585=>"111111111",
  45586=>"000000000",
  45587=>"111111111",
  45588=>"000000000",
  45589=>"010111111",
  45590=>"000000000",
  45591=>"000001100",
  45592=>"111111000",
  45593=>"000111111",
  45594=>"111111001",
  45595=>"111111011",
  45596=>"001101001",
  45597=>"100100100",
  45598=>"011111111",
  45599=>"100100000",
  45600=>"101101001",
  45601=>"010000000",
  45602=>"110101111",
  45603=>"111111111",
  45604=>"001000001",
  45605=>"001001000",
  45606=>"111100000",
  45607=>"000000000",
  45608=>"000000000",
  45609=>"101000000",
  45610=>"000000000",
  45611=>"101000000",
  45612=>"110001000",
  45613=>"111111011",
  45614=>"000101101",
  45615=>"110000000",
  45616=>"011000000",
  45617=>"110111111",
  45618=>"100101111",
  45619=>"000000000",
  45620=>"100100110",
  45621=>"100101111",
  45622=>"000100000",
  45623=>"001000111",
  45624=>"011111111",
  45625=>"000000101",
  45626=>"000000000",
  45627=>"011111111",
  45628=>"110000111",
  45629=>"110010110",
  45630=>"000000000",
  45631=>"000010110",
  45632=>"000000100",
  45633=>"111000000",
  45634=>"001011110",
  45635=>"011010000",
  45636=>"000111111",
  45637=>"001000000",
  45638=>"000101111",
  45639=>"111111111",
  45640=>"111110100",
  45641=>"000000000",
  45642=>"000000000",
  45643=>"101101110",
  45644=>"111111100",
  45645=>"000001011",
  45646=>"001011111",
  45647=>"111111111",
  45648=>"001011011",
  45649=>"111111111",
  45650=>"000000010",
  45651=>"000101111",
  45652=>"110110000",
  45653=>"000000000",
  45654=>"000100000",
  45655=>"000000000",
  45656=>"111111111",
  45657=>"111101100",
  45658=>"000000000",
  45659=>"001000000",
  45660=>"000000011",
  45661=>"000000000",
  45662=>"000111111",
  45663=>"100000100",
  45664=>"110111011",
  45665=>"110111111",
  45666=>"000000000",
  45667=>"111111000",
  45668=>"011011001",
  45669=>"001101101",
  45670=>"111111111",
  45671=>"111101000",
  45672=>"000000111",
  45673=>"010111111",
  45674=>"000100111",
  45675=>"000110001",
  45676=>"000001001",
  45677=>"000000000",
  45678=>"111111111",
  45679=>"000000000",
  45680=>"100111111",
  45681=>"101000000",
  45682=>"000000110",
  45683=>"110111100",
  45684=>"000000100",
  45685=>"000110111",
  45686=>"111111111",
  45687=>"111111110",
  45688=>"100000000",
  45689=>"000100000",
  45690=>"000001101",
  45691=>"000000000",
  45692=>"000000001",
  45693=>"011000011",
  45694=>"000000000",
  45695=>"000000000",
  45696=>"111111111",
  45697=>"100110101",
  45698=>"000000000",
  45699=>"111100000",
  45700=>"001000000",
  45701=>"111111111",
  45702=>"000000000",
  45703=>"111111111",
  45704=>"000100111",
  45705=>"001000000",
  45706=>"111010000",
  45707=>"000000000",
  45708=>"000000000",
  45709=>"000110111",
  45710=>"100100111",
  45711=>"000000010",
  45712=>"111111111",
  45713=>"000000000",
  45714=>"111111111",
  45715=>"000000010",
  45716=>"100100100",
  45717=>"000111111",
  45718=>"000000001",
  45719=>"111111111",
  45720=>"011000111",
  45721=>"000111111",
  45722=>"111110111",
  45723=>"000000000",
  45724=>"100000001",
  45725=>"000101111",
  45726=>"000000001",
  45727=>"111111100",
  45728=>"000110111",
  45729=>"000000000",
  45730=>"000000000",
  45731=>"010000011",
  45732=>"111111111",
  45733=>"110110111",
  45734=>"000000111",
  45735=>"000110110",
  45736=>"000011111",
  45737=>"000001000",
  45738=>"000000000",
  45739=>"000100111",
  45740=>"110111111",
  45741=>"000110100",
  45742=>"111111000",
  45743=>"100000011",
  45744=>"101000000",
  45745=>"111011000",
  45746=>"111111110",
  45747=>"010000001",
  45748=>"111010000",
  45749=>"100000000",
  45750=>"100110110",
  45751=>"111111111",
  45752=>"111000000",
  45753=>"111111111",
  45754=>"000000010",
  45755=>"111101001",
  45756=>"001000000",
  45757=>"011000000",
  45758=>"000000000",
  45759=>"111111101",
  45760=>"000000001",
  45761=>"111111111",
  45762=>"011101111",
  45763=>"111111011",
  45764=>"011001000",
  45765=>"101111111",
  45766=>"101100000",
  45767=>"001000000",
  45768=>"000001111",
  45769=>"000001011",
  45770=>"010011000",
  45771=>"111111001",
  45772=>"000010110",
  45773=>"000110111",
  45774=>"111011000",
  45775=>"000100111",
  45776=>"111111000",
  45777=>"111111111",
  45778=>"101101000",
  45779=>"010111111",
  45780=>"000000111",
  45781=>"111111111",
  45782=>"000000000",
  45783=>"001011000",
  45784=>"000000001",
  45785=>"000000111",
  45786=>"011000100",
  45787=>"000110111",
  45788=>"111111111",
  45789=>"111111111",
  45790=>"111100111",
  45791=>"000000000",
  45792=>"111111111",
  45793=>"011011000",
  45794=>"111111111",
  45795=>"110000011",
  45796=>"000000000",
  45797=>"000001001",
  45798=>"011111111",
  45799=>"000001111",
  45800=>"111111000",
  45801=>"000100111",
  45802=>"110111111",
  45803=>"111111111",
  45804=>"011111111",
  45805=>"111000000",
  45806=>"111111111",
  45807=>"000001000",
  45808=>"111001000",
  45809=>"000000000",
  45810=>"111000111",
  45811=>"101111111",
  45812=>"001001001",
  45813=>"001000001",
  45814=>"000000001",
  45815=>"011001001",
  45816=>"000000000",
  45817=>"011011000",
  45818=>"000000000",
  45819=>"111001011",
  45820=>"011000000",
  45821=>"001001001",
  45822=>"000000000",
  45823=>"000000100",
  45824=>"111110110",
  45825=>"100110110",
  45826=>"000111111",
  45827=>"111111001",
  45828=>"111111111",
  45829=>"101001000",
  45830=>"100000101",
  45831=>"101111111",
  45832=>"000000000",
  45833=>"001000000",
  45834=>"001000000",
  45835=>"011010011",
  45836=>"111111111",
  45837=>"111111111",
  45838=>"111111111",
  45839=>"111111101",
  45840=>"000000000",
  45841=>"111000100",
  45842=>"001000000",
  45843=>"000001111",
  45844=>"000000000",
  45845=>"000001000",
  45846=>"000000111",
  45847=>"000000000",
  45848=>"111111111",
  45849=>"000000000",
  45850=>"001100000",
  45851=>"000110110",
  45852=>"001111111",
  45853=>"000000000",
  45854=>"000000000",
  45855=>"111111111",
  45856=>"000101111",
  45857=>"000101111",
  45858=>"000001011",
  45859=>"101000001",
  45860=>"001000000",
  45861=>"000000000",
  45862=>"111111111",
  45863=>"000001111",
  45864=>"111111111",
  45865=>"010111111",
  45866=>"111000000",
  45867=>"100100000",
  45868=>"111111111",
  45869=>"011011111",
  45870=>"001011001",
  45871=>"011011011",
  45872=>"000000000",
  45873=>"110000011",
  45874=>"101100000",
  45875=>"111011000",
  45876=>"111011000",
  45877=>"100000000",
  45878=>"000000000",
  45879=>"000001011",
  45880=>"000000001",
  45881=>"000001111",
  45882=>"110111111",
  45883=>"111111000",
  45884=>"100110000",
  45885=>"000000000",
  45886=>"000000100",
  45887=>"000111111",
  45888=>"111111111",
  45889=>"111111101",
  45890=>"110000011",
  45891=>"000000000",
  45892=>"110010000",
  45893=>"000110111",
  45894=>"010010000",
  45895=>"111111111",
  45896=>"000000000",
  45897=>"111000000",
  45898=>"000000000",
  45899=>"010111000",
  45900=>"000001000",
  45901=>"000000000",
  45902=>"110111111",
  45903=>"001001001",
  45904=>"000001011",
  45905=>"111110111",
  45906=>"111011000",
  45907=>"111000000",
  45908=>"100000000",
  45909=>"100010010",
  45910=>"011001111",
  45911=>"100100111",
  45912=>"111111111",
  45913=>"000000000",
  45914=>"111010010",
  45915=>"111111111",
  45916=>"000000000",
  45917=>"111000111",
  45918=>"111000000",
  45919=>"000001001",
  45920=>"010000000",
  45921=>"111110111",
  45922=>"100111111",
  45923=>"000000100",
  45924=>"000000100",
  45925=>"000000000",
  45926=>"101000000",
  45927=>"000100111",
  45928=>"000101000",
  45929=>"000000001",
  45930=>"000000000",
  45931=>"110000000",
  45932=>"000000010",
  45933=>"111111111",
  45934=>"000000000",
  45935=>"000011011",
  45936=>"000000100",
  45937=>"000101001",
  45938=>"001001001",
  45939=>"011001011",
  45940=>"000001000",
  45941=>"111111000",
  45942=>"111111111",
  45943=>"000111000",
  45944=>"000000110",
  45945=>"101011011",
  45946=>"000000000",
  45947=>"011111111",
  45948=>"000000001",
  45949=>"101111111",
  45950=>"000000000",
  45951=>"000000000",
  45952=>"001000111",
  45953=>"111111111",
  45954=>"000000000",
  45955=>"000000000",
  45956=>"000100000",
  45957=>"000000111",
  45958=>"000111110",
  45959=>"011000000",
  45960=>"111111010",
  45961=>"000100110",
  45962=>"000000000",
  45963=>"001001001",
  45964=>"111111111",
  45965=>"101111110",
  45966=>"101000000",
  45967=>"000001011",
  45968=>"000000000",
  45969=>"100000000",
  45970=>"001001001",
  45971=>"111011010",
  45972=>"110100111",
  45973=>"110000000",
  45974=>"000000000",
  45975=>"000000000",
  45976=>"111111111",
  45977=>"011011111",
  45978=>"000000111",
  45979=>"000000000",
  45980=>"000111111",
  45981=>"000000000",
  45982=>"111101000",
  45983=>"000000100",
  45984=>"000000000",
  45985=>"100100100",
  45986=>"000000000",
  45987=>"000000000",
  45988=>"111110011",
  45989=>"111010000",
  45990=>"111110000",
  45991=>"000000000",
  45992=>"000000000",
  45993=>"111011000",
  45994=>"100000001",
  45995=>"000000110",
  45996=>"010111010",
  45997=>"000110011",
  45998=>"000001001",
  45999=>"111110111",
  46000=>"011101000",
  46001=>"101101101",
  46002=>"000001111",
  46003=>"101001000",
  46004=>"111111111",
  46005=>"111111111",
  46006=>"111111111",
  46007=>"001000000",
  46008=>"000000011",
  46009=>"111111101",
  46010=>"000000000",
  46011=>"111111111",
  46012=>"000111111",
  46013=>"111111111",
  46014=>"101101111",
  46015=>"111100111",
  46016=>"000110111",
  46017=>"111111111",
  46018=>"111111111",
  46019=>"100111111",
  46020=>"111111011",
  46021=>"100111111",
  46022=>"101000000",
  46023=>"111001001",
  46024=>"101000111",
  46025=>"011111100",
  46026=>"000000000",
  46027=>"111111100",
  46028=>"000110111",
  46029=>"010010111",
  46030=>"100000000",
  46031=>"000000101",
  46032=>"000000001",
  46033=>"111111111",
  46034=>"110000000",
  46035=>"001111111",
  46036=>"000000000",
  46037=>"000000001",
  46038=>"111000000",
  46039=>"111010000",
  46040=>"000000000",
  46041=>"111001001",
  46042=>"001001111",
  46043=>"000000000",
  46044=>"000000000",
  46045=>"000000000",
  46046=>"100000110",
  46047=>"000111110",
  46048=>"111111111",
  46049=>"001011111",
  46050=>"111111000",
  46051=>"100000000",
  46052=>"111111111",
  46053=>"000101101",
  46054=>"110110000",
  46055=>"000010000",
  46056=>"111111111",
  46057=>"000000000",
  46058=>"101000000",
  46059=>"111111111",
  46060=>"000000001",
  46061=>"100100110",
  46062=>"111101100",
  46063=>"001001110",
  46064=>"000010011",
  46065=>"000000000",
  46066=>"111111111",
  46067=>"011111000",
  46068=>"100000111",
  46069=>"111111000",
  46070=>"111111111",
  46071=>"000000000",
  46072=>"111111101",
  46073=>"111001011",
  46074=>"000000000",
  46075=>"000000000",
  46076=>"111011000",
  46077=>"111111101",
  46078=>"000000000",
  46079=>"000000000",
  46080=>"000000000",
  46081=>"110110111",
  46082=>"111111111",
  46083=>"000000101",
  46084=>"000010000",
  46085=>"010011011",
  46086=>"111111111",
  46087=>"000000000",
  46088=>"000000000",
  46089=>"000000000",
  46090=>"000001010",
  46091=>"010111111",
  46092=>"111111111",
  46093=>"110000011",
  46094=>"100100110",
  46095=>"000000000",
  46096=>"000000000",
  46097=>"000000000",
  46098=>"111111111",
  46099=>"000000000",
  46100=>"011011100",
  46101=>"001001000",
  46102=>"111011001",
  46103=>"111110110",
  46104=>"111111111",
  46105=>"000000000",
  46106=>"000000010",
  46107=>"000000000",
  46108=>"000000101",
  46109=>"110000000",
  46110=>"011011001",
  46111=>"000000001",
  46112=>"000111111",
  46113=>"000001001",
  46114=>"110111011",
  46115=>"111111110",
  46116=>"111111111",
  46117=>"111011011",
  46118=>"111111100",
  46119=>"001001001",
  46120=>"100111111",
  46121=>"101111111",
  46122=>"010010000",
  46123=>"000000001",
  46124=>"111111111",
  46125=>"101101111",
  46126=>"100110111",
  46127=>"111111111",
  46128=>"111111111",
  46129=>"110111110",
  46130=>"000000100",
  46131=>"000100000",
  46132=>"101101101",
  46133=>"110000000",
  46134=>"110111001",
  46135=>"010010011",
  46136=>"111111111",
  46137=>"100111111",
  46138=>"111111111",
  46139=>"111011011",
  46140=>"100000000",
  46141=>"111111111",
  46142=>"111111111",
  46143=>"000000000",
  46144=>"111111111",
  46145=>"111111111",
  46146=>"111110000",
  46147=>"111111111",
  46148=>"000000010",
  46149=>"001001000",
  46150=>"111000000",
  46151=>"111111111",
  46152=>"011011010",
  46153=>"000000000",
  46154=>"111111101",
  46155=>"000000000",
  46156=>"000001100",
  46157=>"000010111",
  46158=>"000000000",
  46159=>"100111111",
  46160=>"011011001",
  46161=>"101111101",
  46162=>"000000000",
  46163=>"001001111",
  46164=>"111111111",
  46165=>"000111111",
  46166=>"000000000",
  46167=>"111111111",
  46168=>"100111111",
  46169=>"111111111",
  46170=>"111011111",
  46171=>"111111001",
  46172=>"011000000",
  46173=>"110001101",
  46174=>"010011111",
  46175=>"000000000",
  46176=>"000100111",
  46177=>"010010011",
  46178=>"111111111",
  46179=>"111101111",
  46180=>"100101100",
  46181=>"011111001",
  46182=>"000000000",
  46183=>"001000000",
  46184=>"001101101",
  46185=>"110100000",
  46186=>"100000000",
  46187=>"010010010",
  46188=>"111111000",
  46189=>"111111111",
  46190=>"111111111",
  46191=>"000000110",
  46192=>"001011011",
  46193=>"111111111",
  46194=>"100111111",
  46195=>"000000000",
  46196=>"100000000",
  46197=>"111111111",
  46198=>"111111111",
  46199=>"010000000",
  46200=>"111111111",
  46201=>"000111100",
  46202=>"111111100",
  46203=>"000000000",
  46204=>"000000001",
  46205=>"000111101",
  46206=>"111111000",
  46207=>"011011001",
  46208=>"000000000",
  46209=>"100110111",
  46210=>"111111111",
  46211=>"010110100",
  46212=>"111111001",
  46213=>"111001001",
  46214=>"000000111",
  46215=>"000000011",
  46216=>"000000000",
  46217=>"011001000",
  46218=>"100100101",
  46219=>"000001110",
  46220=>"001111101",
  46221=>"000111000",
  46222=>"111111011",
  46223=>"100100111",
  46224=>"011000000",
  46225=>"000000000",
  46226=>"000000000",
  46227=>"000000000",
  46228=>"001001000",
  46229=>"111111010",
  46230=>"000000000",
  46231=>"111100000",
  46232=>"000001111",
  46233=>"000000000",
  46234=>"110010111",
  46235=>"111111111",
  46236=>"000000000",
  46237=>"110111111",
  46238=>"000000000",
  46239=>"011111111",
  46240=>"000001001",
  46241=>"000000000",
  46242=>"111111111",
  46243=>"111011011",
  46244=>"111111011",
  46245=>"100000000",
  46246=>"000000000",
  46247=>"000100000",
  46248=>"000111000",
  46249=>"000000000",
  46250=>"000000000",
  46251=>"110111111",
  46252=>"000000000",
  46253=>"011110010",
  46254=>"100000000",
  46255=>"111100000",
  46256=>"000100111",
  46257=>"000110000",
  46258=>"111111111",
  46259=>"111000000",
  46260=>"111101100",
  46261=>"000111111",
  46262=>"000000000",
  46263=>"001111000",
  46264=>"111111111",
  46265=>"111111000",
  46266=>"000010000",
  46267=>"010000000",
  46268=>"000110010",
  46269=>"111111111",
  46270=>"111000010",
  46271=>"111111011",
  46272=>"000000000",
  46273=>"111111000",
  46274=>"110110000",
  46275=>"000001111",
  46276=>"111111111",
  46277=>"000000000",
  46278=>"110111011",
  46279=>"010111111",
  46280=>"000000000",
  46281=>"010111110",
  46282=>"011000000",
  46283=>"011001000",
  46284=>"000000000",
  46285=>"000000000",
  46286=>"000000000",
  46287=>"011111001",
  46288=>"111001000",
  46289=>"111001111",
  46290=>"111111111",
  46291=>"010000000",
  46292=>"000000000",
  46293=>"111111010",
  46294=>"111111111",
  46295=>"011000000",
  46296=>"111111111",
  46297=>"000000000",
  46298=>"111111111",
  46299=>"000000111",
  46300=>"000000000",
  46301=>"000100100",
  46302=>"000000000",
  46303=>"111111111",
  46304=>"000000110",
  46305=>"000000000",
  46306=>"111011001",
  46307=>"011001001",
  46308=>"110000000",
  46309=>"010010000",
  46310=>"111111111",
  46311=>"000000000",
  46312=>"111111111",
  46313=>"111111000",
  46314=>"111111110",
  46315=>"110000000",
  46316=>"111111111",
  46317=>"111000000",
  46318=>"000111111",
  46319=>"111111111",
  46320=>"110010011",
  46321=>"010000000",
  46322=>"000000000",
  46323=>"101111101",
  46324=>"000111111",
  46325=>"000000001",
  46326=>"111110111",
  46327=>"011000000",
  46328=>"011011011",
  46329=>"111111111",
  46330=>"000010111",
  46331=>"101110110",
  46332=>"110111111",
  46333=>"111001001",
  46334=>"000100100",
  46335=>"111111111",
  46336=>"010001111",
  46337=>"111011011",
  46338=>"111111111",
  46339=>"010110100",
  46340=>"101111111",
  46341=>"101100100",
  46342=>"111111111",
  46343=>"100101111",
  46344=>"000000000",
  46345=>"000000000",
  46346=>"111111111",
  46347=>"000000000",
  46348=>"111111111",
  46349=>"000000000",
  46350=>"000000011",
  46351=>"111111000",
  46352=>"001000000",
  46353=>"000101001",
  46354=>"110011010",
  46355=>"011110111",
  46356=>"100000000",
  46357=>"111111001",
  46358=>"000000010",
  46359=>"111111111",
  46360=>"111111111",
  46361=>"100110111",
  46362=>"111111111",
  46363=>"111111111",
  46364=>"000000000",
  46365=>"000110110",
  46366=>"111111111",
  46367=>"111111111",
  46368=>"110110111",
  46369=>"100000000",
  46370=>"110111111",
  46371=>"101101101",
  46372=>"000000000",
  46373=>"011011111",
  46374=>"001001000",
  46375=>"100101100",
  46376=>"110110111",
  46377=>"111111000",
  46378=>"111111111",
  46379=>"111111111",
  46380=>"111111111",
  46381=>"111111011",
  46382=>"000000000",
  46383=>"000000000",
  46384=>"110110111",
  46385=>"010000000",
  46386=>"000111000",
  46387=>"111111111",
  46388=>"000000000",
  46389=>"111100000",
  46390=>"100111111",
  46391=>"000011000",
  46392=>"101000000",
  46393=>"000000000",
  46394=>"010111111",
  46395=>"000000000",
  46396=>"000000100",
  46397=>"001000000",
  46398=>"000000100",
  46399=>"110111000",
  46400=>"100111110",
  46401=>"110100000",
  46402=>"000100000",
  46403=>"110000000",
  46404=>"000100000",
  46405=>"000010011",
  46406=>"000000000",
  46407=>"111111111",
  46408=>"000010011",
  46409=>"000011011",
  46410=>"000000011",
  46411=>"110110111",
  46412=>"001111011",
  46413=>"100111111",
  46414=>"110111111",
  46415=>"110111111",
  46416=>"010110100",
  46417=>"000000001",
  46418=>"000000000",
  46419=>"001001111",
  46420=>"111111111",
  46421=>"000010110",
  46422=>"111111111",
  46423=>"000111111",
  46424=>"000000000",
  46425=>"000000101",
  46426=>"100111111",
  46427=>"010000100",
  46428=>"111111111",
  46429=>"111010110",
  46430=>"011000000",
  46431=>"111000000",
  46432=>"000000000",
  46433=>"111000001",
  46434=>"100100100",
  46435=>"000000000",
  46436=>"111111111",
  46437=>"111111111",
  46438=>"111111111",
  46439=>"000000001",
  46440=>"011011111",
  46441=>"111111010",
  46442=>"010010000",
  46443=>"110110111",
  46444=>"101111000",
  46445=>"011111010",
  46446=>"111111111",
  46447=>"111111111",
  46448=>"111111111",
  46449=>"111111111",
  46450=>"011000001",
  46451=>"000010111",
  46452=>"010010101",
  46453=>"101111000",
  46454=>"010000000",
  46455=>"111111111",
  46456=>"000000000",
  46457=>"001000000",
  46458=>"111000000",
  46459=>"000010011",
  46460=>"111100111",
  46461=>"000001001",
  46462=>"101000000",
  46463=>"000000111",
  46464=>"000001011",
  46465=>"000001001",
  46466=>"000000000",
  46467=>"000110111",
  46468=>"111111111",
  46469=>"000000000",
  46470=>"000000001",
  46471=>"000111111",
  46472=>"111011000",
  46473=>"100110110",
  46474=>"111111111",
  46475=>"111111111",
  46476=>"111111111",
  46477=>"011011011",
  46478=>"000001011",
  46479=>"001000000",
  46480=>"000001111",
  46481=>"001111111",
  46482=>"111111111",
  46483=>"010010011",
  46484=>"000000000",
  46485=>"111111000",
  46486=>"110111110",
  46487=>"100000000",
  46488=>"011011111",
  46489=>"010000000",
  46490=>"111111111",
  46491=>"000100110",
  46492=>"000000000",
  46493=>"000000000",
  46494=>"111011001",
  46495=>"000000000",
  46496=>"011111111",
  46497=>"111110110",
  46498=>"111100100",
  46499=>"010111111",
  46500=>"111000000",
  46501=>"000000110",
  46502=>"111011001",
  46503=>"111111111",
  46504=>"000000000",
  46505=>"000011111",
  46506=>"000111111",
  46507=>"111111001",
  46508=>"000000000",
  46509=>"000000000",
  46510=>"011011000",
  46511=>"111111100",
  46512=>"111101111",
  46513=>"011111111",
  46514=>"111100000",
  46515=>"000111000",
  46516=>"000000001",
  46517=>"001001000",
  46518=>"111001001",
  46519=>"000100100",
  46520=>"111111111",
  46521=>"000011001",
  46522=>"111101111",
  46523=>"110000010",
  46524=>"000000000",
  46525=>"000010110",
  46526=>"100111111",
  46527=>"111111111",
  46528=>"100100100",
  46529=>"000000000",
  46530=>"111111111",
  46531=>"111111111",
  46532=>"100000011",
  46533=>"110111011",
  46534=>"001001101",
  46535=>"100100001",
  46536=>"000000111",
  46537=>"111111111",
  46538=>"111101000",
  46539=>"111111111",
  46540=>"101101111",
  46541=>"000000000",
  46542=>"000000011",
  46543=>"000000000",
  46544=>"100100111",
  46545=>"111111111",
  46546=>"111010110",
  46547=>"000000000",
  46548=>"110110110",
  46549=>"111000000",
  46550=>"111111111",
  46551=>"000000100",
  46552=>"000000100",
  46553=>"000110000",
  46554=>"110000000",
  46555=>"010011111",
  46556=>"000000000",
  46557=>"000000111",
  46558=>"101111000",
  46559=>"110000111",
  46560=>"101000000",
  46561=>"111011011",
  46562=>"000000000",
  46563=>"000000000",
  46564=>"000111111",
  46565=>"111100100",
  46566=>"001100000",
  46567=>"111111111",
  46568=>"000000001",
  46569=>"011011001",
  46570=>"110111111",
  46571=>"111111111",
  46572=>"010000011",
  46573=>"000101110",
  46574=>"111111111",
  46575=>"011000000",
  46576=>"011011000",
  46577=>"111111111",
  46578=>"011111110",
  46579=>"111111111",
  46580=>"111111111",
  46581=>"100000100",
  46582=>"111111000",
  46583=>"111010000",
  46584=>"000000000",
  46585=>"000000100",
  46586=>"111110000",
  46587=>"000000000",
  46588=>"111111111",
  46589=>"000111011",
  46590=>"010000000",
  46591=>"000000111",
  46592=>"000011011",
  46593=>"000000000",
  46594=>"111000111",
  46595=>"111111111",
  46596=>"100111111",
  46597=>"111001011",
  46598=>"000000000",
  46599=>"101000000",
  46600=>"001011111",
  46601=>"000000001",
  46602=>"000000000",
  46603=>"100000111",
  46604=>"111111111",
  46605=>"111111111",
  46606=>"010010011",
  46607=>"111111111",
  46608=>"110001001",
  46609=>"110000000",
  46610=>"000000000",
  46611=>"000000000",
  46612=>"000000000",
  46613=>"000111110",
  46614=>"000000000",
  46615=>"111111111",
  46616=>"111111111",
  46617=>"011000000",
  46618=>"100101101",
  46619=>"011111000",
  46620=>"000000000",
  46621=>"001000101",
  46622=>"111111111",
  46623=>"111111111",
  46624=>"111100111",
  46625=>"000000000",
  46626=>"000000000",
  46627=>"000001011",
  46628=>"111111001",
  46629=>"111111111",
  46630=>"111111111",
  46631=>"111111111",
  46632=>"111000000",
  46633=>"000000000",
  46634=>"000000000",
  46635=>"000000000",
  46636=>"111111111",
  46637=>"111111111",
  46638=>"101000111",
  46639=>"000000111",
  46640=>"101111111",
  46641=>"000000000",
  46642=>"111111111",
  46643=>"111111000",
  46644=>"001001000",
  46645=>"100101000",
  46646=>"000100001",
  46647=>"100100000",
  46648=>"000000000",
  46649=>"111111111",
  46650=>"000000000",
  46651=>"111111110",
  46652=>"111100000",
  46653=>"110111111",
  46654=>"011011001",
  46655=>"001000000",
  46656=>"111111111",
  46657=>"110110111",
  46658=>"111111110",
  46659=>"111111111",
  46660=>"111111111",
  46661=>"001000000",
  46662=>"001110111",
  46663=>"000000000",
  46664=>"101101111",
  46665=>"111111111",
  46666=>"011011000",
  46667=>"000000111",
  46668=>"000000000",
  46669=>"111111111",
  46670=>"111111111",
  46671=>"111101001",
  46672=>"110110000",
  46673=>"000000111",
  46674=>"000000000",
  46675=>"001000000",
  46676=>"000100001",
  46677=>"000010111",
  46678=>"110100011",
  46679=>"111101111",
  46680=>"111111110",
  46681=>"000000000",
  46682=>"000000000",
  46683=>"111111111",
  46684=>"000000000",
  46685=>"111111111",
  46686=>"000010111",
  46687=>"111111111",
  46688=>"111110010",
  46689=>"111111000",
  46690=>"011001000",
  46691=>"000000000",
  46692=>"000000001",
  46693=>"111111111",
  46694=>"001000011",
  46695=>"001001111",
  46696=>"000111111",
  46697=>"111111111",
  46698=>"111001000",
  46699=>"111111111",
  46700=>"000000000",
  46701=>"111111111",
  46702=>"111110111",
  46703=>"111111111",
  46704=>"100111111",
  46705=>"000000000",
  46706=>"111111101",
  46707=>"100100000",
  46708=>"000000000",
  46709=>"001011111",
  46710=>"000001011",
  46711=>"000000000",
  46712=>"111111010",
  46713=>"000000000",
  46714=>"000000000",
  46715=>"111111001",
  46716=>"110110100",
  46717=>"111111111",
  46718=>"000010010",
  46719=>"111111110",
  46720=>"101101111",
  46721=>"111111111",
  46722=>"111111010",
  46723=>"111000000",
  46724=>"110100000",
  46725=>"001000000",
  46726=>"000000110",
  46727=>"111111111",
  46728=>"011000000",
  46729=>"111111111",
  46730=>"010010100",
  46731=>"111111111",
  46732=>"000001001",
  46733=>"111111111",
  46734=>"000000010",
  46735=>"000000000",
  46736=>"000000000",
  46737=>"000000000",
  46738=>"100100110",
  46739=>"000101111",
  46740=>"011010111",
  46741=>"111000111",
  46742=>"000100100",
  46743=>"000000000",
  46744=>"111111111",
  46745=>"000000001",
  46746=>"011000000",
  46747=>"000011111",
  46748=>"110000001",
  46749=>"000011011",
  46750=>"110110000",
  46751=>"111100101",
  46752=>"011111001",
  46753=>"000000001",
  46754=>"000000000",
  46755=>"110000000",
  46756=>"000000101",
  46757=>"000000010",
  46758=>"101111001",
  46759=>"111110000",
  46760=>"100000000",
  46761=>"000100100",
  46762=>"001001111",
  46763=>"111111111",
  46764=>"000000000",
  46765=>"001011111",
  46766=>"100111111",
  46767=>"010000000",
  46768=>"111111111",
  46769=>"100011001",
  46770=>"011111111",
  46771=>"111111111",
  46772=>"111001001",
  46773=>"010000001",
  46774=>"100101101",
  46775=>"000000111",
  46776=>"111111111",
  46777=>"000000000",
  46778=>"000111111",
  46779=>"111111011",
  46780=>"111111111",
  46781=>"110000000",
  46782=>"000000000",
  46783=>"111111111",
  46784=>"111100000",
  46785=>"111101001",
  46786=>"111000001",
  46787=>"000011111",
  46788=>"111111111",
  46789=>"100111000",
  46790=>"111111111",
  46791=>"100100000",
  46792=>"001000000",
  46793=>"111111111",
  46794=>"111001101",
  46795=>"000011000",
  46796=>"000010111",
  46797=>"111000000",
  46798=>"000110000",
  46799=>"111111111",
  46800=>"111110110",
  46801=>"111111111",
  46802=>"111111011",
  46803=>"101101000",
  46804=>"000000000",
  46805=>"001001001",
  46806=>"000000111",
  46807=>"000000000",
  46808=>"000000000",
  46809=>"111111000",
  46810=>"000000000",
  46811=>"000000000",
  46812=>"111111101",
  46813=>"111101001",
  46814=>"000001100",
  46815=>"111111000",
  46816=>"000000000",
  46817=>"000000000",
  46818=>"111111111",
  46819=>"100111000",
  46820=>"001000000",
  46821=>"111111111",
  46822=>"000000111",
  46823=>"111111011",
  46824=>"000000111",
  46825=>"101001111",
  46826=>"000000100",
  46827=>"100100111",
  46828=>"111110110",
  46829=>"000000000",
  46830=>"000100111",
  46831=>"011000000",
  46832=>"000000000",
  46833=>"110000000",
  46834=>"100000000",
  46835=>"111110001",
  46836=>"000000000",
  46837=>"111111110",
  46838=>"111000000",
  46839=>"111111000",
  46840=>"111111111",
  46841=>"111111111",
  46842=>"000000000",
  46843=>"000000000",
  46844=>"111111111",
  46845=>"001110111",
  46846=>"000000000",
  46847=>"111111111",
  46848=>"110111111",
  46849=>"111101111",
  46850=>"000000001",
  46851=>"000000000",
  46852=>"001000000",
  46853=>"001000000",
  46854=>"101000000",
  46855=>"000010000",
  46856=>"100111111",
  46857=>"000000000",
  46858=>"111111111",
  46859=>"110110000",
  46860=>"000000000",
  46861=>"000000000",
  46862=>"110100000",
  46863=>"111000111",
  46864=>"100000001",
  46865=>"100100000",
  46866=>"000000000",
  46867=>"111111001",
  46868=>"000000001",
  46869=>"111111111",
  46870=>"001001111",
  46871=>"111111111",
  46872=>"000000000",
  46873=>"000000111",
  46874=>"000000101",
  46875=>"111000000",
  46876=>"111111111",
  46877=>"010000000",
  46878=>"010110110",
  46879=>"111111111",
  46880=>"111001000",
  46881=>"111100111",
  46882=>"001001000",
  46883=>"111101000",
  46884=>"101111111",
  46885=>"000000000",
  46886=>"111110100",
  46887=>"000000000",
  46888=>"111000000",
  46889=>"110111011",
  46890=>"111111111",
  46891=>"111111001",
  46892=>"000010111",
  46893=>"111111111",
  46894=>"111111111",
  46895=>"111111111",
  46896=>"001111001",
  46897=>"100000000",
  46898=>"111111111",
  46899=>"001000000",
  46900=>"111111111",
  46901=>"111111111",
  46902=>"110111111",
  46903=>"000111111",
  46904=>"000000000",
  46905=>"111111111",
  46906=>"000000000",
  46907=>"000000110",
  46908=>"111111011",
  46909=>"001111111",
  46910=>"010001111",
  46911=>"000000000",
  46912=>"111001000",
  46913=>"000000001",
  46914=>"110000000",
  46915=>"000001000",
  46916=>"111111111",
  46917=>"110100000",
  46918=>"100000000",
  46919=>"011011111",
  46920=>"100000000",
  46921=>"110111111",
  46922=>"111111000",
  46923=>"111111111",
  46924=>"111111101",
  46925=>"000000000",
  46926=>"111100111",
  46927=>"011011001",
  46928=>"111001001",
  46929=>"110010110",
  46930=>"111111111",
  46931=>"111111111",
  46932=>"111111111",
  46933=>"011001001",
  46934=>"000011001",
  46935=>"111111011",
  46936=>"111111111",
  46937=>"111111111",
  46938=>"000011111",
  46939=>"111111111",
  46940=>"111111111",
  46941=>"111000000",
  46942=>"100110000",
  46943=>"000000000",
  46944=>"110110111",
  46945=>"110111111",
  46946=>"011010110",
  46947=>"101100111",
  46948=>"100111111",
  46949=>"111100000",
  46950=>"000000100",
  46951=>"101101111",
  46952=>"111110110",
  46953=>"000111111",
  46954=>"000000000",
  46955=>"001000000",
  46956=>"101001101",
  46957=>"000111111",
  46958=>"000000000",
  46959=>"010000000",
  46960=>"000101111",
  46961=>"000000000",
  46962=>"000111110",
  46963=>"001001001",
  46964=>"000000000",
  46965=>"011111111",
  46966=>"111111000",
  46967=>"000110111",
  46968=>"111111111",
  46969=>"111000101",
  46970=>"111111111",
  46971=>"000000000",
  46972=>"000000000",
  46973=>"110000000",
  46974=>"111000111",
  46975=>"000000101",
  46976=>"111111111",
  46977=>"000000000",
  46978=>"000000000",
  46979=>"000000000",
  46980=>"111111111",
  46981=>"111111111",
  46982=>"000110110",
  46983=>"111110100",
  46984=>"000000000",
  46985=>"110100100",
  46986=>"111111111",
  46987=>"111111111",
  46988=>"111111111",
  46989=>"001000000",
  46990=>"000000000",
  46991=>"000000000",
  46992=>"000000000",
  46993=>"111000000",
  46994=>"000000000",
  46995=>"111111111",
  46996=>"111111111",
  46997=>"000000000",
  46998=>"110111111",
  46999=>"101111110",
  47000=>"001011111",
  47001=>"000100111",
  47002=>"000000000",
  47003=>"111111111",
  47004=>"111111111",
  47005=>"111101111",
  47006=>"000000000",
  47007=>"000110010",
  47008=>"000000000",
  47009=>"001010000",
  47010=>"110000000",
  47011=>"000000000",
  47012=>"101101111",
  47013=>"111111011",
  47014=>"111111101",
  47015=>"000000111",
  47016=>"011111111",
  47017=>"110100110",
  47018=>"111011111",
  47019=>"110110000",
  47020=>"111101101",
  47021=>"000000000",
  47022=>"101111111",
  47023=>"000100111",
  47024=>"111111111",
  47025=>"000000111",
  47026=>"111111000",
  47027=>"000000000",
  47028=>"000000000",
  47029=>"000000000",
  47030=>"101001111",
  47031=>"111111111",
  47032=>"000000111",
  47033=>"111111111",
  47034=>"000000000",
  47035=>"111111001",
  47036=>"000000000",
  47037=>"110000110",
  47038=>"111111110",
  47039=>"000000101",
  47040=>"110110110",
  47041=>"111111000",
  47042=>"000111111",
  47043=>"010011011",
  47044=>"111001001",
  47045=>"111111000",
  47046=>"111111010",
  47047=>"000011111",
  47048=>"010110000",
  47049=>"000000000",
  47050=>"110100110",
  47051=>"000000000",
  47052=>"111110110",
  47053=>"000000000",
  47054=>"100100000",
  47055=>"011111000",
  47056=>"111010000",
  47057=>"000000000",
  47058=>"111111111",
  47059=>"111111111",
  47060=>"111110011",
  47061=>"000001111",
  47062=>"000000101",
  47063=>"111110110",
  47064=>"111111001",
  47065=>"000000000",
  47066=>"000000000",
  47067=>"111111111",
  47068=>"000001000",
  47069=>"111110000",
  47070=>"111111111",
  47071=>"100101111",
  47072=>"000100100",
  47073=>"111111111",
  47074=>"000000000",
  47075=>"111111111",
  47076=>"010110111",
  47077=>"111111111",
  47078=>"111000000",
  47079=>"110100111",
  47080=>"111100000",
  47081=>"000011011",
  47082=>"110100000",
  47083=>"100100000",
  47084=>"010010000",
  47085=>"100110110",
  47086=>"000000000",
  47087=>"111111111",
  47088=>"000000011",
  47089=>"110111111",
  47090=>"000000111",
  47091=>"111111111",
  47092=>"000000000",
  47093=>"111111111",
  47094=>"111101001",
  47095=>"111111111",
  47096=>"000000011",
  47097=>"100000000",
  47098=>"110000100",
  47099=>"000001111",
  47100=>"111111111",
  47101=>"000001111",
  47102=>"000000000",
  47103=>"111111010",
  47104=>"110001000",
  47105=>"000000000",
  47106=>"000100101",
  47107=>"000000000",
  47108=>"011011011",
  47109=>"001100100",
  47110=>"111111111",
  47111=>"010000111",
  47112=>"111111101",
  47113=>"111111100",
  47114=>"000000001",
  47115=>"111111111",
  47116=>"010101010",
  47117=>"111111101",
  47118=>"000000000",
  47119=>"110000010",
  47120=>"110100000",
  47121=>"011111111",
  47122=>"111110100",
  47123=>"000111111",
  47124=>"000000000",
  47125=>"111111111",
  47126=>"000000000",
  47127=>"010111011",
  47128=>"111111111",
  47129=>"010000000",
  47130=>"111111111",
  47131=>"111111111",
  47132=>"110000000",
  47133=>"110111001",
  47134=>"100110100",
  47135=>"000011111",
  47136=>"000000000",
  47137=>"111010000",
  47138=>"111001001",
  47139=>"000000000",
  47140=>"101111111",
  47141=>"000001101",
  47142=>"010000000",
  47143=>"000000101",
  47144=>"000000000",
  47145=>"000010111",
  47146=>"011000000",
  47147=>"111100111",
  47148=>"111111100",
  47149=>"100000100",
  47150=>"111111111",
  47151=>"111111001",
  47152=>"110110000",
  47153=>"000000000",
  47154=>"001000000",
  47155=>"011001001",
  47156=>"110110110",
  47157=>"101100010",
  47158=>"111101001",
  47159=>"000000000",
  47160=>"000000000",
  47161=>"000111000",
  47162=>"000000000",
  47163=>"111111111",
  47164=>"000000000",
  47165=>"000100111",
  47166=>"110110110",
  47167=>"001001000",
  47168=>"000000000",
  47169=>"100110110",
  47170=>"111100011",
  47171=>"000000111",
  47172=>"000011011",
  47173=>"010011011",
  47174=>"000111111",
  47175=>"000010110",
  47176=>"000000000",
  47177=>"100111111",
  47178=>"111110100",
  47179=>"111110111",
  47180=>"000000000",
  47181=>"111111111",
  47182=>"000111011",
  47183=>"000000000",
  47184=>"011000000",
  47185=>"111111111",
  47186=>"011011000",
  47187=>"001001000",
  47188=>"000000000",
  47189=>"000000001",
  47190=>"000000001",
  47191=>"111111111",
  47192=>"111011111",
  47193=>"111101101",
  47194=>"000000000",
  47195=>"111111011",
  47196=>"001101111",
  47197=>"000000011",
  47198=>"000110000",
  47199=>"111111111",
  47200=>"100100100",
  47201=>"000000000",
  47202=>"000000111",
  47203=>"000000111",
  47204=>"100000000",
  47205=>"111111101",
  47206=>"000000000",
  47207=>"111111111",
  47208=>"000000000",
  47209=>"010000000",
  47210=>"000000000",
  47211=>"100111111",
  47212=>"001001000",
  47213=>"010000101",
  47214=>"000011111",
  47215=>"111111111",
  47216=>"110110111",
  47217=>"000000000",
  47218=>"111111110",
  47219=>"010111111",
  47220=>"111111101",
  47221=>"000000000",
  47222=>"000000000",
  47223=>"000000001",
  47224=>"000000000",
  47225=>"111100100",
  47226=>"001000000",
  47227=>"011101000",
  47228=>"111111111",
  47229=>"011001001",
  47230=>"111111111",
  47231=>"000000000",
  47232=>"000000001",
  47233=>"111111111",
  47234=>"000100111",
  47235=>"000110011",
  47236=>"001000000",
  47237=>"111000000",
  47238=>"111111010",
  47239=>"000011111",
  47240=>"111111000",
  47241=>"000000000",
  47242=>"000111100",
  47243=>"111111111",
  47244=>"000000000",
  47245=>"111111111",
  47246=>"001000000",
  47247=>"111111000",
  47248=>"111111111",
  47249=>"110110110",
  47250=>"000011111",
  47251=>"111000000",
  47252=>"000111111",
  47253=>"000000011",
  47254=>"111110110",
  47255=>"111000000",
  47256=>"100000101",
  47257=>"101001101",
  47258=>"111000000",
  47259=>"001001001",
  47260=>"000000000",
  47261=>"000000000",
  47262=>"101101001",
  47263=>"000000011",
  47264=>"000100111",
  47265=>"000101111",
  47266=>"111011111",
  47267=>"000011111",
  47268=>"001001001",
  47269=>"111000000",
  47270=>"001101101",
  47271=>"011011011",
  47272=>"000100111",
  47273=>"000000100",
  47274=>"000000111",
  47275=>"111111011",
  47276=>"000000011",
  47277=>"111111011",
  47278=>"111111101",
  47279=>"111111110",
  47280=>"000000001",
  47281=>"111111111",
  47282=>"111111111",
  47283=>"101000000",
  47284=>"001000000",
  47285=>"100000000",
  47286=>"000000110",
  47287=>"000000000",
  47288=>"111011111",
  47289=>"111111111",
  47290=>"001000000",
  47291=>"000000001",
  47292=>"000000000",
  47293=>"000000000",
  47294=>"000000000",
  47295=>"000010111",
  47296=>"000000000",
  47297=>"011110011",
  47298=>"110111110",
  47299=>"000000000",
  47300=>"111111111",
  47301=>"111111111",
  47302=>"000000000",
  47303=>"111111111",
  47304=>"000000000",
  47305=>"000000000",
  47306=>"001000000",
  47307=>"100110110",
  47308=>"000000001",
  47309=>"110111010",
  47310=>"110010000",
  47311=>"000000000",
  47312=>"111111100",
  47313=>"000000000",
  47314=>"000111011",
  47315=>"000000000",
  47316=>"000000000",
  47317=>"001001000",
  47318=>"000000011",
  47319=>"000000100",
  47320=>"000011001",
  47321=>"111001000",
  47322=>"111000001",
  47323=>"111000001",
  47324=>"100110111",
  47325=>"111111111",
  47326=>"000111011",
  47327=>"111001000",
  47328=>"000000000",
  47329=>"110110100",
  47330=>"110111111",
  47331=>"000000000",
  47332=>"001000000",
  47333=>"111000000",
  47334=>"101111001",
  47335=>"111011111",
  47336=>"000000000",
  47337=>"010110110",
  47338=>"100000111",
  47339=>"000000011",
  47340=>"111010000",
  47341=>"000110111",
  47342=>"100100111",
  47343=>"111111111",
  47344=>"100000000",
  47345=>"000010011",
  47346=>"000000000",
  47347=>"000000111",
  47348=>"000100100",
  47349=>"011111111",
  47350=>"000001000",
  47351=>"011001000",
  47352=>"100000100",
  47353=>"000010000",
  47354=>"000101111",
  47355=>"111111010",
  47356=>"000000000",
  47357=>"000000000",
  47358=>"000000000",
  47359=>"111011111",
  47360=>"001001001",
  47361=>"001011011",
  47362=>"000000000",
  47363=>"000001011",
  47364=>"000000000",
  47365=>"110110110",
  47366=>"100100101",
  47367=>"000000000",
  47368=>"010110111",
  47369=>"000000000",
  47370=>"000000001",
  47371=>"000000000",
  47372=>"001001001",
  47373=>"100110110",
  47374=>"111111000",
  47375=>"000000000",
  47376=>"001000000",
  47377=>"000000000",
  47378=>"111000000",
  47379=>"000000111",
  47380=>"000000000",
  47381=>"111111111",
  47382=>"001001001",
  47383=>"111111111",
  47384=>"111111111",
  47385=>"111110000",
  47386=>"011110010",
  47387=>"000111100",
  47388=>"110110110",
  47389=>"001011100",
  47390=>"000000000",
  47391=>"000100110",
  47392=>"000001000",
  47393=>"000000000",
  47394=>"001001001",
  47395=>"111111101",
  47396=>"111100100",
  47397=>"011000000",
  47398=>"100100100",
  47399=>"111111100",
  47400=>"000010000",
  47401=>"100000000",
  47402=>"000000000",
  47403=>"000000000",
  47404=>"000000000",
  47405=>"110111111",
  47406=>"000000000",
  47407=>"000000000",
  47408=>"111111100",
  47409=>"000000000",
  47410=>"100101101",
  47411=>"000111111",
  47412=>"011111011",
  47413=>"000001001",
  47414=>"011000100",
  47415=>"000000000",
  47416=>"000000000",
  47417=>"000000001",
  47418=>"001001011",
  47419=>"100100000",
  47420=>"111111111",
  47421=>"000110110",
  47422=>"001001000",
  47423=>"001001111",
  47424=>"000000011",
  47425=>"000000000",
  47426=>"011011000",
  47427=>"111111111",
  47428=>"101001001",
  47429=>"111000000",
  47430=>"110111111",
  47431=>"111111111",
  47432=>"000000011",
  47433=>"000000000",
  47434=>"111111111",
  47435=>"111111111",
  47436=>"000000000",
  47437=>"111111010",
  47438=>"000100100",
  47439=>"001111111",
  47440=>"111111111",
  47441=>"100000000",
  47442=>"000000000",
  47443=>"010011111",
  47444=>"000000000",
  47445=>"011011011",
  47446=>"111111100",
  47447=>"101000010",
  47448=>"111111111",
  47449=>"000000111",
  47450=>"111000000",
  47451=>"111100111",
  47452=>"111011001",
  47453=>"000110010",
  47454=>"000000000",
  47455=>"110101001",
  47456=>"000000000",
  47457=>"101111111",
  47458=>"110111111",
  47459=>"000000000",
  47460=>"000000000",
  47461=>"000000000",
  47462=>"000110111",
  47463=>"000000000",
  47464=>"111111011",
  47465=>"000000000",
  47466=>"100100110",
  47467=>"111111110",
  47468=>"010000000",
  47469=>"111000000",
  47470=>"000000000",
  47471=>"000010010",
  47472=>"000000111",
  47473=>"000000000",
  47474=>"111000000",
  47475=>"110111111",
  47476=>"111111110",
  47477=>"001000000",
  47478=>"010011111",
  47479=>"001001111",
  47480=>"110110111",
  47481=>"000000111",
  47482=>"111111110",
  47483=>"011000000",
  47484=>"001111010",
  47485=>"101100000",
  47486=>"000000000",
  47487=>"000001111",
  47488=>"110000000",
  47489=>"000000000",
  47490=>"001010110",
  47491=>"001001101",
  47492=>"010011000",
  47493=>"000000000",
  47494=>"011111111",
  47495=>"010000010",
  47496=>"101111111",
  47497=>"100100100",
  47498=>"000101111",
  47499=>"000000000",
  47500=>"101111111",
  47501=>"011011001",
  47502=>"111111101",
  47503=>"111111111",
  47504=>"000000000",
  47505=>"110100100",
  47506=>"100101111",
  47507=>"111111111",
  47508=>"111111000",
  47509=>"000000000",
  47510=>"000000000",
  47511=>"111100001",
  47512=>"000000000",
  47513=>"000000000",
  47514=>"111000000",
  47515=>"111111000",
  47516=>"011000101",
  47517=>"000000000",
  47518=>"111101100",
  47519=>"000000000",
  47520=>"000000001",
  47521=>"000000000",
  47522=>"001000000",
  47523=>"000000000",
  47524=>"000000001",
  47525=>"100000000",
  47526=>"111111111",
  47527=>"101111000",
  47528=>"100110100",
  47529=>"001100100",
  47530=>"111111111",
  47531=>"111111011",
  47532=>"000111100",
  47533=>"110100000",
  47534=>"111110100",
  47535=>"111110000",
  47536=>"000000011",
  47537=>"111110011",
  47538=>"001000000",
  47539=>"111111111",
  47540=>"111111111",
  47541=>"000000000",
  47542=>"111101111",
  47543=>"000110110",
  47544=>"001000000",
  47545=>"000011011",
  47546=>"000000000",
  47547=>"000000000",
  47548=>"000000000",
  47549=>"111001001",
  47550=>"001100000",
  47551=>"011011111",
  47552=>"111111111",
  47553=>"110100010",
  47554=>"000000000",
  47555=>"111111111",
  47556=>"001101101",
  47557=>"000000000",
  47558=>"010011011",
  47559=>"000000000",
  47560=>"111111111",
  47561=>"000000101",
  47562=>"000000000",
  47563=>"011000000",
  47564=>"000000000",
  47565=>"000000000",
  47566=>"100010010",
  47567=>"100100100",
  47568=>"110100000",
  47569=>"000011111",
  47570=>"110000000",
  47571=>"000001111",
  47572=>"000000000",
  47573=>"000000000",
  47574=>"111100000",
  47575=>"111111111",
  47576=>"100111111",
  47577=>"111111111",
  47578=>"111000000",
  47579=>"000000000",
  47580=>"111111000",
  47581=>"111011101",
  47582=>"111111111",
  47583=>"000110110",
  47584=>"000000000",
  47585=>"111111011",
  47586=>"000000000",
  47587=>"000000001",
  47588=>"111111110",
  47589=>"011010010",
  47590=>"000000010",
  47591=>"110111111",
  47592=>"111110111",
  47593=>"110111111",
  47594=>"010010110",
  47595=>"000001000",
  47596=>"111111111",
  47597=>"110110110",
  47598=>"000000000",
  47599=>"111111111",
  47600=>"001111000",
  47601=>"000000000",
  47602=>"111111101",
  47603=>"111111111",
  47604=>"000000000",
  47605=>"100001100",
  47606=>"000000000",
  47607=>"010000000",
  47608=>"111111111",
  47609=>"101101111",
  47610=>"000000000",
  47611=>"101001011",
  47612=>"000100100",
  47613=>"110100101",
  47614=>"000110111",
  47615=>"101000000",
  47616=>"000011001",
  47617=>"111110000",
  47618=>"101000100",
  47619=>"000000000",
  47620=>"000010000",
  47621=>"000000011",
  47622=>"000000000",
  47623=>"000000000",
  47624=>"101111000",
  47625=>"000111111",
  47626=>"000000100",
  47627=>"111111111",
  47628=>"000001110",
  47629=>"111001001",
  47630=>"111111111",
  47631=>"000001000",
  47632=>"000000011",
  47633=>"000000111",
  47634=>"100000000",
  47635=>"000000110",
  47636=>"111111110",
  47637=>"111100000",
  47638=>"010100110",
  47639=>"110111111",
  47640=>"111101001",
  47641=>"011000110",
  47642=>"111111111",
  47643=>"011001000",
  47644=>"001000111",
  47645=>"000001111",
  47646=>"000111111",
  47647=>"000000001",
  47648=>"000001001",
  47649=>"111100100",
  47650=>"110010000",
  47651=>"100111001",
  47652=>"000000000",
  47653=>"111111111",
  47654=>"000111000",
  47655=>"001101111",
  47656=>"000000000",
  47657=>"010111000",
  47658=>"111111000",
  47659=>"000111111",
  47660=>"101101110",
  47661=>"000101111",
  47662=>"111111111",
  47663=>"111111110",
  47664=>"000110111",
  47665=>"000001011",
  47666=>"111111000",
  47667=>"111111111",
  47668=>"000101111",
  47669=>"001011011",
  47670=>"100000110",
  47671=>"000111000",
  47672=>"000001000",
  47673=>"000000110",
  47674=>"000000000",
  47675=>"101000000",
  47676=>"101100101",
  47677=>"001000001",
  47678=>"011111111",
  47679=>"111111001",
  47680=>"110000111",
  47681=>"000000000",
  47682=>"000100111",
  47683=>"000000000",
  47684=>"000110000",
  47685=>"110110110",
  47686=>"111111000",
  47687=>"111111111",
  47688=>"100110010",
  47689=>"000000001",
  47690=>"111101000",
  47691=>"101100111",
  47692=>"010110100",
  47693=>"000111111",
  47694=>"000101111",
  47695=>"111111000",
  47696=>"000000000",
  47697=>"111111011",
  47698=>"001000000",
  47699=>"000000111",
  47700=>"000000111",
  47701=>"000000111",
  47702=>"100000111",
  47703=>"100000000",
  47704=>"111111100",
  47705=>"000000111",
  47706=>"000101111",
  47707=>"110100000",
  47708=>"000000000",
  47709=>"111100110",
  47710=>"111000100",
  47711=>"111111111",
  47712=>"000000000",
  47713=>"000000111",
  47714=>"000000001",
  47715=>"001111111",
  47716=>"000011010",
  47717=>"111100111",
  47718=>"000000000",
  47719=>"000000101",
  47720=>"111111111",
  47721=>"111011111",
  47722=>"111111000",
  47723=>"000000000",
  47724=>"110100000",
  47725=>"111111111",
  47726=>"111101101",
  47727=>"000000111",
  47728=>"000100000",
  47729=>"000000111",
  47730=>"000111111",
  47731=>"111000100",
  47732=>"000000111",
  47733=>"000000000",
  47734=>"000000010",
  47735=>"101001000",
  47736=>"111111011",
  47737=>"000000110",
  47738=>"110110001",
  47739=>"111111001",
  47740=>"110110110",
  47741=>"000000000",
  47742=>"111111111",
  47743=>"111001000",
  47744=>"000000110",
  47745=>"000000111",
  47746=>"000000000",
  47747=>"000000000",
  47748=>"111111111",
  47749=>"111000100",
  47750=>"000111111",
  47751=>"000000000",
  47752=>"000000111",
  47753=>"000000000",
  47754=>"000110000",
  47755=>"000000000",
  47756=>"000000111",
  47757=>"111111111",
  47758=>"000001111",
  47759=>"000000000",
  47760=>"000000111",
  47761=>"000111111",
  47762=>"000000001",
  47763=>"000100000",
  47764=>"110111111",
  47765=>"000000001",
  47766=>"000000000",
  47767=>"001000000",
  47768=>"000000000",
  47769=>"100111101",
  47770=>"110111111",
  47771=>"000001000",
  47772=>"111111111",
  47773=>"111000011",
  47774=>"111111000",
  47775=>"000000111",
  47776=>"111111000",
  47777=>"101000000",
  47778=>"111001111",
  47779=>"000110111",
  47780=>"100111111",
  47781=>"111011111",
  47782=>"111111111",
  47783=>"111111110",
  47784=>"000000101",
  47785=>"101111111",
  47786=>"000000000",
  47787=>"000001111",
  47788=>"001101111",
  47789=>"111111000",
  47790=>"111001000",
  47791=>"100111111",
  47792=>"111000000",
  47793=>"111111110",
  47794=>"100100111",
  47795=>"110000000",
  47796=>"110000000",
  47797=>"000111111",
  47798=>"000000111",
  47799=>"111111111",
  47800=>"111111001",
  47801=>"100000000",
  47802=>"000110111",
  47803=>"000000100",
  47804=>"111111000",
  47805=>"111111111",
  47806=>"100100000",
  47807=>"111111111",
  47808=>"000000000",
  47809=>"111111111",
  47810=>"111001111",
  47811=>"010000000",
  47812=>"100110110",
  47813=>"011111000",
  47814=>"001111111",
  47815=>"010011001",
  47816=>"000000000",
  47817=>"000000000",
  47818=>"000000000",
  47819=>"111000000",
  47820=>"100001001",
  47821=>"100111111",
  47822=>"001111101",
  47823=>"100100111",
  47824=>"111111000",
  47825=>"111111000",
  47826=>"111110000",
  47827=>"000000111",
  47828=>"000111101",
  47829=>"111111111",
  47830=>"000111111",
  47831=>"000110111",
  47832=>"110111000",
  47833=>"111111001",
  47834=>"000000111",
  47835=>"111110000",
  47836=>"000000000",
  47837=>"001000101",
  47838=>"000001001",
  47839=>"001100111",
  47840=>"101111111",
  47841=>"000000111",
  47842=>"110111000",
  47843=>"111111111",
  47844=>"101111111",
  47845=>"011001111",
  47846=>"110000000",
  47847=>"101101000",
  47848=>"011111000",
  47849=>"001001001",
  47850=>"111111011",
  47851=>"111111000",
  47852=>"000000100",
  47853=>"111000000",
  47854=>"110001111",
  47855=>"111110000",
  47856=>"000000000",
  47857=>"011111111",
  47858=>"111100000",
  47859=>"001111111",
  47860=>"001010000",
  47861=>"111111111",
  47862=>"011111100",
  47863=>"000000111",
  47864=>"111111111",
  47865=>"110111000",
  47866=>"111000000",
  47867=>"000111111",
  47868=>"111111000",
  47869=>"010010000",
  47870=>"101000111",
  47871=>"111111111",
  47872=>"000110010",
  47873=>"000111000",
  47874=>"111111000",
  47875=>"110010110",
  47876=>"001101101",
  47877=>"100100110",
  47878=>"111111110",
  47879=>"000111000",
  47880=>"100101111",
  47881=>"000000101",
  47882=>"000000111",
  47883=>"000000001",
  47884=>"000011111",
  47885=>"000000110",
  47886=>"000000111",
  47887=>"001111000",
  47888=>"000000111",
  47889=>"000000000",
  47890=>"000101111",
  47891=>"110111101",
  47892=>"000000000",
  47893=>"111000000",
  47894=>"111110000",
  47895=>"000000111",
  47896=>"000000000",
  47897=>"001000000",
  47898=>"111111111",
  47899=>"000111111",
  47900=>"000111001",
  47901=>"000100110",
  47902=>"111111111",
  47903=>"111101000",
  47904=>"000000000",
  47905=>"011011111",
  47906=>"000000100",
  47907=>"001000000",
  47908=>"000110111",
  47909=>"100111000",
  47910=>"000000010",
  47911=>"111000001",
  47912=>"111110110",
  47913=>"111000000",
  47914=>"101000001",
  47915=>"000000111",
  47916=>"111000000",
  47917=>"001011010",
  47918=>"000000000",
  47919=>"000000111",
  47920=>"110010111",
  47921=>"001000110",
  47922=>"111111111",
  47923=>"000000110",
  47924=>"000000000",
  47925=>"100101101",
  47926=>"000000000",
  47927=>"000000000",
  47928=>"111001001",
  47929=>"111000111",
  47930=>"111101111",
  47931=>"001000000",
  47932=>"110000000",
  47933=>"101000000",
  47934=>"010100111",
  47935=>"111010000",
  47936=>"000000000",
  47937=>"011111111",
  47938=>"111111000",
  47939=>"000000000",
  47940=>"111111111",
  47941=>"111111111",
  47942=>"110111111",
  47943=>"011011000",
  47944=>"101000111",
  47945=>"010111000",
  47946=>"100100100",
  47947=>"011110010",
  47948=>"000000000",
  47949=>"000001111",
  47950=>"101111011",
  47951=>"000001110",
  47952=>"111110111",
  47953=>"000001100",
  47954=>"000001111",
  47955=>"000001000",
  47956=>"000000101",
  47957=>"011011111",
  47958=>"000000000",
  47959=>"011000000",
  47960=>"111111011",
  47961=>"000000111",
  47962=>"011001000",
  47963=>"000001000",
  47964=>"011001101",
  47965=>"001111000",
  47966=>"000000111",
  47967=>"000000000",
  47968=>"001001001",
  47969=>"111111000",
  47970=>"000001001",
  47971=>"001001111",
  47972=>"111111111",
  47973=>"000000000",
  47974=>"111101000",
  47975=>"010000111",
  47976=>"011001000",
  47977=>"000000000",
  47978=>"111111011",
  47979=>"111111111",
  47980=>"110110111",
  47981=>"101101111",
  47982=>"001000110",
  47983=>"000001111",
  47984=>"111111100",
  47985=>"110111111",
  47986=>"000001001",
  47987=>"000000100",
  47988=>"111101000",
  47989=>"000001000",
  47990=>"000100111",
  47991=>"110000110",
  47992=>"111000000",
  47993=>"111111111",
  47994=>"000000000",
  47995=>"111111000",
  47996=>"000111111",
  47997=>"111111000",
  47998=>"000001011",
  47999=>"000000010",
  48000=>"000011011",
  48001=>"000001000",
  48002=>"111011111",
  48003=>"011111000",
  48004=>"111111011",
  48005=>"000000001",
  48006=>"000100111",
  48007=>"000101111",
  48008=>"000000110",
  48009=>"000100101",
  48010=>"000000111",
  48011=>"001000111",
  48012=>"111111111",
  48013=>"001111111",
  48014=>"000001101",
  48015=>"111110000",
  48016=>"110110111",
  48017=>"111111111",
  48018=>"111111101",
  48019=>"111001000",
  48020=>"000000000",
  48021=>"000000000",
  48022=>"000000000",
  48023=>"000000011",
  48024=>"001111111",
  48025=>"000111111",
  48026=>"101111111",
  48027=>"000101000",
  48028=>"111111000",
  48029=>"000101111",
  48030=>"000000111",
  48031=>"000000111",
  48032=>"111111111",
  48033=>"111110000",
  48034=>"100000011",
  48035=>"000000000",
  48036=>"110111111",
  48037=>"000100100",
  48038=>"000010000",
  48039=>"000000011",
  48040=>"000000000",
  48041=>"010000111",
  48042=>"111111110",
  48043=>"000110111",
  48044=>"000111111",
  48045=>"000011111",
  48046=>"111101100",
  48047=>"100100000",
  48048=>"000100110",
  48049=>"000000111",
  48050=>"000000001",
  48051=>"111111000",
  48052=>"111111111",
  48053=>"000000111",
  48054=>"111111111",
  48055=>"000001111",
  48056=>"000000000",
  48057=>"000111111",
  48058=>"101000000",
  48059=>"100000000",
  48060=>"000011111",
  48061=>"111111111",
  48062=>"101000000",
  48063=>"000000010",
  48064=>"000000000",
  48065=>"000000000",
  48066=>"111111111",
  48067=>"001000111",
  48068=>"000011110",
  48069=>"000000000",
  48070=>"011111111",
  48071=>"000000011",
  48072=>"110111000",
  48073=>"111111101",
  48074=>"000000000",
  48075=>"111000000",
  48076=>"000000000",
  48077=>"000000111",
  48078=>"111111110",
  48079=>"111111111",
  48080=>"000000000",
  48081=>"100100000",
  48082=>"000111111",
  48083=>"111111101",
  48084=>"001111111",
  48085=>"000000000",
  48086=>"000000111",
  48087=>"000111111",
  48088=>"100111011",
  48089=>"101001111",
  48090=>"000000000",
  48091=>"000001010",
  48092=>"000111100",
  48093=>"111001101",
  48094=>"000000000",
  48095=>"111011000",
  48096=>"111000000",
  48097=>"010010000",
  48098=>"000000111",
  48099=>"111110111",
  48100=>"110110111",
  48101=>"000000100",
  48102=>"000000000",
  48103=>"000000111",
  48104=>"101000111",
  48105=>"111110111",
  48106=>"010111100",
  48107=>"001001001",
  48108=>"111000000",
  48109=>"011001000",
  48110=>"110111001",
  48111=>"000110111",
  48112=>"000000111",
  48113=>"110111111",
  48114=>"101001000",
  48115=>"011011011",
  48116=>"100000000",
  48117=>"111000000",
  48118=>"000000010",
  48119=>"101111001",
  48120=>"100111101",
  48121=>"110110110",
  48122=>"000000000",
  48123=>"111011000",
  48124=>"011011001",
  48125=>"111111000",
  48126=>"111110110",
  48127=>"101101111",
  48128=>"110111010",
  48129=>"000000000",
  48130=>"000000000",
  48131=>"000000000",
  48132=>"000011111",
  48133=>"000110000",
  48134=>"111111111",
  48135=>"111111111",
  48136=>"111111111",
  48137=>"100100111",
  48138=>"011111111",
  48139=>"011011000",
  48140=>"000100110",
  48141=>"111011011",
  48142=>"000111011",
  48143=>"110111111",
  48144=>"111000000",
  48145=>"010010010",
  48146=>"110111110",
  48147=>"000000000",
  48148=>"111111111",
  48149=>"111111110",
  48150=>"100111111",
  48151=>"011001001",
  48152=>"100000000",
  48153=>"000000111",
  48154=>"111000011",
  48155=>"001001001",
  48156=>"000000000",
  48157=>"100100110",
  48158=>"001001001",
  48159=>"100111110",
  48160=>"000000010",
  48161=>"111100000",
  48162=>"111111001",
  48163=>"000000100",
  48164=>"110000101",
  48165=>"111111111",
  48166=>"000000000",
  48167=>"000000000",
  48168=>"011000011",
  48169=>"000000000",
  48170=>"111111111",
  48171=>"100110111",
  48172=>"100001101",
  48173=>"100000000",
  48174=>"000000100",
  48175=>"110000111",
  48176=>"011111111",
  48177=>"111111111",
  48178=>"011011011",
  48179=>"000000000",
  48180=>"000000101",
  48181=>"000000010",
  48182=>"000000000",
  48183=>"000000101",
  48184=>"001000000",
  48185=>"011000000",
  48186=>"110110000",
  48187=>"011010000",
  48188=>"000000101",
  48189=>"000000000",
  48190=>"000011001",
  48191=>"000000000",
  48192=>"011011011",
  48193=>"001001001",
  48194=>"000000000",
  48195=>"001000000",
  48196=>"000000000",
  48197=>"100100111",
  48198=>"111111110",
  48199=>"111111111",
  48200=>"111011001",
  48201=>"101000000",
  48202=>"111111000",
  48203=>"110100110",
  48204=>"111111111",
  48205=>"001011111",
  48206=>"000000100",
  48207=>"000000111",
  48208=>"110110000",
  48209=>"111001000",
  48210=>"000000001",
  48211=>"011011100",
  48212=>"000010010",
  48213=>"000010000",
  48214=>"000000000",
  48215=>"010000111",
  48216=>"100100000",
  48217=>"000000000",
  48218=>"100110000",
  48219=>"011111111",
  48220=>"011011000",
  48221=>"000111011",
  48222=>"001001111",
  48223=>"000111111",
  48224=>"000100000",
  48225=>"000010110",
  48226=>"000000000",
  48227=>"001001001",
  48228=>"000000000",
  48229=>"000000011",
  48230=>"000110010",
  48231=>"111111111",
  48232=>"000001000",
  48233=>"001001100",
  48234=>"111000000",
  48235=>"011011111",
  48236=>"000000010",
  48237=>"111111000",
  48238=>"010000000",
  48239=>"111111001",
  48240=>"000000000",
  48241=>"000000000",
  48242=>"000100111",
  48243=>"110001001",
  48244=>"000000000",
  48245=>"000010000",
  48246=>"110001000",
  48247=>"111111111",
  48248=>"100100001",
  48249=>"110111100",
  48250=>"000001111",
  48251=>"011111010",
  48252=>"000000010",
  48253=>"101111110",
  48254=>"000000000",
  48255=>"000000000",
  48256=>"110101111",
  48257=>"110000000",
  48258=>"110100000",
  48259=>"111111011",
  48260=>"111111000",
  48261=>"100111111",
  48262=>"111111111",
  48263=>"000000000",
  48264=>"011011110",
  48265=>"000000000",
  48266=>"111111111",
  48267=>"000000000",
  48268=>"111111111",
  48269=>"111111111",
  48270=>"011000000",
  48271=>"111111011",
  48272=>"001011111",
  48273=>"110110110",
  48274=>"111011001",
  48275=>"111111111",
  48276=>"000000000",
  48277=>"111111010",
  48278=>"101000000",
  48279=>"101100000",
  48280=>"100100000",
  48281=>"100111111",
  48282=>"000011111",
  48283=>"000000000",
  48284=>"111111001",
  48285=>"000011010",
  48286=>"000110000",
  48287=>"111100000",
  48288=>"111000000",
  48289=>"000111111",
  48290=>"111111010",
  48291=>"111111000",
  48292=>"000111111",
  48293=>"000000000",
  48294=>"010011011",
  48295=>"010110010",
  48296=>"111110111",
  48297=>"110110111",
  48298=>"000000000",
  48299=>"010011011",
  48300=>"111110000",
  48301=>"001011011",
  48302=>"111111111",
  48303=>"111111101",
  48304=>"000000000",
  48305=>"110110000",
  48306=>"110111011",
  48307=>"000000111",
  48308=>"110111111",
  48309=>"100110111",
  48310=>"000000110",
  48311=>"101111000",
  48312=>"000001000",
  48313=>"100001000",
  48314=>"000000000",
  48315=>"001100110",
  48316=>"001001000",
  48317=>"111111110",
  48318=>"111111111",
  48319=>"111011011",
  48320=>"000000000",
  48321=>"100000000",
  48322=>"011010100",
  48323=>"000000000",
  48324=>"100000000",
  48325=>"111000100",
  48326=>"110100100",
  48327=>"111111011",
  48328=>"110110011",
  48329=>"011000000",
  48330=>"010110110",
  48331=>"111110100",
  48332=>"000001111",
  48333=>"100100100",
  48334=>"000000000",
  48335=>"000010000",
  48336=>"000100110",
  48337=>"111111111",
  48338=>"000011111",
  48339=>"000100000",
  48340=>"011011000",
  48341=>"001000000",
  48342=>"000000111",
  48343=>"000001111",
  48344=>"100000000",
  48345=>"011110100",
  48346=>"110000100",
  48347=>"010010000",
  48348=>"000100111",
  48349=>"100000000",
  48350=>"111111001",
  48351=>"010110000",
  48352=>"001111111",
  48353=>"000001001",
  48354=>"101101101",
  48355=>"111111011",
  48356=>"110110110",
  48357=>"111111101",
  48358=>"001001000",
  48359=>"000000000",
  48360=>"111001110",
  48361=>"110111110",
  48362=>"111111110",
  48363=>"000011011",
  48364=>"000001111",
  48365=>"000000000",
  48366=>"010010111",
  48367=>"000000000",
  48368=>"000000110",
  48369=>"111111111",
  48370=>"110011111",
  48371=>"001001000",
  48372=>"111111111",
  48373=>"001000000",
  48374=>"011101100",
  48375=>"011111011",
  48376=>"111011111",
  48377=>"000000000",
  48378=>"101111111",
  48379=>"000000000",
  48380=>"111111111",
  48381=>"111110110",
  48382=>"110010000",
  48383=>"000000000",
  48384=>"001100000",
  48385=>"000000110",
  48386=>"111111111",
  48387=>"100000000",
  48388=>"000000000",
  48389=>"000000000",
  48390=>"111101111",
  48391=>"000000110",
  48392=>"111111111",
  48393=>"000000000",
  48394=>"100100111",
  48395=>"010011111",
  48396=>"000000000",
  48397=>"000101111",
  48398=>"111111111",
  48399=>"000001111",
  48400=>"000000000",
  48401=>"100000000",
  48402=>"000100110",
  48403=>"000100000",
  48404=>"000000000",
  48405=>"111111111",
  48406=>"001001011",
  48407=>"000000000",
  48408=>"100110011",
  48409=>"110011011",
  48410=>"110110000",
  48411=>"010010000",
  48412=>"100100110",
  48413=>"010011001",
  48414=>"000000000",
  48415=>"000011011",
  48416=>"001010001",
  48417=>"100111111",
  48418=>"111111111",
  48419=>"000000000",
  48420=>"100100111",
  48421=>"011111111",
  48422=>"111111111",
  48423=>"001110000",
  48424=>"110111111",
  48425=>"000000000",
  48426=>"111110110",
  48427=>"000001000",
  48428=>"111011001",
  48429=>"000000000",
  48430=>"000011111",
  48431=>"101111111",
  48432=>"010110111",
  48433=>"000000001",
  48434=>"110010000",
  48435=>"000000000",
  48436=>"111000000",
  48437=>"110111101",
  48438=>"111001001",
  48439=>"111000000",
  48440=>"111010111",
  48441=>"111000000",
  48442=>"000000011",
  48443=>"100111111",
  48444=>"010010111",
  48445=>"100101101",
  48446=>"010011011",
  48447=>"000000110",
  48448=>"000000000",
  48449=>"011001000",
  48450=>"001000000",
  48451=>"111111000",
  48452=>"111111111",
  48453=>"000000000",
  48454=>"110110001",
  48455=>"111111010",
  48456=>"000000000",
  48457=>"100100111",
  48458=>"111111110",
  48459=>"001111101",
  48460=>"000000000",
  48461=>"111111111",
  48462=>"000000010",
  48463=>"001000000",
  48464=>"111111011",
  48465=>"000010010",
  48466=>"110110111",
  48467=>"010010011",
  48468=>"000000000",
  48469=>"001001001",
  48470=>"011111010",
  48471=>"111111111",
  48472=>"000100001",
  48473=>"000000000",
  48474=>"000000011",
  48475=>"111111111",
  48476=>"001001101",
  48477=>"110111111",
  48478=>"001011111",
  48479=>"111111111",
  48480=>"111111100",
  48481=>"111111111",
  48482=>"011111111",
  48483=>"111111100",
  48484=>"000110111",
  48485=>"111111000",
  48486=>"000000000",
  48487=>"011111111",
  48488=>"000011011",
  48489=>"110110100",
  48490=>"000000000",
  48491=>"011001000",
  48492=>"000000000",
  48493=>"001001011",
  48494=>"111111111",
  48495=>"000000001",
  48496=>"111111011",
  48497=>"100101001",
  48498=>"110110000",
  48499=>"110111011",
  48500=>"000000000",
  48501=>"000000000",
  48502=>"111011000",
  48503=>"111111111",
  48504=>"111111111",
  48505=>"111000000",
  48506=>"111111110",
  48507=>"011111010",
  48508=>"100100000",
  48509=>"000000110",
  48510=>"110111111",
  48511=>"000000000",
  48512=>"000000000",
  48513=>"000000000",
  48514=>"001111111",
  48515=>"111111100",
  48516=>"111111000",
  48517=>"000000101",
  48518=>"110110100",
  48519=>"001101001",
  48520=>"000000000",
  48521=>"111111111",
  48522=>"111000000",
  48523=>"100100100",
  48524=>"111111111",
  48525=>"001000001",
  48526=>"000000000",
  48527=>"011111101",
  48528=>"000000000",
  48529=>"111111111",
  48530=>"111110111",
  48531=>"011011011",
  48532=>"000000000",
  48533=>"000010010",
  48534=>"010011011",
  48535=>"001010111",
  48536=>"001001000",
  48537=>"000000011",
  48538=>"111101000",
  48539=>"001000000",
  48540=>"110100111",
  48541=>"000000000",
  48542=>"111101000",
  48543=>"111111111",
  48544=>"111111011",
  48545=>"000010011",
  48546=>"000100111",
  48547=>"101000000",
  48548=>"100000101",
  48549=>"110111000",
  48550=>"000110111",
  48551=>"011110100",
  48552=>"111111111",
  48553=>"111111011",
  48554=>"100110011",
  48555=>"000000000",
  48556=>"000000001",
  48557=>"111111111",
  48558=>"000000000",
  48559=>"000000000",
  48560=>"111111110",
  48561=>"111111111",
  48562=>"000000000",
  48563=>"011011001",
  48564=>"111111001",
  48565=>"111001000",
  48566=>"111111111",
  48567=>"111110110",
  48568=>"111110011",
  48569=>"111111111",
  48570=>"000001001",
  48571=>"100100100",
  48572=>"111110100",
  48573=>"111011111",
  48574=>"111111111",
  48575=>"000010110",
  48576=>"110000000",
  48577=>"001001000",
  48578=>"111111111",
  48579=>"111011111",
  48580=>"000000000",
  48581=>"010011111",
  48582=>"110001011",
  48583=>"000111100",
  48584=>"101100000",
  48585=>"000000111",
  48586=>"101000100",
  48587=>"110111000",
  48588=>"100000000",
  48589=>"100000100",
  48590=>"111101111",
  48591=>"111011010",
  48592=>"000000111",
  48593=>"111111111",
  48594=>"100100000",
  48595=>"011011011",
  48596=>"000010000",
  48597=>"100110000",
  48598=>"000011011",
  48599=>"001011011",
  48600=>"000000000",
  48601=>"000110110",
  48602=>"000000000",
  48603=>"111111111",
  48604=>"001001111",
  48605=>"001010111",
  48606=>"000010011",
  48607=>"010110010",
  48608=>"001011111",
  48609=>"111110111",
  48610=>"100100110",
  48611=>"100001101",
  48612=>"000111111",
  48613=>"111011001",
  48614=>"101100100",
  48615=>"000110000",
  48616=>"111100000",
  48617=>"111111111",
  48618=>"011010000",
  48619=>"001011110",
  48620=>"000001000",
  48621=>"110110110",
  48622=>"000000000",
  48623=>"110110010",
  48624=>"000000000",
  48625=>"000000000",
  48626=>"011011011",
  48627=>"110110110",
  48628=>"000000000",
  48629=>"111000110",
  48630=>"000000011",
  48631=>"110000000",
  48632=>"000100000",
  48633=>"111111101",
  48634=>"000000000",
  48635=>"111010000",
  48636=>"111000000",
  48637=>"111011011",
  48638=>"000000000",
  48639=>"111111001",
  48640=>"001001001",
  48641=>"111101100",
  48642=>"111000000",
  48643=>"000000000",
  48644=>"001000001",
  48645=>"110110111",
  48646=>"111111111",
  48647=>"000000000",
  48648=>"000011000",
  48649=>"110110100",
  48650=>"110111111",
  48651=>"111110110",
  48652=>"111100111",
  48653=>"111111111",
  48654=>"000000000",
  48655=>"111000111",
  48656=>"111111001",
  48657=>"000000000",
  48658=>"000000000",
  48659=>"110111111",
  48660=>"010111001",
  48661=>"111111000",
  48662=>"000001001",
  48663=>"111100110",
  48664=>"111111111",
  48665=>"100000000",
  48666=>"111111111",
  48667=>"111111111",
  48668=>"111111111",
  48669=>"000000000",
  48670=>"011011111",
  48671=>"110110111",
  48672=>"001000110",
  48673=>"111111111",
  48674=>"001011011",
  48675=>"111111111",
  48676=>"001000000",
  48677=>"100100111",
  48678=>"111110111",
  48679=>"011111110",
  48680=>"000000000",
  48681=>"000000100",
  48682=>"111110100",
  48683=>"111111111",
  48684=>"000101110",
  48685=>"000100111",
  48686=>"111111011",
  48687=>"111111100",
  48688=>"001011001",
  48689=>"000000000",
  48690=>"000100110",
  48691=>"011000100",
  48692=>"111010010",
  48693=>"011000000",
  48694=>"111111111",
  48695=>"000000111",
  48696=>"000000000",
  48697=>"000000110",
  48698=>"111000001",
  48699=>"000000000",
  48700=>"110110110",
  48701=>"000000000",
  48702=>"111110110",
  48703=>"000000000",
  48704=>"011111111",
  48705=>"100000100",
  48706=>"110111111",
  48707=>"000000111",
  48708=>"110111111",
  48709=>"000100100",
  48710=>"000000000",
  48711=>"000000001",
  48712=>"000011111",
  48713=>"000000001",
  48714=>"000000000",
  48715=>"001000111",
  48716=>"111111101",
  48717=>"111011011",
  48718=>"010010000",
  48719=>"111111111",
  48720=>"111001000",
  48721=>"010111100",
  48722=>"101000001",
  48723=>"001111111",
  48724=>"111111111",
  48725=>"000110000",
  48726=>"111001000",
  48727=>"111111111",
  48728=>"011000000",
  48729=>"000000101",
  48730=>"000010000",
  48731=>"011011111",
  48732=>"000001000",
  48733=>"000001000",
  48734=>"000000111",
  48735=>"100110011",
  48736=>"001000000",
  48737=>"111011010",
  48738=>"100000000",
  48739=>"000000111",
  48740=>"010001000",
  48741=>"101011111",
  48742=>"000000000",
  48743=>"111111010",
  48744=>"111111111",
  48745=>"000000101",
  48746=>"110000000",
  48747=>"000000000",
  48748=>"011000110",
  48749=>"000000000",
  48750=>"111111000",
  48751=>"000000000",
  48752=>"111111111",
  48753=>"000000111",
  48754=>"000000001",
  48755=>"110111111",
  48756=>"111101111",
  48757=>"001000000",
  48758=>"000000000",
  48759=>"111111111",
  48760=>"001001011",
  48761=>"100000000",
  48762=>"000010100",
  48763=>"000000000",
  48764=>"110011001",
  48765=>"000000000",
  48766=>"001111111",
  48767=>"111111111",
  48768=>"110111111",
  48769=>"000000000",
  48770=>"000000001",
  48771=>"111000000",
  48772=>"000000111",
  48773=>"100000000",
  48774=>"000001011",
  48775=>"000000111",
  48776=>"111110111",
  48777=>"001000110",
  48778=>"000000000",
  48779=>"111101111",
  48780=>"001000000",
  48781=>"111101000",
  48782=>"111111111",
  48783=>"000011111",
  48784=>"110111000",
  48785=>"011011000",
  48786=>"111010000",
  48787=>"011001001",
  48788=>"111000000",
  48789=>"000011011",
  48790=>"111111110",
  48791=>"000001000",
  48792=>"000000001",
  48793=>"111111111",
  48794=>"111111111",
  48795=>"000111111",
  48796=>"111000000",
  48797=>"011011000",
  48798=>"111111011",
  48799=>"111111111",
  48800=>"010000000",
  48801=>"000000000",
  48802=>"011000000",
  48803=>"000000000",
  48804=>"001111111",
  48805=>"111011011",
  48806=>"101001001",
  48807=>"111100100",
  48808=>"110111111",
  48809=>"000000011",
  48810=>"000100100",
  48811=>"000000000",
  48812=>"110111000",
  48813=>"110001000",
  48814=>"001000000",
  48815=>"001000111",
  48816=>"111000000",
  48817=>"111000000",
  48818=>"111111011",
  48819=>"000100110",
  48820=>"000011001",
  48821=>"111111111",
  48822=>"000000001",
  48823=>"111100000",
  48824=>"100000010",
  48825=>"111100111",
  48826=>"000000111",
  48827=>"000000111",
  48828=>"000000000",
  48829=>"111100101",
  48830=>"000001000",
  48831=>"000000000",
  48832=>"000000000",
  48833=>"111010010",
  48834=>"000001101",
  48835=>"111111111",
  48836=>"000000110",
  48837=>"000000000",
  48838=>"100111110",
  48839=>"001101111",
  48840=>"000000111",
  48841=>"111111111",
  48842=>"011000000",
  48843=>"000000000",
  48844=>"111000111",
  48845=>"000111111",
  48846=>"110110111",
  48847=>"111111111",
  48848=>"111111111",
  48849=>"100110110",
  48850=>"111001001",
  48851=>"111111111",
  48852=>"101001001",
  48853=>"111011111",
  48854=>"000010000",
  48855=>"000000001",
  48856=>"000000000",
  48857=>"000100110",
  48858=>"111111111",
  48859=>"111111000",
  48860=>"111111111",
  48861=>"111010000",
  48862=>"000000000",
  48863=>"110110110",
  48864=>"111111111",
  48865=>"000011011",
  48866=>"000000000",
  48867=>"000000100",
  48868=>"000000111",
  48869=>"001100111",
  48870=>"111110111",
  48871=>"100110111",
  48872=>"001000000",
  48873=>"001011001",
  48874=>"111111010",
  48875=>"000000000",
  48876=>"011110110",
  48877=>"000111111",
  48878=>"111111111",
  48879=>"111000000",
  48880=>"111100000",
  48881=>"100000000",
  48882=>"000000111",
  48883=>"001000011",
  48884=>"111111111",
  48885=>"001001000",
  48886=>"111101000",
  48887=>"111011000",
  48888=>"000000000",
  48889=>"000000000",
  48890=>"111000111",
  48891=>"111110000",
  48892=>"111111111",
  48893=>"111111111",
  48894=>"000000100",
  48895=>"000000000",
  48896=>"100000001",
  48897=>"100000111",
  48898=>"000000000",
  48899=>"111111111",
  48900=>"111101111",
  48901=>"111000000",
  48902=>"001001000",
  48903=>"111111000",
  48904=>"000001110",
  48905=>"100000100",
  48906=>"101000000",
  48907=>"011000000",
  48908=>"000011111",
  48909=>"110110111",
  48910=>"110001111",
  48911=>"101001000",
  48912=>"111111000",
  48913=>"111000000",
  48914=>"010010000",
  48915=>"111010001",
  48916=>"110000000",
  48917=>"101001000",
  48918=>"100100111",
  48919=>"111011111",
  48920=>"001000011",
  48921=>"000011111",
  48922=>"111001100",
  48923=>"111110111",
  48924=>"111111111",
  48925=>"111111111",
  48926=>"000000000",
  48927=>"111000000",
  48928=>"111111001",
  48929=>"000000000",
  48930=>"010000111",
  48931=>"111101111",
  48932=>"111111111",
  48933=>"000000111",
  48934=>"111111111",
  48935=>"000101000",
  48936=>"100000110",
  48937=>"111111111",
  48938=>"110000000",
  48939=>"000000110",
  48940=>"111111111",
  48941=>"000000011",
  48942=>"101111010",
  48943=>"101000000",
  48944=>"111110110",
  48945=>"111111111",
  48946=>"000000000",
  48947=>"110110100",
  48948=>"111111111",
  48949=>"111111111",
  48950=>"111000000",
  48951=>"111111011",
  48952=>"011111111",
  48953=>"000000111",
  48954=>"110010000",
  48955=>"111000000",
  48956=>"111000110",
  48957=>"111000000",
  48958=>"000000000",
  48959=>"001111111",
  48960=>"111111111",
  48961=>"000011000",
  48962=>"111111111",
  48963=>"000011111",
  48964=>"010110000",
  48965=>"111111111",
  48966=>"110010011",
  48967=>"111111111",
  48968=>"000000000",
  48969=>"011000000",
  48970=>"111001111",
  48971=>"110110111",
  48972=>"011111111",
  48973=>"000111011",
  48974=>"000000110",
  48975=>"001000000",
  48976=>"011011011",
  48977=>"000110111",
  48978=>"111111011",
  48979=>"000000000",
  48980=>"000000000",
  48981=>"011110110",
  48982=>"111000100",
  48983=>"111011001",
  48984=>"111111111",
  48985=>"011001001",
  48986=>"111111111",
  48987=>"000110110",
  48988=>"000000000",
  48989=>"000000000",
  48990=>"000000000",
  48991=>"110111010",
  48992=>"000000000",
  48993=>"000000011",
  48994=>"000110110",
  48995=>"001011111",
  48996=>"000000000",
  48997=>"111101111",
  48998=>"111000000",
  48999=>"111111000",
  49000=>"111011111",
  49001=>"110100100",
  49002=>"111111111",
  49003=>"010010011",
  49004=>"011011000",
  49005=>"100111110",
  49006=>"111111111",
  49007=>"111110111",
  49008=>"000000000",
  49009=>"111111100",
  49010=>"000000000",
  49011=>"000000100",
  49012=>"000000111",
  49013=>"000000110",
  49014=>"000011011",
  49015=>"111111111",
  49016=>"000000111",
  49017=>"111001111",
  49018=>"000001111",
  49019=>"110010000",
  49020=>"000000101",
  49021=>"111111101",
  49022=>"111011100",
  49023=>"011000000",
  49024=>"100000100",
  49025=>"000100010",
  49026=>"010011001",
  49027=>"000011111",
  49028=>"010000001",
  49029=>"111111111",
  49030=>"000111111",
  49031=>"111111111",
  49032=>"001000101",
  49033=>"111000000",
  49034=>"000000000",
  49035=>"111111110",
  49036=>"111000000",
  49037=>"110001001",
  49038=>"100000000",
  49039=>"111101111",
  49040=>"000000000",
  49041=>"111111011",
  49042=>"010000000",
  49043=>"000000001",
  49044=>"111110000",
  49045=>"110110110",
  49046=>"111101111",
  49047=>"111111111",
  49048=>"111111111",
  49049=>"001000001",
  49050=>"000111111",
  49051=>"111111110",
  49052=>"000000100",
  49053=>"111111111",
  49054=>"000000000",
  49055=>"000000111",
  49056=>"000000000",
  49057=>"111111000",
  49058=>"000111111",
  49059=>"000010000",
  49060=>"000000000",
  49061=>"111111110",
  49062=>"000000000",
  49063=>"000000000",
  49064=>"001001111",
  49065=>"000000110",
  49066=>"101101111",
  49067=>"001001001",
  49068=>"000000001",
  49069=>"111111111",
  49070=>"000000000",
  49071=>"000000001",
  49072=>"111100000",
  49073=>"110000000",
  49074=>"111111111",
  49075=>"111111111",
  49076=>"001001011",
  49077=>"000111111",
  49078=>"000000000",
  49079=>"011111011",
  49080=>"111001001",
  49081=>"100110001",
  49082=>"111111111",
  49083=>"111001000",
  49084=>"000000000",
  49085=>"111111111",
  49086=>"100000000",
  49087=>"100001001",
  49088=>"000000000",
  49089=>"110111111",
  49090=>"000000000",
  49091=>"110110000",
  49092=>"111000000",
  49093=>"111111000",
  49094=>"000101000",
  49095=>"111111111",
  49096=>"111110000",
  49097=>"100110110",
  49098=>"010000110",
  49099=>"001111111",
  49100=>"111101111",
  49101=>"111101100",
  49102=>"100000000",
  49103=>"001000000",
  49104=>"000000110",
  49105=>"100000100",
  49106=>"011000000",
  49107=>"101100111",
  49108=>"100110111",
  49109=>"111111111",
  49110=>"000000010",
  49111=>"110110110",
  49112=>"000100111",
  49113=>"111110100",
  49114=>"111111111",
  49115=>"100100111",
  49116=>"111111111",
  49117=>"011000100",
  49118=>"101101000",
  49119=>"000101111",
  49120=>"111111111",
  49121=>"001001111",
  49122=>"110110100",
  49123=>"001000000",
  49124=>"111111111",
  49125=>"101000000",
  49126=>"000011001",
  49127=>"110010000",
  49128=>"111001000",
  49129=>"111111111",
  49130=>"111111111",
  49131=>"111111111",
  49132=>"011010000",
  49133=>"111101100",
  49134=>"000000001",
  49135=>"000100100",
  49136=>"000000100",
  49137=>"000000000",
  49138=>"000010110",
  49139=>"010111111",
  49140=>"111111101",
  49141=>"111111000",
  49142=>"000000000",
  49143=>"111111010",
  49144=>"100111111",
  49145=>"111011000",
  49146=>"000100100",
  49147=>"000000000",
  49148=>"111111110",
  49149=>"111110110",
  49150=>"111110110",
  49151=>"111011011",
  49152=>"010000000",
  49153=>"111111111",
  49154=>"000000000",
  49155=>"110111111",
  49156=>"000000100",
  49157=>"111111000",
  49158=>"111101001",
  49159=>"111111111",
  49160=>"001111111",
  49161=>"110000000",
  49162=>"001111111",
  49163=>"110100111",
  49164=>"000101111",
  49165=>"000000111",
  49166=>"000000011",
  49167=>"111111111",
  49168=>"000000000",
  49169=>"000001000",
  49170=>"111011001",
  49171=>"100101111",
  49172=>"111111000",
  49173=>"111001111",
  49174=>"000001011",
  49175=>"000100110",
  49176=>"001000000",
  49177=>"101110010",
  49178=>"111111111",
  49179=>"110110110",
  49180=>"000000000",
  49181=>"000000000",
  49182=>"001010010",
  49183=>"111111111",
  49184=>"111111111",
  49185=>"000010110",
  49186=>"100110010",
  49187=>"111000000",
  49188=>"000000001",
  49189=>"000000000",
  49190=>"001001100",
  49191=>"000000000",
  49192=>"101001111",
  49193=>"000000000",
  49194=>"000000000",
  49195=>"011000000",
  49196=>"111111111",
  49197=>"111111000",
  49198=>"111011000",
  49199=>"000000000",
  49200=>"000000000",
  49201=>"100000000",
  49202=>"110110110",
  49203=>"111111111",
  49204=>"000110000",
  49205=>"111001000",
  49206=>"100110000",
  49207=>"101111011",
  49208=>"111100111",
  49209=>"111111111",
  49210=>"000000001",
  49211=>"011011011",
  49212=>"000000000",
  49213=>"011000000",
  49214=>"100000000",
  49215=>"111111111",
  49216=>"000000101",
  49217=>"000100000",
  49218=>"000011111",
  49219=>"000000111",
  49220=>"000110111",
  49221=>"000000000",
  49222=>"000100000",
  49223=>"111111111",
  49224=>"101100100",
  49225=>"101000101",
  49226=>"001000000",
  49227=>"000000000",
  49228=>"111111100",
  49229=>"000100111",
  49230=>"111000000",
  49231=>"111111111",
  49232=>"100100110",
  49233=>"000000000",
  49234=>"000111111",
  49235=>"001001010",
  49236=>"000000001",
  49237=>"111100100",
  49238=>"111011010",
  49239=>"000000000",
  49240=>"100100111",
  49241=>"001000111",
  49242=>"111111001",
  49243=>"111111110",
  49244=>"001000000",
  49245=>"000000000",
  49246=>"111111111",
  49247=>"011011111",
  49248=>"001001111",
  49249=>"111111111",
  49250=>"111111111",
  49251=>"000000000",
  49252=>"001000100",
  49253=>"100000110",
  49254=>"001000000",
  49255=>"011010000",
  49256=>"000000000",
  49257=>"000000000",
  49258=>"111111111",
  49259=>"001001111",
  49260=>"001000000",
  49261=>"101101101",
  49262=>"111110111",
  49263=>"011000000",
  49264=>"111001000",
  49265=>"000000000",
  49266=>"000011111",
  49267=>"101111111",
  49268=>"000000000",
  49269=>"000100100",
  49270=>"111111111",
  49271=>"111111111",
  49272=>"111111111",
  49273=>"000000000",
  49274=>"000000000",
  49275=>"111111111",
  49276=>"111110000",
  49277=>"000000000",
  49278=>"000010000",
  49279=>"000000000",
  49280=>"111111111",
  49281=>"000100000",
  49282=>"111110111",
  49283=>"000000100",
  49284=>"100111111",
  49285=>"000000000",
  49286=>"000000110",
  49287=>"000000001",
  49288=>"001000011",
  49289=>"000100111",
  49290=>"111111111",
  49291=>"000000000",
  49292=>"111100111",
  49293=>"111111111",
  49294=>"111001000",
  49295=>"111111101",
  49296=>"111111111",
  49297=>"100000010",
  49298=>"000000000",
  49299=>"111111111",
  49300=>"010011111",
  49301=>"111011111",
  49302=>"111111111",
  49303=>"101000000",
  49304=>"000000111",
  49305=>"000100000",
  49306=>"000000100",
  49307=>"100000000",
  49308=>"000000000",
  49309=>"101000110",
  49310=>"111111111",
  49311=>"000000000",
  49312=>"111111111",
  49313=>"001000000",
  49314=>"100000110",
  49315=>"000000000",
  49316=>"000000000",
  49317=>"111000100",
  49318=>"001010000",
  49319=>"111111111",
  49320=>"111111111",
  49321=>"111001000",
  49322=>"011000000",
  49323=>"001000111",
  49324=>"111111111",
  49325=>"111111000",
  49326=>"000000110",
  49327=>"000000101",
  49328=>"111011101",
  49329=>"111111111",
  49330=>"001011011",
  49331=>"111100000",
  49332=>"111111111",
  49333=>"000011111",
  49334=>"111111111",
  49335=>"111101111",
  49336=>"000100110",
  49337=>"111111101",
  49338=>"000000000",
  49339=>"000000000",
  49340=>"000111111",
  49341=>"011000000",
  49342=>"000000111",
  49343=>"000000000",
  49344=>"000000000",
  49345=>"111111110",
  49346=>"100000000",
  49347=>"000010010",
  49348=>"111111111",
  49349=>"000000001",
  49350=>"000000000",
  49351=>"000000110",
  49352=>"000000100",
  49353=>"000000000",
  49354=>"100000000",
  49355=>"011001001",
  49356=>"001000000",
  49357=>"000000000",
  49358=>"000000111",
  49359=>"111111111",
  49360=>"111111000",
  49361=>"001000000",
  49362=>"111111111",
  49363=>"000000000",
  49364=>"101100100",
  49365=>"111111111",
  49366=>"000000000",
  49367=>"100100100",
  49368=>"000000011",
  49369=>"111110000",
  49370=>"000000000",
  49371=>"101000111",
  49372=>"000100100",
  49373=>"011111111",
  49374=>"100111001",
  49375=>"101111110",
  49376=>"000010010",
  49377=>"000010010",
  49378=>"000000000",
  49379=>"110000000",
  49380=>"101111000",
  49381=>"111110110",
  49382=>"011001001",
  49383=>"111111111",
  49384=>"000000000",
  49385=>"111111111",
  49386=>"100101111",
  49387=>"111111111",
  49388=>"111111001",
  49389=>"011100000",
  49390=>"111111111",
  49391=>"111101101",
  49392=>"110111111",
  49393=>"101101001",
  49394=>"000000000",
  49395=>"000000000",
  49396=>"000000000",
  49397=>"111100110",
  49398=>"000000000",
  49399=>"000000000",
  49400=>"111111111",
  49401=>"111111111",
  49402=>"100100100",
  49403=>"000000000",
  49404=>"111111111",
  49405=>"111011011",
  49406=>"111110110",
  49407=>"111111111",
  49408=>"111111111",
  49409=>"111111011",
  49410=>"000000000",
  49411=>"111111000",
  49412=>"111000001",
  49413=>"000000001",
  49414=>"110110111",
  49415=>"111111110",
  49416=>"111110111",
  49417=>"000000000",
  49418=>"100000000",
  49419=>"000000000",
  49420=>"001001001",
  49421=>"111111111",
  49422=>"000010111",
  49423=>"010000000",
  49424=>"001000100",
  49425=>"100100111",
  49426=>"111111111",
  49427=>"100100000",
  49428=>"000000000",
  49429=>"111100101",
  49430=>"111001001",
  49431=>"000000000",
  49432=>"111111000",
  49433=>"111111000",
  49434=>"111111101",
  49435=>"000011011",
  49436=>"010110110",
  49437=>"110100100",
  49438=>"111001000",
  49439=>"111111111",
  49440=>"000100110",
  49441=>"110100100",
  49442=>"001000000",
  49443=>"000000101",
  49444=>"101111101",
  49445=>"100000000",
  49446=>"100100100",
  49447=>"000000000",
  49448=>"000000000",
  49449=>"101111111",
  49450=>"000000000",
  49451=>"011000111",
  49452=>"111110110",
  49453=>"000001011",
  49454=>"000111111",
  49455=>"110111010",
  49456=>"000000000",
  49457=>"111111111",
  49458=>"111110111",
  49459=>"000000110",
  49460=>"111101001",
  49461=>"000000010",
  49462=>"000000110",
  49463=>"111111111",
  49464=>"011011001",
  49465=>"000000000",
  49466=>"000000000",
  49467=>"111110111",
  49468=>"000000001",
  49469=>"011001111",
  49470=>"100100000",
  49471=>"110111111",
  49472=>"111111111",
  49473=>"110111000",
  49474=>"100110111",
  49475=>"000000000",
  49476=>"100101000",
  49477=>"000000000",
  49478=>"000101111",
  49479=>"001001011",
  49480=>"110000000",
  49481=>"000111111",
  49482=>"101111111",
  49483=>"111111111",
  49484=>"000000000",
  49485=>"000110111",
  49486=>"111111110",
  49487=>"101001001",
  49488=>"000000000",
  49489=>"100100111",
  49490=>"100000000",
  49491=>"000000000",
  49492=>"000110111",
  49493=>"011011011",
  49494=>"000000000",
  49495=>"111111111",
  49496=>"000000000",
  49497=>"000001001",
  49498=>"000000000",
  49499=>"000000000",
  49500=>"000000000",
  49501=>"000000100",
  49502=>"111101000",
  49503=>"111111000",
  49504=>"100100100",
  49505=>"111111111",
  49506=>"111111101",
  49507=>"000111111",
  49508=>"100011000",
  49509=>"100000010",
  49510=>"000000000",
  49511=>"000000000",
  49512=>"001001111",
  49513=>"010110111",
  49514=>"000000010",
  49515=>"111011001",
  49516=>"000001001",
  49517=>"011111100",
  49518=>"000101111",
  49519=>"101000000",
  49520=>"100100000",
  49521=>"000000100",
  49522=>"110111111",
  49523=>"000000000",
  49524=>"111111101",
  49525=>"111100000",
  49526=>"100000101",
  49527=>"000000101",
  49528=>"000000001",
  49529=>"111111111",
  49530=>"111111111",
  49531=>"111001000",
  49532=>"101110111",
  49533=>"110111111",
  49534=>"000000000",
  49535=>"000110111",
  49536=>"001000110",
  49537=>"000000000",
  49538=>"100100110",
  49539=>"111111111",
  49540=>"111111111",
  49541=>"111111111",
  49542=>"100000000",
  49543=>"001000111",
  49544=>"100100000",
  49545=>"000000011",
  49546=>"000000000",
  49547=>"111111011",
  49548=>"111111111",
  49549=>"000001011",
  49550=>"111111111",
  49551=>"000000010",
  49552=>"000000000",
  49553=>"111111111",
  49554=>"110111111",
  49555=>"011011000",
  49556=>"111001000",
  49557=>"000000000",
  49558=>"100100100",
  49559=>"111000000",
  49560=>"111111111",
  49561=>"100100000",
  49562=>"000000000",
  49563=>"111111010",
  49564=>"000000101",
  49565=>"011000000",
  49566=>"000000000",
  49567=>"000000000",
  49568=>"000100111",
  49569=>"000100000",
  49570=>"111111101",
  49571=>"111101111",
  49572=>"111111111",
  49573=>"111111111",
  49574=>"000000000",
  49575=>"000010010",
  49576=>"100100010",
  49577=>"001000000",
  49578=>"110100101",
  49579=>"000011000",
  49580=>"000000000",
  49581=>"111000111",
  49582=>"001011111",
  49583=>"111111111",
  49584=>"100100111",
  49585=>"000000000",
  49586=>"111111111",
  49587=>"100100010",
  49588=>"000000000",
  49589=>"111111111",
  49590=>"001000000",
  49591=>"111111111",
  49592=>"011000111",
  49593=>"100000000",
  49594=>"111111111",
  49595=>"100100100",
  49596=>"001000000",
  49597=>"110111110",
  49598=>"110000000",
  49599=>"100000100",
  49600=>"111000000",
  49601=>"001000111",
  49602=>"111011111",
  49603=>"000001111",
  49604=>"111111111",
  49605=>"111011111",
  49606=>"000000000",
  49607=>"111011011",
  49608=>"001000100",
  49609=>"000000111",
  49610=>"001000000",
  49611=>"000001000",
  49612=>"111111111",
  49613=>"000011010",
  49614=>"001001000",
  49615=>"111111111",
  49616=>"111000000",
  49617=>"111000000",
  49618=>"000100110",
  49619=>"111111111",
  49620=>"011000000",
  49621=>"111111111",
  49622=>"111111111",
  49623=>"000000110",
  49624=>"111111111",
  49625=>"111001000",
  49626=>"111111111",
  49627=>"111111101",
  49628=>"100111111",
  49629=>"111111111",
  49630=>"000110111",
  49631=>"000001011",
  49632=>"111001001",
  49633=>"000000000",
  49634=>"000101111",
  49635=>"111101000",
  49636=>"111000100",
  49637=>"111111111",
  49638=>"001111111",
  49639=>"000000000",
  49640=>"000000100",
  49641=>"111100111",
  49642=>"111111111",
  49643=>"111111111",
  49644=>"111111110",
  49645=>"111111111",
  49646=>"000000001",
  49647=>"000000000",
  49648=>"000000000",
  49649=>"111111110",
  49650=>"111111101",
  49651=>"000000000",
  49652=>"000000111",
  49653=>"000000000",
  49654=>"111111111",
  49655=>"010000000",
  49656=>"001000000",
  49657=>"000000000",
  49658=>"111111111",
  49659=>"111000000",
  49660=>"001001001",
  49661=>"100000111",
  49662=>"000000000",
  49663=>"000000000",
  49664=>"101100111",
  49665=>"111111111",
  49666=>"111111110",
  49667=>"111111110",
  49668=>"111111111",
  49669=>"110000000",
  49670=>"010010000",
  49671=>"000000000",
  49672=>"001001000",
  49673=>"000000100",
  49674=>"000000000",
  49675=>"110111101",
  49676=>"000010011",
  49677=>"111111110",
  49678=>"000000001",
  49679=>"010111010",
  49680=>"001001111",
  49681=>"000110110",
  49682=>"000000000",
  49683=>"111111110",
  49684=>"111111111",
  49685=>"101101100",
  49686=>"111111111",
  49687=>"101000111",
  49688=>"111110111",
  49689=>"100101100",
  49690=>"100000000",
  49691=>"100000000",
  49692=>"111111011",
  49693=>"111111000",
  49694=>"111111100",
  49695=>"111110010",
  49696=>"011011011",
  49697=>"000000000",
  49698=>"111111111",
  49699=>"000101111",
  49700=>"000010111",
  49701=>"111111111",
  49702=>"100100101",
  49703=>"110111001",
  49704=>"000111110",
  49705=>"111111011",
  49706=>"000000110",
  49707=>"000000011",
  49708=>"000000000",
  49709=>"111100100",
  49710=>"111111111",
  49711=>"111111111",
  49712=>"111001111",
  49713=>"010111011",
  49714=>"111100000",
  49715=>"011101111",
  49716=>"101101111",
  49717=>"101001000",
  49718=>"111111110",
  49719=>"111011011",
  49720=>"001011000",
  49721=>"000000111",
  49722=>"111111111",
  49723=>"111111100",
  49724=>"000000111",
  49725=>"000000100",
  49726=>"001000000",
  49727=>"111001000",
  49728=>"000000000",
  49729=>"000110000",
  49730=>"000000000",
  49731=>"100100110",
  49732=>"111111110",
  49733=>"001111111",
  49734=>"000000000",
  49735=>"101101000",
  49736=>"100101111",
  49737=>"111001111",
  49738=>"000000000",
  49739=>"000000111",
  49740=>"001000000",
  49741=>"000000000",
  49742=>"001100010",
  49743=>"000000110",
  49744=>"111001000",
  49745=>"101000100",
  49746=>"000000000",
  49747=>"000101111",
  49748=>"111101111",
  49749=>"000000000",
  49750=>"111111001",
  49751=>"000000000",
  49752=>"111111000",
  49753=>"111000000",
  49754=>"000000000",
  49755=>"110000000",
  49756=>"111011000",
  49757=>"111000100",
  49758=>"000000111",
  49759=>"011001011",
  49760=>"001111001",
  49761=>"001000001",
  49762=>"000100111",
  49763=>"111000000",
  49764=>"111001000",
  49765=>"111111101",
  49766=>"000000111",
  49767=>"100000011",
  49768=>"000000000",
  49769=>"111110111",
  49770=>"000010011",
  49771=>"011111111",
  49772=>"000000110",
  49773=>"000000000",
  49774=>"000000000",
  49775=>"000000000",
  49776=>"000000000",
  49777=>"001111000",
  49778=>"010010000",
  49779=>"000000110",
  49780=>"001111111",
  49781=>"000000000",
  49782=>"000000000",
  49783=>"000000000",
  49784=>"010111001",
  49785=>"000000000",
  49786=>"101110111",
  49787=>"000100100",
  49788=>"110110110",
  49789=>"000110111",
  49790=>"100100100",
  49791=>"000001001",
  49792=>"000000011",
  49793=>"111111111",
  49794=>"001000110",
  49795=>"001111101",
  49796=>"111100111",
  49797=>"111000100",
  49798=>"001011001",
  49799=>"000000100",
  49800=>"111101111",
  49801=>"000000000",
  49802=>"000111111",
  49803=>"001000001",
  49804=>"111111111",
  49805=>"111111000",
  49806=>"111111000",
  49807=>"000000000",
  49808=>"000000100",
  49809=>"001010110",
  49810=>"001000100",
  49811=>"111111111",
  49812=>"111111011",
  49813=>"111110000",
  49814=>"101000000",
  49815=>"000000111",
  49816=>"000000001",
  49817=>"000000111",
  49818=>"000000000",
  49819=>"111110000",
  49820=>"111111001",
  49821=>"000000000",
  49822=>"111000100",
  49823=>"001001000",
  49824=>"111111011",
  49825=>"000100000",
  49826=>"111100000",
  49827=>"001000000",
  49828=>"010000110",
  49829=>"111110010",
  49830=>"111000100",
  49831=>"110100000",
  49832=>"100111000",
  49833=>"000000000",
  49834=>"001111111",
  49835=>"101100100",
  49836=>"111111111",
  49837=>"100100110",
  49838=>"111111001",
  49839=>"111111000",
  49840=>"000000000",
  49841=>"000100000",
  49842=>"010010010",
  49843=>"111000000",
  49844=>"111111010",
  49845=>"000000001",
  49846=>"000000010",
  49847=>"000010111",
  49848=>"111000001",
  49849=>"111001111",
  49850=>"010110011",
  49851=>"010011011",
  49852=>"011000000",
  49853=>"101000011",
  49854=>"000110110",
  49855=>"111110000",
  49856=>"111111111",
  49857=>"000000111",
  49858=>"111111011",
  49859=>"000000000",
  49860=>"000000111",
  49861=>"000000000",
  49862=>"000000000",
  49863=>"111111011",
  49864=>"111111011",
  49865=>"001111000",
  49866=>"000000000",
  49867=>"011111111",
  49868=>"000000000",
  49869=>"001000000",
  49870=>"111111111",
  49871=>"010010000",
  49872=>"111110110",
  49873=>"111111000",
  49874=>"011000000",
  49875=>"100000001",
  49876=>"001111111",
  49877=>"111110110",
  49878=>"111111110",
  49879=>"000000001",
  49880=>"111111100",
  49881=>"000000000",
  49882=>"100101111",
  49883=>"000111011",
  49884=>"001000000",
  49885=>"001000000",
  49886=>"111111111",
  49887=>"011111011",
  49888=>"000000000",
  49889=>"111111111",
  49890=>"000000010",
  49891=>"000000000",
  49892=>"110010000",
  49893=>"000000000",
  49894=>"111111001",
  49895=>"111111101",
  49896=>"111111111",
  49897=>"000000101",
  49898=>"000000111",
  49899=>"100110111",
  49900=>"111111111",
  49901=>"000000111",
  49902=>"111111111",
  49903=>"111000000",
  49904=>"111111000",
  49905=>"011110110",
  49906=>"000000011",
  49907=>"000000001",
  49908=>"110011011",
  49909=>"111111100",
  49910=>"100110100",
  49911=>"000101111",
  49912=>"111111111",
  49913=>"001000000",
  49914=>"000000000",
  49915=>"111111111",
  49916=>"100000000",
  49917=>"000000000",
  49918=>"111111000",
  49919=>"000011110",
  49920=>"000000001",
  49921=>"101001001",
  49922=>"111111110",
  49923=>"111111000",
  49924=>"000111111",
  49925=>"001110111",
  49926=>"111111111",
  49927=>"101011000",
  49928=>"111111111",
  49929=>"000000000",
  49930=>"011011011",
  49931=>"000000001",
  49932=>"000000110",
  49933=>"111111111",
  49934=>"111111111",
  49935=>"000111111",
  49936=>"011000001",
  49937=>"000101000",
  49938=>"000000100",
  49939=>"000000000",
  49940=>"000000000",
  49941=>"000011000",
  49942=>"100100100",
  49943=>"111101000",
  49944=>"110111111",
  49945=>"111111111",
  49946=>"000000001",
  49947=>"000000000",
  49948=>"010010000",
  49949=>"011011000",
  49950=>"000000000",
  49951=>"000000101",
  49952=>"011011000",
  49953=>"111101111",
  49954=>"000000000",
  49955=>"111111110",
  49956=>"011111011",
  49957=>"110001111",
  49958=>"000001000",
  49959=>"000000101",
  49960=>"111000010",
  49961=>"010111011",
  49962=>"111001001",
  49963=>"011101100",
  49964=>"111111000",
  49965=>"000000001",
  49966=>"000000010",
  49967=>"111111111",
  49968=>"000011111",
  49969=>"111000000",
  49970=>"100000111",
  49971=>"001100111",
  49972=>"111101111",
  49973=>"000000000",
  49974=>"111111001",
  49975=>"000000000",
  49976=>"000000110",
  49977=>"111111111",
  49978=>"010010101",
  49979=>"111111111",
  49980=>"000000001",
  49981=>"111111100",
  49982=>"001011011",
  49983=>"000000000",
  49984=>"000100000",
  49985=>"111100000",
  49986=>"000000001",
  49987=>"000100100",
  49988=>"111111111",
  49989=>"000000001",
  49990=>"111000111",
  49991=>"100111111",
  49992=>"111111001",
  49993=>"000001011",
  49994=>"111101001",
  49995=>"001001001",
  49996=>"111111000",
  49997=>"000000000",
  49998=>"000000000",
  49999=>"101101110",
  50000=>"001001001",
  50001=>"000000110",
  50002=>"111111111",
  50003=>"000000001",
  50004=>"001101000",
  50005=>"001011011",
  50006=>"111111011",
  50007=>"111111111",
  50008=>"000000111",
  50009=>"000000111",
  50010=>"000001011",
  50011=>"111111111",
  50012=>"001000000",
  50013=>"000000111",
  50014=>"000000000",
  50015=>"001111000",
  50016=>"110000011",
  50017=>"000000000",
  50018=>"111001000",
  50019=>"000000111",
  50020=>"000000000",
  50021=>"000001101",
  50022=>"111101101",
  50023=>"001001101",
  50024=>"100110110",
  50025=>"000111111",
  50026=>"000000000",
  50027=>"000111111",
  50028=>"010111111",
  50029=>"001010011",
  50030=>"111111010",
  50031=>"000000000",
  50032=>"111011010",
  50033=>"000011010",
  50034=>"111000000",
  50035=>"000000000",
  50036=>"000010000",
  50037=>"010110000",
  50038=>"001111101",
  50039=>"000000100",
  50040=>"101000000",
  50041=>"111111000",
  50042=>"000000000",
  50043=>"111111011",
  50044=>"000000000",
  50045=>"111111111",
  50046=>"011111100",
  50047=>"000000000",
  50048=>"000011110",
  50049=>"111101110",
  50050=>"111011000",
  50051=>"000000100",
  50052=>"111000000",
  50053=>"110100110",
  50054=>"010110111",
  50055=>"000000000",
  50056=>"000000111",
  50057=>"001001011",
  50058=>"111100111",
  50059=>"100100111",
  50060=>"000111111",
  50061=>"111101100",
  50062=>"111111111",
  50063=>"011111001",
  50064=>"001001001",
  50065=>"111111110",
  50066=>"011000000",
  50067=>"011011011",
  50068=>"011111111",
  50069=>"000000000",
  50070=>"000001000",
  50071=>"100100000",
  50072=>"001001000",
  50073=>"000000000",
  50074=>"000000111",
  50075=>"111111000",
  50076=>"000100101",
  50077=>"000000000",
  50078=>"011111111",
  50079=>"111111111",
  50080=>"001000000",
  50081=>"000000111",
  50082=>"111101111",
  50083=>"111111000",
  50084=>"001101111",
  50085=>"001001111",
  50086=>"111000000",
  50087=>"111011111",
  50088=>"000001000",
  50089=>"000000111",
  50090=>"111111111",
  50091=>"100001100",
  50092=>"111000000",
  50093=>"011111000",
  50094=>"101111111",
  50095=>"111111000",
  50096=>"000000000",
  50097=>"000000000",
  50098=>"111011000",
  50099=>"000000000",
  50100=>"111011001",
  50101=>"100110111",
  50102=>"111111111",
  50103=>"111111111",
  50104=>"000000000",
  50105=>"111111111",
  50106=>"110111111",
  50107=>"000000000",
  50108=>"101111000",
  50109=>"000000100",
  50110=>"111100100",
  50111=>"000000100",
  50112=>"111010000",
  50113=>"001001000",
  50114=>"000000000",
  50115=>"000000000",
  50116=>"000000000",
  50117=>"001000110",
  50118=>"000111000",
  50119=>"001101100",
  50120=>"000000000",
  50121=>"111000000",
  50122=>"000100101",
  50123=>"000111111",
  50124=>"000000000",
  50125=>"101100000",
  50126=>"101100110",
  50127=>"001000000",
  50128=>"011000111",
  50129=>"000000000",
  50130=>"000010111",
  50131=>"111111111",
  50132=>"111111011",
  50133=>"101111011",
  50134=>"000000000",
  50135=>"000110111",
  50136=>"000000111",
  50137=>"111100111",
  50138=>"000000011",
  50139=>"111111000",
  50140=>"011111111",
  50141=>"000000000",
  50142=>"100000000",
  50143=>"011011001",
  50144=>"101000000",
  50145=>"111100000",
  50146=>"011011010",
  50147=>"111111011",
  50148=>"000000111",
  50149=>"000000100",
  50150=>"110000110",
  50151=>"000000000",
  50152=>"101101000",
  50153=>"111111111",
  50154=>"111101111",
  50155=>"000101001",
  50156=>"100000111",
  50157=>"001001001",
  50158=>"111100000",
  50159=>"111111111",
  50160=>"000000111",
  50161=>"111111111",
  50162=>"000111111",
  50163=>"101100110",
  50164=>"001000000",
  50165=>"000000011",
  50166=>"100101111",
  50167=>"110111111",
  50168=>"001001000",
  50169=>"000000000",
  50170=>"000000001",
  50171=>"000000000",
  50172=>"000000000",
  50173=>"111111011",
  50174=>"011110110",
  50175=>"000000111",
  50176=>"111111011",
  50177=>"011111011",
  50178=>"000000000",
  50179=>"111000111",
  50180=>"110000000",
  50181=>"000110110",
  50182=>"000111110",
  50183=>"111111011",
  50184=>"001000011",
  50185=>"011001000",
  50186=>"000000001",
  50187=>"111110110",
  50188=>"110110110",
  50189=>"010011000",
  50190=>"000000101",
  50191=>"000000110",
  50192=>"110100111",
  50193=>"111110010",
  50194=>"110111000",
  50195=>"101100111",
  50196=>"000001111",
  50197=>"111111111",
  50198=>"000111100",
  50199=>"110111111",
  50200=>"000100000",
  50201=>"011011100",
  50202=>"100101101",
  50203=>"111101111",
  50204=>"111111111",
  50205=>"000110111",
  50206=>"000100001",
  50207=>"000000001",
  50208=>"111111111",
  50209=>"001011111",
  50210=>"010000111",
  50211=>"100000100",
  50212=>"100000000",
  50213=>"111110111",
  50214=>"000000000",
  50215=>"000000111",
  50216=>"111111111",
  50217=>"111001000",
  50218=>"000000101",
  50219=>"000001000",
  50220=>"110111000",
  50221=>"000000001",
  50222=>"001000000",
  50223=>"000000111",
  50224=>"110110111",
  50225=>"111000000",
  50226=>"001001100",
  50227=>"101100000",
  50228=>"100000000",
  50229=>"000100110",
  50230=>"000000100",
  50231=>"000110111",
  50232=>"000000000",
  50233=>"110110010",
  50234=>"000111101",
  50235=>"001000000",
  50236=>"101101101",
  50237=>"000000000",
  50238=>"000100111",
  50239=>"000001111",
  50240=>"000110110",
  50241=>"111111010",
  50242=>"010010000",
  50243=>"011111111",
  50244=>"000001111",
  50245=>"001001001",
  50246=>"111000100",
  50247=>"000001000",
  50248=>"001001001",
  50249=>"111111111",
  50250=>"001001111",
  50251=>"001000000",
  50252=>"110110000",
  50253=>"110010000",
  50254=>"011001000",
  50255=>"001001111",
  50256=>"000000000",
  50257=>"110100000",
  50258=>"110110101",
  50259=>"100101001",
  50260=>"111111111",
  50261=>"110111000",
  50262=>"111110010",
  50263=>"000000000",
  50264=>"110110111",
  50265=>"111101000",
  50266=>"000011111",
  50267=>"000000000",
  50268=>"111111111",
  50269=>"111111111",
  50270=>"001001001",
  50271=>"000010110",
  50272=>"000100000",
  50273=>"000000100",
  50274=>"111111111",
  50275=>"010000000",
  50276=>"110111001",
  50277=>"111000000",
  50278=>"000000000",
  50279=>"100111110",
  50280=>"111111111",
  50281=>"111111111",
  50282=>"011010000",
  50283=>"111110111",
  50284=>"001011111",
  50285=>"000001101",
  50286=>"000000000",
  50287=>"001100000",
  50288=>"110100100",
  50289=>"000101111",
  50290=>"010010001",
  50291=>"101101000",
  50292=>"011011000",
  50293=>"000000100",
  50294=>"000000000",
  50295=>"001000000",
  50296=>"111001000",
  50297=>"111111100",
  50298=>"000000000",
  50299=>"000000000",
  50300=>"000000000",
  50301=>"010011000",
  50302=>"010000010",
  50303=>"000000001",
  50304=>"000000001",
  50305=>"111101111",
  50306=>"111000000",
  50307=>"111010000",
  50308=>"000100000",
  50309=>"000000000",
  50310=>"111101000",
  50311=>"000100100",
  50312=>"111111001",
  50313=>"111111111",
  50314=>"011100110",
  50315=>"001001111",
  50316=>"101111111",
  50317=>"111111111",
  50318=>"100110100",
  50319=>"111111111",
  50320=>"000000001",
  50321=>"100000001",
  50322=>"010010111",
  50323=>"000000111",
  50324=>"000000000",
  50325=>"110011011",
  50326=>"001001111",
  50327=>"000000000",
  50328=>"001001111",
  50329=>"101100111",
  50330=>"000000000",
  50331=>"101000000",
  50332=>"110000000",
  50333=>"111111100",
  50334=>"111111101",
  50335=>"000000000",
  50336=>"111111000",
  50337=>"010010000",
  50338=>"010111111",
  50339=>"000000111",
  50340=>"110111101",
  50341=>"000010000",
  50342=>"111111100",
  50343=>"011011010",
  50344=>"000011110",
  50345=>"110100000",
  50346=>"001001111",
  50347=>"000000100",
  50348=>"110100000",
  50349=>"100110011",
  50350=>"000100111",
  50351=>"000111111",
  50352=>"111111111",
  50353=>"000010111",
  50354=>"110111000",
  50355=>"111111111",
  50356=>"000000000",
  50357=>"000011111",
  50358=>"000000000",
  50359=>"001101111",
  50360=>"000001111",
  50361=>"111111110",
  50362=>"111111001",
  50363=>"111000000",
  50364=>"000000000",
  50365=>"110110111",
  50366=>"001001011",
  50367=>"000000000",
  50368=>"111111111",
  50369=>"000000000",
  50370=>"110110010",
  50371=>"110110010",
  50372=>"111110111",
  50373=>"000000101",
  50374=>"111111101",
  50375=>"111111000",
  50376=>"000111111",
  50377=>"110110110",
  50378=>"110110100",
  50379=>"000111000",
  50380=>"111110110",
  50381=>"011011011",
  50382=>"000010001",
  50383=>"111010111",
  50384=>"000011111",
  50385=>"000000111",
  50386=>"000000000",
  50387=>"000000000",
  50388=>"000001111",
  50389=>"111100000",
  50390=>"001100000",
  50391=>"111111110",
  50392=>"000000000",
  50393=>"000000001",
  50394=>"111111111",
  50395=>"110110110",
  50396=>"001001000",
  50397=>"000000001",
  50398=>"100110000",
  50399=>"000000000",
  50400=>"000000111",
  50401=>"001001111",
  50402=>"111111101",
  50403=>"111010011",
  50404=>"000000000",
  50405=>"000000000",
  50406=>"000000100",
  50407=>"000000000",
  50408=>"001111111",
  50409=>"111111111",
  50410=>"000000000",
  50411=>"111101111",
  50412=>"000100101",
  50413=>"011001000",
  50414=>"101001101",
  50415=>"000000000",
  50416=>"000000001",
  50417=>"110111000",
  50418=>"111101101",
  50419=>"000001001",
  50420=>"011001101",
  50421=>"000000000",
  50422=>"111111000",
  50423=>"111111011",
  50424=>"111111111",
  50425=>"111101000",
  50426=>"000000010",
  50427=>"001001001",
  50428=>"011011011",
  50429=>"111111111",
  50430=>"001001000",
  50431=>"000111010",
  50432=>"000001111",
  50433=>"111011010",
  50434=>"100100110",
  50435=>"110111111",
  50436=>"101111111",
  50437=>"000110000",
  50438=>"000110000",
  50439=>"110111000",
  50440=>"000100110",
  50441=>"111100100",
  50442=>"000110111",
  50443=>"010000011",
  50444=>"111110110",
  50445=>"001011111",
  50446=>"000000000",
  50447=>"000000111",
  50448=>"000001001",
  50449=>"000000000",
  50450=>"001001101",
  50451=>"110010010",
  50452=>"100100001",
  50453=>"000100111",
  50454=>"001001110",
  50455=>"000000000",
  50456=>"110110110",
  50457=>"101001001",
  50458=>"000000111",
  50459=>"000011011",
  50460=>"000100000",
  50461=>"000000000",
  50462=>"000000000",
  50463=>"000011111",
  50464=>"011011000",
  50465=>"001000000",
  50466=>"111111010",
  50467=>"000111111",
  50468=>"111111001",
  50469=>"101101111",
  50470=>"111100100",
  50471=>"001001001",
  50472=>"111000000",
  50473=>"111111111",
  50474=>"010110011",
  50475=>"000001000",
  50476=>"111010000",
  50477=>"011000000",
  50478=>"000000000",
  50479=>"000000000",
  50480=>"111111011",
  50481=>"000000101",
  50482=>"111001001",
  50483=>"111111111",
  50484=>"000000000",
  50485=>"100000010",
  50486=>"110110111",
  50487=>"000000000",
  50488=>"000000000",
  50489=>"000001110",
  50490=>"001000100",
  50491=>"001011001",
  50492=>"000000000",
  50493=>"010111000",
  50494=>"111110100",
  50495=>"000000100",
  50496=>"111111101",
  50497=>"000000000",
  50498=>"111111001",
  50499=>"001000100",
  50500=>"000000000",
  50501=>"110011001",
  50502=>"001001000",
  50503=>"000100000",
  50504=>"110000000",
  50505=>"111101011",
  50506=>"111110010",
  50507=>"100100110",
  50508=>"000110111",
  50509=>"111111100",
  50510=>"111111111",
  50511=>"001001000",
  50512=>"000111111",
  50513=>"000010110",
  50514=>"010010100",
  50515=>"111001011",
  50516=>"101000000",
  50517=>"011001001",
  50518=>"111000000",
  50519=>"000000100",
  50520=>"100001001",
  50521=>"011001001",
  50522=>"000000000",
  50523=>"101001111",
  50524=>"011000000",
  50525=>"000100111",
  50526=>"001011000",
  50527=>"001000100",
  50528=>"001000001",
  50529=>"011101111",
  50530=>"000000110",
  50531=>"111001111",
  50532=>"111100000",
  50533=>"000000001",
  50534=>"000000000",
  50535=>"010000100",
  50536=>"011000000",
  50537=>"111110100",
  50538=>"000000000",
  50539=>"111110110",
  50540=>"010010000",
  50541=>"000000001",
  50542=>"001001000",
  50543=>"100000000",
  50544=>"001101000",
  50545=>"011011001",
  50546=>"001111000",
  50547=>"011011111",
  50548=>"100111011",
  50549=>"000000000",
  50550=>"000000000",
  50551=>"000000100",
  50552=>"111111001",
  50553=>"111100000",
  50554=>"000000000",
  50555=>"111111111",
  50556=>"000111111",
  50557=>"000000000",
  50558=>"110000000",
  50559=>"111111111",
  50560=>"111111111",
  50561=>"011111111",
  50562=>"000000100",
  50563=>"000001111",
  50564=>"000000000",
  50565=>"000000111",
  50566=>"000010111",
  50567=>"001011001",
  50568=>"001000001",
  50569=>"000000000",
  50570=>"111111111",
  50571=>"010111111",
  50572=>"111111111",
  50573=>"111111011",
  50574=>"000010011",
  50575=>"000000000",
  50576=>"011110111",
  50577=>"100010111",
  50578=>"110110011",
  50579=>"000000000",
  50580=>"001001111",
  50581=>"001001001",
  50582=>"110110010",
  50583=>"110111000",
  50584=>"111111111",
  50585=>"110000111",
  50586=>"000000001",
  50587=>"000100111",
  50588=>"111011011",
  50589=>"100000000",
  50590=>"001001001",
  50591=>"000010010",
  50592=>"000010000",
  50593=>"100100100",
  50594=>"010110111",
  50595=>"001001100",
  50596=>"110111111",
  50597=>"111111111",
  50598=>"101000000",
  50599=>"111000001",
  50600=>"000000000",
  50601=>"011001111",
  50602=>"000000111",
  50603=>"000000000",
  50604=>"111111100",
  50605=>"111110111",
  50606=>"111001000",
  50607=>"110100100",
  50608=>"101100100",
  50609=>"000000000",
  50610=>"111000000",
  50611=>"011000000",
  50612=>"000100000",
  50613=>"011111111",
  50614=>"111111011",
  50615=>"111111111",
  50616=>"010010000",
  50617=>"110100000",
  50618=>"011011000",
  50619=>"010110011",
  50620=>"000010110",
  50621=>"000000000",
  50622=>"001000001",
  50623=>"000000000",
  50624=>"001001001",
  50625=>"101101110",
  50626=>"001000000",
  50627=>"111001000",
  50628=>"100110111",
  50629=>"000000001",
  50630=>"000000010",
  50631=>"000111111",
  50632=>"001000000",
  50633=>"100001111",
  50634=>"001001001",
  50635=>"001001001",
  50636=>"010000000",
  50637=>"000001111",
  50638=>"010000000",
  50639=>"001111111",
  50640=>"111111000",
  50641=>"111101000",
  50642=>"100111111",
  50643=>"000001000",
  50644=>"101111111",
  50645=>"101000000",
  50646=>"111111110",
  50647=>"111111000",
  50648=>"100111001",
  50649=>"000011111",
  50650=>"000101101",
  50651=>"111000000",
  50652=>"100110110",
  50653=>"000001001",
  50654=>"100000010",
  50655=>"110000000",
  50656=>"100101100",
  50657=>"000000000",
  50658=>"101111111",
  50659=>"111111001",
  50660=>"000100111",
  50661=>"110111011",
  50662=>"101101111",
  50663=>"000000000",
  50664=>"000000000",
  50665=>"111001010",
  50666=>"010110100",
  50667=>"000000000",
  50668=>"001001111",
  50669=>"001010000",
  50670=>"001000101",
  50671=>"000000001",
  50672=>"000111111",
  50673=>"110010000",
  50674=>"111111111",
  50675=>"000100000",
  50676=>"110110111",
  50677=>"000000000",
  50678=>"111111111",
  50679=>"001000000",
  50680=>"011000110",
  50681=>"110010000",
  50682=>"011111111",
  50683=>"001001000",
  50684=>"110100000",
  50685=>"111111111",
  50686=>"111010010",
  50687=>"000000000",
  50688=>"110111011",
  50689=>"100000000",
  50690=>"111001100",
  50691=>"000000100",
  50692=>"000111010",
  50693=>"000000000",
  50694=>"000000000",
  50695=>"111111111",
  50696=>"000000000",
  50697=>"111011011",
  50698=>"000000000",
  50699=>"111111111",
  50700=>"111001001",
  50701=>"000110111",
  50702=>"011011010",
  50703=>"111110000",
  50704=>"100000011",
  50705=>"000000101",
  50706=>"000000000",
  50707=>"111101011",
  50708=>"001100111",
  50709=>"000000111",
  50710=>"110000111",
  50711=>"000110101",
  50712=>"001011111",
  50713=>"110111011",
  50714=>"000000000",
  50715=>"110010001",
  50716=>"001111111",
  50717=>"100111111",
  50718=>"111111001",
  50719=>"000001001",
  50720=>"111111001",
  50721=>"000000100",
  50722=>"100000000",
  50723=>"010001001",
  50724=>"000000000",
  50725=>"100010110",
  50726=>"111000001",
  50727=>"011001000",
  50728=>"000111111",
  50729=>"011011000",
  50730=>"001000000",
  50731=>"111000000",
  50732=>"101000100",
  50733=>"110100000",
  50734=>"000001001",
  50735=>"111111101",
  50736=>"111111001",
  50737=>"110100000",
  50738=>"100110000",
  50739=>"010110100",
  50740=>"000111111",
  50741=>"111011000",
  50742=>"101000110",
  50743=>"000010111",
  50744=>"011101101",
  50745=>"001001001",
  50746=>"000000111",
  50747=>"100110111",
  50748=>"000000000",
  50749=>"111000001",
  50750=>"111000000",
  50751=>"001000000",
  50752=>"001111111",
  50753=>"001001101",
  50754=>"000111111",
  50755=>"000000111",
  50756=>"000000110",
  50757=>"000001111",
  50758=>"000000101",
  50759=>"111100111",
  50760=>"111111111",
  50761=>"111111011",
  50762=>"111100110",
  50763=>"000011111",
  50764=>"110110001",
  50765=>"000000111",
  50766=>"000000111",
  50767=>"011111110",
  50768=>"111101111",
  50769=>"000100100",
  50770=>"110100000",
  50771=>"110111110",
  50772=>"000000111",
  50773=>"001011111",
  50774=>"011011101",
  50775=>"000111111",
  50776=>"000110110",
  50777=>"111111111",
  50778=>"101111111",
  50779=>"000000010",
  50780=>"010000000",
  50781=>"111001000",
  50782=>"001000000",
  50783=>"000111111",
  50784=>"000000000",
  50785=>"011111111",
  50786=>"001111001",
  50787=>"011111111",
  50788=>"000111010",
  50789=>"111111000",
  50790=>"000110000",
  50791=>"111000100",
  50792=>"000111011",
  50793=>"000000000",
  50794=>"000100111",
  50795=>"000000000",
  50796=>"001011111",
  50797=>"001001111",
  50798=>"000000111",
  50799=>"101111000",
  50800=>"000000010",
  50801=>"111111010",
  50802=>"000011000",
  50803=>"111111111",
  50804=>"011000000",
  50805=>"000111111",
  50806=>"111000000",
  50807=>"000000111",
  50808=>"000000011",
  50809=>"111111000",
  50810=>"000000001",
  50811=>"000000111",
  50812=>"110111000",
  50813=>"011111111",
  50814=>"000001000",
  50815=>"111101001",
  50816=>"101111101",
  50817=>"100110111",
  50818=>"000000111",
  50819=>"011011011",
  50820=>"001101111",
  50821=>"000000100",
  50822=>"111111000",
  50823=>"001001001",
  50824=>"000000100",
  50825=>"000000111",
  50826=>"111011011",
  50827=>"011110011",
  50828=>"000000000",
  50829=>"000000000",
  50830=>"100100111",
  50831=>"000010010",
  50832=>"010111111",
  50833=>"100110110",
  50834=>"000000001",
  50835=>"101000110",
  50836=>"111111000",
  50837=>"000000000",
  50838=>"000000111",
  50839=>"101101111",
  50840=>"000000111",
  50841=>"111111111",
  50842=>"111100000",
  50843=>"000011011",
  50844=>"000000000",
  50845=>"000000001",
  50846=>"111111111",
  50847=>"111100111",
  50848=>"000000000",
  50849=>"110100111",
  50850=>"000000000",
  50851=>"000000000",
  50852=>"111000000",
  50853=>"010000000",
  50854=>"010000010",
  50855=>"001011011",
  50856=>"011011111",
  50857=>"000000011",
  50858=>"111000000",
  50859=>"001101000",
  50860=>"100100111",
  50861=>"000001011",
  50862=>"011000000",
  50863=>"100100101",
  50864=>"000000100",
  50865=>"011000000",
  50866=>"111111111",
  50867=>"000011000",
  50868=>"111111001",
  50869=>"111000101",
  50870=>"010100110",
  50871=>"111001011",
  50872=>"001011110",
  50873=>"111111111",
  50874=>"110000001",
  50875=>"110100111",
  50876=>"000000111",
  50877=>"000000111",
  50878=>"000101111",
  50879=>"110000000",
  50880=>"000000100",
  50881=>"001011111",
  50882=>"111110110",
  50883=>"110000000",
  50884=>"101100111",
  50885=>"111111111",
  50886=>"110111111",
  50887=>"111111101",
  50888=>"000000111",
  50889=>"111111101",
  50890=>"010011010",
  50891=>"111111000",
  50892=>"010010000",
  50893=>"110110100",
  50894=>"010011111",
  50895=>"000111011",
  50896=>"001101101",
  50897=>"001101001",
  50898=>"000000111",
  50899=>"011111101",
  50900=>"111111111",
  50901=>"110111111",
  50902=>"000000100",
  50903=>"000000100",
  50904=>"000000000",
  50905=>"011111010",
  50906=>"100111111",
  50907=>"011000111",
  50908=>"110111111",
  50909=>"001100000",
  50910=>"111111011",
  50911=>"110000000",
  50912=>"111111010",
  50913=>"111110100",
  50914=>"000101101",
  50915=>"011011001",
  50916=>"001111110",
  50917=>"100000010",
  50918=>"001011001",
  50919=>"111011001",
  50920=>"111111011",
  50921=>"100101101",
  50922=>"111011001",
  50923=>"000000000",
  50924=>"000000000",
  50925=>"111101100",
  50926=>"111110111",
  50927=>"000000000",
  50928=>"000000000",
  50929=>"001000000",
  50930=>"101111111",
  50931=>"111001000",
  50932=>"111111111",
  50933=>"000001101",
  50934=>"000000000",
  50935=>"101000000",
  50936=>"111111110",
  50937=>"011110100",
  50938=>"000000111",
  50939=>"111111101",
  50940=>"000110110",
  50941=>"111011011",
  50942=>"111000111",
  50943=>"111111000",
  50944=>"000001011",
  50945=>"010010011",
  50946=>"000001111",
  50947=>"000000011",
  50948=>"001000000",
  50949=>"111000010",
  50950=>"100111001",
  50951=>"111000101",
  50952=>"011011111",
  50953=>"010000000",
  50954=>"000000100",
  50955=>"111001111",
  50956=>"100000110",
  50957=>"100000001",
  50958=>"011001000",
  50959=>"001001001",
  50960=>"000111111",
  50961=>"000000010",
  50962=>"001111111",
  50963=>"000000000",
  50964=>"000111010",
  50965=>"000000000",
  50966=>"000011000",
  50967=>"001000000",
  50968=>"110000000",
  50969=>"101111111",
  50970=>"111111111",
  50971=>"000000100",
  50972=>"111111110",
  50973=>"001001000",
  50974=>"111111111",
  50975=>"000000000",
  50976=>"110110001",
  50977=>"111111111",
  50978=>"110111100",
  50979=>"111101000",
  50980=>"100100100",
  50981=>"000111111",
  50982=>"011001000",
  50983=>"111100000",
  50984=>"111101101",
  50985=>"011010110",
  50986=>"000000000",
  50987=>"111110110",
  50988=>"011000011",
  50989=>"011010110",
  50990=>"001111000",
  50991=>"000111011",
  50992=>"001110111",
  50993=>"001001111",
  50994=>"000000111",
  50995=>"111110001",
  50996=>"010000100",
  50997=>"000000011",
  50998=>"000000000",
  50999=>"100000000",
  51000=>"011000111",
  51001=>"101100000",
  51002=>"000000111",
  51003=>"101000101",
  51004=>"011011011",
  51005=>"110000000",
  51006=>"111111111",
  51007=>"110000100",
  51008=>"011111011",
  51009=>"111001001",
  51010=>"010110000",
  51011=>"000000011",
  51012=>"000000111",
  51013=>"000011001",
  51014=>"000000000",
  51015=>"000000000",
  51016=>"000000111",
  51017=>"000000101",
  51018=>"101001011",
  51019=>"111000000",
  51020=>"000000100",
  51021=>"001101000",
  51022=>"000000000",
  51023=>"000000110",
  51024=>"000100000",
  51025=>"000101101",
  51026=>"000000000",
  51027=>"000000111",
  51028=>"110000000",
  51029=>"111111000",
  51030=>"111111111",
  51031=>"100000001",
  51032=>"111111111",
  51033=>"111101000",
  51034=>"000111111",
  51035=>"000000101",
  51036=>"101000000",
  51037=>"000000111",
  51038=>"110000010",
  51039=>"001000000",
  51040=>"001101101",
  51041=>"101000000",
  51042=>"111110000",
  51043=>"000000000",
  51044=>"110110010",
  51045=>"001101001",
  51046=>"000000111",
  51047=>"000000001",
  51048=>"111110000",
  51049=>"000001001",
  51050=>"000110110",
  51051=>"111111101",
  51052=>"011011011",
  51053=>"111000000",
  51054=>"111000000",
  51055=>"000101000",
  51056=>"111111111",
  51057=>"011000000",
  51058=>"111000001",
  51059=>"111011000",
  51060=>"001100111",
  51061=>"011111111",
  51062=>"000001101",
  51063=>"100100001",
  51064=>"000000100",
  51065=>"001101111",
  51066=>"000000111",
  51067=>"111000000",
  51068=>"100000000",
  51069=>"111111111",
  51070=>"000000111",
  51071=>"111000001",
  51072=>"011111110",
  51073=>"111111110",
  51074=>"000110110",
  51075=>"000100111",
  51076=>"110000111",
  51077=>"111111010",
  51078=>"000000011",
  51079=>"111111110",
  51080=>"000000000",
  51081=>"111011011",
  51082=>"000000101",
  51083=>"000000111",
  51084=>"100111000",
  51085=>"111010000",
  51086=>"000011111",
  51087=>"111111111",
  51088=>"100000000",
  51089=>"000110111",
  51090=>"000101111",
  51091=>"110110000",
  51092=>"111000000",
  51093=>"111111110",
  51094=>"111111001",
  51095=>"110100110",
  51096=>"000101111",
  51097=>"101111100",
  51098=>"111111111",
  51099=>"111111011",
  51100=>"111111000",
  51101=>"110100000",
  51102=>"000111010",
  51103=>"111001000",
  51104=>"100000000",
  51105=>"111100000",
  51106=>"111101101",
  51107=>"000000000",
  51108=>"100101101",
  51109=>"100111111",
  51110=>"000111001",
  51111=>"101111010",
  51112=>"100000111",
  51113=>"000001000",
  51114=>"000010111",
  51115=>"111111000",
  51116=>"000000000",
  51117=>"000000011",
  51118=>"111100001",
  51119=>"011111111",
  51120=>"000000000",
  51121=>"000100111",
  51122=>"111111111",
  51123=>"111001001",
  51124=>"111111111",
  51125=>"000000100",
  51126=>"000100111",
  51127=>"111000000",
  51128=>"000000111",
  51129=>"111000000",
  51130=>"111000000",
  51131=>"111111100",
  51132=>"111100111",
  51133=>"011001001",
  51134=>"011000100",
  51135=>"000110111",
  51136=>"000000000",
  51137=>"000111111",
  51138=>"001111010",
  51139=>"000110110",
  51140=>"110100100",
  51141=>"010000000",
  51142=>"111101101",
  51143=>"000111111",
  51144=>"011000100",
  51145=>"111011000",
  51146=>"000000111",
  51147=>"010000010",
  51148=>"000000000",
  51149=>"010110111",
  51150=>"101101101",
  51151=>"000100101",
  51152=>"000000111",
  51153=>"111110000",
  51154=>"000000000",
  51155=>"101111111",
  51156=>"000000000",
  51157=>"001000110",
  51158=>"000000111",
  51159=>"111000110",
  51160=>"111110111",
  51161=>"000000111",
  51162=>"000000001",
  51163=>"100000100",
  51164=>"000011111",
  51165=>"111111001",
  51166=>"000000000",
  51167=>"010000001",
  51168=>"000011111",
  51169=>"111111111",
  51170=>"000000001",
  51171=>"000000000",
  51172=>"111111111",
  51173=>"000001001",
  51174=>"100110110",
  51175=>"111111111",
  51176=>"011000001",
  51177=>"000101100",
  51178=>"101000000",
  51179=>"101100000",
  51180=>"100111111",
  51181=>"010000110",
  51182=>"111011000",
  51183=>"011001001",
  51184=>"000111111",
  51185=>"111111111",
  51186=>"001000000",
  51187=>"000111111",
  51188=>"111001000",
  51189=>"111001101",
  51190=>"101100110",
  51191=>"111011000",
  51192=>"110111111",
  51193=>"011110110",
  51194=>"000000001",
  51195=>"001000111",
  51196=>"111111000",
  51197=>"111111111",
  51198=>"000111111",
  51199=>"000000000",
  51200=>"000000000",
  51201=>"101101100",
  51202=>"111101101",
  51203=>"001001111",
  51204=>"111100100",
  51205=>"111111000",
  51206=>"111111000",
  51207=>"111111001",
  51208=>"111111111",
  51209=>"001001101",
  51210=>"000000011",
  51211=>"110111111",
  51212=>"110110110",
  51213=>"111101110",
  51214=>"100110010",
  51215=>"000000000",
  51216=>"100001111",
  51217=>"110110000",
  51218=>"000000000",
  51219=>"110011001",
  51220=>"111101111",
  51221=>"111001001",
  51222=>"111111101",
  51223=>"111111110",
  51224=>"110111111",
  51225=>"100100000",
  51226=>"000000101",
  51227=>"111010000",
  51228=>"111111111",
  51229=>"000000000",
  51230=>"100110110",
  51231=>"111111110",
  51232=>"110110000",
  51233=>"010111111",
  51234=>"111111000",
  51235=>"000001011",
  51236=>"110000000",
  51237=>"000000000",
  51238=>"111111101",
  51239=>"000100101",
  51240=>"111110010",
  51241=>"110111110",
  51242=>"110110000",
  51243=>"111101111",
  51244=>"000000000",
  51245=>"010011111",
  51246=>"000101000",
  51247=>"000110111",
  51248=>"000000000",
  51249=>"000000000",
  51250=>"001000000",
  51251=>"111111111",
  51252=>"111111111",
  51253=>"001000000",
  51254=>"000000000",
  51255=>"111111111",
  51256=>"000000000",
  51257=>"100101101",
  51258=>"111111111",
  51259=>"000000111",
  51260=>"111101101",
  51261=>"110010000",
  51262=>"111100000",
  51263=>"000001101",
  51264=>"111111011",
  51265=>"000110000",
  51266=>"000000111",
  51267=>"001101111",
  51268=>"110010100",
  51269=>"111111001",
  51270=>"111111000",
  51271=>"000000000",
  51272=>"000101111",
  51273=>"111101000",
  51274=>"111111111",
  51275=>"000000000",
  51276=>"000000111",
  51277=>"011000000",
  51278=>"000110100",
  51279=>"111111111",
  51280=>"000000000",
  51281=>"000000100",
  51282=>"000000110",
  51283=>"111110110",
  51284=>"101000000",
  51285=>"111111000",
  51286=>"000011101",
  51287=>"101101111",
  51288=>"000000000",
  51289=>"101000000",
  51290=>"000011010",
  51291=>"111001100",
  51292=>"000000000",
  51293=>"000000101",
  51294=>"001000000",
  51295=>"011011011",
  51296=>"111111000",
  51297=>"111101101",
  51298=>"111111000",
  51299=>"001101000",
  51300=>"101001101",
  51301=>"111001001",
  51302=>"000001101",
  51303=>"000000001",
  51304=>"111111110",
  51305=>"000000111",
  51306=>"000000001",
  51307=>"001001111",
  51308=>"110110110",
  51309=>"000001001",
  51310=>"000000001",
  51311=>"000000000",
  51312=>"000000000",
  51313=>"000000111",
  51314=>"001011011",
  51315=>"111011000",
  51316=>"000000000",
  51317=>"100000111",
  51318=>"000000101",
  51319=>"011111000",
  51320=>"000110111",
  51321=>"110110110",
  51322=>"000000000",
  51323=>"000000000",
  51324=>"110111110",
  51325=>"111111111",
  51326=>"000000000",
  51327=>"110110000",
  51328=>"000000001",
  51329=>"111111111",
  51330=>"000000000",
  51331=>"001001001",
  51332=>"110110110",
  51333=>"000000000",
  51334=>"111111111",
  51335=>"111000000",
  51336=>"010000000",
  51337=>"100000101",
  51338=>"000000000",
  51339=>"000011011",
  51340=>"101111000",
  51341=>"111011000",
  51342=>"111111111",
  51343=>"000000000",
  51344=>"001001100",
  51345=>"111111111",
  51346=>"000000000",
  51347=>"011111011",
  51348=>"111000000",
  51349=>"111101001",
  51350=>"000000010",
  51351=>"000000010",
  51352=>"000000001",
  51353=>"111111111",
  51354=>"111001000",
  51355=>"011011001",
  51356=>"110000001",
  51357=>"000000111",
  51358=>"111111111",
  51359=>"000000101",
  51360=>"010010011",
  51361=>"000111111",
  51362=>"111111010",
  51363=>"010011111",
  51364=>"000000000",
  51365=>"111111011",
  51366=>"111001000",
  51367=>"100110110",
  51368=>"000000011",
  51369=>"000000101",
  51370=>"000000000",
  51371=>"001111111",
  51372=>"111111111",
  51373=>"001001000",
  51374=>"000000000",
  51375=>"000000010",
  51376=>"000000000",
  51377=>"111111001",
  51378=>"011011010",
  51379=>"001000000",
  51380=>"000100110",
  51381=>"000000001",
  51382=>"111111010",
  51383=>"000011111",
  51384=>"010111000",
  51385=>"000000000",
  51386=>"011011001",
  51387=>"011001011",
  51388=>"001001101",
  51389=>"111111111",
  51390=>"000011000",
  51391=>"100111111",
  51392=>"111111111",
  51393=>"000000000",
  51394=>"000000000",
  51395=>"011010011",
  51396=>"111101101",
  51397=>"000000001",
  51398=>"110111111",
  51399=>"000000000",
  51400=>"000000011",
  51401=>"100101111",
  51402=>"000000000",
  51403=>"000000000",
  51404=>"010110010",
  51405=>"000110000",
  51406=>"001001111",
  51407=>"000100101",
  51408=>"001000000",
  51409=>"000100000",
  51410=>"000000000",
  51411=>"100000010",
  51412=>"001000000",
  51413=>"110010110",
  51414=>"000000001",
  51415=>"111111011",
  51416=>"000000000",
  51417=>"001001001",
  51418=>"111101000",
  51419=>"111111111",
  51420=>"110111011",
  51421=>"100000000",
  51422=>"000000101",
  51423=>"000000000",
  51424=>"111111111",
  51425=>"111011000",
  51426=>"011111111",
  51427=>"111111011",
  51428=>"101111011",
  51429=>"000000000",
  51430=>"111111111",
  51431=>"110111001",
  51432=>"111111001",
  51433=>"011001000",
  51434=>"100000000",
  51435=>"110110000",
  51436=>"011111100",
  51437=>"000111010",
  51438=>"000000110",
  51439=>"111000000",
  51440=>"000000101",
  51441=>"000000001",
  51442=>"001011111",
  51443=>"000100101",
  51444=>"110111010",
  51445=>"100100100",
  51446=>"000011001",
  51447=>"000000000",
  51448=>"100100000",
  51449=>"011111111",
  51450=>"001000111",
  51451=>"111111111",
  51452=>"000000000",
  51453=>"001001001",
  51454=>"111001111",
  51455=>"000000000",
  51456=>"100000000",
  51457=>"101101001",
  51458=>"101111111",
  51459=>"111111010",
  51460=>"000001000",
  51461=>"000011111",
  51462=>"111111101",
  51463=>"111110111",
  51464=>"110111110",
  51465=>"001101111",
  51466=>"111111110",
  51467=>"111110110",
  51468=>"111111111",
  51469=>"111111100",
  51470=>"111111000",
  51471=>"000000110",
  51472=>"100100111",
  51473=>"000000101",
  51474=>"000001111",
  51475=>"000000001",
  51476=>"111101111",
  51477=>"111000000",
  51478=>"001001101",
  51479=>"100100000",
  51480=>"001011111",
  51481=>"001101111",
  51482=>"111111111",
  51483=>"000000000",
  51484=>"000001000",
  51485=>"000000000",
  51486=>"100000000",
  51487=>"000001100",
  51488=>"000000000",
  51489=>"000100001",
  51490=>"011010000",
  51491=>"010001011",
  51492=>"111111000",
  51493=>"111101000",
  51494=>"011000001",
  51495=>"011000000",
  51496=>"000101111",
  51497=>"101101011",
  51498=>"011000000",
  51499=>"111011111",
  51500=>"111111111",
  51501=>"001011001",
  51502=>"000000000",
  51503=>"001000000",
  51504=>"000001111",
  51505=>"001000000",
  51506=>"111011011",
  51507=>"000000010",
  51508=>"011111110",
  51509=>"000000000",
  51510=>"000000000",
  51511=>"000000000",
  51512=>"000000000",
  51513=>"000000111",
  51514=>"111111000",
  51515=>"000000111",
  51516=>"000011000",
  51517=>"111111111",
  51518=>"000000110",
  51519=>"000000000",
  51520=>"000001111",
  51521=>"111111110",
  51522=>"111111010",
  51523=>"111001001",
  51524=>"111101000",
  51525=>"000001111",
  51526=>"011000010",
  51527=>"110110110",
  51528=>"100100100",
  51529=>"010000000",
  51530=>"001001101",
  51531=>"111111111",
  51532=>"010100111",
  51533=>"000010010",
  51534=>"000001001",
  51535=>"011011010",
  51536=>"001001001",
  51537=>"000000100",
  51538=>"110000000",
  51539=>"111000000",
  51540=>"000101111",
  51541=>"011011011",
  51542=>"111111111",
  51543=>"111111111",
  51544=>"000001101",
  51545=>"001000000",
  51546=>"000000000",
  51547=>"000000000",
  51548=>"111111111",
  51549=>"000100111",
  51550=>"000000000",
  51551=>"111111101",
  51552=>"111111001",
  51553=>"001000001",
  51554=>"001101100",
  51555=>"101101111",
  51556=>"000110000",
  51557=>"000000000",
  51558=>"100110111",
  51559=>"100110010",
  51560=>"110111111",
  51561=>"111111111",
  51562=>"001000000",
  51563=>"000000100",
  51564=>"100111110",
  51565=>"011000000",
  51566=>"000000111",
  51567=>"001001001",
  51568=>"000000000",
  51569=>"110000000",
  51570=>"000000111",
  51571=>"011000000",
  51572=>"000000000",
  51573=>"000110110",
  51574=>"001000010",
  51575=>"111111011",
  51576=>"000000000",
  51577=>"000000000",
  51578=>"000000001",
  51579=>"111011011",
  51580=>"111000000",
  51581=>"111111111",
  51582=>"000000000",
  51583=>"000000000",
  51584=>"000000100",
  51585=>"000000000",
  51586=>"111111000",
  51587=>"111111101",
  51588=>"111000000",
  51589=>"111111011",
  51590=>"110111000",
  51591=>"111000000",
  51592=>"101111111",
  51593=>"101101100",
  51594=>"001001100",
  51595=>"011001011",
  51596=>"000000000",
  51597=>"110110000",
  51598=>"000001101",
  51599=>"000000000",
  51600=>"000001001",
  51601=>"111111111",
  51602=>"010000000",
  51603=>"110100000",
  51604=>"011011010",
  51605=>"000010000",
  51606=>"000000000",
  51607=>"011011111",
  51608=>"111111111",
  51609=>"100000000",
  51610=>"000000001",
  51611=>"111111010",
  51612=>"001001001",
  51613=>"111000000",
  51614=>"101111111",
  51615=>"111110000",
  51616=>"000101111",
  51617=>"100000000",
  51618=>"111110010",
  51619=>"000000110",
  51620=>"111111010",
  51621=>"111111111",
  51622=>"111011011",
  51623=>"100111000",
  51624=>"000110111",
  51625=>"000000000",
  51626=>"111111111",
  51627=>"101000100",
  51628=>"111000000",
  51629=>"001111111",
  51630=>"110110000",
  51631=>"000011011",
  51632=>"111110000",
  51633=>"110111111",
  51634=>"000000000",
  51635=>"000000000",
  51636=>"000001001",
  51637=>"110111111",
  51638=>"000000000",
  51639=>"001001111",
  51640=>"000000110",
  51641=>"001000000",
  51642=>"111111111",
  51643=>"111111111",
  51644=>"000000111",
  51645=>"111111111",
  51646=>"011111101",
  51647=>"000100100",
  51648=>"110110010",
  51649=>"111111111",
  51650=>"111111010",
  51651=>"000000101",
  51652=>"000001101",
  51653=>"111111001",
  51654=>"000000101",
  51655=>"111111100",
  51656=>"000000000",
  51657=>"111011011",
  51658=>"000000001",
  51659=>"000000000",
  51660=>"010011111",
  51661=>"000000000",
  51662=>"110101000",
  51663=>"101100101",
  51664=>"000000000",
  51665=>"111111111",
  51666=>"111111111",
  51667=>"111111111",
  51668=>"101100000",
  51669=>"110000000",
  51670=>"000000000",
  51671=>"111111111",
  51672=>"000001101",
  51673=>"000111111",
  51674=>"101111001",
  51675=>"000111111",
  51676=>"110111111",
  51677=>"000000000",
  51678=>"000000100",
  51679=>"111001000",
  51680=>"111100000",
  51681=>"111111111",
  51682=>"000010111",
  51683=>"110101111",
  51684=>"000000000",
  51685=>"111001001",
  51686=>"111000101",
  51687=>"000001001",
  51688=>"101111101",
  51689=>"000000111",
  51690=>"111111110",
  51691=>"000100000",
  51692=>"010000000",
  51693=>"000000001",
  51694=>"101001001",
  51695=>"011111110",
  51696=>"000001011",
  51697=>"101101100",
  51698=>"011000001",
  51699=>"111111111",
  51700=>"111111111",
  51701=>"001000000",
  51702=>"101111001",
  51703=>"000100110",
  51704=>"111111111",
  51705=>"001000000",
  51706=>"100000000",
  51707=>"000000111",
  51708=>"111000000",
  51709=>"111111111",
  51710=>"111111000",
  51711=>"000000000",
  51712=>"000001001",
  51713=>"001000000",
  51714=>"000000000",
  51715=>"111011011",
  51716=>"010010000",
  51717=>"111111111",
  51718=>"111110111",
  51719=>"000000001",
  51720=>"011111111",
  51721=>"111111111",
  51722=>"011000000",
  51723=>"000100000",
  51724=>"011011000",
  51725=>"000100100",
  51726=>"110111011",
  51727=>"001000000",
  51728=>"011011000",
  51729=>"111101111",
  51730=>"111111111",
  51731=>"011000000",
  51732=>"101000000",
  51733=>"111111111",
  51734=>"000000111",
  51735=>"011010010",
  51736=>"000100110",
  51737=>"010000001",
  51738=>"110011111",
  51739=>"000100111",
  51740=>"111111111",
  51741=>"111000000",
  51742=>"100100100",
  51743=>"000000000",
  51744=>"011111111",
  51745=>"000000001",
  51746=>"111111111",
  51747=>"111111111",
  51748=>"000000000",
  51749=>"000000000",
  51750=>"111111111",
  51751=>"111000001",
  51752=>"000000000",
  51753=>"111100000",
  51754=>"001000111",
  51755=>"111110101",
  51756=>"000000000",
  51757=>"000000000",
  51758=>"111111111",
  51759=>"000000100",
  51760=>"000000000",
  51761=>"110110110",
  51762=>"000000000",
  51763=>"000111111",
  51764=>"000000000",
  51765=>"110011001",
  51766=>"000000000",
  51767=>"000100111",
  51768=>"111111000",
  51769=>"000100100",
  51770=>"000000101",
  51771=>"010000000",
  51772=>"000000000",
  51773=>"111111111",
  51774=>"111111111",
  51775=>"111111111",
  51776=>"111111111",
  51777=>"110111111",
  51778=>"111000000",
  51779=>"111110111",
  51780=>"001001000",
  51781=>"000000011",
  51782=>"000000000",
  51783=>"000000000",
  51784=>"110110010",
  51785=>"000110111",
  51786=>"000000000",
  51787=>"000000101",
  51788=>"100000100",
  51789=>"100100000",
  51790=>"111111000",
  51791=>"000111001",
  51792=>"111111111",
  51793=>"000011111",
  51794=>"000010010",
  51795=>"100000000",
  51796=>"000000000",
  51797=>"000000000",
  51798=>"000000100",
  51799=>"111110100",
  51800=>"000011111",
  51801=>"100100100",
  51802=>"001101101",
  51803=>"010010111",
  51804=>"101111111",
  51805=>"001000000",
  51806=>"001000000",
  51807=>"010011000",
  51808=>"111111001",
  51809=>"000100000",
  51810=>"000000000",
  51811=>"000000000",
  51812=>"000001010",
  51813=>"111110110",
  51814=>"110111111",
  51815=>"111000111",
  51816=>"111111011",
  51817=>"000001111",
  51818=>"010000111",
  51819=>"000000010",
  51820=>"111111111",
  51821=>"111111111",
  51822=>"001000000",
  51823=>"000000000",
  51824=>"000000100",
  51825=>"111011111",
  51826=>"001001000",
  51827=>"110011001",
  51828=>"000000100",
  51829=>"111111011",
  51830=>"111000000",
  51831=>"000111100",
  51832=>"100000011",
  51833=>"111111111",
  51834=>"000000000",
  51835=>"000000001",
  51836=>"110110110",
  51837=>"010101000",
  51838=>"011011010",
  51839=>"000000000",
  51840=>"101000100",
  51841=>"000011011",
  51842=>"011110000",
  51843=>"000000000",
  51844=>"000000001",
  51845=>"111011111",
  51846=>"111111111",
  51847=>"000101111",
  51848=>"001111000",
  51849=>"111111000",
  51850=>"110111001",
  51851=>"000000100",
  51852=>"100000000",
  51853=>"000000000",
  51854=>"010111000",
  51855=>"111111000",
  51856=>"001111111",
  51857=>"000000110",
  51858=>"000110110",
  51859=>"111111101",
  51860=>"000000000",
  51861=>"001000000",
  51862=>"001001000",
  51863=>"000000000",
  51864=>"000000000",
  51865=>"111111111",
  51866=>"111111111",
  51867=>"000101011",
  51868=>"011001101",
  51869=>"111111111",
  51870=>"111110111",
  51871=>"100000000",
  51872=>"011000110",
  51873=>"111110110",
  51874=>"000000110",
  51875=>"111000000",
  51876=>"111111111",
  51877=>"001011001",
  51878=>"111000000",
  51879=>"011011011",
  51880=>"110001001",
  51881=>"111111111",
  51882=>"000000001",
  51883=>"001000000",
  51884=>"011010110",
  51885=>"110100100",
  51886=>"000000000",
  51887=>"110010000",
  51888=>"111111111",
  51889=>"000000000",
  51890=>"001011000",
  51891=>"000000000",
  51892=>"111000001",
  51893=>"000000100",
  51894=>"000000000",
  51895=>"000000001",
  51896=>"000000000",
  51897=>"010111111",
  51898=>"011000000",
  51899=>"000000000",
  51900=>"000000000",
  51901=>"111011111",
  51902=>"000000000",
  51903=>"110111000",
  51904=>"111111111",
  51905=>"001001000",
  51906=>"000001000",
  51907=>"111111001",
  51908=>"111001001",
  51909=>"001001000",
  51910=>"100100101",
  51911=>"111111111",
  51912=>"001110111",
  51913=>"000000000",
  51914=>"000000000",
  51915=>"111111111",
  51916=>"011100111",
  51917=>"011111111",
  51918=>"100100100",
  51919=>"000000000",
  51920=>"011111110",
  51921=>"000000100",
  51922=>"000000100",
  51923=>"111111111",
  51924=>"111111111",
  51925=>"000000000",
  51926=>"000000000",
  51927=>"000000000",
  51928=>"000000110",
  51929=>"111110000",
  51930=>"111111111",
  51931=>"111000110",
  51932=>"000100111",
  51933=>"000000000",
  51934=>"111000000",
  51935=>"111111000",
  51936=>"111111001",
  51937=>"000000000",
  51938=>"011111000",
  51939=>"000100000",
  51940=>"000001011",
  51941=>"001011111",
  51942=>"011000110",
  51943=>"000000000",
  51944=>"000000000",
  51945=>"111111110",
  51946=>"000000001",
  51947=>"001000000",
  51948=>"000000000",
  51949=>"111011111",
  51950=>"000111111",
  51951=>"011111000",
  51952=>"101111111",
  51953=>"111000011",
  51954=>"111111111",
  51955=>"011110111",
  51956=>"111001001",
  51957=>"111110010",
  51958=>"000001001",
  51959=>"111111011",
  51960=>"111001000",
  51961=>"111111111",
  51962=>"000100111",
  51963=>"000000000",
  51964=>"111111001",
  51965=>"111111111",
  51966=>"001000000",
  51967=>"111111110",
  51968=>"111111111",
  51969=>"000001011",
  51970=>"000000011",
  51971=>"101100111",
  51972=>"000000000",
  51973=>"000000101",
  51974=>"000000000",
  51975=>"111011000",
  51976=>"100100000",
  51977=>"000000000",
  51978=>"111101000",
  51979=>"110001001",
  51980=>"000000000",
  51981=>"000100111",
  51982=>"000000000",
  51983=>"010111111",
  51984=>"000000000",
  51985=>"000110110",
  51986=>"001101111",
  51987=>"111111111",
  51988=>"000000100",
  51989=>"100110000",
  51990=>"110111111",
  51991=>"100111111",
  51992=>"111010000",
  51993=>"111111011",
  51994=>"000000101",
  51995=>"010000111",
  51996=>"111111111",
  51997=>"000000111",
  51998=>"000000000",
  51999=>"000010110",
  52000=>"010001011",
  52001=>"111111111",
  52002=>"000000110",
  52003=>"000000000",
  52004=>"110000000",
  52005=>"000000000",
  52006=>"111111111",
  52007=>"111111111",
  52008=>"000000000",
  52009=>"001001000",
  52010=>"110110100",
  52011=>"011011001",
  52012=>"000000111",
  52013=>"000000000",
  52014=>"111001110",
  52015=>"000100000",
  52016=>"000000111",
  52017=>"000000001",
  52018=>"111111111",
  52019=>"111000000",
  52020=>"110110110",
  52021=>"100000000",
  52022=>"111111111",
  52023=>"000000000",
  52024=>"111111000",
  52025=>"111111111",
  52026=>"000000000",
  52027=>"011001000",
  52028=>"111111111",
  52029=>"100100110",
  52030=>"110011011",
  52031=>"011000000",
  52032=>"111111011",
  52033=>"000011000",
  52034=>"111111111",
  52035=>"111010111",
  52036=>"110110110",
  52037=>"111100001",
  52038=>"110110110",
  52039=>"110110110",
  52040=>"000000000",
  52041=>"000110000",
  52042=>"100000000",
  52043=>"110100110",
  52044=>"101101111",
  52045=>"110111110",
  52046=>"111100111",
  52047=>"000000010",
  52048=>"111101100",
  52049=>"000000001",
  52050=>"000000000",
  52051=>"111100100",
  52052=>"000000000",
  52053=>"011011111",
  52054=>"000000011",
  52055=>"000000000",
  52056=>"000000000",
  52057=>"101111000",
  52058=>"100100000",
  52059=>"100000000",
  52060=>"111010011",
  52061=>"110110111",
  52062=>"000000000",
  52063=>"010000000",
  52064=>"010000000",
  52065=>"111111111",
  52066=>"000110011",
  52067=>"000000000",
  52068=>"111111111",
  52069=>"000000000",
  52070=>"000000010",
  52071=>"000000000",
  52072=>"011011111",
  52073=>"000001111",
  52074=>"111000000",
  52075=>"000111000",
  52076=>"110110110",
  52077=>"011100100",
  52078=>"110100000",
  52079=>"010000000",
  52080=>"010111111",
  52081=>"111111111",
  52082=>"101101110",
  52083=>"111110010",
  52084=>"000110111",
  52085=>"001000110",
  52086=>"100101111",
  52087=>"000000000",
  52088=>"111111111",
  52089=>"011011010",
  52090=>"111101100",
  52091=>"000000100",
  52092=>"100111111",
  52093=>"111110100",
  52094=>"000000000",
  52095=>"100000000",
  52096=>"000000000",
  52097=>"111110100",
  52098=>"010000000",
  52099=>"101101100",
  52100=>"111111000",
  52101=>"110110110",
  52102=>"111000100",
  52103=>"000000000",
  52104=>"000010101",
  52105=>"000000111",
  52106=>"001000000",
  52107=>"000010111",
  52108=>"001100101",
  52109=>"110110110",
  52110=>"100000001",
  52111=>"100110111",
  52112=>"000000000",
  52113=>"000000000",
  52114=>"000001111",
  52115=>"110000011",
  52116=>"111111011",
  52117=>"000001010",
  52118=>"001011011",
  52119=>"111111111",
  52120=>"011111111",
  52121=>"011000100",
  52122=>"110000000",
  52123=>"000000001",
  52124=>"111110110",
  52125=>"000000000",
  52126=>"001000000",
  52127=>"010011111",
  52128=>"101000000",
  52129=>"000001001",
  52130=>"111111111",
  52131=>"001000000",
  52132=>"111110111",
  52133=>"011011011",
  52134=>"000111111",
  52135=>"111111110",
  52136=>"001000001",
  52137=>"110100001",
  52138=>"000000001",
  52139=>"011001000",
  52140=>"111111111",
  52141=>"001000111",
  52142=>"111011011",
  52143=>"111010000",
  52144=>"000000010",
  52145=>"000000000",
  52146=>"000000000",
  52147=>"000100100",
  52148=>"100110110",
  52149=>"000000000",
  52150=>"000000000",
  52151=>"000001001",
  52152=>"001111111",
  52153=>"001011011",
  52154=>"100000111",
  52155=>"111111110",
  52156=>"011001000",
  52157=>"000000000",
  52158=>"111110000",
  52159=>"001100110",
  52160=>"110111011",
  52161=>"111111111",
  52162=>"000000000",
  52163=>"000000110",
  52164=>"110110111",
  52165=>"110000000",
  52166=>"000000111",
  52167=>"111001001",
  52168=>"111110111",
  52169=>"000110111",
  52170=>"110100100",
  52171=>"110000000",
  52172=>"001101000",
  52173=>"000000000",
  52174=>"101100100",
  52175=>"001000110",
  52176=>"011000000",
  52177=>"011110111",
  52178=>"111111111",
  52179=>"000000000",
  52180=>"000000000",
  52181=>"000000001",
  52182=>"011000000",
  52183=>"110111011",
  52184=>"111111111",
  52185=>"001000000",
  52186=>"000000000",
  52187=>"111111111",
  52188=>"111111111",
  52189=>"111111001",
  52190=>"000000000",
  52191=>"000000000",
  52192=>"011111110",
  52193=>"111111000",
  52194=>"111111001",
  52195=>"000010000",
  52196=>"111111111",
  52197=>"001001001",
  52198=>"000000000",
  52199=>"111100000",
  52200=>"000000000",
  52201=>"000000000",
  52202=>"001001011",
  52203=>"110110111",
  52204=>"011000000",
  52205=>"111111111",
  52206=>"011011000",
  52207=>"000000000",
  52208=>"000000000",
  52209=>"000000001",
  52210=>"111111111",
  52211=>"000000000",
  52212=>"011111110",
  52213=>"000000000",
  52214=>"000000000",
  52215=>"011011000",
  52216=>"010010010",
  52217=>"111111111",
  52218=>"000000000",
  52219=>"000000000",
  52220=>"000000111",
  52221=>"000000000",
  52222=>"111100100",
  52223=>"000000000",
  52224=>"110111110",
  52225=>"010001001",
  52226=>"001000111",
  52227=>"000000000",
  52228=>"111111110",
  52229=>"100000000",
  52230=>"000000111",
  52231=>"111000000",
  52232=>"010000001",
  52233=>"111110000",
  52234=>"111111100",
  52235=>"111111111",
  52236=>"000000110",
  52237=>"111111000",
  52238=>"111011011",
  52239=>"111111100",
  52240=>"000001111",
  52241=>"000111111",
  52242=>"111111000",
  52243=>"111000000",
  52244=>"011111111",
  52245=>"111001001",
  52246=>"000111111",
  52247=>"000000111",
  52248=>"000000111",
  52249=>"000100110",
  52250=>"111111111",
  52251=>"111101100",
  52252=>"111111111",
  52253=>"000000000",
  52254=>"101000000",
  52255=>"000010000",
  52256=>"000001101",
  52257=>"100000000",
  52258=>"111111001",
  52259=>"000000111",
  52260=>"000011100",
  52261=>"000011011",
  52262=>"000000000",
  52263=>"111111000",
  52264=>"111001000",
  52265=>"000000111",
  52266=>"000100000",
  52267=>"111111111",
  52268=>"000000000",
  52269=>"111111111",
  52270=>"111111100",
  52271=>"000111111",
  52272=>"111101101",
  52273=>"111000000",
  52274=>"000001111",
  52275=>"100111011",
  52276=>"111000001",
  52277=>"000000111",
  52278=>"000000000",
  52279=>"011001000",
  52280=>"000011111",
  52281=>"111111101",
  52282=>"000000001",
  52283=>"111000000",
  52284=>"000000111",
  52285=>"000000000",
  52286=>"111011100",
  52287=>"000111111",
  52288=>"011111110",
  52289=>"000000000",
  52290=>"001011000",
  52291=>"000000000",
  52292=>"011100111",
  52293=>"111100100",
  52294=>"111010000",
  52295=>"111111000",
  52296=>"111111011",
  52297=>"000000111",
  52298=>"111111111",
  52299=>"110101101",
  52300=>"111111000",
  52301=>"000111111",
  52302=>"000000111",
  52303=>"000000001",
  52304=>"110111111",
  52305=>"101000000",
  52306=>"000000000",
  52307=>"110110111",
  52308=>"000000000",
  52309=>"111111111",
  52310=>"111100000",
  52311=>"000101111",
  52312=>"000111111",
  52313=>"000000000",
  52314=>"000000000",
  52315=>"111000000",
  52316=>"000111111",
  52317=>"111001000",
  52318=>"110100000",
  52319=>"000000100",
  52320=>"101000000",
  52321=>"100000000",
  52322=>"111111111",
  52323=>"010000000",
  52324=>"000000010",
  52325=>"000000111",
  52326=>"111110000",
  52327=>"000000000",
  52328=>"011000000",
  52329=>"111111000",
  52330=>"111000000",
  52331=>"111010000",
  52332=>"111111001",
  52333=>"000110111",
  52334=>"111000000",
  52335=>"111000000",
  52336=>"000000000",
  52337=>"000001011",
  52338=>"111111000",
  52339=>"001000001",
  52340=>"011000101",
  52341=>"000111111",
  52342=>"111000111",
  52343=>"111011111",
  52344=>"000000000",
  52345=>"000000101",
  52346=>"110111111",
  52347=>"111000001",
  52348=>"110110000",
  52349=>"100000000",
  52350=>"000111111",
  52351=>"100111001",
  52352=>"001000000",
  52353=>"000111111",
  52354=>"000000000",
  52355=>"000000111",
  52356=>"000000000",
  52357=>"000000011",
  52358=>"111000000",
  52359=>"000000000",
  52360=>"000000000",
  52361=>"000000000",
  52362=>"100111111",
  52363=>"111111111",
  52364=>"011000011",
  52365=>"000000000",
  52366=>"000000111",
  52367=>"000011000",
  52368=>"000000111",
  52369=>"000110110",
  52370=>"111110000",
  52371=>"100110110",
  52372=>"000000000",
  52373=>"000000000",
  52374=>"001011111",
  52375=>"111000000",
  52376=>"000000101",
  52377=>"000000000",
  52378=>"001111000",
  52379=>"001000001",
  52380=>"111110111",
  52381=>"111111101",
  52382=>"000111111",
  52383=>"110111110",
  52384=>"001000001",
  52385=>"100000010",
  52386=>"000000000",
  52387=>"000000001",
  52388=>"000011111",
  52389=>"000111111",
  52390=>"111111111",
  52391=>"000010010",
  52392=>"111111101",
  52393=>"000000000",
  52394=>"111000000",
  52395=>"111110100",
  52396=>"110100100",
  52397=>"000011111",
  52398=>"111000100",
  52399=>"111111111",
  52400=>"111111111",
  52401=>"000010011",
  52402=>"111111101",
  52403=>"010101111",
  52404=>"111111000",
  52405=>"000001000",
  52406=>"111111000",
  52407=>"111111100",
  52408=>"001000100",
  52409=>"111111111",
  52410=>"000000011",
  52411=>"001001001",
  52412=>"111001000",
  52413=>"111000001",
  52414=>"111111000",
  52415=>"111110000",
  52416=>"000000000",
  52417=>"110110111",
  52418=>"111111111",
  52419=>"111110001",
  52420=>"111000000",
  52421=>"000100001",
  52422=>"000000110",
  52423=>"000000000",
  52424=>"111011000",
  52425=>"111000000",
  52426=>"001000111",
  52427=>"111001000",
  52428=>"111111000",
  52429=>"010111000",
  52430=>"000010110",
  52431=>"000000111",
  52432=>"000000000",
  52433=>"000000000",
  52434=>"011001101",
  52435=>"000000000",
  52436=>"000000000",
  52437=>"100111111",
  52438=>"111111011",
  52439=>"111000000",
  52440=>"101110000",
  52441=>"111111000",
  52442=>"101000000",
  52443=>"001000000",
  52444=>"111111111",
  52445=>"000000001",
  52446=>"111111111",
  52447=>"000000000",
  52448=>"110110010",
  52449=>"000000000",
  52450=>"000111000",
  52451=>"000000000",
  52452=>"000001111",
  52453=>"111010000",
  52454=>"000100111",
  52455=>"111111111",
  52456=>"011011111",
  52457=>"111100000",
  52458=>"111111110",
  52459=>"100111000",
  52460=>"000000011",
  52461=>"000111000",
  52462=>"100100011",
  52463=>"000000111",
  52464=>"000000000",
  52465=>"000011111",
  52466=>"111101110",
  52467=>"001111111",
  52468=>"111000000",
  52469=>"110100110",
  52470=>"100100101",
  52471=>"001001111",
  52472=>"110111111",
  52473=>"000000000",
  52474=>"111110000",
  52475=>"011000000",
  52476=>"001001000",
  52477=>"101001111",
  52478=>"000000111",
  52479=>"000000000",
  52480=>"000000001",
  52481=>"000000001",
  52482=>"010000000",
  52483=>"011111111",
  52484=>"100000000",
  52485=>"000100000",
  52486=>"111111000",
  52487=>"000000000",
  52488=>"000000111",
  52489=>"000000111",
  52490=>"000000000",
  52491=>"000011000",
  52492=>"101100111",
  52493=>"000010000",
  52494=>"001001000",
  52495=>"000000111",
  52496=>"000000111",
  52497=>"111011111",
  52498=>"000000000",
  52499=>"101000000",
  52500=>"000100111",
  52501=>"000100000",
  52502=>"111100001",
  52503=>"000000000",
  52504=>"111111011",
  52505=>"000000000",
  52506=>"100100000",
  52507=>"000000000",
  52508=>"110110110",
  52509=>"000000111",
  52510=>"111110000",
  52511=>"010111010",
  52512=>"111111000",
  52513=>"111111000",
  52514=>"110001000",
  52515=>"111111001",
  52516=>"111000000",
  52517=>"111111111",
  52518=>"000111011",
  52519=>"111000001",
  52520=>"111111111",
  52521=>"110111010",
  52522=>"000011111",
  52523=>"111111111",
  52524=>"111011000",
  52525=>"000101100",
  52526=>"000111001",
  52527=>"000000000",
  52528=>"100000000",
  52529=>"111111111",
  52530=>"000000000",
  52531=>"111011111",
  52532=>"110100000",
  52533=>"010010011",
  52534=>"100110001",
  52535=>"111101111",
  52536=>"000000000",
  52537=>"111001111",
  52538=>"000000111",
  52539=>"111111010",
  52540=>"111110000",
  52541=>"101000011",
  52542=>"000100010",
  52543=>"011000000",
  52544=>"000101111",
  52545=>"000111100",
  52546=>"000000110",
  52547=>"110110111",
  52548=>"110111000",
  52549=>"101000000",
  52550=>"000111111",
  52551=>"101111111",
  52552=>"111010000",
  52553=>"000000000",
  52554=>"110110000",
  52555=>"001110100",
  52556=>"011000111",
  52557=>"001111111",
  52558=>"000101101",
  52559=>"100001111",
  52560=>"000000001",
  52561=>"001011000",
  52562=>"000101111",
  52563=>"000101111",
  52564=>"000000001",
  52565=>"011011011",
  52566=>"001111111",
  52567=>"001000001",
  52568=>"111011011",
  52569=>"111000001",
  52570=>"101111111",
  52571=>"010111110",
  52572=>"111000000",
  52573=>"001000000",
  52574=>"000000111",
  52575=>"111010111",
  52576=>"000000000",
  52577=>"111000001",
  52578=>"000000100",
  52579=>"000000101",
  52580=>"100000000",
  52581=>"100110001",
  52582=>"000000000",
  52583=>"000111001",
  52584=>"000100100",
  52585=>"111000000",
  52586=>"000111111",
  52587=>"001111111",
  52588=>"000000000",
  52589=>"000011111",
  52590=>"000000000",
  52591=>"000000000",
  52592=>"101100000",
  52593=>"100000111",
  52594=>"000111111",
  52595=>"111111001",
  52596=>"000000000",
  52597=>"000100100",
  52598=>"111111111",
  52599=>"111111101",
  52600=>"000000000",
  52601=>"111111000",
  52602=>"000000111",
  52603=>"000111111",
  52604=>"111111111",
  52605=>"111111001",
  52606=>"111101001",
  52607=>"111010110",
  52608=>"110011111",
  52609=>"111111111",
  52610=>"111001111",
  52611=>"111111111",
  52612=>"111011001",
  52613=>"110110000",
  52614=>"011011000",
  52615=>"111111000",
  52616=>"000000111",
  52617=>"011011000",
  52618=>"101111111",
  52619=>"000111111",
  52620=>"111100111",
  52621=>"110100000",
  52622=>"111111111",
  52623=>"110111001",
  52624=>"100111111",
  52625=>"111001000",
  52626=>"111011001",
  52627=>"111100000",
  52628=>"000001100",
  52629=>"000000000",
  52630=>"011111111",
  52631=>"010001000",
  52632=>"101001011",
  52633=>"000000001",
  52634=>"111111011",
  52635=>"000001111",
  52636=>"001000100",
  52637=>"111111000",
  52638=>"000100000",
  52639=>"000000000",
  52640=>"111100000",
  52641=>"111111111",
  52642=>"000010000",
  52643=>"000000000",
  52644=>"111110101",
  52645=>"000000000",
  52646=>"000000011",
  52647=>"111111100",
  52648=>"111000111",
  52649=>"110110000",
  52650=>"111111111",
  52651=>"000000000",
  52652=>"000110100",
  52653=>"101111111",
  52654=>"111111111",
  52655=>"111101101",
  52656=>"000111111",
  52657=>"111111111",
  52658=>"000111111",
  52659=>"011000011",
  52660=>"111111111",
  52661=>"111111110",
  52662=>"011011001",
  52663=>"111111111",
  52664=>"000000001",
  52665=>"000111111",
  52666=>"000000000",
  52667=>"000000000",
  52668=>"101011101",
  52669=>"111000000",
  52670=>"000000111",
  52671=>"100100111",
  52672=>"111111111",
  52673=>"111111101",
  52674=>"111100000",
  52675=>"000000000",
  52676=>"000000000",
  52677=>"101101111",
  52678=>"110111000",
  52679=>"000000000",
  52680=>"000000001",
  52681=>"111111000",
  52682=>"000000000",
  52683=>"111000000",
  52684=>"111111000",
  52685=>"111111001",
  52686=>"111100100",
  52687=>"011111100",
  52688=>"000000111",
  52689=>"001111111",
  52690=>"001001111",
  52691=>"011011111",
  52692=>"000100100",
  52693=>"111000000",
  52694=>"000111111",
  52695=>"000111001",
  52696=>"000000111",
  52697=>"111111000",
  52698=>"000000000",
  52699=>"111001000",
  52700=>"000000000",
  52701=>"111000001",
  52702=>"000110111",
  52703=>"001000001",
  52704=>"111111111",
  52705=>"000000000",
  52706=>"000000000",
  52707=>"011000000",
  52708=>"000001011",
  52709=>"000000000",
  52710=>"100111000",
  52711=>"000010110",
  52712=>"000000111",
  52713=>"111110111",
  52714=>"000000010",
  52715=>"101010000",
  52716=>"111111111",
  52717=>"000110000",
  52718=>"000000000",
  52719=>"000000000",
  52720=>"000111111",
  52721=>"000111001",
  52722=>"111100000",
  52723=>"000111000",
  52724=>"111111011",
  52725=>"011011111",
  52726=>"000000110",
  52727=>"111001011",
  52728=>"000111111",
  52729=>"111111011",
  52730=>"001000000",
  52731=>"111000000",
  52732=>"111111111",
  52733=>"001100111",
  52734=>"100000000",
  52735=>"000111111",
  52736=>"000000000",
  52737=>"000000011",
  52738=>"000000001",
  52739=>"111111111",
  52740=>"111111111",
  52741=>"111000100",
  52742=>"111111110",
  52743=>"000000000",
  52744=>"111111111",
  52745=>"110010010",
  52746=>"111101111",
  52747=>"011010111",
  52748=>"111101101",
  52749=>"111111001",
  52750=>"000000001",
  52751=>"111111111",
  52752=>"111111111",
  52753=>"111101100",
  52754=>"100000000",
  52755=>"111111101",
  52756=>"000111111",
  52757=>"000011010",
  52758=>"100111110",
  52759=>"000000000",
  52760=>"001001001",
  52761=>"000000001",
  52762=>"000000000",
  52763=>"000000000",
  52764=>"000000000",
  52765=>"000001001",
  52766=>"000000000",
  52767=>"111111111",
  52768=>"111110111",
  52769=>"001011111",
  52770=>"001111000",
  52771=>"011001111",
  52772=>"000010111",
  52773=>"000000101",
  52774=>"001000000",
  52775=>"000000001",
  52776=>"000000001",
  52777=>"000000111",
  52778=>"000000101",
  52779=>"000000000",
  52780=>"111101111",
  52781=>"000000110",
  52782=>"111111111",
  52783=>"011110000",
  52784=>"111111111",
  52785=>"111000000",
  52786=>"111111111",
  52787=>"000001001",
  52788=>"110110010",
  52789=>"110000000",
  52790=>"110110110",
  52791=>"001000001",
  52792=>"111111101",
  52793=>"100100111",
  52794=>"111111111",
  52795=>"000000110",
  52796=>"000000111",
  52797=>"100000000",
  52798=>"011011001",
  52799=>"111111111",
  52800=>"111111111",
  52801=>"111111111",
  52802=>"111111111",
  52803=>"000100110",
  52804=>"111101100",
  52805=>"000000000",
  52806=>"000000000",
  52807=>"111111111",
  52808=>"111111111",
  52809=>"000000000",
  52810=>"000000000",
  52811=>"111000000",
  52812=>"000000000",
  52813=>"000000111",
  52814=>"000000011",
  52815=>"000000000",
  52816=>"110000000",
  52817=>"110010001",
  52818=>"010011000",
  52819=>"000000000",
  52820=>"000100111",
  52821=>"001111110",
  52822=>"111111111",
  52823=>"000000000",
  52824=>"000000000",
  52825=>"000000000",
  52826=>"111111111",
  52827=>"001011111",
  52828=>"000000010",
  52829=>"111000111",
  52830=>"001101111",
  52831=>"010111011",
  52832=>"111000010",
  52833=>"000000000",
  52834=>"101111111",
  52835=>"111101111",
  52836=>"100000000",
  52837=>"111111111",
  52838=>"111111111",
  52839=>"000100000",
  52840=>"000000000",
  52841=>"111101111",
  52842=>"000000000",
  52843=>"010111111",
  52844=>"010110000",
  52845=>"001001111",
  52846=>"000000111",
  52847=>"000000000",
  52848=>"000000111",
  52849=>"000010000",
  52850=>"111011011",
  52851=>"111111110",
  52852=>"000000000",
  52853=>"000000000",
  52854=>"111111010",
  52855=>"000000000",
  52856=>"100000000",
  52857=>"100000111",
  52858=>"000000000",
  52859=>"000000000",
  52860=>"000000001",
  52861=>"010000000",
  52862=>"110000000",
  52863=>"111000000",
  52864=>"111111011",
  52865=>"111111111",
  52866=>"011010110",
  52867=>"001000100",
  52868=>"010000000",
  52869=>"000100000",
  52870=>"111111111",
  52871=>"110111111",
  52872=>"000001011",
  52873=>"111111000",
  52874=>"111111111",
  52875=>"100100111",
  52876=>"100000111",
  52877=>"111111110",
  52878=>"111111111",
  52879=>"101111101",
  52880=>"011111001",
  52881=>"000000000",
  52882=>"111010000",
  52883=>"111111011",
  52884=>"000011000",
  52885=>"110100100",
  52886=>"001000000",
  52887=>"000001111",
  52888=>"000000000",
  52889=>"000000010",
  52890=>"011111111",
  52891=>"111111111",
  52892=>"000000000",
  52893=>"101001001",
  52894=>"100111111",
  52895=>"000111111",
  52896=>"000000000",
  52897=>"111111111",
  52898=>"110110100",
  52899=>"000000101",
  52900=>"000100000",
  52901=>"101111001",
  52902=>"000001001",
  52903=>"111111100",
  52904=>"011111111",
  52905=>"001000000",
  52906=>"100000000",
  52907=>"111111111",
  52908=>"111111111",
  52909=>"000000000",
  52910=>"000010000",
  52911=>"000000111",
  52912=>"011000000",
  52913=>"100110000",
  52914=>"111111111",
  52915=>"000111000",
  52916=>"000110110",
  52917=>"001111011",
  52918=>"111111110",
  52919=>"111000000",
  52920=>"111001000",
  52921=>"011001011",
  52922=>"100100100",
  52923=>"111001011",
  52924=>"000000000",
  52925=>"001000000",
  52926=>"000110111",
  52927=>"111111011",
  52928=>"111111101",
  52929=>"000000000",
  52930=>"000000111",
  52931=>"011111111",
  52932=>"111111111",
  52933=>"000000000",
  52934=>"001011000",
  52935=>"111111111",
  52936=>"111111111",
  52937=>"000000000",
  52938=>"001101101",
  52939=>"000010010",
  52940=>"111111111",
  52941=>"110110000",
  52942=>"010000111",
  52943=>"100100110",
  52944=>"111011001",
  52945=>"000000111",
  52946=>"000000001",
  52947=>"111101111",
  52948=>"000010000",
  52949=>"000100000",
  52950=>"000000000",
  52951=>"111111111",
  52952=>"000000000",
  52953=>"111111011",
  52954=>"000000000",
  52955=>"000010010",
  52956=>"110000010",
  52957=>"001000101",
  52958=>"000011000",
  52959=>"100100000",
  52960=>"000001011",
  52961=>"000011000",
  52962=>"000111111",
  52963=>"000000000",
  52964=>"110111001",
  52965=>"100100110",
  52966=>"011001111",
  52967=>"000001111",
  52968=>"111100100",
  52969=>"000000011",
  52970=>"000000011",
  52971=>"100000000",
  52972=>"111111011",
  52973=>"000000011",
  52974=>"010000100",
  52975=>"000001111",
  52976=>"000000000",
  52977=>"000100110",
  52978=>"100000110",
  52979=>"000000000",
  52980=>"000000000",
  52981=>"111111111",
  52982=>"001011110",
  52983=>"111111111",
  52984=>"111000000",
  52985=>"110100111",
  52986=>"111111111",
  52987=>"111000000",
  52988=>"000000000",
  52989=>"111111111",
  52990=>"111111110",
  52991=>"111111111",
  52992=>"111111001",
  52993=>"011001000",
  52994=>"000000000",
  52995=>"111111111",
  52996=>"000000000",
  52997=>"110111111",
  52998=>"000000000",
  52999=>"011111111",
  53000=>"010010000",
  53001=>"111111101",
  53002=>"110100101",
  53003=>"000000001",
  53004=>"111101001",
  53005=>"010000111",
  53006=>"000000001",
  53007=>"001001000",
  53008=>"101101111",
  53009=>"100000000",
  53010=>"001000000",
  53011=>"000000000",
  53012=>"000000001",
  53013=>"000000111",
  53014=>"001011100",
  53015=>"000000000",
  53016=>"111111010",
  53017=>"111111000",
  53018=>"110110100",
  53019=>"111111111",
  53020=>"111111111",
  53021=>"000000110",
  53022=>"000000000",
  53023=>"110011011",
  53024=>"000000000",
  53025=>"011111111",
  53026=>"000000101",
  53027=>"010000000",
  53028=>"001000000",
  53029=>"000000000",
  53030=>"100011000",
  53031=>"001000100",
  53032=>"000000100",
  53033=>"111111111",
  53034=>"000000110",
  53035=>"000000011",
  53036=>"111111011",
  53037=>"011000000",
  53038=>"111010001",
  53039=>"111111111",
  53040=>"111001001",
  53041=>"000000111",
  53042=>"111111111",
  53043=>"111111111",
  53044=>"110000111",
  53045=>"010011000",
  53046=>"000000000",
  53047=>"110110111",
  53048=>"000000000",
  53049=>"000000001",
  53050=>"100000000",
  53051=>"100000000",
  53052=>"000000000",
  53053=>"000000000",
  53054=>"111100100",
  53055=>"101000000",
  53056=>"111101000",
  53057=>"111011000",
  53058=>"100000000",
  53059=>"001001100",
  53060=>"111111111",
  53061=>"111001001",
  53062=>"000000101",
  53063=>"000000000",
  53064=>"100000000",
  53065=>"011111111",
  53066=>"000111000",
  53067=>"110110110",
  53068=>"111111000",
  53069=>"000000000",
  53070=>"100000000",
  53071=>"111110000",
  53072=>"110110100",
  53073=>"000000001",
  53074=>"000000100",
  53075=>"111110111",
  53076=>"011001111",
  53077=>"111111111",
  53078=>"011000111",
  53079=>"111111111",
  53080=>"111111111",
  53081=>"111111111",
  53082=>"111111111",
  53083=>"100000111",
  53084=>"011001001",
  53085=>"111110010",
  53086=>"000110111",
  53087=>"000111111",
  53088=>"000000000",
  53089=>"000000000",
  53090=>"001000000",
  53091=>"111001001",
  53092=>"111111011",
  53093=>"000000000",
  53094=>"110100110",
  53095=>"000000100",
  53096=>"001111111",
  53097=>"000000111",
  53098=>"000000100",
  53099=>"111111011",
  53100=>"000000000",
  53101=>"011111000",
  53102=>"111000000",
  53103=>"111111111",
  53104=>"000000000",
  53105=>"000000000",
  53106=>"000000010",
  53107=>"111111100",
  53108=>"101111100",
  53109=>"000000110",
  53110=>"110000000",
  53111=>"000000111",
  53112=>"101001111",
  53113=>"000000000",
  53114=>"011000000",
  53115=>"001111111",
  53116=>"000111111",
  53117=>"000000000",
  53118=>"111111111",
  53119=>"000100100",
  53120=>"001001011",
  53121=>"100110000",
  53122=>"000000001",
  53123=>"111000000",
  53124=>"000111111",
  53125=>"011000000",
  53126=>"001000000",
  53127=>"111111111",
  53128=>"001000001",
  53129=>"111111111",
  53130=>"111111111",
  53131=>"001111111",
  53132=>"111111111",
  53133=>"101100100",
  53134=>"000000000",
  53135=>"111111111",
  53136=>"000000000",
  53137=>"111111111",
  53138=>"000000001",
  53139=>"000000100",
  53140=>"000000011",
  53141=>"000000000",
  53142=>"111111111",
  53143=>"111010000",
  53144=>"000111111",
  53145=>"101100101",
  53146=>"111111111",
  53147=>"110111111",
  53148=>"001010111",
  53149=>"111111010",
  53150=>"011000000",
  53151=>"111100110",
  53152=>"111111111",
  53153=>"000001001",
  53154=>"101000001",
  53155=>"000000000",
  53156=>"000011111",
  53157=>"010010000",
  53158=>"000000111",
  53159=>"000000000",
  53160=>"000000000",
  53161=>"000001011",
  53162=>"111001111",
  53163=>"011011010",
  53164=>"000000000",
  53165=>"000000000",
  53166=>"111100101",
  53167=>"100101101",
  53168=>"100000101",
  53169=>"000000101",
  53170=>"000010000",
  53171=>"000010111",
  53172=>"000000000",
  53173=>"000000100",
  53174=>"111111111",
  53175=>"111111111",
  53176=>"000110111",
  53177=>"111001000",
  53178=>"000100000",
  53179=>"100100100",
  53180=>"000000000",
  53181=>"110000000",
  53182=>"000000001",
  53183=>"111111011",
  53184=>"000010000",
  53185=>"000001000",
  53186=>"111000011",
  53187=>"111111010",
  53188=>"111111010",
  53189=>"111111111",
  53190=>"000011000",
  53191=>"011011011",
  53192=>"000000000",
  53193=>"111111000",
  53194=>"011110111",
  53195=>"110110110",
  53196=>"000111000",
  53197=>"000000000",
  53198=>"000010000",
  53199=>"100101000",
  53200=>"000001011",
  53201=>"001101100",
  53202=>"111111111",
  53203=>"000000000",
  53204=>"111111111",
  53205=>"001000001",
  53206=>"000000101",
  53207=>"111001000",
  53208=>"000000000",
  53209=>"111111111",
  53210=>"001000111",
  53211=>"111111111",
  53212=>"111111100",
  53213=>"000010011",
  53214=>"000000011",
  53215=>"000000100",
  53216=>"001011010",
  53217=>"011001100",
  53218=>"111111011",
  53219=>"000000001",
  53220=>"000000000",
  53221=>"111000000",
  53222=>"001011000",
  53223=>"000000000",
  53224=>"111111111",
  53225=>"111111110",
  53226=>"000000000",
  53227=>"111111101",
  53228=>"000000000",
  53229=>"110110110",
  53230=>"000000101",
  53231=>"111111111",
  53232=>"000000100",
  53233=>"111010010",
  53234=>"000000001",
  53235=>"111111111",
  53236=>"000010011",
  53237=>"000111000",
  53238=>"000100110",
  53239=>"100100000",
  53240=>"001000000",
  53241=>"111111111",
  53242=>"011011111",
  53243=>"000000000",
  53244=>"000000100",
  53245=>"011111111",
  53246=>"000111110",
  53247=>"111111111",
  53248=>"000000001",
  53249=>"110000111",
  53250=>"001000000",
  53251=>"011001000",
  53252=>"100010000",
  53253=>"000000001",
  53254=>"111000101",
  53255=>"000000000",
  53256=>"000000001",
  53257=>"111111111",
  53258=>"111111110",
  53259=>"111111111",
  53260=>"101001111",
  53261=>"111000000",
  53262=>"011001001",
  53263=>"110110110",
  53264=>"000111111",
  53265=>"001001101",
  53266=>"110111111",
  53267=>"000000000",
  53268=>"111110011",
  53269=>"000000000",
  53270=>"000000000",
  53271=>"100110111",
  53272=>"111111111",
  53273=>"111110000",
  53274=>"100000000",
  53275=>"101111110",
  53276=>"110100000",
  53277=>"000000100",
  53278=>"000000000",
  53279=>"000000000",
  53280=>"100000100",
  53281=>"111111000",
  53282=>"000110110",
  53283=>"000000001",
  53284=>"111111111",
  53285=>"101100111",
  53286=>"111110110",
  53287=>"110100000",
  53288=>"101110111",
  53289=>"000000000",
  53290=>"111101001",
  53291=>"000000100",
  53292=>"111111111",
  53293=>"000000000",
  53294=>"000000001",
  53295=>"111111000",
  53296=>"100000000",
  53297=>"111111000",
  53298=>"000000000",
  53299=>"010000101",
  53300=>"000000000",
  53301=>"111110100",
  53302=>"100101111",
  53303=>"001001000",
  53304=>"001001111",
  53305=>"000101111",
  53306=>"110110000",
  53307=>"000000000",
  53308=>"000000000",
  53309=>"110110110",
  53310=>"000000001",
  53311=>"111111000",
  53312=>"111111101",
  53313=>"010011000",
  53314=>"010010000",
  53315=>"111111001",
  53316=>"111111111",
  53317=>"111111110",
  53318=>"000000000",
  53319=>"001000111",
  53320=>"101000001",
  53321=>"001001111",
  53322=>"000000000",
  53323=>"011111111",
  53324=>"000000000",
  53325=>"001000000",
  53326=>"101000001",
  53327=>"100110110",
  53328=>"111001000",
  53329=>"000000010",
  53330=>"111110000",
  53331=>"110110111",
  53332=>"000000000",
  53333=>"111111111",
  53334=>"101111111",
  53335=>"111111100",
  53336=>"000011111",
  53337=>"000000000",
  53338=>"111111100",
  53339=>"111111110",
  53340=>"011011111",
  53341=>"111111111",
  53342=>"111111001",
  53343=>"111100000",
  53344=>"000000000",
  53345=>"001001001",
  53346=>"101000000",
  53347=>"100000000",
  53348=>"111110110",
  53349=>"111001000",
  53350=>"111111111",
  53351=>"011001000",
  53352=>"000000000",
  53353=>"010111111",
  53354=>"111111000",
  53355=>"111111000",
  53356=>"000000000",
  53357=>"000000101",
  53358=>"000000000",
  53359=>"111100000",
  53360=>"011000001",
  53361=>"000000111",
  53362=>"100000101",
  53363=>"001001011",
  53364=>"010010000",
  53365=>"001011111",
  53366=>"000000000",
  53367=>"001111111",
  53368=>"100000100",
  53369=>"111100000",
  53370=>"001000001",
  53371=>"000000000",
  53372=>"110110110",
  53373=>"111111000",
  53374=>"001000000",
  53375=>"001000011",
  53376=>"111101000",
  53377=>"111111111",
  53378=>"111100000",
  53379=>"000100000",
  53380=>"000000000",
  53381=>"111111111",
  53382=>"000000000",
  53383=>"000000010",
  53384=>"111111111",
  53385=>"001000100",
  53386=>"111110110",
  53387=>"000000001",
  53388=>"011111111",
  53389=>"000011011",
  53390=>"111110000",
  53391=>"111111111",
  53392=>"000011000",
  53393=>"000010000",
  53394=>"111111000",
  53395=>"111111111",
  53396=>"000000000",
  53397=>"111111110",
  53398=>"111111111",
  53399=>"000000000",
  53400=>"000000000",
  53401=>"111111111",
  53402=>"111111111",
  53403=>"000000000",
  53404=>"111000000",
  53405=>"000000111",
  53406=>"111110111",
  53407=>"011111111",
  53408=>"000000000",
  53409=>"111001011",
  53410=>"000000111",
  53411=>"111111111",
  53412=>"011001111",
  53413=>"111110110",
  53414=>"001111000",
  53415=>"111011000",
  53416=>"111111011",
  53417=>"111101111",
  53418=>"111111111",
  53419=>"000000000",
  53420=>"110111000",
  53421=>"110100100",
  53422=>"001011011",
  53423=>"110011111",
  53424=>"000111111",
  53425=>"110110111",
  53426=>"000110000",
  53427=>"111111101",
  53428=>"111010000",
  53429=>"111111111",
  53430=>"000000000",
  53431=>"000001001",
  53432=>"100100101",
  53433=>"011111111",
  53434=>"011000000",
  53435=>"001000000",
  53436=>"111111111",
  53437=>"111111111",
  53438=>"011000111",
  53439=>"111111111",
  53440=>"000000000",
  53441=>"000000000",
  53442=>"000011111",
  53443=>"000010000",
  53444=>"010111111",
  53445=>"000000000",
  53446=>"001000000",
  53447=>"111111111",
  53448=>"000000000",
  53449=>"111111111",
  53450=>"000000000",
  53451=>"111111110",
  53452=>"101101111",
  53453=>"000111010",
  53454=>"111111111",
  53455=>"111000101",
  53456=>"000001001",
  53457=>"000000110",
  53458=>"100110110",
  53459=>"111101001",
  53460=>"000111011",
  53461=>"111111111",
  53462=>"000000000",
  53463=>"000000111",
  53464=>"111111011",
  53465=>"010010100",
  53466=>"000000111",
  53467=>"000000000",
  53468=>"101111111",
  53469=>"101000111",
  53470=>"000000000",
  53471=>"111111100",
  53472=>"000000000",
  53473=>"111011011",
  53474=>"111111000",
  53475=>"011011001",
  53476=>"000000001",
  53477=>"011010000",
  53478=>"000111111",
  53479=>"111111111",
  53480=>"000000000",
  53481=>"000000000",
  53482=>"000000000",
  53483=>"111111111",
  53484=>"111111100",
  53485=>"000011010",
  53486=>"111111111",
  53487=>"110110111",
  53488=>"000000000",
  53489=>"111111111",
  53490=>"111111111",
  53491=>"011000000",
  53492=>"000000000",
  53493=>"110110110",
  53494=>"001000000",
  53495=>"000001101",
  53496=>"011001000",
  53497=>"000000000",
  53498=>"000000000",
  53499=>"000000000",
  53500=>"000000000",
  53501=>"000100100",
  53502=>"010110111",
  53503=>"011111111",
  53504=>"000000000",
  53505=>"111101111",
  53506=>"110000111",
  53507=>"111010010",
  53508=>"110111111",
  53509=>"000000000",
  53510=>"001001111",
  53511=>"111111111",
  53512=>"000000001",
  53513=>"000000000",
  53514=>"000000000",
  53515=>"011000101",
  53516=>"100000000",
  53517=>"100001001",
  53518=>"111100111",
  53519=>"111111111",
  53520=>"111001101",
  53521=>"000000000",
  53522=>"000000001",
  53523=>"000000111",
  53524=>"111000000",
  53525=>"001111111",
  53526=>"101101111",
  53527=>"110110111",
  53528=>"000000000",
  53529=>"111111011",
  53530=>"000000000",
  53531=>"010010011",
  53532=>"111111111",
  53533=>"010000000",
  53534=>"000000000",
  53535=>"001000010",
  53536=>"000000000",
  53537=>"000110001",
  53538=>"111000100",
  53539=>"111111011",
  53540=>"110100100",
  53541=>"001001111",
  53542=>"110110111",
  53543=>"010000111",
  53544=>"101000000",
  53545=>"000001000",
  53546=>"000010111",
  53547=>"111000000",
  53548=>"000001101",
  53549=>"100100100",
  53550=>"111110111",
  53551=>"000000000",
  53552=>"111111110",
  53553=>"001001001",
  53554=>"110100110",
  53555=>"111001000",
  53556=>"111111000",
  53557=>"000000000",
  53558=>"111000000",
  53559=>"001000111",
  53560=>"000000000",
  53561=>"001001011",
  53562=>"111111110",
  53563=>"000000000",
  53564=>"000000000",
  53565=>"000111110",
  53566=>"110110000",
  53567=>"000000000",
  53568=>"111111111",
  53569=>"000000000",
  53570=>"111111111",
  53571=>"111111111",
  53572=>"000000111",
  53573=>"000110110",
  53574=>"000000000",
  53575=>"000110110",
  53576=>"000000100",
  53577=>"000110111",
  53578=>"011000100",
  53579=>"010010100",
  53580=>"000000100",
  53581=>"111111011",
  53582=>"000100110",
  53583=>"110010000",
  53584=>"010010000",
  53585=>"100100000",
  53586=>"111001101",
  53587=>"110000000",
  53588=>"111111100",
  53589=>"001001000",
  53590=>"000000000",
  53591=>"101111000",
  53592=>"000101111",
  53593=>"100110100",
  53594=>"111111011",
  53595=>"111111111",
  53596=>"110110110",
  53597=>"111111001",
  53598=>"000000000",
  53599=>"101100100",
  53600=>"000000011",
  53601=>"111111111",
  53602=>"000000000",
  53603=>"110110111",
  53604=>"111111100",
  53605=>"001111000",
  53606=>"000000111",
  53607=>"111110111",
  53608=>"111111111",
  53609=>"010011111",
  53610=>"110110100",
  53611=>"000000000",
  53612=>"111111111",
  53613=>"001001000",
  53614=>"111010000",
  53615=>"000000000",
  53616=>"000000000",
  53617=>"011001111",
  53618=>"001000001",
  53619=>"111111111",
  53620=>"111111001",
  53621=>"000010111",
  53622=>"001000100",
  53623=>"111111111",
  53624=>"111111001",
  53625=>"000000000",
  53626=>"000000000",
  53627=>"111111110",
  53628=>"000000111",
  53629=>"101111110",
  53630=>"111101111",
  53631=>"111111111",
  53632=>"000000110",
  53633=>"111011111",
  53634=>"111111000",
  53635=>"000001011",
  53636=>"000000111",
  53637=>"000000000",
  53638=>"000000101",
  53639=>"110100100",
  53640=>"000000000",
  53641=>"000000000",
  53642=>"111011001",
  53643=>"011001011",
  53644=>"111110111",
  53645=>"111111111",
  53646=>"000111111",
  53647=>"111111111",
  53648=>"000000000",
  53649=>"110000000",
  53650=>"000000000",
  53651=>"000000000",
  53652=>"111111111",
  53653=>"000000000",
  53654=>"101000000",
  53655=>"101111000",
  53656=>"001001011",
  53657=>"011111111",
  53658=>"111111111",
  53659=>"111001111",
  53660=>"000000000",
  53661=>"100000011",
  53662=>"000000000",
  53663=>"111000000",
  53664=>"111111001",
  53665=>"101000000",
  53666=>"000000100",
  53667=>"011011001",
  53668=>"001000001",
  53669=>"111111111",
  53670=>"000000000",
  53671=>"000000101",
  53672=>"000001001",
  53673=>"110110110",
  53674=>"100000000",
  53675=>"001001000",
  53676=>"000000000",
  53677=>"001011111",
  53678=>"000000000",
  53679=>"000000111",
  53680=>"000000111",
  53681=>"011111011",
  53682=>"101011111",
  53683=>"111000000",
  53684=>"000000000",
  53685=>"000000010",
  53686=>"000000111",
  53687=>"000000000",
  53688=>"001000000",
  53689=>"000000100",
  53690=>"110000000",
  53691=>"000000000",
  53692=>"000000000",
  53693=>"000001111",
  53694=>"111111111",
  53695=>"100111101",
  53696=>"110111011",
  53697=>"000000000",
  53698=>"111111111",
  53699=>"111111111",
  53700=>"000000111",
  53701=>"000000000",
  53702=>"001000000",
  53703=>"000000111",
  53704=>"000000000",
  53705=>"011111000",
  53706=>"111111111",
  53707=>"000000111",
  53708=>"000001000",
  53709=>"000000000",
  53710=>"011101100",
  53711=>"011001111",
  53712=>"011011111",
  53713=>"000000000",
  53714=>"001101000",
  53715=>"000000000",
  53716=>"011011001",
  53717=>"000000000",
  53718=>"000000111",
  53719=>"000000000",
  53720=>"000011001",
  53721=>"000000000",
  53722=>"010111111",
  53723=>"000000000",
  53724=>"000000000",
  53725=>"111111111",
  53726=>"111111111",
  53727=>"111100100",
  53728=>"100100000",
  53729=>"011111010",
  53730=>"110111000",
  53731=>"000001001",
  53732=>"111111000",
  53733=>"000000000",
  53734=>"000000001",
  53735=>"111111000",
  53736=>"011000000",
  53737=>"111111111",
  53738=>"010000000",
  53739=>"111110010",
  53740=>"111111111",
  53741=>"011011100",
  53742=>"100000000",
  53743=>"000001111",
  53744=>"100110000",
  53745=>"001000111",
  53746=>"111011001",
  53747=>"010111110",
  53748=>"111111110",
  53749=>"000010011",
  53750=>"111111111",
  53751=>"110000111",
  53752=>"010111100",
  53753=>"000010000",
  53754=>"111111111",
  53755=>"000000000",
  53756=>"110100000",
  53757=>"111111111",
  53758=>"001011111",
  53759=>"111111111",
  53760=>"111111111",
  53761=>"111111111",
  53762=>"111111111",
  53763=>"100000100",
  53764=>"000111111",
  53765=>"001001001",
  53766=>"000000000",
  53767=>"000000000",
  53768=>"000100100",
  53769=>"111111111",
  53770=>"000000000",
  53771=>"000000110",
  53772=>"100010000",
  53773=>"111001000",
  53774=>"000000000",
  53775=>"000000000",
  53776=>"000000000",
  53777=>"000000111",
  53778=>"000000111",
  53779=>"000111111",
  53780=>"000000000",
  53781=>"000000001",
  53782=>"111001001",
  53783=>"011011001",
  53784=>"011011001",
  53785=>"110100111",
  53786=>"000011011",
  53787=>"000000100",
  53788=>"000000000",
  53789=>"001000001",
  53790=>"111111000",
  53791=>"111111111",
  53792=>"110010111",
  53793=>"100111111",
  53794=>"011001000",
  53795=>"000000011",
  53796=>"000001010",
  53797=>"000101111",
  53798=>"010111111",
  53799=>"000001000",
  53800=>"101100000",
  53801=>"000000111",
  53802=>"110111111",
  53803=>"111100111",
  53804=>"011001001",
  53805=>"011000000",
  53806=>"000000000",
  53807=>"010000000",
  53808=>"000000001",
  53809=>"110011010",
  53810=>"110000000",
  53811=>"000000110",
  53812=>"001000000",
  53813=>"111001101",
  53814=>"110111111",
  53815=>"001001000",
  53816=>"000000010",
  53817=>"111111011",
  53818=>"000000100",
  53819=>"111111000",
  53820=>"011111111",
  53821=>"000101111",
  53822=>"000000001",
  53823=>"100100110",
  53824=>"001101111",
  53825=>"111111000",
  53826=>"011011111",
  53827=>"000100111",
  53828=>"111111010",
  53829=>"000000000",
  53830=>"101111111",
  53831=>"111100110",
  53832=>"111111111",
  53833=>"001000101",
  53834=>"000000010",
  53835=>"000000000",
  53836=>"000011011",
  53837=>"101001111",
  53838=>"110000000",
  53839=>"111111111",
  53840=>"000000000",
  53841=>"000110111",
  53842=>"111000000",
  53843=>"000111111",
  53844=>"111101001",
  53845=>"000011111",
  53846=>"000000000",
  53847=>"000000111",
  53848=>"000000000",
  53849=>"000000000",
  53850=>"000000000",
  53851=>"110000111",
  53852=>"000000000",
  53853=>"000100111",
  53854=>"000000110",
  53855=>"111110100",
  53856=>"100000000",
  53857=>"000000000",
  53858=>"111111000",
  53859=>"000000111",
  53860=>"001000000",
  53861=>"001001000",
  53862=>"111111101",
  53863=>"111111111",
  53864=>"000001001",
  53865=>"000000000",
  53866=>"000010110",
  53867=>"000000000",
  53868=>"000000100",
  53869=>"000000000",
  53870=>"000000000",
  53871=>"000001110",
  53872=>"000010111",
  53873=>"111111101",
  53874=>"101111010",
  53875=>"000000000",
  53876=>"111100000",
  53877=>"011011000",
  53878=>"000000000",
  53879=>"001001011",
  53880=>"000000000",
  53881=>"100100100",
  53882=>"000000000",
  53883=>"110000000",
  53884=>"010011010",
  53885=>"011111111",
  53886=>"110011000",
  53887=>"000000000",
  53888=>"001111111",
  53889=>"110110111",
  53890=>"111000001",
  53891=>"000111111",
  53892=>"111111111",
  53893=>"101111111",
  53894=>"100100000",
  53895=>"001000000",
  53896=>"000000011",
  53897=>"111011000",
  53898=>"001111011",
  53899=>"000000000",
  53900=>"111000000",
  53901=>"000111111",
  53902=>"110100000",
  53903=>"101100110",
  53904=>"111111010",
  53905=>"111111111",
  53906=>"000000111",
  53907=>"111111111",
  53908=>"111111111",
  53909=>"111100001",
  53910=>"001001001",
  53911=>"100101100",
  53912=>"000000000",
  53913=>"001001111",
  53914=>"000010000",
  53915=>"101100100",
  53916=>"000100110",
  53917=>"000100000",
  53918=>"111101111",
  53919=>"000000000",
  53920=>"111111111",
  53921=>"100100101",
  53922=>"100000001",
  53923=>"001000000",
  53924=>"110000100",
  53925=>"111111111",
  53926=>"011111011",
  53927=>"001000010",
  53928=>"001000011",
  53929=>"111100100",
  53930=>"111111111",
  53931=>"111111000",
  53932=>"001001000",
  53933=>"100111100",
  53934=>"110000000",
  53935=>"000000000",
  53936=>"111111101",
  53937=>"000100100",
  53938=>"110110110",
  53939=>"000001001",
  53940=>"000100000",
  53941=>"000001011",
  53942=>"111111111",
  53943=>"111100000",
  53944=>"111111111",
  53945=>"111001110",
  53946=>"111000000",
  53947=>"111111110",
  53948=>"011000000",
  53949=>"111111000",
  53950=>"000111001",
  53951=>"000000000",
  53952=>"000000000",
  53953=>"000000111",
  53954=>"111110110",
  53955=>"111111011",
  53956=>"111000001",
  53957=>"111111111",
  53958=>"000111001",
  53959=>"111111111",
  53960=>"000000000",
  53961=>"000000101",
  53962=>"110000000",
  53963=>"111000110",
  53964=>"000001101",
  53965=>"000000000",
  53966=>"010000000",
  53967=>"011110000",
  53968=>"001001111",
  53969=>"011111111",
  53970=>"111001000",
  53971=>"000000000",
  53972=>"111111011",
  53973=>"110000000",
  53974=>"001011011",
  53975=>"111111000",
  53976=>"111111111",
  53977=>"000100000",
  53978=>"000000000",
  53979=>"111111111",
  53980=>"111111111",
  53981=>"111111111",
  53982=>"111110111",
  53983=>"001001011",
  53984=>"101000000",
  53985=>"000000111",
  53986=>"001001000",
  53987=>"101111111",
  53988=>"000001001",
  53989=>"000100110",
  53990=>"011110111",
  53991=>"110111000",
  53992=>"000100111",
  53993=>"111110111",
  53994=>"110110001",
  53995=>"010000000",
  53996=>"000000000",
  53997=>"001001111",
  53998=>"110000000",
  53999=>"000000000",
  54000=>"000000000",
  54001=>"111111111",
  54002=>"100110000",
  54003=>"011001111",
  54004=>"001001100",
  54005=>"111001001",
  54006=>"111100100",
  54007=>"000000001",
  54008=>"100111111",
  54009=>"111111000",
  54010=>"001000000",
  54011=>"000000001",
  54012=>"000000000",
  54013=>"001000000",
  54014=>"111100110",
  54015=>"000000100",
  54016=>"000000000",
  54017=>"011011000",
  54018=>"010000000",
  54019=>"000000000",
  54020=>"100011000",
  54021=>"111101100",
  54022=>"000100110",
  54023=>"000100111",
  54024=>"000000111",
  54025=>"111111101",
  54026=>"000001101",
  54027=>"000000110",
  54028=>"110000000",
  54029=>"100111111",
  54030=>"000111111",
  54031=>"000111011",
  54032=>"111111000",
  54033=>"111111000",
  54034=>"111000111",
  54035=>"000001000",
  54036=>"001001000",
  54037=>"111111011",
  54038=>"111111000",
  54039=>"000000101",
  54040=>"111111111",
  54041=>"001001011",
  54042=>"001000111",
  54043=>"001001000",
  54044=>"000111101",
  54045=>"100000111",
  54046=>"101001111",
  54047=>"100100101",
  54048=>"101101101",
  54049=>"010111110",
  54050=>"000011000",
  54051=>"111111010",
  54052=>"111111111",
  54053=>"000000111",
  54054=>"001010111",
  54055=>"001001001",
  54056=>"111111101",
  54057=>"010010001",
  54058=>"110111111",
  54059=>"000000000",
  54060=>"100001111",
  54061=>"010001010",
  54062=>"000001111",
  54063=>"000001111",
  54064=>"111111111",
  54065=>"001001001",
  54066=>"111111111",
  54067=>"000111110",
  54068=>"000100000",
  54069=>"000001011",
  54070=>"111111100",
  54071=>"000000000",
  54072=>"000001001",
  54073=>"101000001",
  54074=>"010000000",
  54075=>"000000001",
  54076=>"011111000",
  54077=>"111000100",
  54078=>"110111000",
  54079=>"011111010",
  54080=>"100001001",
  54081=>"111000011",
  54082=>"111111111",
  54083=>"000000000",
  54084=>"101101111",
  54085=>"000000000",
  54086=>"111000111",
  54087=>"001000001",
  54088=>"111111010",
  54089=>"000001000",
  54090=>"000000000",
  54091=>"001011011",
  54092=>"111001000",
  54093=>"000000101",
  54094=>"000000001",
  54095=>"000110100",
  54096=>"000100111",
  54097=>"000000001",
  54098=>"000000111",
  54099=>"011000000",
  54100=>"000000000",
  54101=>"000101011",
  54102=>"000000111",
  54103=>"111011111",
  54104=>"111111111",
  54105=>"111111101",
  54106=>"111111111",
  54107=>"011111111",
  54108=>"000111111",
  54109=>"110111111",
  54110=>"111000001",
  54111=>"000001111",
  54112=>"000000111",
  54113=>"000000011",
  54114=>"110111000",
  54115=>"101111001",
  54116=>"110110110",
  54117=>"001001111",
  54118=>"000000000",
  54119=>"000000001",
  54120=>"111100111",
  54121=>"000000100",
  54122=>"001101111",
  54123=>"100100000",
  54124=>"000011011",
  54125=>"111001111",
  54126=>"000000100",
  54127=>"100000000",
  54128=>"011111110",
  54129=>"000111110",
  54130=>"111111111",
  54131=>"111111011",
  54132=>"000000110",
  54133=>"000000000",
  54134=>"000000000",
  54135=>"000000111",
  54136=>"000000000",
  54137=>"000000000",
  54138=>"000000010",
  54139=>"111000001",
  54140=>"111101101",
  54141=>"111111110",
  54142=>"111111110",
  54143=>"100100100",
  54144=>"000000110",
  54145=>"111001111",
  54146=>"100000000",
  54147=>"111111111",
  54148=>"000001001",
  54149=>"000100000",
  54150=>"001000000",
  54151=>"000000010",
  54152=>"000000000",
  54153=>"111111111",
  54154=>"000000000",
  54155=>"001001001",
  54156=>"111111100",
  54157=>"111011111",
  54158=>"000011111",
  54159=>"000000000",
  54160=>"111100100",
  54161=>"000000000",
  54162=>"011000000",
  54163=>"111111110",
  54164=>"100111011",
  54165=>"001000000",
  54166=>"000100100",
  54167=>"110011111",
  54168=>"000000111",
  54169=>"001000000",
  54170=>"111000000",
  54171=>"000000011",
  54172=>"010111111",
  54173=>"111111100",
  54174=>"111111111",
  54175=>"000000000",
  54176=>"001000001",
  54177=>"000111011",
  54178=>"001001100",
  54179=>"001001000",
  54180=>"101001101",
  54181=>"111111111",
  54182=>"000000011",
  54183=>"010111111",
  54184=>"000000000",
  54185=>"000001111",
  54186=>"000011000",
  54187=>"111101100",
  54188=>"111111111",
  54189=>"111111001",
  54190=>"000000111",
  54191=>"111101101",
  54192=>"000001000",
  54193=>"111111111",
  54194=>"111000111",
  54195=>"000000010",
  54196=>"111110111",
  54197=>"101000000",
  54198=>"100100000",
  54199=>"000000111",
  54200=>"000000010",
  54201=>"000000111",
  54202=>"000000001",
  54203=>"111111111",
  54204=>"001011111",
  54205=>"111111111",
  54206=>"011000000",
  54207=>"110000000",
  54208=>"000000000",
  54209=>"011111111",
  54210=>"000000000",
  54211=>"000001011",
  54212=>"000100100",
  54213=>"110000001",
  54214=>"110111111",
  54215=>"111111111",
  54216=>"000000000",
  54217=>"111111100",
  54218=>"000000000",
  54219=>"000000000",
  54220=>"100000000",
  54221=>"000111111",
  54222=>"000000010",
  54223=>"000000001",
  54224=>"000000000",
  54225=>"011111000",
  54226=>"011001010",
  54227=>"000110111",
  54228=>"111111000",
  54229=>"000111100",
  54230=>"000000000",
  54231=>"000000000",
  54232=>"000011111",
  54233=>"101001111",
  54234=>"000000001",
  54235=>"011100100",
  54236=>"101101111",
  54237=>"111000100",
  54238=>"110100111",
  54239=>"110000000",
  54240=>"000000011",
  54241=>"111101111",
  54242=>"010000001",
  54243=>"000000001",
  54244=>"111111111",
  54245=>"111001000",
  54246=>"111111000",
  54247=>"001000001",
  54248=>"000000111",
  54249=>"111111111",
  54250=>"010110110",
  54251=>"001001110",
  54252=>"000100101",
  54253=>"011011001",
  54254=>"000110110",
  54255=>"000011111",
  54256=>"111111110",
  54257=>"111000011",
  54258=>"111111011",
  54259=>"000011111",
  54260=>"111111000",
  54261=>"101000001",
  54262=>"111111001",
  54263=>"000000100",
  54264=>"000100111",
  54265=>"111100100",
  54266=>"001000101",
  54267=>"000000000",
  54268=>"101101101",
  54269=>"110101001",
  54270=>"001111110",
  54271=>"000100100",
  54272=>"111111111",
  54273=>"000010010",
  54274=>"111111111",
  54275=>"011111111",
  54276=>"100000000",
  54277=>"010000000",
  54278=>"000100100",
  54279=>"110110110",
  54280=>"111101000",
  54281=>"110000000",
  54282=>"000000000",
  54283=>"111011111",
  54284=>"011111111",
  54285=>"001001000",
  54286=>"000000111",
  54287=>"111011000",
  54288=>"110100000",
  54289=>"010000000",
  54290=>"001101110",
  54291=>"111110111",
  54292=>"000111001",
  54293=>"000000000",
  54294=>"111111111",
  54295=>"100110001",
  54296=>"100000000",
  54297=>"111111111",
  54298=>"000000001",
  54299=>"001001000",
  54300=>"000001000",
  54301=>"111101001",
  54302=>"000000010",
  54303=>"111111100",
  54304=>"100110001",
  54305=>"110111111",
  54306=>"110110110",
  54307=>"101111111",
  54308=>"000000000",
  54309=>"001011001",
  54310=>"000000000",
  54311=>"000000000",
  54312=>"100101001",
  54313=>"100111000",
  54314=>"000000000",
  54315=>"111111110",
  54316=>"000000000",
  54317=>"001000111",
  54318=>"110111111",
  54319=>"111111111",
  54320=>"100110000",
  54321=>"100000000",
  54322=>"001111111",
  54323=>"100111111",
  54324=>"000100111",
  54325=>"000110111",
  54326=>"101101000",
  54327=>"100100100",
  54328=>"000000000",
  54329=>"000001000",
  54330=>"000000000",
  54331=>"001011010",
  54332=>"101000000",
  54333=>"111111011",
  54334=>"111000000",
  54335=>"000000110",
  54336=>"011111110",
  54337=>"000000000",
  54338=>"000100110",
  54339=>"111111111",
  54340=>"000000110",
  54341=>"110011011",
  54342=>"111000000",
  54343=>"111111111",
  54344=>"111111000",
  54345=>"000000000",
  54346=>"111001001",
  54347=>"000000111",
  54348=>"111111100",
  54349=>"000010000",
  54350=>"100110110",
  54351=>"111001111",
  54352=>"000000110",
  54353=>"001000000",
  54354=>"111111000",
  54355=>"011011000",
  54356=>"111111000",
  54357=>"000010010",
  54358=>"000000111",
  54359=>"000000000",
  54360=>"111111111",
  54361=>"000000111",
  54362=>"000101100",
  54363=>"001001001",
  54364=>"100101111",
  54365=>"000000111",
  54366=>"001110110",
  54367=>"111111111",
  54368=>"000100000",
  54369=>"111010110",
  54370=>"111111011",
  54371=>"000000111",
  54372=>"000100100",
  54373=>"111111111",
  54374=>"000100111",
  54375=>"000000111",
  54376=>"100000000",
  54377=>"111111111",
  54378=>"000000000",
  54379=>"001001000",
  54380=>"000001111",
  54381=>"110111111",
  54382=>"000001000",
  54383=>"000000000",
  54384=>"000000111",
  54385=>"001000000",
  54386=>"110000000",
  54387=>"010000000",
  54388=>"011011001",
  54389=>"001000000",
  54390=>"111111000",
  54391=>"000000000",
  54392=>"000000100",
  54393=>"000000000",
  54394=>"100111111",
  54395=>"000000000",
  54396=>"000100100",
  54397=>"000000000",
  54398=>"000000000",
  54399=>"011111110",
  54400=>"000000000",
  54401=>"110010110",
  54402=>"110000011",
  54403=>"111110000",
  54404=>"000000001",
  54405=>"101001000",
  54406=>"001111111",
  54407=>"111111111",
  54408=>"001001101",
  54409=>"000000000",
  54410=>"100100000",
  54411=>"110111111",
  54412=>"000000101",
  54413=>"001011011",
  54414=>"111110110",
  54415=>"000100110",
  54416=>"011000000",
  54417=>"000000000",
  54418=>"011000000",
  54419=>"111111011",
  54420=>"000010000",
  54421=>"000000000",
  54422=>"000000001",
  54423=>"111111111",
  54424=>"100111111",
  54425=>"100000101",
  54426=>"101111111",
  54427=>"000001011",
  54428=>"111111111",
  54429=>"111111111",
  54430=>"100000101",
  54431=>"111110000",
  54432=>"111111111",
  54433=>"000100111",
  54434=>"000000111",
  54435=>"111111001",
  54436=>"000110111",
  54437=>"111011000",
  54438=>"110111111",
  54439=>"011011010",
  54440=>"001111111",
  54441=>"111011111",
  54442=>"111000000",
  54443=>"011111111",
  54444=>"011010000",
  54445=>"000000000",
  54446=>"000000000",
  54447=>"111111111",
  54448=>"000000000",
  54449=>"110100000",
  54450=>"111110110",
  54451=>"111101101",
  54452=>"111111111",
  54453=>"100100000",
  54454=>"000000000",
  54455=>"000000000",
  54456=>"111111111",
  54457=>"000000111",
  54458=>"000000111",
  54459=>"111110100",
  54460=>"011011000",
  54461=>"111111001",
  54462=>"000000000",
  54463=>"001101001",
  54464=>"111111111",
  54465=>"000000111",
  54466=>"100100101",
  54467=>"111111111",
  54468=>"000000000",
  54469=>"000000111",
  54470=>"000111111",
  54471=>"010010100",
  54472=>"100000000",
  54473=>"111111111",
  54474=>"111001001",
  54475=>"000000000",
  54476=>"000000000",
  54477=>"111111111",
  54478=>"111100110",
  54479=>"111111111",
  54480=>"111011011",
  54481=>"000110111",
  54482=>"111111011",
  54483=>"000000000",
  54484=>"000000000",
  54485=>"111000000",
  54486=>"111110100",
  54487=>"010010110",
  54488=>"010010000",
  54489=>"100110110",
  54490=>"111111000",
  54491=>"111111111",
  54492=>"111011001",
  54493=>"000111111",
  54494=>"010010010",
  54495=>"000000000",
  54496=>"000001111",
  54497=>"111111111",
  54498=>"000000000",
  54499=>"111110000",
  54500=>"111111111",
  54501=>"100010010",
  54502=>"111111111",
  54503=>"000111111",
  54504=>"111111000",
  54505=>"111111111",
  54506=>"000100100",
  54507=>"011011111",
  54508=>"000000000",
  54509=>"011111011",
  54510=>"111010111",
  54511=>"000000111",
  54512=>"100100110",
  54513=>"100000000",
  54514=>"100100101",
  54515=>"001011111",
  54516=>"001011100",
  54517=>"111011011",
  54518=>"110110100",
  54519=>"111111000",
  54520=>"000000000",
  54521=>"111011011",
  54522=>"111111111",
  54523=>"100000000",
  54524=>"001000000",
  54525=>"111111111",
  54526=>"001000000",
  54527=>"001111111",
  54528=>"111110100",
  54529=>"011011011",
  54530=>"111110110",
  54531=>"011011111",
  54532=>"000100100",
  54533=>"000000000",
  54534=>"111111111",
  54535=>"001001100",
  54536=>"000000000",
  54537=>"000110000",
  54538=>"100000000",
  54539=>"101111111",
  54540=>"111101111",
  54541=>"000000111",
  54542=>"111111111",
  54543=>"011001111",
  54544=>"011111011",
  54545=>"100100000",
  54546=>"011000101",
  54547=>"000100100",
  54548=>"111111110",
  54549=>"010010100",
  54550=>"011011001",
  54551=>"000000000",
  54552=>"111111110",
  54553=>"000000000",
  54554=>"010010010",
  54555=>"111110100",
  54556=>"000000110",
  54557=>"000000000",
  54558=>"111111000",
  54559=>"000000000",
  54560=>"001100000",
  54561=>"000000000",
  54562=>"111111000",
  54563=>"111111100",
  54564=>"111111111",
  54565=>"110111000",
  54566=>"110110110",
  54567=>"101111111",
  54568=>"000000000",
  54569=>"000000110",
  54570=>"100110110",
  54571=>"111111111",
  54572=>"111000000",
  54573=>"000000000",
  54574=>"000001000",
  54575=>"000000001",
  54576=>"010000000",
  54577=>"111011111",
  54578=>"000010000",
  54579=>"111111111",
  54580=>"001001100",
  54581=>"111000000",
  54582=>"111111000",
  54583=>"000000000",
  54584=>"000000110",
  54585=>"001000101",
  54586=>"111001001",
  54587=>"111101111",
  54588=>"000000000",
  54589=>"111101101",
  54590=>"000000010",
  54591=>"111100111",
  54592=>"000000011",
  54593=>"111111111",
  54594=>"000000000",
  54595=>"000000000",
  54596=>"110110111",
  54597=>"111111111",
  54598=>"111111001",
  54599=>"101101100",
  54600=>"011011111",
  54601=>"000111111",
  54602=>"100111111",
  54603=>"000000100",
  54604=>"111010010",
  54605=>"000010111",
  54606=>"000000011",
  54607=>"101111111",
  54608=>"100100100",
  54609=>"000100111",
  54610=>"111111111",
  54611=>"100111000",
  54612=>"000000000",
  54613=>"011011011",
  54614=>"001001000",
  54615=>"011001011",
  54616=>"111100101",
  54617=>"000001111",
  54618=>"111111011",
  54619=>"111111111",
  54620=>"111111111",
  54621=>"111000000",
  54622=>"001011111",
  54623=>"111000111",
  54624=>"000000000",
  54625=>"111011111",
  54626=>"101001000",
  54627=>"100100100",
  54628=>"100100110",
  54629=>"000001000",
  54630=>"001001000",
  54631=>"111111111",
  54632=>"000000011",
  54633=>"111111001",
  54634=>"000000000",
  54635=>"111101111",
  54636=>"100000010",
  54637=>"000000111",
  54638=>"000010010",
  54639=>"111111111",
  54640=>"000000000",
  54641=>"001000000",
  54642=>"111101011",
  54643=>"011011111",
  54644=>"111100000",
  54645=>"111111111",
  54646=>"000000100",
  54647=>"111011010",
  54648=>"000000000",
  54649=>"000000000",
  54650=>"111000000",
  54651=>"001011010",
  54652=>"111111111",
  54653=>"010111111",
  54654=>"000011111",
  54655=>"000100110",
  54656=>"000000000",
  54657=>"000000011",
  54658=>"001000100",
  54659=>"000001011",
  54660=>"000000000",
  54661=>"100100111",
  54662=>"111011011",
  54663=>"100000000",
  54664=>"010010111",
  54665=>"111001100",
  54666=>"111111111",
  54667=>"000000000",
  54668=>"111111111",
  54669=>"001000001",
  54670=>"000111111",
  54671=>"111111000",
  54672=>"111000000",
  54673=>"001000000",
  54674=>"000000000",
  54675=>"000000000",
  54676=>"111000000",
  54677=>"000000000",
  54678=>"110111111",
  54679=>"110110001",
  54680=>"000100000",
  54681=>"011011000",
  54682=>"010010110",
  54683=>"000000000",
  54684=>"011010000",
  54685=>"011011000",
  54686=>"110111111",
  54687=>"000000000",
  54688=>"100110100",
  54689=>"110110110",
  54690=>"000000100",
  54691=>"111111111",
  54692=>"111111111",
  54693=>"000000000",
  54694=>"111111111",
  54695=>"110010010",
  54696=>"111111111",
  54697=>"111000000",
  54698=>"111001111",
  54699=>"000000000",
  54700=>"000100100",
  54701=>"000000110",
  54702=>"111111111",
  54703=>"111111111",
  54704=>"000111111",
  54705=>"111111010",
  54706=>"101101000",
  54707=>"111111111",
  54708=>"110111111",
  54709=>"111111101",
  54710=>"111110111",
  54711=>"111111011",
  54712=>"000110100",
  54713=>"111111111",
  54714=>"100111111",
  54715=>"000000111",
  54716=>"111111111",
  54717=>"101001111",
  54718=>"110100111",
  54719=>"111111011",
  54720=>"111111111",
  54721=>"111101000",
  54722=>"111111111",
  54723=>"000000000",
  54724=>"100000001",
  54725=>"111111100",
  54726=>"110010110",
  54727=>"111110111",
  54728=>"100100100",
  54729=>"101000000",
  54730=>"111001111",
  54731=>"000000000",
  54732=>"111110000",
  54733=>"111010000",
  54734=>"010010011",
  54735=>"011011010",
  54736=>"000000110",
  54737=>"100100110",
  54738=>"000100110",
  54739=>"111111100",
  54740=>"011001010",
  54741=>"111111111",
  54742=>"011111111",
  54743=>"110111111",
  54744=>"110100000",
  54745=>"100000000",
  54746=>"000001000",
  54747=>"111111111",
  54748=>"000111011",
  54749=>"001001001",
  54750=>"001111111",
  54751=>"001000000",
  54752=>"110011111",
  54753=>"000000010",
  54754=>"110111100",
  54755=>"000000111",
  54756=>"111111111",
  54757=>"011011011",
  54758=>"111000000",
  54759=>"011010000",
  54760=>"100000000",
  54761=>"110100000",
  54762=>"000000000",
  54763=>"000100110",
  54764=>"100110110",
  54765=>"011000000",
  54766=>"000000000",
  54767=>"100000000",
  54768=>"001011011",
  54769=>"000000000",
  54770=>"001100010",
  54771=>"000000000",
  54772=>"000000000",
  54773=>"100000010",
  54774=>"111010011",
  54775=>"011111111",
  54776=>"100100100",
  54777=>"100100100",
  54778=>"100000000",
  54779=>"111111111",
  54780=>"111110011",
  54781=>"110010000",
  54782=>"100000111",
  54783=>"000000100",
  54784=>"001110000",
  54785=>"111000111",
  54786=>"111000101",
  54787=>"000100111",
  54788=>"101000000",
  54789=>"111000000",
  54790=>"000010111",
  54791=>"111000000",
  54792=>"111111011",
  54793=>"000000000",
  54794=>"111111111",
  54795=>"000001111",
  54796=>"000110111",
  54797=>"111111111",
  54798=>"111111001",
  54799=>"111111010",
  54800=>"110111111",
  54801=>"000000111",
  54802=>"010110111",
  54803=>"111000000",
  54804=>"111011000",
  54805=>"101100000",
  54806=>"111111110",
  54807=>"000111111",
  54808=>"100000000",
  54809=>"001000110",
  54810=>"000000000",
  54811=>"000000110",
  54812=>"110100000",
  54813=>"111111001",
  54814=>"000000000",
  54815=>"111111000",
  54816=>"011011111",
  54817=>"110111000",
  54818=>"111000000",
  54819=>"101001111",
  54820=>"000000000",
  54821=>"100000000",
  54822=>"101110110",
  54823=>"101111111",
  54824=>"100000111",
  54825=>"000111000",
  54826=>"111111110",
  54827=>"111111111",
  54828=>"000000111",
  54829=>"111000111",
  54830=>"000111111",
  54831=>"001111111",
  54832=>"111100000",
  54833=>"000000000",
  54834=>"000111000",
  54835=>"111100000",
  54836=>"000101000",
  54837=>"010011110",
  54838=>"111100110",
  54839=>"111110110",
  54840=>"001011001",
  54841=>"111111001",
  54842=>"111111111",
  54843=>"000001011",
  54844=>"111000000",
  54845=>"111111110",
  54846=>"000001101",
  54847=>"111111000",
  54848=>"100111010",
  54849=>"100111000",
  54850=>"000000111",
  54851=>"111111000",
  54852=>"111111010",
  54853=>"001000110",
  54854=>"000001000",
  54855=>"011000000",
  54856=>"000111111",
  54857=>"111001111",
  54858=>"111001111",
  54859=>"111000000",
  54860=>"111110100",
  54861=>"100100000",
  54862=>"111000000",
  54863=>"111111111",
  54864=>"101110110",
  54865=>"001001111",
  54866=>"000001001",
  54867=>"111110111",
  54868=>"110000000",
  54869=>"111110111",
  54870=>"100100110",
  54871=>"010111010",
  54872=>"111000111",
  54873=>"000000000",
  54874=>"111111001",
  54875=>"000001111",
  54876=>"000000000",
  54877=>"111111111",
  54878=>"101000001",
  54879=>"011011011",
  54880=>"111000000",
  54881=>"111100000",
  54882=>"100000111",
  54883=>"000000000",
  54884=>"110100100",
  54885=>"000000011",
  54886=>"111111111",
  54887=>"110100101",
  54888=>"111000000",
  54889=>"111000000",
  54890=>"111010000",
  54891=>"000001111",
  54892=>"011010010",
  54893=>"111011010",
  54894=>"100000111",
  54895=>"000000000",
  54896=>"111000010",
  54897=>"101000111",
  54898=>"001001000",
  54899=>"111100111",
  54900=>"000000001",
  54901=>"111100000",
  54902=>"111000000",
  54903=>"000010110",
  54904=>"000111000",
  54905=>"011000000",
  54906=>"000000000",
  54907=>"000000001",
  54908=>"110111000",
  54909=>"000000001",
  54910=>"000000000",
  54911=>"111111111",
  54912=>"001000011",
  54913=>"111001010",
  54914=>"010010110",
  54915=>"101011111",
  54916=>"000111111",
  54917=>"100000000",
  54918=>"111000001",
  54919=>"111010111",
  54920=>"111110110",
  54921=>"000000001",
  54922=>"111111011",
  54923=>"110000111",
  54924=>"000001111",
  54925=>"001000001",
  54926=>"111111101",
  54927=>"000000000",
  54928=>"000000111",
  54929=>"000000000",
  54930=>"100111000",
  54931=>"001110111",
  54932=>"111111000",
  54933=>"000100111",
  54934=>"111101111",
  54935=>"001000111",
  54936=>"011000111",
  54937=>"111111100",
  54938=>"100110111",
  54939=>"110011000",
  54940=>"111110000",
  54941=>"001000000",
  54942=>"111111111",
  54943=>"111001000",
  54944=>"110110100",
  54945=>"000000111",
  54946=>"011000111",
  54947=>"111111001",
  54948=>"000000000",
  54949=>"111000001",
  54950=>"110000000",
  54951=>"000111111",
  54952=>"000000001",
  54953=>"000000000",
  54954=>"100100000",
  54955=>"111000111",
  54956=>"110111111",
  54957=>"100111000",
  54958=>"000000110",
  54959=>"000001111",
  54960=>"111111001",
  54961=>"000001011",
  54962=>"010010011",
  54963=>"000000000",
  54964=>"000000111",
  54965=>"000000000",
  54966=>"111111000",
  54967=>"111111111",
  54968=>"111000000",
  54969=>"111110111",
  54970=>"000010010",
  54971=>"000000000",
  54972=>"000110111",
  54973=>"010000000",
  54974=>"111111110",
  54975=>"001011011",
  54976=>"000000000",
  54977=>"111111000",
  54978=>"011000011",
  54979=>"111111011",
  54980=>"111111111",
  54981=>"010100000",
  54982=>"011111110",
  54983=>"011111110",
  54984=>"010110111",
  54985=>"000000000",
  54986=>"110110000",
  54987=>"000111000",
  54988=>"101111101",
  54989=>"000000111",
  54990=>"000001110",
  54991=>"000100000",
  54992=>"101011111",
  54993=>"000110111",
  54994=>"000000111",
  54995=>"000100101",
  54996=>"000111111",
  54997=>"111111111",
  54998=>"000000111",
  54999=>"111011111",
  55000=>"111111000",
  55001=>"001000011",
  55002=>"000000100",
  55003=>"111001111",
  55004=>"111111100",
  55005=>"111111011",
  55006=>"111000111",
  55007=>"000000010",
  55008=>"000000000",
  55009=>"000110111",
  55010=>"111100100",
  55011=>"101000000",
  55012=>"000000000",
  55013=>"001001001",
  55014=>"111111111",
  55015=>"100110111",
  55016=>"111000000",
  55017=>"111111111",
  55018=>"111111010",
  55019=>"010111110",
  55020=>"000001001",
  55021=>"000100111",
  55022=>"000000011",
  55023=>"111000000",
  55024=>"000010000",
  55025=>"000000000",
  55026=>"111111111",
  55027=>"000010110",
  55028=>"001001001",
  55029=>"000110100",
  55030=>"010011010",
  55031=>"111100101",
  55032=>"111111111",
  55033=>"010111101",
  55034=>"111011000",
  55035=>"000111110",
  55036=>"000111111",
  55037=>"111110110",
  55038=>"111000000",
  55039=>"100111111",
  55040=>"111000010",
  55041=>"000111111",
  55042=>"111101110",
  55043=>"000111101",
  55044=>"101111000",
  55045=>"000000000",
  55046=>"111111111",
  55047=>"111000000",
  55048=>"000110110",
  55049=>"111111011",
  55050=>"001000101",
  55051=>"110100111",
  55052=>"011111000",
  55053=>"001000110",
  55054=>"000000001",
  55055=>"000001001",
  55056=>"000000111",
  55057=>"000000011",
  55058=>"111010111",
  55059=>"000000011",
  55060=>"000000111",
  55061=>"111111100",
  55062=>"100111111",
  55063=>"000000101",
  55064=>"111111010",
  55065=>"111001001",
  55066=>"000110111",
  55067=>"111000000",
  55068=>"000111010",
  55069=>"000000001",
  55070=>"000000000",
  55071=>"111001000",
  55072=>"100010000",
  55073=>"000010111",
  55074=>"011000000",
  55075=>"000000000",
  55076=>"000111111",
  55077=>"100110100",
  55078=>"100000011",
  55079=>"101000010",
  55080=>"011100111",
  55081=>"000000010",
  55082=>"101000110",
  55083=>"100000001",
  55084=>"111000000",
  55085=>"001011011",
  55086=>"000100111",
  55087=>"000000000",
  55088=>"000110110",
  55089=>"111100000",
  55090=>"001100111",
  55091=>"000010100",
  55092=>"111000111",
  55093=>"000100000",
  55094=>"000111111",
  55095=>"011000111",
  55096=>"000001000",
  55097=>"111001001",
  55098=>"000000000",
  55099=>"111000111",
  55100=>"000011000",
  55101=>"000111001",
  55102=>"000100110",
  55103=>"100000000",
  55104=>"111000000",
  55105=>"111111110",
  55106=>"000000111",
  55107=>"001011000",
  55108=>"111111101",
  55109=>"100110000",
  55110=>"000000000",
  55111=>"001111111",
  55112=>"000000000",
  55113=>"000010111",
  55114=>"101100100",
  55115=>"000110000",
  55116=>"110110111",
  55117=>"111111101",
  55118=>"111100110",
  55119=>"000011000",
  55120=>"000011000",
  55121=>"111111000",
  55122=>"111110110",
  55123=>"000000000",
  55124=>"000000111",
  55125=>"001011011",
  55126=>"111111110",
  55127=>"101000011",
  55128=>"111111111",
  55129=>"010100000",
  55130=>"110100000",
  55131=>"001000000",
  55132=>"111111101",
  55133=>"011001111",
  55134=>"111001000",
  55135=>"101111001",
  55136=>"000000000",
  55137=>"001001111",
  55138=>"111001100",
  55139=>"111111111",
  55140=>"010111111",
  55141=>"000000000",
  55142=>"111111111",
  55143=>"111111111",
  55144=>"101111000",
  55145=>"101111001",
  55146=>"000000000",
  55147=>"011000100",
  55148=>"000011011",
  55149=>"001101001",
  55150=>"100111001",
  55151=>"001000001",
  55152=>"000010011",
  55153=>"010000110",
  55154=>"000000111",
  55155=>"001011001",
  55156=>"000000000",
  55157=>"011000000",
  55158=>"110111000",
  55159=>"100101001",
  55160=>"111111111",
  55161=>"111000111",
  55162=>"111111111",
  55163=>"000110000",
  55164=>"100000111",
  55165=>"101000101",
  55166=>"001000101",
  55167=>"000000011",
  55168=>"100110100",
  55169=>"101110110",
  55170=>"000000011",
  55171=>"001000000",
  55172=>"001111011",
  55173=>"000000000",
  55174=>"000000000",
  55175=>"000111111",
  55176=>"000000100",
  55177=>"000000000",
  55178=>"011011011",
  55179=>"000111111",
  55180=>"111101111",
  55181=>"100100100",
  55182=>"111100000",
  55183=>"001000000",
  55184=>"000000000",
  55185=>"111111111",
  55186=>"111110111",
  55187=>"000110111",
  55188=>"111111111",
  55189=>"000001000",
  55190=>"110100100",
  55191=>"000010010",
  55192=>"111000011",
  55193=>"000110000",
  55194=>"111111000",
  55195=>"011110000",
  55196=>"111111011",
  55197=>"000000011",
  55198=>"111000000",
  55199=>"000100111",
  55200=>"000000011",
  55201=>"010110001",
  55202=>"111111111",
  55203=>"111100000",
  55204=>"111111100",
  55205=>"111000000",
  55206=>"111000111",
  55207=>"011001011",
  55208=>"000001000",
  55209=>"100100111",
  55210=>"111111111",
  55211=>"001000000",
  55212=>"000000000",
  55213=>"000110111",
  55214=>"110110000",
  55215=>"000000000",
  55216=>"000000110",
  55217=>"000111110",
  55218=>"111110000",
  55219=>"111111110",
  55220=>"000111111",
  55221=>"111000111",
  55222=>"111110000",
  55223=>"000000000",
  55224=>"111110000",
  55225=>"000000000",
  55226=>"000001111",
  55227=>"000010111",
  55228=>"000000011",
  55229=>"111111101",
  55230=>"101001000",
  55231=>"100111000",
  55232=>"001101000",
  55233=>"000000000",
  55234=>"111011111",
  55235=>"000000000",
  55236=>"001000100",
  55237=>"111111000",
  55238=>"101000011",
  55239=>"111000000",
  55240=>"000100111",
  55241=>"111110000",
  55242=>"111001000",
  55243=>"000000100",
  55244=>"111111001",
  55245=>"111111000",
  55246=>"001111111",
  55247=>"101111111",
  55248=>"111101000",
  55249=>"011111000",
  55250=>"000011111",
  55251=>"111111111",
  55252=>"111001001",
  55253=>"000100101",
  55254=>"001000011",
  55255=>"000001010",
  55256=>"100100001",
  55257=>"111111000",
  55258=>"111000111",
  55259=>"111011001",
  55260=>"011011110",
  55261=>"001101110",
  55262=>"011000000",
  55263=>"111111000",
  55264=>"000100000",
  55265=>"111110111",
  55266=>"101000000",
  55267=>"000000000",
  55268=>"000111110",
  55269=>"000000111",
  55270=>"000100110",
  55271=>"111001111",
  55272=>"001001000",
  55273=>"111000111",
  55274=>"110110111",
  55275=>"011011011",
  55276=>"001000000",
  55277=>"000011000",
  55278=>"000110111",
  55279=>"011001111",
  55280=>"000000000",
  55281=>"000010000",
  55282=>"000111111",
  55283=>"001000000",
  55284=>"101000000",
  55285=>"000101111",
  55286=>"000000100",
  55287=>"000000000",
  55288=>"000111001",
  55289=>"000111111",
  55290=>"111100000",
  55291=>"001000000",
  55292=>"111100001",
  55293=>"110111111",
  55294=>"000000000",
  55295=>"000000111",
  55296=>"111100100",
  55297=>"000000000",
  55298=>"111111111",
  55299=>"000010111",
  55300=>"001100000",
  55301=>"111011111",
  55302=>"111111111",
  55303=>"111111111",
  55304=>"111111110",
  55305=>"111100000",
  55306=>"000000111",
  55307=>"000110111",
  55308=>"001001011",
  55309=>"000000000",
  55310=>"000100111",
  55311=>"111000000",
  55312=>"110111111",
  55313=>"000111111",
  55314=>"000010111",
  55315=>"110100000",
  55316=>"111111001",
  55317=>"110110000",
  55318=>"011111111",
  55319=>"111111111",
  55320=>"111111100",
  55321=>"011011010",
  55322=>"111011111",
  55323=>"000000101",
  55324=>"000100111",
  55325=>"001001101",
  55326=>"010110110",
  55327=>"000000000",
  55328=>"000000000",
  55329=>"000000000",
  55330=>"111111111",
  55331=>"010011111",
  55332=>"000000000",
  55333=>"111100000",
  55334=>"000000111",
  55335=>"010000000",
  55336=>"001000000",
  55337=>"010111111",
  55338=>"001000000",
  55339=>"001111111",
  55340=>"100011000",
  55341=>"010111111",
  55342=>"100000000",
  55343=>"111111111",
  55344=>"111000000",
  55345=>"100100111",
  55346=>"010111100",
  55347=>"010001111",
  55348=>"111111011",
  55349=>"000000000",
  55350=>"101000111",
  55351=>"110110011",
  55352=>"000111110",
  55353=>"100000000",
  55354=>"111111111",
  55355=>"111001001",
  55356=>"111111111",
  55357=>"000000000",
  55358=>"011000000",
  55359=>"111111100",
  55360=>"000000000",
  55361=>"011111111",
  55362=>"000000000",
  55363=>"111111111",
  55364=>"001001000",
  55365=>"111111111",
  55366=>"111111000",
  55367=>"110110000",
  55368=>"100110100",
  55369=>"000000111",
  55370=>"000001111",
  55371=>"111010110",
  55372=>"000100000",
  55373=>"110000000",
  55374=>"111100100",
  55375=>"111111111",
  55376=>"000000000",
  55377=>"000101111",
  55378=>"101000000",
  55379=>"001001111",
  55380=>"000000000",
  55381=>"111111111",
  55382=>"000000111",
  55383=>"111111000",
  55384=>"000000110",
  55385=>"000000100",
  55386=>"001001000",
  55387=>"001001001",
  55388=>"010110000",
  55389=>"111111110",
  55390=>"111111111",
  55391=>"000000000",
  55392=>"000010000",
  55393=>"001001111",
  55394=>"111111111",
  55395=>"000111111",
  55396=>"001001001",
  55397=>"111100100",
  55398=>"000000001",
  55399=>"000101000",
  55400=>"111110101",
  55401=>"000000000",
  55402=>"010010000",
  55403=>"111111111",
  55404=>"111000100",
  55405=>"111101000",
  55406=>"111111111",
  55407=>"111110010",
  55408=>"110111111",
  55409=>"011111111",
  55410=>"110110111",
  55411=>"000000000",
  55412=>"000000111",
  55413=>"111111100",
  55414=>"111111000",
  55415=>"110110111",
  55416=>"111001000",
  55417=>"111111111",
  55418=>"000000011",
  55419=>"000000000",
  55420=>"100110110",
  55421=>"111111000",
  55422=>"000000000",
  55423=>"110111110",
  55424=>"000000000",
  55425=>"001000100",
  55426=>"111100011",
  55427=>"010000010",
  55428=>"110111011",
  55429=>"111100000",
  55430=>"001001111",
  55431=>"000000000",
  55432=>"000011111",
  55433=>"100110111",
  55434=>"000111111",
  55435=>"111111110",
  55436=>"111111010",
  55437=>"010111011",
  55438=>"001000111",
  55439=>"111111111",
  55440=>"100100111",
  55441=>"000000000",
  55442=>"111000111",
  55443=>"001000000",
  55444=>"111111000",
  55445=>"001001000",
  55446=>"111101111",
  55447=>"000000111",
  55448=>"111111111",
  55449=>"111010110",
  55450=>"010011010",
  55451=>"101100110",
  55452=>"000000111",
  55453=>"111000000",
  55454=>"111111111",
  55455=>"110111010",
  55456=>"111111010",
  55457=>"000000000",
  55458=>"000000000",
  55459=>"000111111",
  55460=>"000000000",
  55461=>"000000000",
  55462=>"000111111",
  55463=>"001011000",
  55464=>"000100100",
  55465=>"000000001",
  55466=>"001011000",
  55467=>"000000001",
  55468=>"111101011",
  55469=>"000110100",
  55470=>"111111000",
  55471=>"000000100",
  55472=>"111111111",
  55473=>"001000000",
  55474=>"110111111",
  55475=>"011111110",
  55476=>"101000000",
  55477=>"110101000",
  55478=>"000000000",
  55479=>"111111001",
  55480=>"101101001",
  55481=>"001000000",
  55482=>"100000111",
  55483=>"000000000",
  55484=>"111011000",
  55485=>"111111100",
  55486=>"011001111",
  55487=>"111000000",
  55488=>"001000000",
  55489=>"001001111",
  55490=>"110111100",
  55491=>"010111110",
  55492=>"000000000",
  55493=>"111111111",
  55494=>"000000000",
  55495=>"000010000",
  55496=>"000000000",
  55497=>"000000001",
  55498=>"111111111",
  55499=>"000000010",
  55500=>"001000111",
  55501=>"100000000",
  55502=>"111011000",
  55503=>"110110110",
  55504=>"000000011",
  55505=>"000010111",
  55506=>"000010011",
  55507=>"000000000",
  55508=>"111111000",
  55509=>"111111110",
  55510=>"111111111",
  55511=>"111111111",
  55512=>"111111000",
  55513=>"111111111",
  55514=>"000000000",
  55515=>"111111111",
  55516=>"111111000",
  55517=>"101001000",
  55518=>"111111111",
  55519=>"111111111",
  55520=>"000000000",
  55521=>"011111111",
  55522=>"111010011",
  55523=>"000111111",
  55524=>"111111111",
  55525=>"100000100",
  55526=>"010000000",
  55527=>"000000100",
  55528=>"000000100",
  55529=>"010000110",
  55530=>"000111111",
  55531=>"111011111",
  55532=>"001000111",
  55533=>"111111111",
  55534=>"100001111",
  55535=>"111011111",
  55536=>"000000000",
  55537=>"111111111",
  55538=>"111000000",
  55539=>"000000001",
  55540=>"111110000",
  55541=>"000000000",
  55542=>"111111110",
  55543=>"000111000",
  55544=>"000000000",
  55545=>"000000011",
  55546=>"000000000",
  55547=>"000000000",
  55548=>"000000011",
  55549=>"000000001",
  55550=>"000000000",
  55551=>"111111010",
  55552=>"111111111",
  55553=>"000111111",
  55554=>"011111101",
  55555=>"000000101",
  55556=>"001000000",
  55557=>"111000000",
  55558=>"110111111",
  55559=>"000110111",
  55560=>"000101100",
  55561=>"111001001",
  55562=>"101100101",
  55563=>"000100110",
  55564=>"001011111",
  55565=>"000011101",
  55566=>"110000000",
  55567=>"110111111",
  55568=>"001000000",
  55569=>"100111000",
  55570=>"111000000",
  55571=>"000000010",
  55572=>"000111111",
  55573=>"000000001",
  55574=>"001110110",
  55575=>"000000111",
  55576=>"100000000",
  55577=>"111111111",
  55578=>"110110010",
  55579=>"111000000",
  55580=>"111111111",
  55581=>"011111111",
  55582=>"000010000",
  55583=>"011111111",
  55584=>"000101001",
  55585=>"101101000",
  55586=>"000100111",
  55587=>"000001111",
  55588=>"111111111",
  55589=>"111001000",
  55590=>"000111111",
  55591=>"000000000",
  55592=>"101011000",
  55593=>"000000000",
  55594=>"000000000",
  55595=>"000101111",
  55596=>"101000111",
  55597=>"111111011",
  55598=>"111101000",
  55599=>"000000000",
  55600=>"011110110",
  55601=>"000000000",
  55602=>"111111111",
  55603=>"010000000",
  55604=>"111000000",
  55605=>"111000000",
  55606=>"000011111",
  55607=>"100001111",
  55608=>"000000000",
  55609=>"000001000",
  55610=>"001001101",
  55611=>"000000000",
  55612=>"111111100",
  55613=>"001000000",
  55614=>"001000111",
  55615=>"111000000",
  55616=>"111000000",
  55617=>"111000000",
  55618=>"100010010",
  55619=>"001000101",
  55620=>"100110111",
  55621=>"111110111",
  55622=>"111111111",
  55623=>"111101000",
  55624=>"110111110",
  55625=>"010000000",
  55626=>"011000000",
  55627=>"001101111",
  55628=>"100111000",
  55629=>"000000000",
  55630=>"111011111",
  55631=>"101111111",
  55632=>"111111100",
  55633=>"111111100",
  55634=>"000000011",
  55635=>"000000101",
  55636=>"000011111",
  55637=>"011011011",
  55638=>"111111000",
  55639=>"100000000",
  55640=>"111111111",
  55641=>"111111111",
  55642=>"001000000",
  55643=>"000000000",
  55644=>"010010000",
  55645=>"001000000",
  55646=>"110000000",
  55647=>"111111111",
  55648=>"110110100",
  55649=>"000000000",
  55650=>"111111111",
  55651=>"111111111",
  55652=>"000000110",
  55653=>"000000000",
  55654=>"111111111",
  55655=>"111111110",
  55656=>"110111111",
  55657=>"101110111",
  55658=>"000000111",
  55659=>"100000000",
  55660=>"110111111",
  55661=>"111111111",
  55662=>"000000000",
  55663=>"000000101",
  55664=>"110111110",
  55665=>"000000000",
  55666=>"000010000",
  55667=>"011010000",
  55668=>"001000000",
  55669=>"000000000",
  55670=>"111100000",
  55671=>"000000111",
  55672=>"111000000",
  55673=>"000000011",
  55674=>"011011001",
  55675=>"111111000",
  55676=>"000100111",
  55677=>"000011000",
  55678=>"011011111",
  55679=>"000000101",
  55680=>"111100100",
  55681=>"001001100",
  55682=>"111111011",
  55683=>"000000000",
  55684=>"011000101",
  55685=>"000000000",
  55686=>"000000000",
  55687=>"110000101",
  55688=>"000000000",
  55689=>"111111111",
  55690=>"111111111",
  55691=>"100100100",
  55692=>"111111111",
  55693=>"011111111",
  55694=>"111111110",
  55695=>"111111111",
  55696=>"111100000",
  55697=>"000000000",
  55698=>"000000000",
  55699=>"111111001",
  55700=>"000110111",
  55701=>"000000000",
  55702=>"000000000",
  55703=>"001001111",
  55704=>"000000000",
  55705=>"111101111",
  55706=>"111111010",
  55707=>"000100111",
  55708=>"011111111",
  55709=>"110110000",
  55710=>"101101101",
  55711=>"001101111",
  55712=>"011011000",
  55713=>"111111111",
  55714=>"000000000",
  55715=>"001000000",
  55716=>"100111100",
  55717=>"001011000",
  55718=>"110101111",
  55719=>"111011111",
  55720=>"100000011",
  55721=>"010011111",
  55722=>"111111000",
  55723=>"111111111",
  55724=>"000000000",
  55725=>"011111100",
  55726=>"111111111",
  55727=>"000000100",
  55728=>"011000000",
  55729=>"000110000",
  55730=>"111101101",
  55731=>"111111111",
  55732=>"101001001",
  55733=>"111111111",
  55734=>"110000000",
  55735=>"000000001",
  55736=>"000000000",
  55737=>"111111111",
  55738=>"000000111",
  55739=>"111000000",
  55740=>"101011000",
  55741=>"111001000",
  55742=>"111111111",
  55743=>"111101001",
  55744=>"111111111",
  55745=>"111000000",
  55746=>"000000000",
  55747=>"111100000",
  55748=>"110100101",
  55749=>"111111111",
  55750=>"111111010",
  55751=>"000101100",
  55752=>"111111101",
  55753=>"111110000",
  55754=>"000000100",
  55755=>"010110111",
  55756=>"111000001",
  55757=>"111111110",
  55758=>"111111111",
  55759=>"000000000",
  55760=>"111111111",
  55761=>"100100100",
  55762=>"111111010",
  55763=>"100111111",
  55764=>"011111011",
  55765=>"111111000",
  55766=>"000000110",
  55767=>"000000010",
  55768=>"111110011",
  55769=>"000000000",
  55770=>"011011011",
  55771=>"111111111",
  55772=>"110110111",
  55773=>"001000000",
  55774=>"111100000",
  55775=>"111001001",
  55776=>"011000000",
  55777=>"111101111",
  55778=>"001000000",
  55779=>"010110000",
  55780=>"000000001",
  55781=>"010010010",
  55782=>"101000101",
  55783=>"111111111",
  55784=>"101111111",
  55785=>"111000111",
  55786=>"000001111",
  55787=>"000000000",
  55788=>"111101001",
  55789=>"100000000",
  55790=>"000000000",
  55791=>"111111011",
  55792=>"100100111",
  55793=>"100111111",
  55794=>"000000000",
  55795=>"000000000",
  55796=>"001000000",
  55797=>"000000000",
  55798=>"001000000",
  55799=>"111111111",
  55800=>"000111111",
  55801=>"111111111",
  55802=>"111111000",
  55803=>"111010000",
  55804=>"000000000",
  55805=>"001111100",
  55806=>"111010000",
  55807=>"111111111",
  55808=>"110110000",
  55809=>"001001001",
  55810=>"001000000",
  55811=>"000000000",
  55812=>"010000010",
  55813=>"111000001",
  55814=>"111011111",
  55815=>"100111100",
  55816=>"000000000",
  55817=>"011000111",
  55818=>"000001001",
  55819=>"000000000",
  55820=>"001110100",
  55821=>"001000001",
  55822=>"100000000",
  55823=>"101100100",
  55824=>"000100000",
  55825=>"010110111",
  55826=>"111100101",
  55827=>"111111010",
  55828=>"000000000",
  55829=>"111001000",
  55830=>"000011010",
  55831=>"011011000",
  55832=>"110110000",
  55833=>"111111100",
  55834=>"101000011",
  55835=>"000101101",
  55836=>"111100101",
  55837=>"110000000",
  55838=>"011001001",
  55839=>"001000110",
  55840=>"000000011",
  55841=>"111111111",
  55842=>"011011001",
  55843=>"111111111",
  55844=>"110110011",
  55845=>"000000000",
  55846=>"100111111",
  55847=>"100000101",
  55848=>"110111111",
  55849=>"000000000",
  55850=>"000000111",
  55851=>"010110000",
  55852=>"000010000",
  55853=>"010010010",
  55854=>"101101101",
  55855=>"001100101",
  55856=>"010110000",
  55857=>"111000001",
  55858=>"000000000",
  55859=>"000000000",
  55860=>"000010110",
  55861=>"001001001",
  55862=>"000100111",
  55863=>"000000000",
  55864=>"110111111",
  55865=>"000110000",
  55866=>"101001011",
  55867=>"101101000",
  55868=>"111100000",
  55869=>"000001011",
  55870=>"111101011",
  55871=>"111000001",
  55872=>"000000000",
  55873=>"001001000",
  55874=>"000000001",
  55875=>"010101111",
  55876=>"001000100",
  55877=>"110100111",
  55878=>"001011011",
  55879=>"000110111",
  55880=>"011011011",
  55881=>"001100111",
  55882=>"111001101",
  55883=>"110110100",
  55884=>"000000000",
  55885=>"001001000",
  55886=>"000010111",
  55887=>"000000111",
  55888=>"101111111",
  55889=>"010010000",
  55890=>"111001001",
  55891=>"100100100",
  55892=>"010011000",
  55893=>"110111110",
  55894=>"101111111",
  55895=>"000111111",
  55896=>"111000000",
  55897=>"100000111",
  55898=>"000010000",
  55899=>"000100101",
  55900=>"000000111",
  55901=>"000001011",
  55902=>"001001111",
  55903=>"000001001",
  55904=>"000101111",
  55905=>"110110010",
  55906=>"111111011",
  55907=>"000101111",
  55908=>"110110100",
  55909=>"111111110",
  55910=>"010000010",
  55911=>"111001000",
  55912=>"000000111",
  55913=>"111111001",
  55914=>"000001111",
  55915=>"000000010",
  55916=>"111110110",
  55917=>"111110000",
  55918=>"111111111",
  55919=>"000000000",
  55920=>"111000000",
  55921=>"000000001",
  55922=>"100000100",
  55923=>"110111111",
  55924=>"010010010",
  55925=>"001001111",
  55926=>"010000001",
  55927=>"101101111",
  55928=>"110001111",
  55929=>"001000011",
  55930=>"111000000",
  55931=>"010000000",
  55932=>"100100100",
  55933=>"000101001",
  55934=>"000000000",
  55935=>"000000001",
  55936=>"101101101",
  55937=>"100101000",
  55938=>"000000100",
  55939=>"011011000",
  55940=>"111111111",
  55941=>"111000000",
  55942=>"001000011",
  55943=>"000000000",
  55944=>"000000000",
  55945=>"100111111",
  55946=>"000000000",
  55947=>"011010011",
  55948=>"111110000",
  55949=>"100101100",
  55950=>"011000000",
  55951=>"111111111",
  55952=>"000000000",
  55953=>"110111010",
  55954=>"010110110",
  55955=>"001000101",
  55956=>"111111010",
  55957=>"111000000",
  55958=>"000001001",
  55959=>"111111000",
  55960=>"001001001",
  55961=>"111110001",
  55962=>"111011111",
  55963=>"000000000",
  55964=>"011001000",
  55965=>"111110000",
  55966=>"110000000",
  55967=>"000101101",
  55968=>"111111001",
  55969=>"000100101",
  55970=>"110010000",
  55971=>"001111111",
  55972=>"000000000",
  55973=>"111111111",
  55974=>"000000000",
  55975=>"011100111",
  55976=>"000000111",
  55977=>"000000000",
  55978=>"000000100",
  55979=>"110110010",
  55980=>"001101000",
  55981=>"110110000",
  55982=>"000001111",
  55983=>"111111000",
  55984=>"010010000",
  55985=>"111111011",
  55986=>"111111111",
  55987=>"010111110",
  55988=>"100000001",
  55989=>"000100111",
  55990=>"111101001",
  55991=>"000000011",
  55992=>"000001111",
  55993=>"101001111",
  55994=>"101001001",
  55995=>"011111111",
  55996=>"000000000",
  55997=>"111111111",
  55998=>"000000001",
  55999=>"111111000",
  56000=>"100110111",
  56001=>"000000000",
  56002=>"000010110",
  56003=>"110111110",
  56004=>"001001111",
  56005=>"101101001",
  56006=>"001000110",
  56007=>"110110101",
  56008=>"111111010",
  56009=>"010100000",
  56010=>"001000101",
  56011=>"101001101",
  56012=>"111111101",
  56013=>"001011111",
  56014=>"000010110",
  56015=>"010010011",
  56016=>"000000111",
  56017=>"000000001",
  56018=>"111111111",
  56019=>"101000001",
  56020=>"111100101",
  56021=>"000000000",
  56022=>"100000000",
  56023=>"110110111",
  56024=>"110110011",
  56025=>"000000000",
  56026=>"000000111",
  56027=>"101101000",
  56028=>"111001001",
  56029=>"000000000",
  56030=>"010110010",
  56031=>"001101111",
  56032=>"000000000",
  56033=>"000000000",
  56034=>"111111000",
  56035=>"001000000",
  56036=>"010100111",
  56037=>"111111111",
  56038=>"000010000",
  56039=>"001001111",
  56040=>"111111011",
  56041=>"111111110",
  56042=>"111111110",
  56043=>"111110100",
  56044=>"111111111",
  56045=>"000000000",
  56046=>"011011101",
  56047=>"111101101",
  56048=>"000011111",
  56049=>"111111010",
  56050=>"110010000",
  56051=>"000000000",
  56052=>"100111111",
  56053=>"110000000",
  56054=>"001001001",
  56055=>"010110010",
  56056=>"101000001",
  56057=>"011110000",
  56058=>"000001001",
  56059=>"000000111",
  56060=>"001001000",
  56061=>"110110110",
  56062=>"001000000",
  56063=>"000000100",
  56064=>"000000000",
  56065=>"000000101",
  56066=>"111111111",
  56067=>"111111000",
  56068=>"000000000",
  56069=>"110110111",
  56070=>"111111111",
  56071=>"111000101",
  56072=>"111111010",
  56073=>"111100000",
  56074=>"000001101",
  56075=>"111111010",
  56076=>"001000100",
  56077=>"010010010",
  56078=>"011001101",
  56079=>"111101100",
  56080=>"000011000",
  56081=>"000000000",
  56082=>"000000011",
  56083=>"010110110",
  56084=>"111011111",
  56085=>"101000111",
  56086=>"000100111",
  56087=>"010110010",
  56088=>"110110110",
  56089=>"111111111",
  56090=>"000111111",
  56091=>"101101111",
  56092=>"101101101",
  56093=>"111111111",
  56094=>"000000010",
  56095=>"111110100",
  56096=>"011011010",
  56097=>"000110110",
  56098=>"111111011",
  56099=>"001000001",
  56100=>"001001000",
  56101=>"111111010",
  56102=>"000000000",
  56103=>"010011111",
  56104=>"101100111",
  56105=>"000000111",
  56106=>"010010000",
  56107=>"000000000",
  56108=>"111111110",
  56109=>"110110110",
  56110=>"000000111",
  56111=>"100000100",
  56112=>"110110110",
  56113=>"010011010",
  56114=>"111111111",
  56115=>"000010011",
  56116=>"010010000",
  56117=>"101111111",
  56118=>"100000001",
  56119=>"111101101",
  56120=>"000000000",
  56121=>"000000101",
  56122=>"001001000",
  56123=>"000000000",
  56124=>"010010011",
  56125=>"010000000",
  56126=>"000111111",
  56127=>"001101101",
  56128=>"000000110",
  56129=>"100111110",
  56130=>"000000000",
  56131=>"001000000",
  56132=>"111100000",
  56133=>"111100000",
  56134=>"111000111",
  56135=>"111111111",
  56136=>"001100110",
  56137=>"000000001",
  56138=>"111100000",
  56139=>"000000000",
  56140=>"000110111",
  56141=>"100000000",
  56142=>"010001101",
  56143=>"100111001",
  56144=>"000000000",
  56145=>"001000000",
  56146=>"010000000",
  56147=>"000000001",
  56148=>"011011001",
  56149=>"001001001",
  56150=>"111011011",
  56151=>"001001111",
  56152=>"111001001",
  56153=>"000000001",
  56154=>"111000000",
  56155=>"101000001",
  56156=>"010010000",
  56157=>"000001111",
  56158=>"111000111",
  56159=>"000000000",
  56160=>"101000001",
  56161=>"010010111",
  56162=>"101111011",
  56163=>"101000000",
  56164=>"001001001",
  56165=>"000000000",
  56166=>"111110110",
  56167=>"110111010",
  56168=>"010000100",
  56169=>"001000100",
  56170=>"000000000",
  56171=>"011010110",
  56172=>"110110100",
  56173=>"000001101",
  56174=>"001000001",
  56175=>"000000111",
  56176=>"000100111",
  56177=>"000000000",
  56178=>"101100111",
  56179=>"111111110",
  56180=>"110111000",
  56181=>"000101111",
  56182=>"000000000",
  56183=>"000000000",
  56184=>"101001000",
  56185=>"000000000",
  56186=>"000101111",
  56187=>"000000000",
  56188=>"100000000",
  56189=>"111110111",
  56190=>"001111110",
  56191=>"000101111",
  56192=>"101101000",
  56193=>"111111101",
  56194=>"001001111",
  56195=>"000010000",
  56196=>"001101101",
  56197=>"010011110",
  56198=>"000000111",
  56199=>"101001001",
  56200=>"001000100",
  56201=>"000111101",
  56202=>"111111001",
  56203=>"000001000",
  56204=>"011010111",
  56205=>"001001000",
  56206=>"100010011",
  56207=>"000000000",
  56208=>"010000000",
  56209=>"111111001",
  56210=>"111110111",
  56211=>"010100110",
  56212=>"110111111",
  56213=>"010010000",
  56214=>"001000000",
  56215=>"000010001",
  56216=>"111000010",
  56217=>"000001000",
  56218=>"111111111",
  56219=>"000000000",
  56220=>"000101100",
  56221=>"010111111",
  56222=>"101001101",
  56223=>"000000111",
  56224=>"111111111",
  56225=>"001111111",
  56226=>"000110110",
  56227=>"111001000",
  56228=>"000000011",
  56229=>"010010010",
  56230=>"111010111",
  56231=>"011110111",
  56232=>"000000000",
  56233=>"011011110",
  56234=>"001011100",
  56235=>"000000000",
  56236=>"000000001",
  56237=>"000000000",
  56238=>"000010000",
  56239=>"010010000",
  56240=>"000000000",
  56241=>"000000101",
  56242=>"000000100",
  56243=>"000001000",
  56244=>"010110111",
  56245=>"001000101",
  56246=>"110111111",
  56247=>"010010010",
  56248=>"110110111",
  56249=>"010010010",
  56250=>"110000000",
  56251=>"101111111",
  56252=>"000000000",
  56253=>"001001000",
  56254=>"000000000",
  56255=>"000100110",
  56256=>"001001000",
  56257=>"100100111",
  56258=>"001111001",
  56259=>"111111111",
  56260=>"111110010",
  56261=>"111111011",
  56262=>"011010000",
  56263=>"111101100",
  56264=>"000000100",
  56265=>"000000001",
  56266=>"000000001",
  56267=>"100110110",
  56268=>"111110010",
  56269=>"000000001",
  56270=>"101000000",
  56271=>"111000101",
  56272=>"000000111",
  56273=>"000000100",
  56274=>"110111101",
  56275=>"001111111",
  56276=>"101111111",
  56277=>"110000000",
  56278=>"101001000",
  56279=>"100010011",
  56280=>"000000000",
  56281=>"110111110",
  56282=>"000000011",
  56283=>"110111011",
  56284=>"000000000",
  56285=>"011000101",
  56286=>"101111011",
  56287=>"000100110",
  56288=>"000000000",
  56289=>"100000001",
  56290=>"111111100",
  56291=>"000100101",
  56292=>"111111111",
  56293=>"001000000",
  56294=>"111010000",
  56295=>"000000000",
  56296=>"110110010",
  56297=>"010100000",
  56298=>"110110010",
  56299=>"000000000",
  56300=>"100111111",
  56301=>"011111000",
  56302=>"000001111",
  56303=>"000010111",
  56304=>"100000111",
  56305=>"001000000",
  56306=>"011111010",
  56307=>"000000100",
  56308=>"000000100",
  56309=>"010000000",
  56310=>"101111111",
  56311=>"001011111",
  56312=>"111111000",
  56313=>"000001000",
  56314=>"010110010",
  56315=>"000000100",
  56316=>"110110100",
  56317=>"000000000",
  56318=>"000111111",
  56319=>"000111111",
  56320=>"000000000",
  56321=>"001011100",
  56322=>"000100111",
  56323=>"111111111",
  56324=>"110111110",
  56325=>"100000111",
  56326=>"101111111",
  56327=>"100000000",
  56328=>"111111111",
  56329=>"111111011",
  56330=>"010000000",
  56331=>"000100100",
  56332=>"111111001",
  56333=>"000000101",
  56334=>"111111001",
  56335=>"111111000",
  56336=>"011111111",
  56337=>"011111011",
  56338=>"000100100",
  56339=>"000000111",
  56340=>"000000100",
  56341=>"111111110",
  56342=>"000000000",
  56343=>"110100100",
  56344=>"011011010",
  56345=>"000000000",
  56346=>"111001000",
  56347=>"011011011",
  56348=>"000000000",
  56349=>"000011111",
  56350=>"000100011",
  56351=>"000110110",
  56352=>"001011111",
  56353=>"110110110",
  56354=>"000000000",
  56355=>"110111000",
  56356=>"111111001",
  56357=>"110100100",
  56358=>"110100000",
  56359=>"000000111",
  56360=>"111111100",
  56361=>"011111111",
  56362=>"001000000",
  56363=>"000110110",
  56364=>"000000000",
  56365=>"000000000",
  56366=>"000000011",
  56367=>"111111111",
  56368=>"111111100",
  56369=>"110111001",
  56370=>"000000000",
  56371=>"000000001",
  56372=>"000010000",
  56373=>"100000000",
  56374=>"001000000",
  56375=>"000000000",
  56376=>"000011010",
  56377=>"000101110",
  56378=>"001101111",
  56379=>"111010111",
  56380=>"000100100",
  56381=>"000000000",
  56382=>"111011011",
  56383=>"000000000",
  56384=>"010011011",
  56385=>"010000000",
  56386=>"111100000",
  56387=>"110110000",
  56388=>"000000011",
  56389=>"000000110",
  56390=>"000001000",
  56391=>"100000000",
  56392=>"011011011",
  56393=>"111001001",
  56394=>"100111111",
  56395=>"000000000",
  56396=>"111111111",
  56397=>"000000000",
  56398=>"111111101",
  56399=>"111000000",
  56400=>"000000000",
  56401=>"010110001",
  56402=>"000000000",
  56403=>"111111000",
  56404=>"000010111",
  56405=>"000000001",
  56406=>"111100100",
  56407=>"000000101",
  56408=>"000000111",
  56409=>"111101001",
  56410=>"111111011",
  56411=>"000001010",
  56412=>"000000110",
  56413=>"001101011",
  56414=>"011001001",
  56415=>"001111110",
  56416=>"111111111",
  56417=>"111101001",
  56418=>"111111101",
  56419=>"111111111",
  56420=>"000000000",
  56421=>"010000000",
  56422=>"110000000",
  56423=>"011111101",
  56424=>"111111000",
  56425=>"000000000",
  56426=>"000101111",
  56427=>"101100100",
  56428=>"000100111",
  56429=>"000000111",
  56430=>"111000000",
  56431=>"111101000",
  56432=>"111111000",
  56433=>"110010000",
  56434=>"011111111",
  56435=>"000000000",
  56436=>"000001101",
  56437=>"100111111",
  56438=>"011001001",
  56439=>"000010111",
  56440=>"011001000",
  56441=>"000000000",
  56442=>"000111101",
  56443=>"111111101",
  56444=>"111010111",
  56445=>"111111000",
  56446=>"010111111",
  56447=>"000000000",
  56448=>"000100111",
  56449=>"100100000",
  56450=>"100111100",
  56451=>"111111000",
  56452=>"111111101",
  56453=>"000000000",
  56454=>"001000011",
  56455=>"111110000",
  56456=>"000000100",
  56457=>"000000001",
  56458=>"111110000",
  56459=>"000000111",
  56460=>"011001001",
  56461=>"000000110",
  56462=>"000000100",
  56463=>"000000111",
  56464=>"100111111",
  56465=>"000000000",
  56466=>"111111001",
  56467=>"001001101",
  56468=>"100111111",
  56469=>"000100110",
  56470=>"111101000",
  56471=>"000000000",
  56472=>"111001000",
  56473=>"000000000",
  56474=>"000010110",
  56475=>"011010111",
  56476=>"110100000",
  56477=>"111000000",
  56478=>"000000000",
  56479=>"000111001",
  56480=>"100100111",
  56481=>"000011111",
  56482=>"000111111",
  56483=>"000001111",
  56484=>"110111111",
  56485=>"000000001",
  56486=>"000111111",
  56487=>"000011011",
  56488=>"110111111",
  56489=>"000000000",
  56490=>"000000001",
  56491=>"000000000",
  56492=>"110110011",
  56493=>"100001011",
  56494=>"110111011",
  56495=>"110010000",
  56496=>"111111111",
  56497=>"000000000",
  56498=>"010110011",
  56499=>"111111010",
  56500=>"011000001",
  56501=>"100110110",
  56502=>"000100111",
  56503=>"111000000",
  56504=>"100000000",
  56505=>"000001011",
  56506=>"011110000",
  56507=>"111111111",
  56508=>"000000100",
  56509=>"111111000",
  56510=>"100111111",
  56511=>"111111001",
  56512=>"000001001",
  56513=>"111111111",
  56514=>"111001011",
  56515=>"000111001",
  56516=>"111011111",
  56517=>"000000000",
  56518=>"111111010",
  56519=>"111011011",
  56520=>"000000000",
  56521=>"101000111",
  56522=>"011111101",
  56523=>"000011111",
  56524=>"000000111",
  56525=>"111111110",
  56526=>"101111001",
  56527=>"111100000",
  56528=>"000000100",
  56529=>"001000000",
  56530=>"001000110",
  56531=>"000001111",
  56532=>"111111101",
  56533=>"111110000",
  56534=>"111101000",
  56535=>"011111100",
  56536=>"111111111",
  56537=>"000000000",
  56538=>"111111111",
  56539=>"000000000",
  56540=>"000100111",
  56541=>"000000000",
  56542=>"011110000",
  56543=>"000000111",
  56544=>"111011000",
  56545=>"111111000",
  56546=>"000111110",
  56547=>"111111111",
  56548=>"000000000",
  56549=>"000110100",
  56550=>"000111000",
  56551=>"000000000",
  56552=>"101000011",
  56553=>"000011000",
  56554=>"111111101",
  56555=>"000000000",
  56556=>"000000111",
  56557=>"111111111",
  56558=>"000000000",
  56559=>"011001111",
  56560=>"011000000",
  56561=>"000000000",
  56562=>"111100100",
  56563=>"110110010",
  56564=>"111111111",
  56565=>"000001001",
  56566=>"010001001",
  56567=>"000000000",
  56568=>"111111111",
  56569=>"001111101",
  56570=>"000000000",
  56571=>"000000000",
  56572=>"000000000",
  56573=>"001111111",
  56574=>"100110111",
  56575=>"001000000",
  56576=>"111111000",
  56577=>"001001011",
  56578=>"000000000",
  56579=>"010100111",
  56580=>"000000111",
  56581=>"111111111",
  56582=>"111111111",
  56583=>"000000000",
  56584=>"110010011",
  56585=>"000000000",
  56586=>"111111111",
  56587=>"111111000",
  56588=>"001000000",
  56589=>"000000101",
  56590=>"000000000",
  56591=>"000000011",
  56592=>"001111111",
  56593=>"000110111",
  56594=>"111111111",
  56595=>"000001000",
  56596=>"111111111",
  56597=>"111111111",
  56598=>"000000000",
  56599=>"100000000",
  56600=>"011010110",
  56601=>"000000000",
  56602=>"111111111",
  56603=>"000011010",
  56604=>"100000110",
  56605=>"111111011",
  56606=>"011000000",
  56607=>"111111111",
  56608=>"000100001",
  56609=>"110111010",
  56610=>"000100111",
  56611=>"111111100",
  56612=>"111111111",
  56613=>"110111111",
  56614=>"011111111",
  56615=>"000000011",
  56616=>"111100101",
  56617=>"000000111",
  56618=>"111111000",
  56619=>"111111001",
  56620=>"000100100",
  56621=>"001011111",
  56622=>"111110100",
  56623=>"101111111",
  56624=>"000000100",
  56625=>"111111111",
  56626=>"111111100",
  56627=>"000000100",
  56628=>"111110000",
  56629=>"100000000",
  56630=>"111101111",
  56631=>"011001001",
  56632=>"000001000",
  56633=>"111000000",
  56634=>"111111111",
  56635=>"110110111",
  56636=>"000100100",
  56637=>"100110111",
  56638=>"000000000",
  56639=>"100000100",
  56640=>"100111111",
  56641=>"000000111",
  56642=>"111000000",
  56643=>"001000000",
  56644=>"011011000",
  56645=>"111000000",
  56646=>"111111100",
  56647=>"000000001",
  56648=>"000000000",
  56649=>"111111111",
  56650=>"011000000",
  56651=>"011000000",
  56652=>"001101100",
  56653=>"100111111",
  56654=>"100000000",
  56655=>"111011111",
  56656=>"000000100",
  56657=>"010010110",
  56658=>"000100100",
  56659=>"111011111",
  56660=>"000011000",
  56661=>"001111100",
  56662=>"111100000",
  56663=>"100100110",
  56664=>"000001111",
  56665=>"111111101",
  56666=>"110110100",
  56667=>"000000001",
  56668=>"110111111",
  56669=>"000110111",
  56670=>"000000000",
  56671=>"000000000",
  56672=>"111111001",
  56673=>"001111111",
  56674=>"000000110",
  56675=>"000000000",
  56676=>"000001111",
  56677=>"000000111",
  56678=>"000000001",
  56679=>"001001111",
  56680=>"011001001",
  56681=>"011111111",
  56682=>"000001000",
  56683=>"011001001",
  56684=>"111111111",
  56685=>"111110100",
  56686=>"001111111",
  56687=>"100000000",
  56688=>"010000000",
  56689=>"000000000",
  56690=>"111111111",
  56691=>"000110000",
  56692=>"001101111",
  56693=>"000000000",
  56694=>"110000000",
  56695=>"111111111",
  56696=>"000000001",
  56697=>"001011111",
  56698=>"000111111",
  56699=>"001001111",
  56700=>"111111111",
  56701=>"110110010",
  56702=>"111000101",
  56703=>"000000000",
  56704=>"001001001",
  56705=>"000000000",
  56706=>"111000100",
  56707=>"000011111",
  56708=>"000000111",
  56709=>"110111100",
  56710=>"001011111",
  56711=>"111000000",
  56712=>"111101101",
  56713=>"101111111",
  56714=>"000000000",
  56715=>"001001101",
  56716=>"111101000",
  56717=>"110111111",
  56718=>"000000000",
  56719=>"100110111",
  56720=>"000010000",
  56721=>"000000100",
  56722=>"111110100",
  56723=>"100000000",
  56724=>"111001000",
  56725=>"001011111",
  56726=>"001001001",
  56727=>"000000110",
  56728=>"000000111",
  56729=>"000011001",
  56730=>"000000000",
  56731=>"000000000",
  56732=>"111100100",
  56733=>"111111110",
  56734=>"001110100",
  56735=>"010100000",
  56736=>"000000001",
  56737=>"110110100",
  56738=>"110100000",
  56739=>"000001101",
  56740=>"110110100",
  56741=>"000000010",
  56742=>"111001010",
  56743=>"111000111",
  56744=>"100000010",
  56745=>"111111001",
  56746=>"111111111",
  56747=>"000000100",
  56748=>"101100111",
  56749=>"001001111",
  56750=>"111000001",
  56751=>"001110111",
  56752=>"101111111",
  56753=>"111011000",
  56754=>"000000000",
  56755=>"111111000",
  56756=>"100000000",
  56757=>"000000111",
  56758=>"000000111",
  56759=>"111111110",
  56760=>"000000111",
  56761=>"000000000",
  56762=>"000000011",
  56763=>"010111111",
  56764=>"001000000",
  56765=>"111111001",
  56766=>"111001000",
  56767=>"011011011",
  56768=>"111111010",
  56769=>"111111111",
  56770=>"000000000",
  56771=>"010000010",
  56772=>"111111111",
  56773=>"000010111",
  56774=>"000000011",
  56775=>"000001011",
  56776=>"111110000",
  56777=>"001000111",
  56778=>"000000001",
  56779=>"000000111",
  56780=>"000011001",
  56781=>"110110010",
  56782=>"111111111",
  56783=>"111111111",
  56784=>"111111110",
  56785=>"111111111",
  56786=>"000001001",
  56787=>"111000100",
  56788=>"000100111",
  56789=>"100111111",
  56790=>"100100101",
  56791=>"110110000",
  56792=>"111111100",
  56793=>"000000000",
  56794=>"111111100",
  56795=>"110110110",
  56796=>"101111111",
  56797=>"111100000",
  56798=>"000000010",
  56799=>"001011111",
  56800=>"000001000",
  56801=>"000100111",
  56802=>"111110110",
  56803=>"010000001",
  56804=>"110100100",
  56805=>"111111111",
  56806=>"000111111",
  56807=>"111101101",
  56808=>"011000000",
  56809=>"111100010",
  56810=>"000000000",
  56811=>"100110010",
  56812=>"000000110",
  56813=>"000000110",
  56814=>"111111111",
  56815=>"000000000",
  56816=>"110110100",
  56817=>"000000000",
  56818=>"000000111",
  56819=>"101000010",
  56820=>"111111111",
  56821=>"111000000",
  56822=>"000000000",
  56823=>"000000000",
  56824=>"011111010",
  56825=>"000111110",
  56826=>"001011011",
  56827=>"101111011",
  56828=>"000000100",
  56829=>"011111000",
  56830=>"111111011",
  56831=>"000001100",
  56832=>"000000000",
  56833=>"100100000",
  56834=>"101000000",
  56835=>"000001111",
  56836=>"000110111",
  56837=>"101000000",
  56838=>"000000000",
  56839=>"000000000",
  56840=>"111111111",
  56841=>"011111111",
  56842=>"000000000",
  56843=>"111101101",
  56844=>"110000000",
  56845=>"111100101",
  56846=>"011101000",
  56847=>"000000001",
  56848=>"110000000",
  56849=>"000110101",
  56850=>"111111111",
  56851=>"000000010",
  56852=>"000000100",
  56853=>"101111000",
  56854=>"011011110",
  56855=>"000000000",
  56856=>"000000000",
  56857=>"110000000",
  56858=>"000000001",
  56859=>"110000011",
  56860=>"101001101",
  56861=>"111110110",
  56862=>"101111001",
  56863=>"111110111",
  56864=>"000010000",
  56865=>"011100000",
  56866=>"100000000",
  56867=>"111111111",
  56868=>"000000111",
  56869=>"000000100",
  56870=>"010011001",
  56871=>"110110111",
  56872=>"000100111",
  56873=>"111101000",
  56874=>"111111111",
  56875=>"000000000",
  56876=>"101000000",
  56877=>"010111110",
  56878=>"000111011",
  56879=>"010000000",
  56880=>"100000001",
  56881=>"111111111",
  56882=>"111100011",
  56883=>"001101101",
  56884=>"001111111",
  56885=>"111111111",
  56886=>"001000000",
  56887=>"001111111",
  56888=>"000000000",
  56889=>"100000110",
  56890=>"111111111",
  56891=>"011000000",
  56892=>"000000000",
  56893=>"000011111",
  56894=>"110110111",
  56895=>"000111111",
  56896=>"111001000",
  56897=>"110110110",
  56898=>"111111111",
  56899=>"111111111",
  56900=>"010010000",
  56901=>"001001001",
  56902=>"111100000",
  56903=>"111111000",
  56904=>"011011011",
  56905=>"000000000",
  56906=>"100000000",
  56907=>"011001011",
  56908=>"111111111",
  56909=>"111000000",
  56910=>"000101101",
  56911=>"000000000",
  56912=>"000000000",
  56913=>"000000010",
  56914=>"111111001",
  56915=>"000000000",
  56916=>"000000000",
  56917=>"111110111",
  56918=>"111101000",
  56919=>"001011101",
  56920=>"100000000",
  56921=>"000000111",
  56922=>"011000000",
  56923=>"000000000",
  56924=>"000000000",
  56925=>"000000000",
  56926=>"111111111",
  56927=>"111111111",
  56928=>"100100000",
  56929=>"101000001",
  56930=>"101101111",
  56931=>"100100000",
  56932=>"000010010",
  56933=>"000000100",
  56934=>"101000111",
  56935=>"111111111",
  56936=>"000000000",
  56937=>"101000000",
  56938=>"001000000",
  56939=>"111111111",
  56940=>"111111111",
  56941=>"000000000",
  56942=>"100100100",
  56943=>"000000000",
  56944=>"000010111",
  56945=>"000000000",
  56946=>"111111111",
  56947=>"000000000",
  56948=>"011111111",
  56949=>"000110110",
  56950=>"000000000",
  56951=>"000000000",
  56952=>"011111100",
  56953=>"000110100",
  56954=>"111111100",
  56955=>"000000000",
  56956=>"100000110",
  56957=>"000000000",
  56958=>"111010100",
  56959=>"001001111",
  56960=>"101111111",
  56961=>"111100100",
  56962=>"111111110",
  56963=>"111111011",
  56964=>"100111000",
  56965=>"000000011",
  56966=>"110111111",
  56967=>"000000000",
  56968=>"111100000",
  56969=>"000111011",
  56970=>"000000110",
  56971=>"111111111",
  56972=>"111111111",
  56973=>"111001000",
  56974=>"011001110",
  56975=>"000000000",
  56976=>"000000000",
  56977=>"000010010",
  56978=>"111111000",
  56979=>"001000000",
  56980=>"000100111",
  56981=>"000100110",
  56982=>"000100000",
  56983=>"000000000",
  56984=>"110010010",
  56985=>"101111111",
  56986=>"100100101",
  56987=>"011011010",
  56988=>"000000110",
  56989=>"000000000",
  56990=>"000001111",
  56991=>"000000001",
  56992=>"000000000",
  56993=>"100100101",
  56994=>"000000010",
  56995=>"000000000",
  56996=>"111110000",
  56997=>"110110111",
  56998=>"101000111",
  56999=>"111011011",
  57000=>"001101111",
  57001=>"100111011",
  57002=>"110000000",
  57003=>"000000011",
  57004=>"000111111",
  57005=>"111001110",
  57006=>"110111111",
  57007=>"000000000",
  57008=>"001000000",
  57009=>"011011111",
  57010=>"111111111",
  57011=>"001000111",
  57012=>"000111111",
  57013=>"000000000",
  57014=>"111111111",
  57015=>"010010100",
  57016=>"100111111",
  57017=>"111111100",
  57018=>"111101001",
  57019=>"111111011",
  57020=>"100110110",
  57021=>"000000000",
  57022=>"110110111",
  57023=>"000000110",
  57024=>"100000000",
  57025=>"000000100",
  57026=>"000000111",
  57027=>"000000000",
  57028=>"000000100",
  57029=>"111100001",
  57030=>"000100111",
  57031=>"000000111",
  57032=>"111111111",
  57033=>"000000000",
  57034=>"000000001",
  57035=>"110000100",
  57036=>"100000001",
  57037=>"110000011",
  57038=>"100100011",
  57039=>"111111111",
  57040=>"010111111",
  57041=>"000010000",
  57042=>"000000000",
  57043=>"000000000",
  57044=>"111111111",
  57045=>"000000110",
  57046=>"111000000",
  57047=>"111111111",
  57048=>"101000000",
  57049=>"000100111",
  57050=>"001000000",
  57051=>"000000100",
  57052=>"110110111",
  57053=>"110111111",
  57054=>"101101111",
  57055=>"000000000",
  57056=>"011000000",
  57057=>"110111110",
  57058=>"000000111",
  57059=>"000000000",
  57060=>"001011011",
  57061=>"011110000",
  57062=>"111111111",
  57063=>"100111111",
  57064=>"000000000",
  57065=>"110110000",
  57066=>"000000000",
  57067=>"000000000",
  57068=>"101001001",
  57069=>"100110111",
  57070=>"110110100",
  57071=>"111111111",
  57072=>"111100100",
  57073=>"000000000",
  57074=>"000011011",
  57075=>"111001001",
  57076=>"010110100",
  57077=>"111111111",
  57078=>"100111011",
  57079=>"111111111",
  57080=>"011000000",
  57081=>"111000000",
  57082=>"100100110",
  57083=>"000011111",
  57084=>"010000000",
  57085=>"111111111",
  57086=>"111110111",
  57087=>"110111111",
  57088=>"011001011",
  57089=>"001001001",
  57090=>"111111111",
  57091=>"000000000",
  57092=>"111100100",
  57093=>"111111011",
  57094=>"000000011",
  57095=>"100000000",
  57096=>"100000100",
  57097=>"000000000",
  57098=>"111111111",
  57099=>"000000100",
  57100=>"001000001",
  57101=>"011011111",
  57102=>"000000000",
  57103=>"111111111",
  57104=>"000000000",
  57105=>"111011011",
  57106=>"111111111",
  57107=>"100000000",
  57108=>"011111111",
  57109=>"000001011",
  57110=>"000001001",
  57111=>"000110111",
  57112=>"111111111",
  57113=>"111110000",
  57114=>"011111000",
  57115=>"000110111",
  57116=>"111011111",
  57117=>"111111111",
  57118=>"000011111",
  57119=>"101001000",
  57120=>"111100001",
  57121=>"111111111",
  57122=>"010011111",
  57123=>"000000001",
  57124=>"111111001",
  57125=>"101111111",
  57126=>"001011001",
  57127=>"000000000",
  57128=>"000000000",
  57129=>"111111111",
  57130=>"100101011",
  57131=>"000000111",
  57132=>"000100110",
  57133=>"011011011",
  57134=>"000000000",
  57135=>"000000011",
  57136=>"000000000",
  57137=>"001001111",
  57138=>"111111111",
  57139=>"100111111",
  57140=>"101000000",
  57141=>"100100000",
  57142=>"000000000",
  57143=>"000000000",
  57144=>"011000000",
  57145=>"111111001",
  57146=>"001000000",
  57147=>"111111111",
  57148=>"000000000",
  57149=>"000000111",
  57150=>"000000011",
  57151=>"111101111",
  57152=>"111111111",
  57153=>"111111111",
  57154=>"000010000",
  57155=>"000000000",
  57156=>"111001000",
  57157=>"111111111",
  57158=>"000000000",
  57159=>"110111111",
  57160=>"110000000",
  57161=>"110110000",
  57162=>"111101001",
  57163=>"111111111",
  57164=>"000000000",
  57165=>"000000000",
  57166=>"111111100",
  57167=>"111111111",
  57168=>"001100100",
  57169=>"100000111",
  57170=>"001000000",
  57171=>"111111111",
  57172=>"000000000",
  57173=>"001011011",
  57174=>"111111100",
  57175=>"111111111",
  57176=>"000000000",
  57177=>"110110000",
  57178=>"100100011",
  57179=>"000000000",
  57180=>"000000000",
  57181=>"000000011",
  57182=>"000000000",
  57183=>"100000001",
  57184=>"100000000",
  57185=>"100000111",
  57186=>"110111011",
  57187=>"111111111",
  57188=>"000000000",
  57189=>"000000001",
  57190=>"111101110",
  57191=>"111111110",
  57192=>"111001101",
  57193=>"111111111",
  57194=>"011000000",
  57195=>"110110000",
  57196=>"110110110",
  57197=>"111001111",
  57198=>"111111111",
  57199=>"000000110",
  57200=>"110011000",
  57201=>"110100000",
  57202=>"110110010",
  57203=>"111111011",
  57204=>"000000000",
  57205=>"111111110",
  57206=>"111011011",
  57207=>"100110110",
  57208=>"001000011",
  57209=>"111000000",
  57210=>"001101101",
  57211=>"111111111",
  57212=>"001001001",
  57213=>"000000000",
  57214=>"111111001",
  57215=>"111111111",
  57216=>"111111111",
  57217=>"000110111",
  57218=>"110011010",
  57219=>"001000000",
  57220=>"000000111",
  57221=>"000000111",
  57222=>"000000000",
  57223=>"000000001",
  57224=>"001001111",
  57225=>"011100111",
  57226=>"111111111",
  57227=>"000011111",
  57228=>"101101111",
  57229=>"000110000",
  57230=>"100000010",
  57231=>"001000000",
  57232=>"000000000",
  57233=>"111000000",
  57234=>"100111111",
  57235=>"011000000",
  57236=>"111111011",
  57237=>"000100000",
  57238=>"001001011",
  57239=>"111001000",
  57240=>"001111111",
  57241=>"111000000",
  57242=>"111111111",
  57243=>"111111111",
  57244=>"111111111",
  57245=>"100100110",
  57246=>"111100111",
  57247=>"111111111",
  57248=>"001011000",
  57249=>"000111111",
  57250=>"011001111",
  57251=>"111111111",
  57252=>"000000000",
  57253=>"000000000",
  57254=>"111101111",
  57255=>"000000000",
  57256=>"010110100",
  57257=>"000000100",
  57258=>"000000000",
  57259=>"011111111",
  57260=>"101000000",
  57261=>"100000001",
  57262=>"111111111",
  57263=>"111111111",
  57264=>"111111111",
  57265=>"000110111",
  57266=>"111111111",
  57267=>"111111111",
  57268=>"100100000",
  57269=>"000000100",
  57270=>"000000110",
  57271=>"000111111",
  57272=>"000000011",
  57273=>"000000001",
  57274=>"100110011",
  57275=>"010111111",
  57276=>"111111111",
  57277=>"000111111",
  57278=>"000000000",
  57279=>"110100100",
  57280=>"111110011",
  57281=>"000000000",
  57282=>"111111111",
  57283=>"111111110",
  57284=>"101110000",
  57285=>"011001111",
  57286=>"110000000",
  57287=>"010010000",
  57288=>"011010111",
  57289=>"111111001",
  57290=>"011111100",
  57291=>"111111111",
  57292=>"101111000",
  57293=>"101000000",
  57294=>"000000001",
  57295=>"010111111",
  57296=>"000011001",
  57297=>"000000000",
  57298=>"101100000",
  57299=>"111110100",
  57300=>"111000000",
  57301=>"111101111",
  57302=>"000000100",
  57303=>"000000001",
  57304=>"000000000",
  57305=>"000000000",
  57306=>"000000000",
  57307=>"101101001",
  57308=>"001001001",
  57309=>"111110110",
  57310=>"000001000",
  57311=>"001011111",
  57312=>"111011001",
  57313=>"000100000",
  57314=>"000000000",
  57315=>"111101111",
  57316=>"000000010",
  57317=>"111111110",
  57318=>"111111111",
  57319=>"111111111",
  57320=>"000001001",
  57321=>"100100100",
  57322=>"000000000",
  57323=>"100000001",
  57324=>"111111001",
  57325=>"000000000",
  57326=>"000000100",
  57327=>"011111111",
  57328=>"111111100",
  57329=>"000001111",
  57330=>"000001000",
  57331=>"011000000",
  57332=>"111111111",
  57333=>"111111111",
  57334=>"111011000",
  57335=>"111111110",
  57336=>"000111111",
  57337=>"101001001",
  57338=>"000000110",
  57339=>"101001111",
  57340=>"011111111",
  57341=>"100000000",
  57342=>"110100000",
  57343=>"111111111",
  57344=>"111100000",
  57345=>"011011000",
  57346=>"101101111",
  57347=>"111111111",
  57348=>"011110000",
  57349=>"000000111",
  57350=>"111111011",
  57351=>"000100000",
  57352=>"011111111",
  57353=>"111100100",
  57354=>"000000000",
  57355=>"111001100",
  57356=>"111111001",
  57357=>"010000000",
  57358=>"000000000",
  57359=>"111111111",
  57360=>"100000001",
  57361=>"111110110",
  57362=>"111111001",
  57363=>"000000111",
  57364=>"000011000",
  57365=>"000110000",
  57366=>"000101111",
  57367=>"110110110",
  57368=>"011011111",
  57369=>"001111111",
  57370=>"010111110",
  57371=>"100111111",
  57372=>"011000100",
  57373=>"111111111",
  57374=>"000001000",
  57375=>"000101111",
  57376=>"111000001",
  57377=>"000000000",
  57378=>"111111111",
  57379=>"111000101",
  57380=>"000000000",
  57381=>"100100100",
  57382=>"000000000",
  57383=>"000101111",
  57384=>"000000111",
  57385=>"111011000",
  57386=>"000000000",
  57387=>"000000000",
  57388=>"000000000",
  57389=>"000101000",
  57390=>"001001001",
  57391=>"100000000",
  57392=>"000111111",
  57393=>"011111011",
  57394=>"000011111",
  57395=>"000000000",
  57396=>"111001001",
  57397=>"110010110",
  57398=>"000000100",
  57399=>"011000000",
  57400=>"000001001",
  57401=>"000001000",
  57402=>"010000000",
  57403=>"111000000",
  57404=>"101000111",
  57405=>"111111110",
  57406=>"111111000",
  57407=>"111111011",
  57408=>"100110110",
  57409=>"001001100",
  57410=>"011110000",
  57411=>"000000000",
  57412=>"000000000",
  57413=>"011111111",
  57414=>"000000100",
  57415=>"110000000",
  57416=>"110110000",
  57417=>"111111100",
  57418=>"000000000",
  57419=>"111111111",
  57420=>"101001001",
  57421=>"110100000",
  57422=>"111011000",
  57423=>"110100111",
  57424=>"111111111",
  57425=>"100111111",
  57426=>"000000000",
  57427=>"111110100",
  57428=>"111111011",
  57429=>"000000111",
  57430=>"110110111",
  57431=>"111111110",
  57432=>"111001111",
  57433=>"000000101",
  57434=>"000000001",
  57435=>"010110000",
  57436=>"010000110",
  57437=>"100000000",
  57438=>"000000000",
  57439=>"010010011",
  57440=>"000000000",
  57441=>"000000000",
  57442=>"000000000",
  57443=>"000000000",
  57444=>"000000000",
  57445=>"000000000",
  57446=>"001111111",
  57447=>"111111111",
  57448=>"111111111",
  57449=>"111110110",
  57450=>"000000010",
  57451=>"111110000",
  57452=>"111001111",
  57453=>"000001111",
  57454=>"100000100",
  57455=>"101101000",
  57456=>"000111111",
  57457=>"100000000",
  57458=>"010000000",
  57459=>"100110000",
  57460=>"011011011",
  57461=>"000100111",
  57462=>"001000000",
  57463=>"000000000",
  57464=>"000000011",
  57465=>"000101111",
  57466=>"010000110",
  57467=>"100000100",
  57468=>"001001001",
  57469=>"011111001",
  57470=>"010000000",
  57471=>"000111111",
  57472=>"111111111",
  57473=>"000000111",
  57474=>"000011111",
  57475=>"111001001",
  57476=>"011111111",
  57477=>"111110111",
  57478=>"100100000",
  57479=>"111000000",
  57480=>"111111111",
  57481=>"100000001",
  57482=>"111111111",
  57483=>"011111011",
  57484=>"000111111",
  57485=>"111110111",
  57486=>"000001111",
  57487=>"111001011",
  57488=>"000000000",
  57489=>"101000000",
  57490=>"001111111",
  57491=>"001001011",
  57492=>"010010110",
  57493=>"111011001",
  57494=>"111111111",
  57495=>"000101001",
  57496=>"101000000",
  57497=>"000000110",
  57498=>"111111111",
  57499=>"001000000",
  57500=>"010111111",
  57501=>"100110000",
  57502=>"111000101",
  57503=>"010000000",
  57504=>"000011011",
  57505=>"111000000",
  57506=>"001000111",
  57507=>"100111111",
  57508=>"110000000",
  57509=>"001000000",
  57510=>"110110000",
  57511=>"000000000",
  57512=>"100111111",
  57513=>"000001111",
  57514=>"111111111",
  57515=>"000000000",
  57516=>"000111111",
  57517=>"001111111",
  57518=>"100000100",
  57519=>"000001000",
  57520=>"001000000",
  57521=>"010010011",
  57522=>"111111010",
  57523=>"000001101",
  57524=>"111111001",
  57525=>"000000001",
  57526=>"000001001",
  57527=>"111111111",
  57528=>"100000000",
  57529=>"111111111",
  57530=>"111000110",
  57531=>"100000001",
  57532=>"000000100",
  57533=>"110111010",
  57534=>"000000101",
  57535=>"011001000",
  57536=>"100000000",
  57537=>"001000001",
  57538=>"101000110",
  57539=>"111100111",
  57540=>"111111000",
  57541=>"000000111",
  57542=>"000000111",
  57543=>"111111111",
  57544=>"110111111",
  57545=>"000111110",
  57546=>"100000111",
  57547=>"100100111",
  57548=>"111001111",
  57549=>"000000000",
  57550=>"010001000",
  57551=>"011011001",
  57552=>"000001001",
  57553=>"111111011",
  57554=>"000000010",
  57555=>"000001111",
  57556=>"111111111",
  57557=>"100000000",
  57558=>"000000000",
  57559=>"000100110",
  57560=>"111111000",
  57561=>"000000100",
  57562=>"111111111",
  57563=>"111001001",
  57564=>"111111111",
  57565=>"000000000",
  57566=>"110111011",
  57567=>"000000000",
  57568=>"101000000",
  57569=>"110110100",
  57570=>"000000110",
  57571=>"111111010",
  57572=>"000001001",
  57573=>"011111000",
  57574=>"000000110",
  57575=>"000000000",
  57576=>"010010010",
  57577=>"010111010",
  57578=>"101111110",
  57579=>"000000101",
  57580=>"001000001",
  57581=>"111111111",
  57582=>"000001011",
  57583=>"111111110",
  57584=>"000000111",
  57585=>"010111011",
  57586=>"000000000",
  57587=>"110101101",
  57588=>"111111111",
  57589=>"001000000",
  57590=>"110111111",
  57591=>"111111111",
  57592=>"000011111",
  57593=>"111111000",
  57594=>"000000001",
  57595=>"111001001",
  57596=>"001000011",
  57597=>"000000101",
  57598=>"000000000",
  57599=>"111101101",
  57600=>"100110111",
  57601=>"000110111",
  57602=>"111001111",
  57603=>"111111111",
  57604=>"000111111",
  57605=>"000000000",
  57606=>"111111111",
  57607=>"100111111",
  57608=>"000111111",
  57609=>"111110111",
  57610=>"111111111",
  57611=>"111111000",
  57612=>"010010000",
  57613=>"111111111",
  57614=>"110111111",
  57615=>"011111110",
  57616=>"001111111",
  57617=>"111000000",
  57618=>"000000111",
  57619=>"000000111",
  57620=>"000100111",
  57621=>"111101000",
  57622=>"111111011",
  57623=>"001010100",
  57624=>"011111111",
  57625=>"011001000",
  57626=>"110010000",
  57627=>"000011011",
  57628=>"111111011",
  57629=>"111111000",
  57630=>"011000000",
  57631=>"001011000",
  57632=>"111111111",
  57633=>"000111111",
  57634=>"011001001",
  57635=>"111111111",
  57636=>"101101100",
  57637=>"000110111",
  57638=>"010011111",
  57639=>"111110000",
  57640=>"000010000",
  57641=>"011001011",
  57642=>"001000010",
  57643=>"111101111",
  57644=>"111111001",
  57645=>"011111110",
  57646=>"000110000",
  57647=>"101111000",
  57648=>"000000101",
  57649=>"111110111",
  57650=>"111011111",
  57651=>"011111000",
  57652=>"110010100",
  57653=>"111111111",
  57654=>"000000000",
  57655=>"110011001",
  57656=>"001000000",
  57657=>"001000000",
  57658=>"000010010",
  57659=>"111000101",
  57660=>"111110111",
  57661=>"011011000",
  57662=>"011001011",
  57663=>"001000111",
  57664=>"111111111",
  57665=>"111110111",
  57666=>"000000101",
  57667=>"111111111",
  57668=>"000000000",
  57669=>"000111000",
  57670=>"111111111",
  57671=>"101000000",
  57672=>"000000000",
  57673=>"000000000",
  57674=>"001110111",
  57675=>"100110110",
  57676=>"111100100",
  57677=>"011110000",
  57678=>"100000000",
  57679=>"000000100",
  57680=>"001000000",
  57681=>"011001111",
  57682=>"010000110",
  57683=>"000001011",
  57684=>"000000000",
  57685=>"011001111",
  57686=>"111010000",
  57687=>"000000001",
  57688=>"111111001",
  57689=>"000000000",
  57690=>"000111011",
  57691=>"110111001",
  57692=>"000000000",
  57693=>"111111111",
  57694=>"000010111",
  57695=>"000000111",
  57696=>"001111000",
  57697=>"000000000",
  57698=>"100110110",
  57699=>"000111111",
  57700=>"111110110",
  57701=>"111101111",
  57702=>"110000111",
  57703=>"001000000",
  57704=>"001001001",
  57705=>"111111111",
  57706=>"011000001",
  57707=>"000000000",
  57708=>"001010000",
  57709=>"111000111",
  57710=>"011111110",
  57711=>"000000101",
  57712=>"101101001",
  57713=>"000011111",
  57714=>"111111000",
  57715=>"011011011",
  57716=>"010011010",
  57717=>"000000011",
  57718=>"000100100",
  57719=>"000110000",
  57720=>"001111011",
  57721=>"100111000",
  57722=>"001000000",
  57723=>"100000000",
  57724=>"000000000",
  57725=>"111111111",
  57726=>"000000111",
  57727=>"100110000",
  57728=>"011000010",
  57729=>"111000110",
  57730=>"000011000",
  57731=>"000000001",
  57732=>"000010001",
  57733=>"110000100",
  57734=>"000010110",
  57735=>"001000001",
  57736=>"000011000",
  57737=>"111000000",
  57738=>"000000000",
  57739=>"111110100",
  57740=>"111011101",
  57741=>"110100000",
  57742=>"000000111",
  57743=>"100100000",
  57744=>"000000000",
  57745=>"001001001",
  57746=>"111111111",
  57747=>"001011011",
  57748=>"011001001",
  57749=>"001001001",
  57750=>"100000100",
  57751=>"111110000",
  57752=>"111011000",
  57753=>"011001011",
  57754=>"111111000",
  57755=>"110100111",
  57756=>"111111111",
  57757=>"111110000",
  57758=>"001000111",
  57759=>"000000111",
  57760=>"001000000",
  57761=>"000000000",
  57762=>"111111000",
  57763=>"111100000",
  57764=>"100000110",
  57765=>"111111101",
  57766=>"000000100",
  57767=>"000000010",
  57768=>"111111000",
  57769=>"000000100",
  57770=>"111111111",
  57771=>"101000000",
  57772=>"101011000",
  57773=>"011000000",
  57774=>"000000000",
  57775=>"001011010",
  57776=>"011000111",
  57777=>"111111111",
  57778=>"000000000",
  57779=>"000000000",
  57780=>"111101101",
  57781=>"000000111",
  57782=>"000000111",
  57783=>"011010010",
  57784=>"000001000",
  57785=>"011001000",
  57786=>"001001111",
  57787=>"010000001",
  57788=>"001001000",
  57789=>"011000110",
  57790=>"101101001",
  57791=>"110011001",
  57792=>"000111011",
  57793=>"000001001",
  57794=>"010011000",
  57795=>"000111000",
  57796=>"111000101",
  57797=>"000000100",
  57798=>"000010000",
  57799=>"001001001",
  57800=>"110110000",
  57801=>"001000000",
  57802=>"001000000",
  57803=>"000111000",
  57804=>"000111000",
  57805=>"111110111",
  57806=>"111001000",
  57807=>"001101111",
  57808=>"111111000",
  57809=>"111111111",
  57810=>"011111011",
  57811=>"011111111",
  57812=>"111001101",
  57813=>"100000001",
  57814=>"000000100",
  57815=>"111111011",
  57816=>"001111111",
  57817=>"101000111",
  57818=>"101100000",
  57819=>"101101001",
  57820=>"010111111",
  57821=>"000000110",
  57822=>"011111111",
  57823=>"100110110",
  57824=>"110111110",
  57825=>"001000000",
  57826=>"001000001",
  57827=>"111000000",
  57828=>"111111111",
  57829=>"111111010",
  57830=>"100100000",
  57831=>"111100000",
  57832=>"111101100",
  57833=>"000101001",
  57834=>"111111111",
  57835=>"000000011",
  57836=>"001000000",
  57837=>"111111001",
  57838=>"100100000",
  57839=>"010111110",
  57840=>"000000011",
  57841=>"111000010",
  57842=>"110000000",
  57843=>"000001011",
  57844=>"110101111",
  57845=>"111101111",
  57846=>"111000000",
  57847=>"000011110",
  57848=>"000010111",
  57849=>"010010000",
  57850=>"000010110",
  57851=>"000000000",
  57852=>"000000000",
  57853=>"111101101",
  57854=>"011001001",
  57855=>"111101101",
  57856=>"010000110",
  57857=>"011011010",
  57858=>"000000000",
  57859=>"111111111",
  57860=>"000000000",
  57861=>"110110111",
  57862=>"001000000",
  57863=>"000000000",
  57864=>"111000000",
  57865=>"111111001",
  57866=>"000000000",
  57867=>"110000000",
  57868=>"111111111",
  57869=>"110111111",
  57870=>"000000000",
  57871=>"111111111",
  57872=>"000000000",
  57873=>"000011111",
  57874=>"111101001",
  57875=>"111010111",
  57876=>"010000001",
  57877=>"111011100",
  57878=>"111111111",
  57879=>"111111111",
  57880=>"111111111",
  57881=>"110110000",
  57882=>"111111101",
  57883=>"000000001",
  57884=>"111111111",
  57885=>"000000000",
  57886=>"110100100",
  57887=>"111111011",
  57888=>"000000000",
  57889=>"111111111",
  57890=>"000111111",
  57891=>"111111111",
  57892=>"011001000",
  57893=>"001000000",
  57894=>"000100111",
  57895=>"101111111",
  57896=>"111111000",
  57897=>"111100111",
  57898=>"111111111",
  57899=>"001000011",
  57900=>"111111111",
  57901=>"110111111",
  57902=>"000000000",
  57903=>"111111111",
  57904=>"010111100",
  57905=>"111111111",
  57906=>"000011000",
  57907=>"111111111",
  57908=>"111111111",
  57909=>"000000000",
  57910=>"101000100",
  57911=>"000000000",
  57912=>"110010000",
  57913=>"110000000",
  57914=>"111111111",
  57915=>"100000000",
  57916=>"000000111",
  57917=>"000000000",
  57918=>"000000000",
  57919=>"000000000",
  57920=>"100000000",
  57921=>"000000000",
  57922=>"000000000",
  57923=>"111111111",
  57924=>"000001101",
  57925=>"110110110",
  57926=>"111011011",
  57927=>"000000110",
  57928=>"110100100",
  57929=>"111111111",
  57930=>"111111111",
  57931=>"111111110",
  57932=>"000000111",
  57933=>"110110100",
  57934=>"000001001",
  57935=>"000000000",
  57936=>"000000000",
  57937=>"000001001",
  57938=>"111111111",
  57939=>"100100000",
  57940=>"000000000",
  57941=>"111111000",
  57942=>"111100000",
  57943=>"101111111",
  57944=>"001001001",
  57945=>"001001001",
  57946=>"000000000",
  57947=>"111111111",
  57948=>"111111000",
  57949=>"000000000",
  57950=>"100000000",
  57951=>"100000000",
  57952=>"111111111",
  57953=>"110111111",
  57954=>"111111111",
  57955=>"101100111",
  57956=>"111111001",
  57957=>"110010000",
  57958=>"111111000",
  57959=>"111110000",
  57960=>"000101101",
  57961=>"110111111",
  57962=>"111001000",
  57963=>"000000000",
  57964=>"000000000",
  57965=>"000000000",
  57966=>"000011101",
  57967=>"000000000",
  57968=>"000000110",
  57969=>"000100000",
  57970=>"100100100",
  57971=>"100101111",
  57972=>"111000111",
  57973=>"011001001",
  57974=>"001011111",
  57975=>"111111111",
  57976=>"100010011",
  57977=>"110100100",
  57978=>"000000000",
  57979=>"111111011",
  57980=>"100110111",
  57981=>"001111111",
  57982=>"111111100",
  57983=>"000111110",
  57984=>"000000000",
  57985=>"000000100",
  57986=>"000001000",
  57987=>"111110000",
  57988=>"111111111",
  57989=>"111001111",
  57990=>"011011011",
  57991=>"000000000",
  57992=>"101111111",
  57993=>"111111111",
  57994=>"111111111",
  57995=>"011011111",
  57996=>"000000100",
  57997=>"101101111",
  57998=>"100101111",
  57999=>"011011000",
  58000=>"000000111",
  58001=>"000000000",
  58002=>"001000000",
  58003=>"000000100",
  58004=>"111111100",
  58005=>"010010010",
  58006=>"000000000",
  58007=>"000000000",
  58008=>"000000000",
  58009=>"111111111",
  58010=>"111111111",
  58011=>"000000000",
  58012=>"111001001",
  58013=>"111010000",
  58014=>"001011111",
  58015=>"110010111",
  58016=>"111000000",
  58017=>"000000000",
  58018=>"000001100",
  58019=>"111111010",
  58020=>"111100100",
  58021=>"000000000",
  58022=>"100000000",
  58023=>"010000000",
  58024=>"111111111",
  58025=>"000000000",
  58026=>"111111111",
  58027=>"010111110",
  58028=>"111111111",
  58029=>"110101101",
  58030=>"011111101",
  58031=>"000010001",
  58032=>"111111111",
  58033=>"000010000",
  58034=>"110111111",
  58035=>"100100100",
  58036=>"011101000",
  58037=>"110110001",
  58038=>"111000000",
  58039=>"000000000",
  58040=>"001101111",
  58041=>"000000000",
  58042=>"001011000",
  58043=>"000000000",
  58044=>"000000001",
  58045=>"100100111",
  58046=>"111111111",
  58047=>"111100111",
  58048=>"111100111",
  58049=>"111000000",
  58050=>"000111110",
  58051=>"000100000",
  58052=>"111111111",
  58053=>"000000000",
  58054=>"111001000",
  58055=>"111111111",
  58056=>"000000000",
  58057=>"111011011",
  58058=>"000000000",
  58059=>"001001111",
  58060=>"000000110",
  58061=>"000010111",
  58062=>"100101000",
  58063=>"000000000",
  58064=>"001111111",
  58065=>"000011111",
  58066=>"111000111",
  58067=>"000001000",
  58068=>"000000000",
  58069=>"000000000",
  58070=>"011011011",
  58071=>"000000000",
  58072=>"111111111",
  58073=>"000000000",
  58074=>"100000000",
  58075=>"011111111",
  58076=>"111111011",
  58077=>"000000000",
  58078=>"111010100",
  58079=>"111111011",
  58080=>"000000000",
  58081=>"000000110",
  58082=>"001011001",
  58083=>"000000000",
  58084=>"011011111",
  58085=>"111111110",
  58086=>"001000000",
  58087=>"001001001",
  58088=>"000000000",
  58089=>"111111111",
  58090=>"111111111",
  58091=>"000010000",
  58092=>"100111111",
  58093=>"000000100",
  58094=>"100000111",
  58095=>"111111111",
  58096=>"000000000",
  58097=>"111111111",
  58098=>"111111111",
  58099=>"100100100",
  58100=>"111111111",
  58101=>"001011111",
  58102=>"001101111",
  58103=>"111111110",
  58104=>"000000000",
  58105=>"100101111",
  58106=>"000000000",
  58107=>"110110111",
  58108=>"111111111",
  58109=>"000000001",
  58110=>"111011111",
  58111=>"011011111",
  58112=>"000000000",
  58113=>"111011011",
  58114=>"100100111",
  58115=>"000000101",
  58116=>"000000000",
  58117=>"000000000",
  58118=>"001001001",
  58119=>"001000100",
  58120=>"011000001",
  58121=>"111000100",
  58122=>"111110010",
  58123=>"000001001",
  58124=>"111011111",
  58125=>"000000000",
  58126=>"000000001",
  58127=>"000001001",
  58128=>"101010111",
  58129=>"000000000",
  58130=>"000000000",
  58131=>"111111111",
  58132=>"000000000",
  58133=>"000000000",
  58134=>"111001011",
  58135=>"111001001",
  58136=>"000000000",
  58137=>"110111111",
  58138=>"111111111",
  58139=>"100111101",
  58140=>"111111111",
  58141=>"000000000",
  58142=>"000000000",
  58143=>"111111111",
  58144=>"111111111",
  58145=>"000000000",
  58146=>"000000000",
  58147=>"000000101",
  58148=>"111111111",
  58149=>"111111111",
  58150=>"111111111",
  58151=>"010100100",
  58152=>"000010110",
  58153=>"111000000",
  58154=>"111111111",
  58155=>"000000000",
  58156=>"010010110",
  58157=>"000111001",
  58158=>"111110000",
  58159=>"001001111",
  58160=>"000000000",
  58161=>"001000000",
  58162=>"111111111",
  58163=>"000000000",
  58164=>"011000000",
  58165=>"111011011",
  58166=>"111100100",
  58167=>"101111111",
  58168=>"001001101",
  58169=>"000000000",
  58170=>"000000111",
  58171=>"000000011",
  58172=>"000001001",
  58173=>"101111100",
  58174=>"000000000",
  58175=>"111001011",
  58176=>"110111111",
  58177=>"111111111",
  58178=>"111111011",
  58179=>"111111111",
  58180=>"000100000",
  58181=>"000011011",
  58182=>"000100100",
  58183=>"001001001",
  58184=>"111111111",
  58185=>"100000000",
  58186=>"000100111",
  58187=>"100111111",
  58188=>"111111111",
  58189=>"101101000",
  58190=>"110000001",
  58191=>"011011011",
  58192=>"000000000",
  58193=>"000000000",
  58194=>"100100111",
  58195=>"000010111",
  58196=>"000110110",
  58197=>"011011111",
  58198=>"111111111",
  58199=>"111001101",
  58200=>"000000000",
  58201=>"110111111",
  58202=>"110110100",
  58203=>"000000000",
  58204=>"100101100",
  58205=>"011011111",
  58206=>"000000000",
  58207=>"000000110",
  58208=>"000000000",
  58209=>"111111111",
  58210=>"001100111",
  58211=>"001011000",
  58212=>"000011111",
  58213=>"000000000",
  58214=>"000000111",
  58215=>"011111111",
  58216=>"111100100",
  58217=>"111111011",
  58218=>"000010000",
  58219=>"111110110",
  58220=>"110110111",
  58221=>"011001101",
  58222=>"010000100",
  58223=>"111111010",
  58224=>"111000000",
  58225=>"010001011",
  58226=>"000000111",
  58227=>"010110100",
  58228=>"111111000",
  58229=>"011001001",
  58230=>"000000000",
  58231=>"111111111",
  58232=>"111111111",
  58233=>"100010111",
  58234=>"011101111",
  58235=>"010000000",
  58236=>"000000000",
  58237=>"010110010",
  58238=>"000000111",
  58239=>"111111111",
  58240=>"111111111",
  58241=>"111111111",
  58242=>"111111111",
  58243=>"111101111",
  58244=>"000010111",
  58245=>"111111111",
  58246=>"000000111",
  58247=>"001001111",
  58248=>"000101111",
  58249=>"101100111",
  58250=>"000000000",
  58251=>"001001011",
  58252=>"111111111",
  58253=>"011111111",
  58254=>"000000000",
  58255=>"111111100",
  58256=>"101100111",
  58257=>"111111111",
  58258=>"000000000",
  58259=>"111110111",
  58260=>"000000000",
  58261=>"000000000",
  58262=>"111110100",
  58263=>"110100000",
  58264=>"001001000",
  58265=>"111011011",
  58266=>"111111111",
  58267=>"000000111",
  58268=>"001000000",
  58269=>"100111111",
  58270=>"000000001",
  58271=>"000000000",
  58272=>"000000000",
  58273=>"110010000",
  58274=>"000000000",
  58275=>"000000000",
  58276=>"000001001",
  58277=>"110111111",
  58278=>"100111011",
  58279=>"000000011",
  58280=>"100100011",
  58281=>"000000100",
  58282=>"000000000",
  58283=>"000000000",
  58284=>"000000000",
  58285=>"111111011",
  58286=>"011011001",
  58287=>"111111111",
  58288=>"100000000",
  58289=>"000000111",
  58290=>"001001000",
  58291=>"000000111",
  58292=>"111110011",
  58293=>"101100100",
  58294=>"111111001",
  58295=>"111111111",
  58296=>"000000000",
  58297=>"000110111",
  58298=>"111111111",
  58299=>"100000000",
  58300=>"000111111",
  58301=>"000000000",
  58302=>"000111111",
  58303=>"001000000",
  58304=>"000000000",
  58305=>"111111000",
  58306=>"000000000",
  58307=>"111111111",
  58308=>"111100000",
  58309=>"001000100",
  58310=>"111111111",
  58311=>"111011011",
  58312=>"111100001",
  58313=>"111010000",
  58314=>"000000100",
  58315=>"111111111",
  58316=>"110100000",
  58317=>"111000000",
  58318=>"001010110",
  58319=>"000000000",
  58320=>"001000001",
  58321=>"000000000",
  58322=>"110000000",
  58323=>"111111000",
  58324=>"110111111",
  58325=>"111110010",
  58326=>"000000001",
  58327=>"011011111",
  58328=>"000000000",
  58329=>"000000000",
  58330=>"000000000",
  58331=>"100000000",
  58332=>"011100100",
  58333=>"000100100",
  58334=>"000000100",
  58335=>"000000101",
  58336=>"111111111",
  58337=>"000000000",
  58338=>"000000000",
  58339=>"111111110",
  58340=>"000000000",
  58341=>"010111111",
  58342=>"001000000",
  58343=>"111111111",
  58344=>"111111111",
  58345=>"101111111",
  58346=>"011011000",
  58347=>"111111010",
  58348=>"110111001",
  58349=>"001000000",
  58350=>"001000000",
  58351=>"001000101",
  58352=>"000000000",
  58353=>"111111111",
  58354=>"000000000",
  58355=>"111111111",
  58356=>"100100000",
  58357=>"000000000",
  58358=>"111111111",
  58359=>"010010110",
  58360=>"000100001",
  58361=>"001101101",
  58362=>"000101111",
  58363=>"100000110",
  58364=>"111111000",
  58365=>"111111111",
  58366=>"111111111",
  58367=>"111000000",
  58368=>"111011100",
  58369=>"000000000",
  58370=>"000000111",
  58371=>"000000000",
  58372=>"000110111",
  58373=>"000000000",
  58374=>"101101101",
  58375=>"111111111",
  58376=>"111100000",
  58377=>"111111111",
  58378=>"000000011",
  58379=>"101101001",
  58380=>"011111111",
  58381=>"000000000",
  58382=>"111111000",
  58383=>"101111111",
  58384=>"110110111",
  58385=>"000000001",
  58386=>"111000000",
  58387=>"000000111",
  58388=>"000000000",
  58389=>"111111110",
  58390=>"110111111",
  58391=>"111111000",
  58392=>"111110100",
  58393=>"001001011",
  58394=>"001000010",
  58395=>"111101001",
  58396=>"111111111",
  58397=>"111111011",
  58398=>"111111110",
  58399=>"101100000",
  58400=>"100111101",
  58401=>"111111111",
  58402=>"111111011",
  58403=>"110111000",
  58404=>"000111111",
  58405=>"000111111",
  58406=>"000001111",
  58407=>"001001001",
  58408=>"000010111",
  58409=>"000000000",
  58410=>"000000101",
  58411=>"110110111",
  58412=>"100000111",
  58413=>"110111111",
  58414=>"111111111",
  58415=>"111111011",
  58416=>"011111111",
  58417=>"100000001",
  58418=>"011011001",
  58419=>"000000000",
  58420=>"000000111",
  58421=>"001001000",
  58422=>"000000101",
  58423=>"111011000",
  58424=>"000000000",
  58425=>"001011110",
  58426=>"001000001",
  58427=>"111110111",
  58428=>"000001111",
  58429=>"000000000",
  58430=>"111010000",
  58431=>"111011000",
  58432=>"111100000",
  58433=>"000000111",
  58434=>"101000011",
  58435=>"101111001",
  58436=>"111011111",
  58437=>"111100000",
  58438=>"101000000",
  58439=>"111111111",
  58440=>"100000000",
  58441=>"000000111",
  58442=>"111111010",
  58443=>"111111111",
  58444=>"000000000",
  58445=>"111011011",
  58446=>"000000000",
  58447=>"110011110",
  58448=>"111111111",
  58449=>"100010000",
  58450=>"100100000",
  58451=>"000000000",
  58452=>"111111111",
  58453=>"001111000",
  58454=>"011111111",
  58455=>"000000001",
  58456=>"011100000",
  58457=>"000001111",
  58458=>"111110010",
  58459=>"110110110",
  58460=>"000000000",
  58461=>"011111001",
  58462=>"111111000",
  58463=>"111111111",
  58464=>"100000000",
  58465=>"000000000",
  58466=>"010000010",
  58467=>"110110110",
  58468=>"010010101",
  58469=>"010001001",
  58470=>"000000000",
  58471=>"000000000",
  58472=>"000000000",
  58473=>"111111110",
  58474=>"000000000",
  58475=>"000011111",
  58476=>"111111100",
  58477=>"000110111",
  58478=>"000000000",
  58479=>"000000000",
  58480=>"000111000",
  58481=>"000000000",
  58482=>"100100110",
  58483=>"001000000",
  58484=>"100001111",
  58485=>"111001001",
  58486=>"000000000",
  58487=>"111001001",
  58488=>"111111111",
  58489=>"111111011",
  58490=>"111111010",
  58491=>"010000011",
  58492=>"011111001",
  58493=>"001001111",
  58494=>"100010011",
  58495=>"111111000",
  58496=>"011000111",
  58497=>"111011000",
  58498=>"111000111",
  58499=>"000000000",
  58500=>"111111111",
  58501=>"101000000",
  58502=>"111010100",
  58503=>"111010000",
  58504=>"011011011",
  58505=>"111000000",
  58506=>"011000000",
  58507=>"000000000",
  58508=>"000100000",
  58509=>"101100100",
  58510=>"000000010",
  58511=>"000111111",
  58512=>"000000110",
  58513=>"000000111",
  58514=>"110111000",
  58515=>"111100000",
  58516=>"011111111",
  58517=>"111001001",
  58518=>"111000000",
  58519=>"011000000",
  58520=>"111011001",
  58521=>"001001101",
  58522=>"000000000",
  58523=>"000000000",
  58524=>"111111000",
  58525=>"111111000",
  58526=>"111111111",
  58527=>"101111111",
  58528=>"111111010",
  58529=>"100100000",
  58530=>"000001111",
  58531=>"000011000",
  58532=>"000000101",
  58533=>"100100000",
  58534=>"111111111",
  58535=>"110100110",
  58536=>"001001011",
  58537=>"010000100",
  58538=>"001000000",
  58539=>"001001001",
  58540=>"111111110",
  58541=>"111111000",
  58542=>"111111111",
  58543=>"111111111",
  58544=>"001000001",
  58545=>"100111111",
  58546=>"110110110",
  58547=>"000000010",
  58548=>"000001001",
  58549=>"111111111",
  58550=>"111001111",
  58551=>"111111111",
  58552=>"000000100",
  58553=>"110111111",
  58554=>"100100000",
  58555=>"011011000",
  58556=>"010010000",
  58557=>"111010000",
  58558=>"111000000",
  58559=>"000000001",
  58560=>"000000010",
  58561=>"111111111",
  58562=>"000011010",
  58563=>"000000000",
  58564=>"111101111",
  58565=>"111111000",
  58566=>"101000100",
  58567=>"000000000",
  58568=>"111111111",
  58569=>"101000111",
  58570=>"101011000",
  58571=>"111111101",
  58572=>"000000000",
  58573=>"110110111",
  58574=>"000011011",
  58575=>"001011011",
  58576=>"011111001",
  58577=>"000000000",
  58578=>"011001111",
  58579=>"000000011",
  58580=>"000000000",
  58581=>"001001001",
  58582=>"000111000",
  58583=>"000000000",
  58584=>"001000000",
  58585=>"000000000",
  58586=>"111011000",
  58587=>"000000101",
  58588=>"001001000",
  58589=>"000000111",
  58590=>"000000101",
  58591=>"011101110",
  58592=>"000000011",
  58593=>"000000000",
  58594=>"111111001",
  58595=>"111111110",
  58596=>"111111011",
  58597=>"110000001",
  58598=>"100000010",
  58599=>"111111000",
  58600=>"111111111",
  58601=>"111111111",
  58602=>"011011011",
  58603=>"000000000",
  58604=>"100000100",
  58605=>"010110110",
  58606=>"011111111",
  58607=>"000000000",
  58608=>"111111100",
  58609=>"000001000",
  58610=>"000110100",
  58611=>"000111011",
  58612=>"111111100",
  58613=>"111011110",
  58614=>"000000000",
  58615=>"011000011",
  58616=>"000100111",
  58617=>"000000010",
  58618=>"001001111",
  58619=>"111101111",
  58620=>"111011001",
  58621=>"111111010",
  58622=>"111111000",
  58623=>"101100000",
  58624=>"011011000",
  58625=>"001001111",
  58626=>"001011111",
  58627=>"000000111",
  58628=>"111110100",
  58629=>"000000000",
  58630=>"001001111",
  58631=>"011001000",
  58632=>"111111111",
  58633=>"000000000",
  58634=>"110000000",
  58635=>"000001111",
  58636=>"000000111",
  58637=>"111100110",
  58638=>"100000000",
  58639=>"000111001",
  58640=>"010111111",
  58641=>"000001111",
  58642=>"001000000",
  58643=>"111111001",
  58644=>"000000100",
  58645=>"111111011",
  58646=>"111111110",
  58647=>"100000000",
  58648=>"000000000",
  58649=>"000000000",
  58650=>"000001000",
  58651=>"111111000",
  58652=>"100110000",
  58653=>"000111111",
  58654=>"111111111",
  58655=>"000000001",
  58656=>"001000000",
  58657=>"000000111",
  58658=>"011111000",
  58659=>"000000000",
  58660=>"111010110",
  58661=>"110110111",
  58662=>"000000000",
  58663=>"000000000",
  58664=>"000000000",
  58665=>"111001001",
  58666=>"100000000",
  58667=>"000000000",
  58668=>"111000001",
  58669=>"001011100",
  58670=>"111111011",
  58671=>"000100100",
  58672=>"111111111",
  58673=>"111111111",
  58674=>"110111100",
  58675=>"000000000",
  58676=>"001000000",
  58677=>"111111101",
  58678=>"011111011",
  58679=>"111100000",
  58680=>"111111000",
  58681=>"111000111",
  58682=>"111100100",
  58683=>"000001111",
  58684=>"000001001",
  58685=>"101111111",
  58686=>"000000100",
  58687=>"001011000",
  58688=>"110110000",
  58689=>"100111111",
  58690=>"010010010",
  58691=>"111111000",
  58692=>"000000110",
  58693=>"000011111",
  58694=>"111100000",
  58695=>"011001111",
  58696=>"111111111",
  58697=>"111011000",
  58698=>"111110000",
  58699=>"111110010",
  58700=>"100000000",
  58701=>"111110000",
  58702=>"000000001",
  58703=>"000000011",
  58704=>"011001011",
  58705=>"001001000",
  58706=>"000011111",
  58707=>"111111111",
  58708=>"000000111",
  58709=>"011011001",
  58710=>"000000000",
  58711=>"000111111",
  58712=>"100000000",
  58713=>"000000000",
  58714=>"000111000",
  58715=>"010110000",
  58716=>"011111111",
  58717=>"111001111",
  58718=>"111111001",
  58719=>"011011000",
  58720=>"000111111",
  58721=>"000000111",
  58722=>"111111011",
  58723=>"000000100",
  58724=>"111111011",
  58725=>"100000000",
  58726=>"111000000",
  58727=>"111111111",
  58728=>"111111000",
  58729=>"011111000",
  58730=>"110111110",
  58731=>"001001011",
  58732=>"100110110",
  58733=>"101111111",
  58734=>"000101111",
  58735=>"000111111",
  58736=>"011000000",
  58737=>"111111100",
  58738=>"010111111",
  58739=>"110110110",
  58740=>"111111000",
  58741=>"000000100",
  58742=>"000000000",
  58743=>"010000000",
  58744=>"011111111",
  58745=>"111111011",
  58746=>"000000011",
  58747=>"111111001",
  58748=>"000000000",
  58749=>"110110111",
  58750=>"111111111",
  58751=>"111111011",
  58752=>"000010000",
  58753=>"011000101",
  58754=>"111011011",
  58755=>"110110110",
  58756=>"101001111",
  58757=>"000000100",
  58758=>"011000110",
  58759=>"101011011",
  58760=>"010110110",
  58761=>"001001100",
  58762=>"111111000",
  58763=>"111010000",
  58764=>"000000111",
  58765=>"000001000",
  58766=>"000011001",
  58767=>"100100000",
  58768=>"010111000",
  58769=>"110111111",
  58770=>"000000001",
  58771=>"110110100",
  58772=>"000111111",
  58773=>"000111111",
  58774=>"000111111",
  58775=>"111111111",
  58776=>"101101000",
  58777=>"111000000",
  58778=>"001011111",
  58779=>"111111111",
  58780=>"111111000",
  58781=>"100110010",
  58782=>"000011111",
  58783=>"010110000",
  58784=>"111011001",
  58785=>"011011011",
  58786=>"000110110",
  58787=>"000000000",
  58788=>"010000000",
  58789=>"110100101",
  58790=>"111111000",
  58791=>"111111111",
  58792=>"110000000",
  58793=>"000000000",
  58794=>"011111111",
  58795=>"001001000",
  58796=>"000000000",
  58797=>"011100100",
  58798=>"000000110",
  58799=>"000000111",
  58800=>"000000110",
  58801=>"101001000",
  58802=>"000000100",
  58803=>"010001001",
  58804=>"000000011",
  58805=>"001001100",
  58806=>"100000000",
  58807=>"001000000",
  58808=>"000011111",
  58809=>"010111111",
  58810=>"000000000",
  58811=>"111111111",
  58812=>"000000000",
  58813=>"100000111",
  58814=>"111000000",
  58815=>"000000011",
  58816=>"111011011",
  58817=>"000110100",
  58818=>"111111111",
  58819=>"111111000",
  58820=>"010111100",
  58821=>"100001111",
  58822=>"000000000",
  58823=>"100111111",
  58824=>"000000000",
  58825=>"000000000",
  58826=>"000110110",
  58827=>"000110000",
  58828=>"111000000",
  58829=>"100100000",
  58830=>"111111000",
  58831=>"111110000",
  58832=>"110100000",
  58833=>"110111111",
  58834=>"000000000",
  58835=>"001000101",
  58836=>"111111011",
  58837=>"111010000",
  58838=>"000100000",
  58839=>"110110001",
  58840=>"000011011",
  58841=>"111001101",
  58842=>"100000110",
  58843=>"011010000",
  58844=>"111110000",
  58845=>"111110011",
  58846=>"000000001",
  58847=>"000000100",
  58848=>"110100000",
  58849=>"111111111",
  58850=>"000000000",
  58851=>"000000000",
  58852=>"000000001",
  58853=>"001101111",
  58854=>"001000000",
  58855=>"000000001",
  58856=>"000000001",
  58857=>"011111110",
  58858=>"111001001",
  58859=>"011010011",
  58860=>"000000110",
  58861=>"101100000",
  58862=>"000000101",
  58863=>"100111100",
  58864=>"001000000",
  58865=>"011110110",
  58866=>"101101001",
  58867=>"010010000",
  58868=>"000010011",
  58869=>"111001000",
  58870=>"111110010",
  58871=>"111111110",
  58872=>"000101111",
  58873=>"000000000",
  58874=>"000000000",
  58875=>"111111000",
  58876=>"000000100",
  58877=>"111000101",
  58878=>"000100110",
  58879=>"000000100",
  58880=>"111111111",
  58881=>"001000111",
  58882=>"000000000",
  58883=>"110000000",
  58884=>"000000000",
  58885=>"110000000",
  58886=>"000000000",
  58887=>"111111111",
  58888=>"011001101",
  58889=>"000000000",
  58890=>"000000000",
  58891=>"000110111",
  58892=>"000110110",
  58893=>"011000000",
  58894=>"111111111",
  58895=>"100101000",
  58896=>"111111111",
  58897=>"100000000",
  58898=>"111111111",
  58899=>"000000000",
  58900=>"110110100",
  58901=>"111111111",
  58902=>"111001000",
  58903=>"011011001",
  58904=>"110110110",
  58905=>"110000000",
  58906=>"111111111",
  58907=>"111001111",
  58908=>"000000000",
  58909=>"000000000",
  58910=>"111111001",
  58911=>"100110111",
  58912=>"001011011",
  58913=>"000001001",
  58914=>"111111011",
  58915=>"001111111",
  58916=>"110010010",
  58917=>"000001001",
  58918=>"000011011",
  58919=>"000000011",
  58920=>"000000000",
  58921=>"000111111",
  58922=>"000000100",
  58923=>"111011000",
  58924=>"100100111",
  58925=>"111001000",
  58926=>"000011111",
  58927=>"011010111",
  58928=>"000000100",
  58929=>"100000000",
  58930=>"001001001",
  58931=>"111011011",
  58932=>"000000000",
  58933=>"000000100",
  58934=>"000000000",
  58935=>"100100100",
  58936=>"111111111",
  58937=>"100100100",
  58938=>"000000000",
  58939=>"001001011",
  58940=>"000000000",
  58941=>"000000000",
  58942=>"000110000",
  58943=>"111111011",
  58944=>"000000000",
  58945=>"110110000",
  58946=>"000001011",
  58947=>"000110110",
  58948=>"000010111",
  58949=>"000000000",
  58950=>"000000000",
  58951=>"111111111",
  58952=>"001001000",
  58953=>"111100100",
  58954=>"011111011",
  58955=>"111000000",
  58956=>"000000000",
  58957=>"000000000",
  58958=>"000110110",
  58959=>"111111111",
  58960=>"111111111",
  58961=>"000000000",
  58962=>"000000000",
  58963=>"111111001",
  58964=>"000000000",
  58965=>"000010110",
  58966=>"000100111",
  58967=>"000000001",
  58968=>"000000010",
  58969=>"000000000",
  58970=>"111111111",
  58971=>"001000000",
  58972=>"111110000",
  58973=>"111001010",
  58974=>"000000000",
  58975=>"010110110",
  58976=>"000000000",
  58977=>"000000100",
  58978=>"000000000",
  58979=>"111111111",
  58980=>"100001000",
  58981=>"000000110",
  58982=>"110000000",
  58983=>"111110100",
  58984=>"000000000",
  58985=>"000111111",
  58986=>"000000000",
  58987=>"000000000",
  58988=>"000100000",
  58989=>"111111111",
  58990=>"000111110",
  58991=>"000000000",
  58992=>"000000000",
  58993=>"000000000",
  58994=>"011111111",
  58995=>"111111111",
  58996=>"110110100",
  58997=>"111111111",
  58998=>"111111011",
  58999=>"011011011",
  59000=>"010000000",
  59001=>"000000000",
  59002=>"100100001",
  59003=>"000001001",
  59004=>"110000000",
  59005=>"011111111",
  59006=>"000000000",
  59007=>"000011000",
  59008=>"000000000",
  59009=>"000001011",
  59010=>"111111111",
  59011=>"000001000",
  59012=>"011010101",
  59013=>"101111111",
  59014=>"000110111",
  59015=>"000110000",
  59016=>"000000110",
  59017=>"000000000",
  59018=>"100110000",
  59019=>"000000001",
  59020=>"000001011",
  59021=>"000000000",
  59022=>"000100000",
  59023=>"000010111",
  59024=>"000001011",
  59025=>"011001110",
  59026=>"000000000",
  59027=>"010001101",
  59028=>"000000000",
  59029=>"000000000",
  59030=>"111001001",
  59031=>"000000000",
  59032=>"011111110",
  59033=>"100000000",
  59034=>"111111111",
  59035=>"011011011",
  59036=>"000110000",
  59037=>"000000000",
  59038=>"111111111",
  59039=>"000111011",
  59040=>"100000000",
  59041=>"111111011",
  59042=>"011011000",
  59043=>"000010110",
  59044=>"000000001",
  59045=>"110111111",
  59046=>"111111111",
  59047=>"011011011",
  59048=>"000000010",
  59049=>"000000000",
  59050=>"000000000",
  59051=>"001011111",
  59052=>"100000000",
  59053=>"001001001",
  59054=>"110110010",
  59055=>"000011011",
  59056=>"000011000",
  59057=>"011010010",
  59058=>"000000000",
  59059=>"000000000",
  59060=>"110000000",
  59061=>"000000011",
  59062=>"001011011",
  59063=>"111111010",
  59064=>"001011010",
  59065=>"000000111",
  59066=>"000000000",
  59067=>"101111111",
  59068=>"000000000",
  59069=>"000000010",
  59070=>"000000010",
  59071=>"111111011",
  59072=>"111111111",
  59073=>"100111111",
  59074=>"011111010",
  59075=>"000000000",
  59076=>"001000000",
  59077=>"000010111",
  59078=>"111111111",
  59079=>"000011000",
  59080=>"000000000",
  59081=>"001101001",
  59082=>"000000000",
  59083=>"001001000",
  59084=>"111111111",
  59085=>"100001011",
  59086=>"111000000",
  59087=>"110010010",
  59088=>"001011111",
  59089=>"011011110",
  59090=>"000000000",
  59091=>"000000000",
  59092=>"000111111",
  59093=>"001001000",
  59094=>"111001111",
  59095=>"000010000",
  59096=>"001000100",
  59097=>"010010001",
  59098=>"000000111",
  59099=>"111011011",
  59100=>"000000011",
  59101=>"000011111",
  59102=>"001000000",
  59103=>"111111000",
  59104=>"000000001",
  59105=>"011101000",
  59106=>"110111100",
  59107=>"001111111",
  59108=>"100100111",
  59109=>"111111101",
  59110=>"000100000",
  59111=>"111111111",
  59112=>"111001000",
  59113=>"010111111",
  59114=>"111111111",
  59115=>"000110110",
  59116=>"100111100",
  59117=>"000000100",
  59118=>"110000011",
  59119=>"111111111",
  59120=>"001000000",
  59121=>"111111100",
  59122=>"111111111",
  59123=>"111111011",
  59124=>"111010100",
  59125=>"001000000",
  59126=>"011101101",
  59127=>"000000100",
  59128=>"000000000",
  59129=>"000000000",
  59130=>"000000000",
  59131=>"000000000",
  59132=>"111111000",
  59133=>"000000000",
  59134=>"000000101",
  59135=>"101111011",
  59136=>"000000000",
  59137=>"100100000",
  59138=>"000000000",
  59139=>"100111111",
  59140=>"100000111",
  59141=>"111111111",
  59142=>"011111011",
  59143=>"111111110",
  59144=>"100110111",
  59145=>"000000000",
  59146=>"000000000",
  59147=>"111110011",
  59148=>"111111111",
  59149=>"000000000",
  59150=>"111111111",
  59151=>"110111111",
  59152=>"110111111",
  59153=>"011111111",
  59154=>"000000111",
  59155=>"000000001",
  59156=>"000000010",
  59157=>"100110000",
  59158=>"011011001",
  59159=>"000000000",
  59160=>"111011000",
  59161=>"111111111",
  59162=>"001001000",
  59163=>"000001011",
  59164=>"000000110",
  59165=>"100110111",
  59166=>"000000000",
  59167=>"111111111",
  59168=>"111111000",
  59169=>"110111111",
  59170=>"000000000",
  59171=>"111111111",
  59172=>"011011000",
  59173=>"111111111",
  59174=>"111111111",
  59175=>"111000000",
  59176=>"111111100",
  59177=>"000000000",
  59178=>"111111010",
  59179=>"000000000",
  59180=>"000000000",
  59181=>"111111000",
  59182=>"000111000",
  59183=>"100100000",
  59184=>"100000100",
  59185=>"000000000",
  59186=>"011111001",
  59187=>"001001110",
  59188=>"111111110",
  59189=>"110111110",
  59190=>"111110100",
  59191=>"000000001",
  59192=>"001001000",
  59193=>"000000000",
  59194=>"000000110",
  59195=>"110011011",
  59196=>"101111110",
  59197=>"000111000",
  59198=>"100101101",
  59199=>"000000000",
  59200=>"110000000",
  59201=>"000010000",
  59202=>"011110010",
  59203=>"111111111",
  59204=>"111111110",
  59205=>"110100100",
  59206=>"100100000",
  59207=>"111111110",
  59208=>"111111111",
  59209=>"100000111",
  59210=>"111111110",
  59211=>"111111111",
  59212=>"111011101",
  59213=>"000000111",
  59214=>"000000000",
  59215=>"111011001",
  59216=>"001000000",
  59217=>"110110111",
  59218=>"111111111",
  59219=>"000000000",
  59220=>"111001111",
  59221=>"001001001",
  59222=>"000000000",
  59223=>"010000010",
  59224=>"111111011",
  59225=>"111011000",
  59226=>"100000001",
  59227=>"000000000",
  59228=>"010011011",
  59229=>"111111000",
  59230=>"000000110",
  59231=>"111111111",
  59232=>"001011011",
  59233=>"111100100",
  59234=>"110110010",
  59235=>"001111111",
  59236=>"000000000",
  59237=>"000100100",
  59238=>"111100100",
  59239=>"001101001",
  59240=>"001001001",
  59241=>"010000000",
  59242=>"100101101",
  59243=>"111111111",
  59244=>"000110110",
  59245=>"001000100",
  59246=>"010010000",
  59247=>"000000000",
  59248=>"111111110",
  59249=>"000000000",
  59250=>"011110010",
  59251=>"111111001",
  59252=>"111111111",
  59253=>"111100110",
  59254=>"000110111",
  59255=>"000110000",
  59256=>"101101111",
  59257=>"111001000",
  59258=>"111111111",
  59259=>"000000000",
  59260=>"000010000",
  59261=>"111111001",
  59262=>"011111111",
  59263=>"010000000",
  59264=>"010010010",
  59265=>"101101111",
  59266=>"000000000",
  59267=>"100000000",
  59268=>"110100111",
  59269=>"000000000",
  59270=>"001000000",
  59271=>"001000100",
  59272=>"100100000",
  59273=>"111111111",
  59274=>"111111111",
  59275=>"010010010",
  59276=>"111111111",
  59277=>"000000000",
  59278=>"000010011",
  59279=>"110000000",
  59280=>"000000000",
  59281=>"111111111",
  59282=>"010011000",
  59283=>"000000000",
  59284=>"111000000",
  59285=>"000000000",
  59286=>"000000000",
  59287=>"111100000",
  59288=>"000001111",
  59289=>"000001001",
  59290=>"111111111",
  59291=>"011111001",
  59292=>"000000110",
  59293=>"000000000",
  59294=>"000000000",
  59295=>"100000000",
  59296=>"111111011",
  59297=>"111111001",
  59298=>"000000000",
  59299=>"011000000",
  59300=>"001111111",
  59301=>"000000000",
  59302=>"111111111",
  59303=>"000001111",
  59304=>"100111111",
  59305=>"111111100",
  59306=>"010110111",
  59307=>"011000000",
  59308=>"100000110",
  59309=>"000100100",
  59310=>"000000000",
  59311=>"011000000",
  59312=>"001000000",
  59313=>"001001000",
  59314=>"011011011",
  59315=>"101111111",
  59316=>"000000000",
  59317=>"000000111",
  59318=>"000111111",
  59319=>"000010000",
  59320=>"111111111",
  59321=>"000000001",
  59322=>"110000000",
  59323=>"000011111",
  59324=>"000011111",
  59325=>"111011011",
  59326=>"111111011",
  59327=>"000001000",
  59328=>"000000000",
  59329=>"000000000",
  59330=>"111111111",
  59331=>"000000000",
  59332=>"000000011",
  59333=>"110100000",
  59334=>"111000000",
  59335=>"011011011",
  59336=>"000000000",
  59337=>"111110110",
  59338=>"000001000",
  59339=>"110100000",
  59340=>"000000000",
  59341=>"000000000",
  59342=>"001011110",
  59343=>"100100100",
  59344=>"000000000",
  59345=>"001011011",
  59346=>"000000001",
  59347=>"111111110",
  59348=>"110110000",
  59349=>"110111111",
  59350=>"000000100",
  59351=>"100100001",
  59352=>"111111111",
  59353=>"000100000",
  59354=>"000100111",
  59355=>"111111110",
  59356=>"111000111",
  59357=>"001011000",
  59358=>"000000000",
  59359=>"000000000",
  59360=>"011000000",
  59361=>"011011110",
  59362=>"000101111",
  59363=>"011110000",
  59364=>"000100111",
  59365=>"000000000",
  59366=>"000000000",
  59367=>"100110100",
  59368=>"101010000",
  59369=>"110111111",
  59370=>"011111111",
  59371=>"011011011",
  59372=>"000000000",
  59373=>"111111011",
  59374=>"001001111",
  59375=>"111111101",
  59376=>"000110100",
  59377=>"110111111",
  59378=>"001000000",
  59379=>"000000000",
  59380=>"001111011",
  59381=>"100100001",
  59382=>"001001111",
  59383=>"001001001",
  59384=>"111111011",
  59385=>"001000000",
  59386=>"000000000",
  59387=>"000000000",
  59388=>"000000000",
  59389=>"000101001",
  59390=>"000000011",
  59391=>"111111111",
  59392=>"001001111",
  59393=>"110111111",
  59394=>"010000111",
  59395=>"010010010",
  59396=>"000000000",
  59397=>"001000001",
  59398=>"001000000",
  59399=>"111111111",
  59400=>"000000000",
  59401=>"111110100",
  59402=>"110110110",
  59403=>"000000111",
  59404=>"111000000",
  59405=>"111111111",
  59406=>"000001001",
  59407=>"001001001",
  59408=>"110000110",
  59409=>"111001001",
  59410=>"011001101",
  59411=>"010000000",
  59412=>"000111111",
  59413=>"000000110",
  59414=>"110110110",
  59415=>"011111111",
  59416=>"110110110",
  59417=>"110000010",
  59418=>"111101101",
  59419=>"111000000",
  59420=>"000000000",
  59421=>"000000111",
  59422=>"011011110",
  59423=>"000000111",
  59424=>"111000100",
  59425=>"000111111",
  59426=>"000000000",
  59427=>"000000000",
  59428=>"100000111",
  59429=>"011111111",
  59430=>"111111111",
  59431=>"000000000",
  59432=>"000000011",
  59433=>"111001000",
  59434=>"000000000",
  59435=>"111000000",
  59436=>"001000100",
  59437=>"111001000",
  59438=>"110000000",
  59439=>"000000000",
  59440=>"001101100",
  59441=>"001000000",
  59442=>"000011011",
  59443=>"000000000",
  59444=>"111000000",
  59445=>"111011001",
  59446=>"000000000",
  59447=>"001000000",
  59448=>"000110111",
  59449=>"001001111",
  59450=>"000011010",
  59451=>"000000000",
  59452=>"101001101",
  59453=>"000011111",
  59454=>"011000001",
  59455=>"011111111",
  59456=>"111110000",
  59457=>"110110000",
  59458=>"000000001",
  59459=>"000000000",
  59460=>"100110110",
  59461=>"110110100",
  59462=>"110000000",
  59463=>"100100100",
  59464=>"011111011",
  59465=>"000000000",
  59466=>"000010011",
  59467=>"001001010",
  59468=>"110110110",
  59469=>"110000111",
  59470=>"000000111",
  59471=>"000001001",
  59472=>"111000000",
  59473=>"111110000",
  59474=>"001000000",
  59475=>"011011011",
  59476=>"000100000",
  59477=>"000001111",
  59478=>"000000000",
  59479=>"111111010",
  59480=>"001111111",
  59481=>"111000000",
  59482=>"111111000",
  59483=>"000111111",
  59484=>"000000001",
  59485=>"111000000",
  59486=>"000000111",
  59487=>"000011111",
  59488=>"001000101",
  59489=>"011111110",
  59490=>"000110110",
  59491=>"000000100",
  59492=>"111110000",
  59493=>"111000000",
  59494=>"111111000",
  59495=>"111110111",
  59496=>"001001001",
  59497=>"000000011",
  59498=>"111110100",
  59499=>"000000100",
  59500=>"001000011",
  59501=>"111111111",
  59502=>"111111000",
  59503=>"110000101",
  59504=>"111011011",
  59505=>"000001011",
  59506=>"111111001",
  59507=>"000111111",
  59508=>"000000000",
  59509=>"000001111",
  59510=>"110111110",
  59511=>"001000000",
  59512=>"111101000",
  59513=>"111000000",
  59514=>"111111111",
  59515=>"000000010",
  59516=>"110100110",
  59517=>"000000010",
  59518=>"111111110",
  59519=>"010110010",
  59520=>"000000111",
  59521=>"011011010",
  59522=>"110110111",
  59523=>"100000100",
  59524=>"111100111",
  59525=>"110000000",
  59526=>"000000110",
  59527=>"110011000",
  59528=>"110000110",
  59529=>"111000000",
  59530=>"000001111",
  59531=>"100111111",
  59532=>"111101001",
  59533=>"111111111",
  59534=>"110111011",
  59535=>"100111111",
  59536=>"000000000",
  59537=>"111101101",
  59538=>"100000000",
  59539=>"000000000",
  59540=>"001001001",
  59541=>"111111110",
  59542=>"111000001",
  59543=>"000000110",
  59544=>"111111111",
  59545=>"111001000",
  59546=>"000110000",
  59547=>"111000000",
  59548=>"000000100",
  59549=>"111000110",
  59550=>"011111011",
  59551=>"000000000",
  59552=>"000000000",
  59553=>"111011001",
  59554=>"111011001",
  59555=>"111111100",
  59556=>"011001001",
  59557=>"000000000",
  59558=>"111111101",
  59559=>"011111011",
  59560=>"001000110",
  59561=>"001001001",
  59562=>"111000000",
  59563=>"110111111",
  59564=>"111100000",
  59565=>"000110110",
  59566=>"000100111",
  59567=>"000001111",
  59568=>"111010000",
  59569=>"111010000",
  59570=>"111111111",
  59571=>"111111111",
  59572=>"111110110",
  59573=>"000010110",
  59574=>"000111110",
  59575=>"111111001",
  59576=>"111111111",
  59577=>"001000001",
  59578=>"111000000",
  59579=>"000000011",
  59580=>"110000100",
  59581=>"000001001",
  59582=>"111111111",
  59583=>"010010010",
  59584=>"101001001",
  59585=>"111000000",
  59586=>"111000000",
  59587=>"000000000",
  59588=>"000000000",
  59589=>"111010000",
  59590=>"000000000",
  59591=>"100000000",
  59592=>"111011000",
  59593=>"010010010",
  59594=>"011000000",
  59595=>"111000100",
  59596=>"000101111",
  59597=>"100011011",
  59598=>"100000011",
  59599=>"010000000",
  59600=>"111111011",
  59601=>"100000000",
  59602=>"111000011",
  59603=>"111001000",
  59604=>"100000000",
  59605=>"111000000",
  59606=>"100000000",
  59607=>"111011101",
  59608=>"010111111",
  59609=>"000110111",
  59610=>"011000000",
  59611=>"011000000",
  59612=>"110011000",
  59613=>"010000000",
  59614=>"000000000",
  59615=>"001000001",
  59616=>"001000000",
  59617=>"001001010",
  59618=>"100000100",
  59619=>"011000100",
  59620=>"000111111",
  59621=>"110111110",
  59622=>"000000001",
  59623=>"001000000",
  59624=>"000000000",
  59625=>"111111011",
  59626=>"000000111",
  59627=>"111100000",
  59628=>"111111011",
  59629=>"000000000",
  59630=>"111000000",
  59631=>"001111110",
  59632=>"100000011",
  59633=>"000111111",
  59634=>"111110111",
  59635=>"001000000",
  59636=>"000000000",
  59637=>"001111111",
  59638=>"000000111",
  59639=>"111010010",
  59640=>"000000000",
  59641=>"110001001",
  59642=>"001000000",
  59643=>"000000000",
  59644=>"110110000",
  59645=>"100100111",
  59646=>"010010000",
  59647=>"111000011",
  59648=>"000000000",
  59649=>"111111010",
  59650=>"111111111",
  59651=>"111111111",
  59652=>"000000011",
  59653=>"000000000",
  59654=>"001001111",
  59655=>"000000000",
  59656=>"001001000",
  59657=>"101001001",
  59658=>"111111100",
  59659=>"111111111",
  59660=>"111001001",
  59661=>"010110010",
  59662=>"110110111",
  59663=>"100110110",
  59664=>"001000001",
  59665=>"000000001",
  59666=>"010010000",
  59667=>"101010010",
  59668=>"000000000",
  59669=>"101101111",
  59670=>"110100000",
  59671=>"101000000",
  59672=>"011011001",
  59673=>"000110111",
  59674=>"000000000",
  59675=>"111111110",
  59676=>"100110100",
  59677=>"000000000",
  59678=>"111000001",
  59679=>"111001000",
  59680=>"011111000",
  59681=>"000000000",
  59682=>"000110111",
  59683=>"111111111",
  59684=>"001000000",
  59685=>"010000000",
  59686=>"111100000",
  59687=>"001011000",
  59688=>"010110000",
  59689=>"000111111",
  59690=>"111110110",
  59691=>"100000110",
  59692=>"000000000",
  59693=>"110110000",
  59694=>"011000111",
  59695=>"101001101",
  59696=>"101000000",
  59697=>"000110110",
  59698=>"111111110",
  59699=>"110110110",
  59700=>"110110000",
  59701=>"111111000",
  59702=>"000001001",
  59703=>"111001001",
  59704=>"001000001",
  59705=>"101000000",
  59706=>"010000000",
  59707=>"110000010",
  59708=>"000000000",
  59709=>"100001000",
  59710=>"111001001",
  59711=>"011111111",
  59712=>"111001000",
  59713=>"100100011",
  59714=>"000000001",
  59715=>"000000111",
  59716=>"111111010",
  59717=>"001011111",
  59718=>"000101101",
  59719=>"000000110",
  59720=>"011000000",
  59721=>"001001111",
  59722=>"111111001",
  59723=>"111111001",
  59724=>"000000111",
  59725=>"000001111",
  59726=>"101100000",
  59727=>"111111110",
  59728=>"110001000",
  59729=>"111111111",
  59730=>"111000000",
  59731=>"100000110",
  59732=>"000000000",
  59733=>"001011001",
  59734=>"110000110",
  59735=>"010111111",
  59736=>"000000001",
  59737=>"000010001",
  59738=>"000000001",
  59739=>"001001111",
  59740=>"111110000",
  59741=>"011111111",
  59742=>"011001000",
  59743=>"000000000",
  59744=>"111111111",
  59745=>"110000000",
  59746=>"000111011",
  59747=>"101000000",
  59748=>"000011011",
  59749=>"111101111",
  59750=>"111111111",
  59751=>"111010110",
  59752=>"110000000",
  59753=>"000101111",
  59754=>"111111000",
  59755=>"001000110",
  59756=>"000000000",
  59757=>"110000000",
  59758=>"101001011",
  59759=>"010000000",
  59760=>"011000000",
  59761=>"110000111",
  59762=>"110000000",
  59763=>"100100100",
  59764=>"000000000",
  59765=>"010110111",
  59766=>"111000000",
  59767=>"000011011",
  59768=>"101000000",
  59769=>"111011000",
  59770=>"000000111",
  59771=>"000000000",
  59772=>"000101111",
  59773=>"110110111",
  59774=>"111001000",
  59775=>"101001101",
  59776=>"011001001",
  59777=>"101110110",
  59778=>"000111011",
  59779=>"000000000",
  59780=>"000000000",
  59781=>"011111011",
  59782=>"111111111",
  59783=>"111010100",
  59784=>"001001111",
  59785=>"000101101",
  59786=>"011111111",
  59787=>"000100000",
  59788=>"111110111",
  59789=>"111111111",
  59790=>"000000110",
  59791=>"000010010",
  59792=>"111111101",
  59793=>"111010000",
  59794=>"001000000",
  59795=>"001001011",
  59796=>"111110000",
  59797=>"110010000",
  59798=>"111001001",
  59799=>"111111110",
  59800=>"000010110",
  59801=>"001000110",
  59802=>"111111111",
  59803=>"000101111",
  59804=>"000000000",
  59805=>"110110010",
  59806=>"111001001",
  59807=>"100000000",
  59808=>"111111000",
  59809=>"110111011",
  59810=>"000000111",
  59811=>"111111111",
  59812=>"000011111",
  59813=>"100000000",
  59814=>"111101101",
  59815=>"000010111",
  59816=>"110000000",
  59817=>"110111111",
  59818=>"111110111",
  59819=>"111000001",
  59820=>"111111000",
  59821=>"000000000",
  59822=>"111101000",
  59823=>"011001010",
  59824=>"011000111",
  59825=>"100000000",
  59826=>"111111100",
  59827=>"111101100",
  59828=>"111101001",
  59829=>"000000000",
  59830=>"110000110",
  59831=>"100111101",
  59832=>"000000000",
  59833=>"000110111",
  59834=>"111001000",
  59835=>"111111100",
  59836=>"100110000",
  59837=>"001101101",
  59838=>"101101111",
  59839=>"001000001",
  59840=>"010111011",
  59841=>"111110110",
  59842=>"001001001",
  59843=>"010010000",
  59844=>"100000110",
  59845=>"111011000",
  59846=>"111100001",
  59847=>"111000000",
  59848=>"110100100",
  59849=>"000011011",
  59850=>"001000001",
  59851=>"111100000",
  59852=>"111111100",
  59853=>"000111111",
  59854=>"111110011",
  59855=>"110000011",
  59856=>"111000100",
  59857=>"111111111",
  59858=>"111000000",
  59859=>"110000001",
  59860=>"001001001",
  59861=>"010000111",
  59862=>"011000000",
  59863=>"100000000",
  59864=>"000000001",
  59865=>"000010011",
  59866=>"101100101",
  59867=>"111000000",
  59868=>"010010000",
  59869=>"001001111",
  59870=>"111111010",
  59871=>"000000000",
  59872=>"101001111",
  59873=>"001111111",
  59874=>"000100111",
  59875=>"111011111",
  59876=>"001001111",
  59877=>"111010111",
  59878=>"000111100",
  59879=>"111111111",
  59880=>"001000000",
  59881=>"000000000",
  59882=>"111001000",
  59883=>"010000000",
  59884=>"101000001",
  59885=>"100111111",
  59886=>"111101111",
  59887=>"111101000",
  59888=>"111101100",
  59889=>"000001111",
  59890=>"001111111",
  59891=>"111001000",
  59892=>"000000110",
  59893=>"000101111",
  59894=>"010011111",
  59895=>"111111111",
  59896=>"110010000",
  59897=>"111101000",
  59898=>"011111111",
  59899=>"000110111",
  59900=>"111111000",
  59901=>"000000000",
  59902=>"111011010",
  59903=>"111011111",
  59904=>"000000000",
  59905=>"000011111",
  59906=>"000000000",
  59907=>"000000000",
  59908=>"111101111",
  59909=>"001000100",
  59910=>"000000000",
  59911=>"111001001",
  59912=>"000111101",
  59913=>"000111111",
  59914=>"111011111",
  59915=>"100000000",
  59916=>"000000000",
  59917=>"011010010",
  59918=>"000100111",
  59919=>"000000000",
  59920=>"110111110",
  59921=>"001001001",
  59922=>"000100010",
  59923=>"000000000",
  59924=>"111111111",
  59925=>"100000111",
  59926=>"111111111",
  59927=>"111111001",
  59928=>"000101110",
  59929=>"111111111",
  59930=>"001000000",
  59931=>"011000000",
  59932=>"111111111",
  59933=>"000000000",
  59934=>"000000111",
  59935=>"001111111",
  59936=>"111111111",
  59937=>"001001000",
  59938=>"000000000",
  59939=>"000000000",
  59940=>"001111000",
  59941=>"111111111",
  59942=>"001101101",
  59943=>"000000000",
  59944=>"100000100",
  59945=>"000000001",
  59946=>"000111111",
  59947=>"111111111",
  59948=>"011111111",
  59949=>"111110001",
  59950=>"001001000",
  59951=>"000000100",
  59952=>"000000000",
  59953=>"000000000",
  59954=>"001001001",
  59955=>"000111111",
  59956=>"011111111",
  59957=>"001000110",
  59958=>"111100000",
  59959=>"000000110",
  59960=>"110100000",
  59961=>"111111111",
  59962=>"000000000",
  59963=>"110100111",
  59964=>"000000101",
  59965=>"000000000",
  59966=>"000000000",
  59967=>"100000000",
  59968=>"001000000",
  59969=>"111101111",
  59970=>"111111111",
  59971=>"111111111",
  59972=>"111111000",
  59973=>"111111111",
  59974=>"000000011",
  59975=>"000000000",
  59976=>"011001011",
  59977=>"111101111",
  59978=>"000000000",
  59979=>"111111111",
  59980=>"111000000",
  59981=>"000001000",
  59982=>"000000000",
  59983=>"000000000",
  59984=>"000000001",
  59985=>"000010000",
  59986=>"111111111",
  59987=>"000000000",
  59988=>"010100100",
  59989=>"000000000",
  59990=>"001111111",
  59991=>"101101111",
  59992=>"000000110",
  59993=>"000000000",
  59994=>"101111111",
  59995=>"110100111",
  59996=>"000000111",
  59997=>"000000111",
  59998=>"000111111",
  59999=>"011111111",
  60000=>"111111000",
  60001=>"000000000",
  60002=>"111111111",
  60003=>"010011111",
  60004=>"000000000",
  60005=>"101000111",
  60006=>"111011010",
  60007=>"100001101",
  60008=>"111111000",
  60009=>"111111111",
  60010=>"000000011",
  60011=>"000110000",
  60012=>"100000000",
  60013=>"000000000",
  60014=>"111111110",
  60015=>"001000000",
  60016=>"011001011",
  60017=>"111111111",
  60018=>"011000000",
  60019=>"000001001",
  60020=>"001111111",
  60021=>"000000000",
  60022=>"000000000",
  60023=>"000000000",
  60024=>"001000001",
  60025=>"111111111",
  60026=>"101000000",
  60027=>"101000000",
  60028=>"000000000",
  60029=>"000000001",
  60030=>"001000110",
  60031=>"111111111",
  60032=>"000000000",
  60033=>"111111111",
  60034=>"000000000",
  60035=>"000000000",
  60036=>"000001111",
  60037=>"000000100",
  60038=>"000100100",
  60039=>"111011111",
  60040=>"110010000",
  60041=>"100100110",
  60042=>"000000000",
  60043=>"110110010",
  60044=>"111110111",
  60045=>"111110000",
  60046=>"111001001",
  60047=>"000000000",
  60048=>"000000000",
  60049=>"011111111",
  60050=>"100000000",
  60051=>"111101000",
  60052=>"011010111",
  60053=>"000000000",
  60054=>"000000000",
  60055=>"000000000",
  60056=>"000000000",
  60057=>"000111111",
  60058=>"111111111",
  60059=>"001001000",
  60060=>"001011000",
  60061=>"001001001",
  60062=>"000000000",
  60063=>"101001101",
  60064=>"001001111",
  60065=>"111011001",
  60066=>"111111111",
  60067=>"000100111",
  60068=>"101001000",
  60069=>"111111111",
  60070=>"111111110",
  60071=>"100110000",
  60072=>"001000000",
  60073=>"111111111",
  60074=>"000000000",
  60075=>"000000000",
  60076=>"000001100",
  60077=>"111100111",
  60078=>"111111100",
  60079=>"111111111",
  60080=>"111111010",
  60081=>"111111111",
  60082=>"111111011",
  60083=>"111111001",
  60084=>"110111111",
  60085=>"111111000",
  60086=>"000000000",
  60087=>"100000000",
  60088=>"000000110",
  60089=>"000000011",
  60090=>"111111111",
  60091=>"000001111",
  60092=>"111111111",
  60093=>"000000000",
  60094=>"000000000",
  60095=>"001001111",
  60096=>"000000111",
  60097=>"000001111",
  60098=>"111101111",
  60099=>"111111111",
  60100=>"000000111",
  60101=>"101001111",
  60102=>"001000000",
  60103=>"001111111",
  60104=>"111111111",
  60105=>"000110000",
  60106=>"000000000",
  60107=>"000000000",
  60108=>"111001111",
  60109=>"011111011",
  60110=>"111110111",
  60111=>"111000111",
  60112=>"000011111",
  60113=>"001001111",
  60114=>"111011111",
  60115=>"000000000",
  60116=>"000000000",
  60117=>"000001011",
  60118=>"000000110",
  60119=>"100000000",
  60120=>"101000100",
  60121=>"001011001",
  60122=>"111111111",
  60123=>"111111000",
  60124=>"111111111",
  60125=>"000000000",
  60126=>"111111111",
  60127=>"000000100",
  60128=>"010001111",
  60129=>"111011011",
  60130=>"011111111",
  60131=>"100100110",
  60132=>"000000000",
  60133=>"111111111",
  60134=>"011111111",
  60135=>"000000000",
  60136=>"100111110",
  60137=>"110110111",
  60138=>"000000000",
  60139=>"011011011",
  60140=>"111111110",
  60141=>"111111111",
  60142=>"111111111",
  60143=>"000000000",
  60144=>"111000001",
  60145=>"011010011",
  60146=>"111111100",
  60147=>"000000100",
  60148=>"000000000",
  60149=>"000100110",
  60150=>"100100110",
  60151=>"111111111",
  60152=>"111111001",
  60153=>"001001111",
  60154=>"000000011",
  60155=>"000000000",
  60156=>"001001111",
  60157=>"000000000",
  60158=>"000001100",
  60159=>"000000000",
  60160=>"101111111",
  60161=>"001000100",
  60162=>"000000001",
  60163=>"000000001",
  60164=>"000000100",
  60165=>"000000001",
  60166=>"101100100",
  60167=>"000000000",
  60168=>"000000000",
  60169=>"000000001",
  60170=>"111111111",
  60171=>"010110000",
  60172=>"100101111",
  60173=>"000000000",
  60174=>"000100111",
  60175=>"100000000",
  60176=>"111111000",
  60177=>"110000000",
  60178=>"000000000",
  60179=>"111111001",
  60180=>"100100000",
  60181=>"111111000",
  60182=>"111001111",
  60183=>"000000000",
  60184=>"110110110",
  60185=>"000000000",
  60186=>"000000110",
  60187=>"111111101",
  60188=>"111000110",
  60189=>"110110000",
  60190=>"111111111",
  60191=>"000000000",
  60192=>"110000000",
  60193=>"110111111",
  60194=>"000000110",
  60195=>"110100110",
  60196=>"001011011",
  60197=>"000000000",
  60198=>"000000000",
  60199=>"110100000",
  60200=>"101001111",
  60201=>"000111111",
  60202=>"011110000",
  60203=>"111111111",
  60204=>"000000111",
  60205=>"000000000",
  60206=>"111111111",
  60207=>"101000000",
  60208=>"001001000",
  60209=>"000000000",
  60210=>"111011001",
  60211=>"000000000",
  60212=>"000100111",
  60213=>"000000000",
  60214=>"000001111",
  60215=>"000000100",
  60216=>"000000000",
  60217=>"111100000",
  60218=>"000000000",
  60219=>"101111110",
  60220=>"111111111",
  60221=>"111111110",
  60222=>"010111110",
  60223=>"111110000",
  60224=>"111100000",
  60225=>"001000000",
  60226=>"000000111",
  60227=>"111111111",
  60228=>"111111111",
  60229=>"111111111",
  60230=>"001001000",
  60231=>"000000000",
  60232=>"000000000",
  60233=>"000000111",
  60234=>"111011100",
  60235=>"001001101",
  60236=>"110100110",
  60237=>"111111110",
  60238=>"110111000",
  60239=>"111111111",
  60240=>"000000100",
  60241=>"000100111",
  60242=>"111111111",
  60243=>"000000000",
  60244=>"111101000",
  60245=>"011011000",
  60246=>"110110100",
  60247=>"111111110",
  60248=>"111111100",
  60249=>"111111111",
  60250=>"011010010",
  60251=>"000000000",
  60252=>"111111111",
  60253=>"000000000",
  60254=>"000000000",
  60255=>"000000111",
  60256=>"110110111",
  60257=>"000111111",
  60258=>"101001001",
  60259=>"100000000",
  60260=>"001000000",
  60261=>"010111111",
  60262=>"110110110",
  60263=>"001001111",
  60264=>"000100100",
  60265=>"000000000",
  60266=>"001011011",
  60267=>"011111100",
  60268=>"110111001",
  60269=>"000000000",
  60270=>"000000000",
  60271=>"000011000",
  60272=>"111001000",
  60273=>"111111110",
  60274=>"011000000",
  60275=>"110000000",
  60276=>"000000000",
  60277=>"001111111",
  60278=>"111111111",
  60279=>"000000000",
  60280=>"111111111",
  60281=>"000000111",
  60282=>"000000000",
  60283=>"110111111",
  60284=>"100100000",
  60285=>"111111110",
  60286=>"111111111",
  60287=>"111111111",
  60288=>"011111110",
  60289=>"110111111",
  60290=>"111111111",
  60291=>"000000000",
  60292=>"000000000",
  60293=>"000000000",
  60294=>"111011001",
  60295=>"111011011",
  60296=>"011101111",
  60297=>"000111111",
  60298=>"101001000",
  60299=>"100000000",
  60300=>"000110111",
  60301=>"111101101",
  60302=>"100100100",
  60303=>"000000000",
  60304=>"111111111",
  60305=>"011000111",
  60306=>"111111111",
  60307=>"111111110",
  60308=>"000000000",
  60309=>"000000000",
  60310=>"011011111",
  60311=>"000000000",
  60312=>"000000000",
  60313=>"111111111",
  60314=>"000000000",
  60315=>"000000101",
  60316=>"000000000",
  60317=>"111000000",
  60318=>"000000000",
  60319=>"100000000",
  60320=>"111111111",
  60321=>"111111001",
  60322=>"111110110",
  60323=>"010110000",
  60324=>"000100000",
  60325=>"000011001",
  60326=>"000000000",
  60327=>"000111111",
  60328=>"111111111",
  60329=>"100110100",
  60330=>"111111111",
  60331=>"000000000",
  60332=>"000001001",
  60333=>"011111111",
  60334=>"000000100",
  60335=>"000000000",
  60336=>"000000000",
  60337=>"111111111",
  60338=>"000000000",
  60339=>"111111111",
  60340=>"111111111",
  60341=>"000000000",
  60342=>"111111101",
  60343=>"000000000",
  60344=>"010110000",
  60345=>"010000000",
  60346=>"000000000",
  60347=>"110011001",
  60348=>"000000000",
  60349=>"000000100",
  60350=>"000000000",
  60351=>"001000000",
  60352=>"000010000",
  60353=>"000111011",
  60354=>"111111111",
  60355=>"000011111",
  60356=>"111111101",
  60357=>"000000000",
  60358=>"111111111",
  60359=>"111111110",
  60360=>"000000110",
  60361=>"001001000",
  60362=>"100101101",
  60363=>"000000111",
  60364=>"000000000",
  60365=>"111111111",
  60366=>"000100111",
  60367=>"000110000",
  60368=>"000000000",
  60369=>"000101010",
  60370=>"000011111",
  60371=>"011001001",
  60372=>"001111110",
  60373=>"000000000",
  60374=>"001011011",
  60375=>"000000000",
  60376=>"000000001",
  60377=>"000000000",
  60378=>"000010000",
  60379=>"100010111",
  60380=>"000000001",
  60381=>"111111111",
  60382=>"001001111",
  60383=>"111111111",
  60384=>"111000000",
  60385=>"000000111",
  60386=>"111111111",
  60387=>"000000000",
  60388=>"111011010",
  60389=>"001000000",
  60390=>"000000000",
  60391=>"000000000",
  60392=>"101101111",
  60393=>"001111111",
  60394=>"000001011",
  60395=>"111111111",
  60396=>"111010000",
  60397=>"000000000",
  60398=>"111111111",
  60399=>"110111111",
  60400=>"111111010",
  60401=>"101111111",
  60402=>"111011001",
  60403=>"001001011",
  60404=>"000000000",
  60405=>"001000000",
  60406=>"001111001",
  60407=>"111111111",
  60408=>"001000101",
  60409=>"000000100",
  60410=>"000000011",
  60411=>"000000000",
  60412=>"000000000",
  60413=>"000000000",
  60414=>"011111111",
  60415=>"111100111",
  60416=>"001111111",
  60417=>"000000000",
  60418=>"001111111",
  60419=>"000100000",
  60420=>"101111111",
  60421=>"000000000",
  60422=>"111111111",
  60423=>"000001111",
  60424=>"110100111",
  60425=>"010010010",
  60426=>"000000000",
  60427=>"001000000",
  60428=>"000110110",
  60429=>"000010000",
  60430=>"000100000",
  60431=>"100111001",
  60432=>"111011000",
  60433=>"000000000",
  60434=>"000000010",
  60435=>"000000000",
  60436=>"111111111",
  60437=>"100100100",
  60438=>"111100110",
  60439=>"000000000",
  60440=>"111100000",
  60441=>"111111011",
  60442=>"111001001",
  60443=>"100100000",
  60444=>"111001110",
  60445=>"010011000",
  60446=>"100100000",
  60447=>"110000000",
  60448=>"110110111",
  60449=>"100100000",
  60450=>"000000000",
  60451=>"111111111",
  60452=>"111111111",
  60453=>"111011011",
  60454=>"110111111",
  60455=>"111111001",
  60456=>"110111111",
  60457=>"000000000",
  60458=>"101101111",
  60459=>"000000000",
  60460=>"111111111",
  60461=>"000011111",
  60462=>"100000000",
  60463=>"111111111",
  60464=>"101101001",
  60465=>"111111111",
  60466=>"000000001",
  60467=>"000000000",
  60468=>"010010010",
  60469=>"000000000",
  60470=>"000111111",
  60471=>"000110110",
  60472=>"111101101",
  60473=>"000001000",
  60474=>"001100100",
  60475=>"001001111",
  60476=>"111111111",
  60477=>"011000011",
  60478=>"000001101",
  60479=>"000000101",
  60480=>"000100100",
  60481=>"011111111",
  60482=>"111110010",
  60483=>"111011111",
  60484=>"001000000",
  60485=>"100100000",
  60486=>"000000110",
  60487=>"001000000",
  60488=>"001011011",
  60489=>"000000000",
  60490=>"001000000",
  60491=>"110111000",
  60492=>"111111111",
  60493=>"011101000",
  60494=>"000000000",
  60495=>"111111111",
  60496=>"111110000",
  60497=>"000001000",
  60498=>"000000000",
  60499=>"111110110",
  60500=>"000000011",
  60501=>"111111111",
  60502=>"000100111",
  60503=>"000000000",
  60504=>"111111011",
  60505=>"000000101",
  60506=>"111111111",
  60507=>"100011111",
  60508=>"111111101",
  60509=>"001001111",
  60510=>"001100000",
  60511=>"101111000",
  60512=>"111111111",
  60513=>"000010010",
  60514=>"000000000",
  60515=>"110110111",
  60516=>"100100000",
  60517=>"000000000",
  60518=>"111111011",
  60519=>"111111000",
  60520=>"000000000",
  60521=>"000000000",
  60522=>"111011111",
  60523=>"111110110",
  60524=>"010000000",
  60525=>"000100000",
  60526=>"001011111",
  60527=>"000000000",
  60528=>"010110111",
  60529=>"000010000",
  60530=>"100110100",
  60531=>"011001001",
  60532=>"000000000",
  60533=>"000000010",
  60534=>"111110010",
  60535=>"111100100",
  60536=>"000000011",
  60537=>"111000011",
  60538=>"000000001",
  60539=>"111111111",
  60540=>"000100100",
  60541=>"000000000",
  60542=>"000010111",
  60543=>"100100000",
  60544=>"111111111",
  60545=>"000011111",
  60546=>"111111110",
  60547=>"111111011",
  60548=>"111111100",
  60549=>"100110111",
  60550=>"111011001",
  60551=>"000111100",
  60552=>"110111111",
  60553=>"111111111",
  60554=>"111101111",
  60555=>"111011010",
  60556=>"111111111",
  60557=>"001001111",
  60558=>"111001000",
  60559=>"111111111",
  60560=>"001111111",
  60561=>"111111111",
  60562=>"010010110",
  60563=>"111100100",
  60564=>"111111000",
  60565=>"000000010",
  60566=>"001000000",
  60567=>"000000000",
  60568=>"001001001",
  60569=>"000000111",
  60570=>"000000000",
  60571=>"000000000",
  60572=>"000000000",
  60573=>"000000010",
  60574=>"111111111",
  60575=>"110110111",
  60576=>"110110110",
  60577=>"101001000",
  60578=>"111111111",
  60579=>"001000000",
  60580=>"011001010",
  60581=>"111000011",
  60582=>"000000111",
  60583=>"111011011",
  60584=>"101100000",
  60585=>"000000001",
  60586=>"000000000",
  60587=>"000000000",
  60588=>"111111110",
  60589=>"110110000",
  60590=>"000100111",
  60591=>"000000000",
  60592=>"000000110",
  60593=>"001111100",
  60594=>"111111110",
  60595=>"000001010",
  60596=>"111110011",
  60597=>"000001111",
  60598=>"110111111",
  60599=>"000000000",
  60600=>"111111011",
  60601=>"110010000",
  60602=>"111000000",
  60603=>"001001011",
  60604=>"101001111",
  60605=>"000000111",
  60606=>"000110111",
  60607=>"011000100",
  60608=>"000000100",
  60609=>"000001001",
  60610=>"000000000",
  60611=>"111111111",
  60612=>"111111111",
  60613=>"000111111",
  60614=>"000000110",
  60615=>"111111111",
  60616=>"000010001",
  60617=>"101101111",
  60618=>"000000000",
  60619=>"111001000",
  60620=>"000101101",
  60621=>"101101000",
  60622=>"000000000",
  60623=>"000000100",
  60624=>"000000000",
  60625=>"000000000",
  60626=>"000000000",
  60627=>"000000000",
  60628=>"110111111",
  60629=>"001000111",
  60630=>"000111111",
  60631=>"000000000",
  60632=>"111111100",
  60633=>"100111111",
  60634=>"000110111",
  60635=>"000111111",
  60636=>"100010000",
  60637=>"111111111",
  60638=>"111111111",
  60639=>"011000000",
  60640=>"111111111",
  60641=>"000000110",
  60642=>"000000000",
  60643=>"111110110",
  60644=>"111111111",
  60645=>"111111111",
  60646=>"010010000",
  60647=>"000001111",
  60648=>"000000000",
  60649=>"111011011",
  60650=>"000000000",
  60651=>"111001101",
  60652=>"101111111",
  60653=>"100011001",
  60654=>"111001000",
  60655=>"000000000",
  60656=>"010000000",
  60657=>"001111111",
  60658=>"011000000",
  60659=>"001000000",
  60660=>"000000000",
  60661=>"111011110",
  60662=>"001001001",
  60663=>"000000000",
  60664=>"111111111",
  60665=>"111110100",
  60666=>"001000000",
  60667=>"000100110",
  60668=>"000111111",
  60669=>"001000000",
  60670=>"101001000",
  60671=>"000110110",
  60672=>"001000001",
  60673=>"111101101",
  60674=>"111111111",
  60675=>"000000000",
  60676=>"111111111",
  60677=>"000000000",
  60678=>"111111010",
  60679=>"111111011",
  60680=>"111111100",
  60681=>"111111111",
  60682=>"111111101",
  60683=>"111111111",
  60684=>"000000000",
  60685=>"000111011",
  60686=>"000000001",
  60687=>"011000000",
  60688=>"000000000",
  60689=>"000000000",
  60690=>"000000000",
  60691=>"000000000",
  60692=>"110111100",
  60693=>"001000000",
  60694=>"110111110",
  60695=>"001111111",
  60696=>"101000000",
  60697=>"000111111",
  60698=>"011011001",
  60699=>"111000011",
  60700=>"000101101",
  60701=>"000000000",
  60702=>"000000000",
  60703=>"000101100",
  60704=>"000000000",
  60705=>"101101111",
  60706=>"000000000",
  60707=>"011100110",
  60708=>"000000000",
  60709=>"000000101",
  60710=>"111111111",
  60711=>"011000000",
  60712=>"101100100",
  60713=>"101100000",
  60714=>"000000100",
  60715=>"000100100",
  60716=>"001001001",
  60717=>"100100110",
  60718=>"111111000",
  60719=>"111111111",
  60720=>"001001000",
  60721=>"000011011",
  60722=>"111110111",
  60723=>"000000111",
  60724=>"111111000",
  60725=>"000000001",
  60726=>"010010000",
  60727=>"111011000",
  60728=>"111010000",
  60729=>"111111110",
  60730=>"111000000",
  60731=>"000000000",
  60732=>"100100110",
  60733=>"111111001",
  60734=>"101101101",
  60735=>"000000111",
  60736=>"111111100",
  60737=>"100001101",
  60738=>"000000001",
  60739=>"000000001",
  60740=>"101111000",
  60741=>"100110000",
  60742=>"111111011",
  60743=>"000000000",
  60744=>"000000000",
  60745=>"000000000",
  60746=>"111111111",
  60747=>"000100100",
  60748=>"000000000",
  60749=>"001001110",
  60750=>"111001001",
  60751=>"001001000",
  60752=>"001100111",
  60753=>"111110111",
  60754=>"111111110",
  60755=>"111101101",
  60756=>"000001000",
  60757=>"001011011",
  60758=>"011111010",
  60759=>"100111111",
  60760=>"000000000",
  60761=>"111111110",
  60762=>"001100110",
  60763=>"000000010",
  60764=>"010111111",
  60765=>"000000100",
  60766=>"000000011",
  60767=>"011000110",
  60768=>"111111110",
  60769=>"100101100",
  60770=>"001001001",
  60771=>"111111111",
  60772=>"000000000",
  60773=>"000000000",
  60774=>"000011000",
  60775=>"111111111",
  60776=>"100100100",
  60777=>"000111000",
  60778=>"101111111",
  60779=>"111111101",
  60780=>"100000100",
  60781=>"111111111",
  60782=>"000010000",
  60783=>"111100111",
  60784=>"111000000",
  60785=>"111000000",
  60786=>"000111111",
  60787=>"100100100",
  60788=>"000000000",
  60789=>"000000000",
  60790=>"000100110",
  60791=>"111111100",
  60792=>"111000001",
  60793=>"111110111",
  60794=>"111111111",
  60795=>"111100111",
  60796=>"111111000",
  60797=>"011110111",
  60798=>"111011011",
  60799=>"101100100",
  60800=>"000100100",
  60801=>"101101111",
  60802=>"001001000",
  60803=>"110101111",
  60804=>"000000011",
  60805=>"011111010",
  60806=>"010011111",
  60807=>"011100000",
  60808=>"111011111",
  60809=>"111111001",
  60810=>"111000010",
  60811=>"000000000",
  60812=>"110110111",
  60813=>"110110110",
  60814=>"000000101",
  60815=>"000000000",
  60816=>"110000000",
  60817=>"001101001",
  60818=>"010011011",
  60819=>"001000011",
  60820=>"001001011",
  60821=>"000010010",
  60822=>"000000000",
  60823=>"001011001",
  60824=>"111101000",
  60825=>"111100000",
  60826=>"111111001",
  60827=>"000001000",
  60828=>"001010000",
  60829=>"111111111",
  60830=>"001001000",
  60831=>"111111111",
  60832=>"000000000",
  60833=>"001000000",
  60834=>"000000010",
  60835=>"000000111",
  60836=>"000000001",
  60837=>"111011000",
  60838=>"111111111",
  60839=>"000000000",
  60840=>"111111111",
  60841=>"000000000",
  60842=>"000000000",
  60843=>"000110111",
  60844=>"000000000",
  60845=>"000001001",
  60846=>"111000100",
  60847=>"000100100",
  60848=>"110000100",
  60849=>"001001001",
  60850=>"111111111",
  60851=>"000000000",
  60852=>"100111001",
  60853=>"000000000",
  60854=>"111111101",
  60855=>"111111010",
  60856=>"111111111",
  60857=>"101000000",
  60858=>"000111101",
  60859=>"011111111",
  60860=>"000000001",
  60861=>"111111111",
  60862=>"000000000",
  60863=>"001001111",
  60864=>"000000001",
  60865=>"111111111",
  60866=>"011000000",
  60867=>"111111000",
  60868=>"111111110",
  60869=>"001001001",
  60870=>"000010000",
  60871=>"000110111",
  60872=>"000000000",
  60873=>"000100110",
  60874=>"001000000",
  60875=>"000000000",
  60876=>"111000000",
  60877=>"111111111",
  60878=>"111111000",
  60879=>"000000111",
  60880=>"101110111",
  60881=>"000000000",
  60882=>"000000100",
  60883=>"000010011",
  60884=>"000001011",
  60885=>"111111111",
  60886=>"000000000",
  60887=>"000000100",
  60888=>"110100101",
  60889=>"000111111",
  60890=>"001100000",
  60891=>"111110000",
  60892=>"101001110",
  60893=>"000000010",
  60894=>"111111111",
  60895=>"111001001",
  60896=>"110101111",
  60897=>"110100000",
  60898=>"010000000",
  60899=>"000011011",
  60900=>"101111100",
  60901=>"011010000",
  60902=>"101111111",
  60903=>"111000000",
  60904=>"011001000",
  60905=>"010010000",
  60906=>"000100000",
  60907=>"101100001",
  60908=>"010111111",
  60909=>"001000000",
  60910=>"111111111",
  60911=>"111000000",
  60912=>"111110010",
  60913=>"000000000",
  60914=>"111111001",
  60915=>"100110110",
  60916=>"000000001",
  60917=>"110110111",
  60918=>"000001110",
  60919=>"000101101",
  60920=>"100111111",
  60921=>"111011011",
  60922=>"000000000",
  60923=>"111000000",
  60924=>"000000000",
  60925=>"000000101",
  60926=>"000000000",
  60927=>"110110111",
  60928=>"001000000",
  60929=>"111111111",
  60930=>"000000001",
  60931=>"111000000",
  60932=>"001000111",
  60933=>"000000000",
  60934=>"000000000",
  60935=>"111000000",
  60936=>"111111111",
  60937=>"111111100",
  60938=>"000000000",
  60939=>"000001001",
  60940=>"001001001",
  60941=>"111101100",
  60942=>"000100111",
  60943=>"000000000",
  60944=>"110000000",
  60945=>"000000000",
  60946=>"001000000",
  60947=>"000000000",
  60948=>"111111111",
  60949=>"110110111",
  60950=>"101100000",
  60951=>"010010000",
  60952=>"111010000",
  60953=>"000000000",
  60954=>"001000111",
  60955=>"111110110",
  60956=>"000000110",
  60957=>"000111111",
  60958=>"010011011",
  60959=>"011011111",
  60960=>"100111111",
  60961=>"110110110",
  60962=>"000000100",
  60963=>"000000001",
  60964=>"000000000",
  60965=>"100110000",
  60966=>"000000000",
  60967=>"001000100",
  60968=>"110101100",
  60969=>"110111110",
  60970=>"001011011",
  60971=>"000000000",
  60972=>"111111101",
  60973=>"000000000",
  60974=>"111111111",
  60975=>"111000000",
  60976=>"101111100",
  60977=>"100111111",
  60978=>"110110000",
  60979=>"110000100",
  60980=>"000001000",
  60981=>"000110111",
  60982=>"000000000",
  60983=>"000110111",
  60984=>"111111111",
  60985=>"111111000",
  60986=>"111111111",
  60987=>"000010011",
  60988=>"111111111",
  60989=>"000011111",
  60990=>"110111111",
  60991=>"000000000",
  60992=>"111000011",
  60993=>"111000000",
  60994=>"111111111",
  60995=>"001000000",
  60996=>"000011111",
  60997=>"011111110",
  60998=>"111110110",
  60999=>"111111111",
  61000=>"111111111",
  61001=>"111111111",
  61002=>"111101100",
  61003=>"000000111",
  61004=>"111111111",
  61005=>"100000000",
  61006=>"011011111",
  61007=>"000111111",
  61008=>"111111111",
  61009=>"001000111",
  61010=>"100000000",
  61011=>"000001001",
  61012=>"000000000",
  61013=>"101001111",
  61014=>"001111111",
  61015=>"100001011",
  61016=>"000111111",
  61017=>"000000000",
  61018=>"111111000",
  61019=>"111111111",
  61020=>"000000001",
  61021=>"111111111",
  61022=>"111111111",
  61023=>"111111110",
  61024=>"111111111",
  61025=>"000000000",
  61026=>"111000000",
  61027=>"101000000",
  61028=>"010110111",
  61029=>"000000110",
  61030=>"000000000",
  61031=>"000000000",
  61032=>"111111100",
  61033=>"000000000",
  61034=>"111111111",
  61035=>"000000000",
  61036=>"011010110",
  61037=>"111111111",
  61038=>"000000000",
  61039=>"001001000",
  61040=>"001000000",
  61041=>"111111111",
  61042=>"000100100",
  61043=>"001000000",
  61044=>"111111111",
  61045=>"000000000",
  61046=>"011111011",
  61047=>"100111111",
  61048=>"000000111",
  61049=>"000000000",
  61050=>"000000000",
  61051=>"000000111",
  61052=>"000100110",
  61053=>"111110001",
  61054=>"000000000",
  61055=>"000000000",
  61056=>"111101110",
  61057=>"000000000",
  61058=>"111011111",
  61059=>"000000111",
  61060=>"000000111",
  61061=>"110000111",
  61062=>"000000110",
  61063=>"000100100",
  61064=>"111001111",
  61065=>"100000000",
  61066=>"000000000",
  61067=>"111111111",
  61068=>"111111111",
  61069=>"111111111",
  61070=>"111111011",
  61071=>"100111101",
  61072=>"000000000",
  61073=>"000000110",
  61074=>"101000000",
  61075=>"111110111",
  61076=>"111100101",
  61077=>"000000000",
  61078=>"000000000",
  61079=>"011011111",
  61080=>"000001001",
  61081=>"000000111",
  61082=>"000000000",
  61083=>"000000000",
  61084=>"011011111",
  61085=>"111101100",
  61086=>"001111111",
  61087=>"111111111",
  61088=>"111111000",
  61089=>"111111111",
  61090=>"000110111",
  61091=>"101001011",
  61092=>"000000100",
  61093=>"111111011",
  61094=>"111111111",
  61095=>"101111111",
  61096=>"001111111",
  61097=>"000100101",
  61098=>"000000000",
  61099=>"101100100",
  61100=>"000000000",
  61101=>"000001001",
  61102=>"000000111",
  61103=>"000000100",
  61104=>"111111000",
  61105=>"111111111",
  61106=>"100111111",
  61107=>"111011000",
  61108=>"111100000",
  61109=>"000000000",
  61110=>"111111110",
  61111=>"111111100",
  61112=>"111111001",
  61113=>"000000000",
  61114=>"000000100",
  61115=>"111111111",
  61116=>"000110111",
  61117=>"000000100",
  61118=>"000000000",
  61119=>"000000111",
  61120=>"111111111",
  61121=>"001001000",
  61122=>"000000000",
  61123=>"111111111",
  61124=>"000000000",
  61125=>"000000000",
  61126=>"010110111",
  61127=>"111111111",
  61128=>"110000000",
  61129=>"111111110",
  61130=>"101110110",
  61131=>"111111111",
  61132=>"000001111",
  61133=>"000000000",
  61134=>"000000101",
  61135=>"000100110",
  61136=>"100111010",
  61137=>"111000000",
  61138=>"000000000",
  61139=>"111000000",
  61140=>"000100111",
  61141=>"100110111",
  61142=>"111000000",
  61143=>"000000000",
  61144=>"110110111",
  61145=>"100100100",
  61146=>"000000000",
  61147=>"100111111",
  61148=>"111111111",
  61149=>"111111111",
  61150=>"011000000",
  61151=>"000011111",
  61152=>"111110000",
  61153=>"110111111",
  61154=>"111111111",
  61155=>"111011111",
  61156=>"000000001",
  61157=>"111111111",
  61158=>"111111111",
  61159=>"111111111",
  61160=>"111000000",
  61161=>"100000000",
  61162=>"000000100",
  61163=>"110000010",
  61164=>"111111000",
  61165=>"101000000",
  61166=>"000100100",
  61167=>"100111111",
  61168=>"111111110",
  61169=>"000000000",
  61170=>"000000000",
  61171=>"000000111",
  61172=>"010000000",
  61173=>"100110111",
  61174=>"000000000",
  61175=>"100110111",
  61176=>"111001000",
  61177=>"001001011",
  61178=>"001000100",
  61179=>"111111110",
  61180=>"110111111",
  61181=>"111110110",
  61182=>"111111111",
  61183=>"111101101",
  61184=>"000001111",
  61185=>"001000000",
  61186=>"000100000",
  61187=>"000000000",
  61188=>"111111001",
  61189=>"000101111",
  61190=>"000000100",
  61191=>"111111111",
  61192=>"100001001",
  61193=>"000000000",
  61194=>"111111111",
  61195=>"111111111",
  61196=>"000111111",
  61197=>"000011111",
  61198=>"000000000",
  61199=>"111000011",
  61200=>"110010000",
  61201=>"100110100",
  61202=>"100000100",
  61203=>"000001001",
  61204=>"111111111",
  61205=>"100000000",
  61206=>"111101111",
  61207=>"000000001",
  61208=>"101101111",
  61209=>"101001100",
  61210=>"000000000",
  61211=>"111111111",
  61212=>"111111111",
  61213=>"000000111",
  61214=>"000000001",
  61215=>"111111111",
  61216=>"011011000",
  61217=>"111111111",
  61218=>"000000000",
  61219=>"111101100",
  61220=>"100000000",
  61221=>"000000000",
  61222=>"100100100",
  61223=>"111111011",
  61224=>"111111111",
  61225=>"000000100",
  61226=>"000000000",
  61227=>"000010010",
  61228=>"100111111",
  61229=>"000000100",
  61230=>"000010000",
  61231=>"110000000",
  61232=>"001001011",
  61233=>"000010000",
  61234=>"111111111",
  61235=>"000000000",
  61236=>"000000000",
  61237=>"000000111",
  61238=>"001111011",
  61239=>"000000000",
  61240=>"000000000",
  61241=>"111111011",
  61242=>"100000111",
  61243=>"110000111",
  61244=>"010110110",
  61245=>"001100110",
  61246=>"000010000",
  61247=>"100111111",
  61248=>"111111000",
  61249=>"111111111",
  61250=>"000000110",
  61251=>"111111111",
  61252=>"100110110",
  61253=>"001000100",
  61254=>"101101000",
  61255=>"001001101",
  61256=>"110100000",
  61257=>"000110111",
  61258=>"011001001",
  61259=>"111111111",
  61260=>"111011000",
  61261=>"001110000",
  61262=>"101001001",
  61263=>"111001000",
  61264=>"111111111",
  61265=>"000000000",
  61266=>"111111111",
  61267=>"000000000",
  61268=>"000000000",
  61269=>"001001001",
  61270=>"000000111",
  61271=>"111111111",
  61272=>"011111011",
  61273=>"000111111",
  61274=>"000000000",
  61275=>"000001100",
  61276=>"001001001",
  61277=>"111111111",
  61278=>"000000111",
  61279=>"111111111",
  61280=>"001000000",
  61281=>"000000000",
  61282=>"011111111",
  61283=>"000000000",
  61284=>"111111111",
  61285=>"111111111",
  61286=>"000000000",
  61287=>"100100111",
  61288=>"111111111",
  61289=>"110000000",
  61290=>"000111111",
  61291=>"111111111",
  61292=>"011001011",
  61293=>"000000001",
  61294=>"111111111",
  61295=>"111111111",
  61296=>"111111111",
  61297=>"000001001",
  61298=>"000000000",
  61299=>"110110110",
  61300=>"000000000",
  61301=>"100001001",
  61302=>"100001000",
  61303=>"111110110",
  61304=>"001000000",
  61305=>"111111010",
  61306=>"111111111",
  61307=>"000110111",
  61308=>"000000110",
  61309=>"111000111",
  61310=>"000000000",
  61311=>"111000000",
  61312=>"111011111",
  61313=>"000010100",
  61314=>"110110110",
  61315=>"000111111",
  61316=>"000100101",
  61317=>"000000100",
  61318=>"000000111",
  61319=>"111111111",
  61320=>"111111110",
  61321=>"000000000",
  61322=>"101100000",
  61323=>"010111111",
  61324=>"111111111",
  61325=>"000000000",
  61326=>"101001001",
  61327=>"110100000",
  61328=>"001101111",
  61329=>"111011000",
  61330=>"001000111",
  61331=>"001001111",
  61332=>"000000000",
  61333=>"000010000",
  61334=>"011010111",
  61335=>"000000111",
  61336=>"011000011",
  61337=>"100100100",
  61338=>"100100100",
  61339=>"000000000",
  61340=>"000000000",
  61341=>"011110110",
  61342=>"000000000",
  61343=>"111111000",
  61344=>"111110111",
  61345=>"011110000",
  61346=>"101111110",
  61347=>"001000000",
  61348=>"101101111",
  61349=>"000000000",
  61350=>"111111110",
  61351=>"111111111",
  61352=>"100000000",
  61353=>"110111111",
  61354=>"000000000",
  61355=>"000100100",
  61356=>"000000000",
  61357=>"000011001",
  61358=>"000000000",
  61359=>"000000000",
  61360=>"000000000",
  61361=>"000000000",
  61362=>"111111111",
  61363=>"000000000",
  61364=>"000000000",
  61365=>"000000000",
  61366=>"111111111",
  61367=>"110000000",
  61368=>"000000010",
  61369=>"001000000",
  61370=>"111000000",
  61371=>"101100000",
  61372=>"111111111",
  61373=>"000000000",
  61374=>"001000001",
  61375=>"111101100",
  61376=>"111111111",
  61377=>"000000000",
  61378=>"000000000",
  61379=>"111111111",
  61380=>"000110111",
  61381=>"111000110",
  61382=>"011001000",
  61383=>"011011011",
  61384=>"101101100",
  61385=>"111111111",
  61386=>"111000000",
  61387=>"001001000",
  61388=>"111111111",
  61389=>"011001000",
  61390=>"001000000",
  61391=>"111111111",
  61392=>"101001111",
  61393=>"101000000",
  61394=>"111011111",
  61395=>"000000000",
  61396=>"001000010",
  61397=>"100111111",
  61398=>"100000000",
  61399=>"100000000",
  61400=>"111001000",
  61401=>"101101111",
  61402=>"111000000",
  61403=>"011011000",
  61404=>"111111111",
  61405=>"000100100",
  61406=>"110111111",
  61407=>"011110110",
  61408=>"111111100",
  61409=>"111001000",
  61410=>"000000100",
  61411=>"111111100",
  61412=>"000110111",
  61413=>"010000000",
  61414=>"000111100",
  61415=>"000000000",
  61416=>"000000000",
  61417=>"111100111",
  61418=>"000000010",
  61419=>"000100000",
  61420=>"000110111",
  61421=>"000100111",
  61422=>"000000000",
  61423=>"000110111",
  61424=>"000000000",
  61425=>"000001001",
  61426=>"111001001",
  61427=>"001011111",
  61428=>"101111000",
  61429=>"001001100",
  61430=>"000000000",
  61431=>"110011000",
  61432=>"000000000",
  61433=>"001001011",
  61434=>"110110110",
  61435=>"111000000",
  61436=>"001111111",
  61437=>"111111011",
  61438=>"111111111",
  61439=>"000000110",
  61440=>"111111111",
  61441=>"000000000",
  61442=>"111101000",
  61443=>"000000111",
  61444=>"101000010",
  61445=>"111001000",
  61446=>"000000100",
  61447=>"000101111",
  61448=>"111000000",
  61449=>"000111000",
  61450=>"111111000",
  61451=>"110111111",
  61452=>"110110110",
  61453=>"000000111",
  61454=>"100100110",
  61455=>"000110111",
  61456=>"000000000",
  61457=>"000000000",
  61458=>"111000111",
  61459=>"000111100",
  61460=>"000000111",
  61461=>"111000000",
  61462=>"111010101",
  61463=>"000011111",
  61464=>"111111111",
  61465=>"000100101",
  61466=>"011011011",
  61467=>"100111111",
  61468=>"111100100",
  61469=>"100000000",
  61470=>"100000101",
  61471=>"000101111",
  61472=>"000010111",
  61473=>"100110111",
  61474=>"111111000",
  61475=>"110111000",
  61476=>"000000111",
  61477=>"100111111",
  61478=>"100100000",
  61479=>"000000111",
  61480=>"100111111",
  61481=>"111111000",
  61482=>"111111111",
  61483=>"111000000",
  61484=>"100000000",
  61485=>"111111000",
  61486=>"000000000",
  61487=>"000001011",
  61488=>"000000000",
  61489=>"110111111",
  61490=>"011011001",
  61491=>"111011000",
  61492=>"000111111",
  61493=>"011111111",
  61494=>"111111110",
  61495=>"000110111",
  61496=>"110100000",
  61497=>"111111000",
  61498=>"111111111",
  61499=>"111001011",
  61500=>"111111001",
  61501=>"111111011",
  61502=>"000011111",
  61503=>"000000100",
  61504=>"111000000",
  61505=>"010011011",
  61506=>"100010000",
  61507=>"101000000",
  61508=>"001111111",
  61509=>"000000000",
  61510=>"000000000",
  61511=>"000000000",
  61512=>"000000111",
  61513=>"111111111",
  61514=>"111111111",
  61515=>"000000000",
  61516=>"001001000",
  61517=>"110111000",
  61518=>"000001111",
  61519=>"101000001",
  61520=>"101000000",
  61521=>"011011000",
  61522=>"111001001",
  61523=>"101111111",
  61524=>"000000001",
  61525=>"000110100",
  61526=>"000000101",
  61527=>"000000111",
  61528=>"001001000",
  61529=>"111101101",
  61530=>"011000000",
  61531=>"111000000",
  61532=>"000000000",
  61533=>"000111111",
  61534=>"111000000",
  61535=>"000011011",
  61536=>"000000000",
  61537=>"000111111",
  61538=>"000000000",
  61539=>"111111000",
  61540=>"111110000",
  61541=>"011000100",
  61542=>"000000000",
  61543=>"111111111",
  61544=>"111011000",
  61545=>"111100111",
  61546=>"111011111",
  61547=>"000010111",
  61548=>"001011000",
  61549=>"111001011",
  61550=>"111100000",
  61551=>"000000000",
  61552=>"111000000",
  61553=>"101111111",
  61554=>"111111111",
  61555=>"101101001",
  61556=>"111111111",
  61557=>"111111110",
  61558=>"111111000",
  61559=>"011111100",
  61560=>"000000001",
  61561=>"000000111",
  61562=>"111111000",
  61563=>"111111111",
  61564=>"100110000",
  61565=>"000000110",
  61566=>"000000111",
  61567=>"000000000",
  61568=>"000100111",
  61569=>"101001000",
  61570=>"000000000",
  61571=>"011111111",
  61572=>"111001011",
  61573=>"100000000",
  61574=>"111111111",
  61575=>"001000000",
  61576=>"000101111",
  61577=>"010010000",
  61578=>"000000000",
  61579=>"000001111",
  61580=>"011000110",
  61581=>"011111000",
  61582=>"001000101",
  61583=>"111000000",
  61584=>"001000100",
  61585=>"000000100",
  61586=>"010010000",
  61587=>"000111111",
  61588=>"111110001",
  61589=>"000000010",
  61590=>"111000000",
  61591=>"111000001",
  61592=>"000000000",
  61593=>"111111000",
  61594=>"111111000",
  61595=>"001000000",
  61596=>"000110111",
  61597=>"111111111",
  61598=>"100000000",
  61599=>"110100000",
  61600=>"000001110",
  61601=>"111011011",
  61602=>"111100111",
  61603=>"000000000",
  61604=>"111111111",
  61605=>"100110110",
  61606=>"111111111",
  61607=>"100111111",
  61608=>"000101001",
  61609=>"000000000",
  61610=>"000001111",
  61611=>"111111111",
  61612=>"111111000",
  61613=>"100000000",
  61614=>"101000000",
  61615=>"000000000",
  61616=>"111001000",
  61617=>"100111111",
  61618=>"101111010",
  61619=>"100000011",
  61620=>"000000000",
  61621=>"000011010",
  61622=>"000000000",
  61623=>"000000111",
  61624=>"001101111",
  61625=>"111111000",
  61626=>"100000100",
  61627=>"110110010",
  61628=>"111100111",
  61629=>"000000111",
  61630=>"100111100",
  61631=>"000100111",
  61632=>"100000100",
  61633=>"001001111",
  61634=>"000111111",
  61635=>"110111100",
  61636=>"010000111",
  61637=>"000000000",
  61638=>"010100110",
  61639=>"111111111",
  61640=>"111111000",
  61641=>"100100000",
  61642=>"000111010",
  61643=>"111111000",
  61644=>"000101111",
  61645=>"100000111",
  61646=>"000000000",
  61647=>"000011111",
  61648=>"111101000",
  61649=>"011001010",
  61650=>"000000111",
  61651=>"111111000",
  61652=>"111111111",
  61653=>"101111110",
  61654=>"000000000",
  61655=>"000000000",
  61656=>"000001000",
  61657=>"111111000",
  61658=>"111101000",
  61659=>"010111101",
  61660=>"111111000",
  61661=>"101001111",
  61662=>"111111000",
  61663=>"000111111",
  61664=>"111000001",
  61665=>"000000000",
  61666=>"000010110",
  61667=>"111000000",
  61668=>"111110000",
  61669=>"111000000",
  61670=>"010011000",
  61671=>"000000111",
  61672=>"000011111",
  61673=>"101001111",
  61674=>"000111111",
  61675=>"000000000",
  61676=>"000000100",
  61677=>"000011111",
  61678=>"000000000",
  61679=>"000101110",
  61680=>"111111000",
  61681=>"000000000",
  61682=>"000000000",
  61683=>"101100111",
  61684=>"000000111",
  61685=>"000000110",
  61686=>"000000000",
  61687=>"111101001",
  61688=>"011010000",
  61689=>"000000000",
  61690=>"111111000",
  61691=>"111001001",
  61692=>"000000001",
  61693=>"111111111",
  61694=>"111111111",
  61695=>"111111000",
  61696=>"011000000",
  61697=>"000100000",
  61698=>"111101100",
  61699=>"000000111",
  61700=>"111011000",
  61701=>"001000111",
  61702=>"101111111",
  61703=>"111111000",
  61704=>"111110000",
  61705=>"000000000",
  61706=>"111000000",
  61707=>"000000000",
  61708=>"111100101",
  61709=>"111111000",
  61710=>"100000000",
  61711=>"000000000",
  61712=>"000100100",
  61713=>"000000000",
  61714=>"111000001",
  61715=>"000000111",
  61716=>"000000000",
  61717=>"001111111",
  61718=>"011111100",
  61719=>"011000000",
  61720=>"000111111",
  61721=>"111001001",
  61722=>"000000000",
  61723=>"000000000",
  61724=>"111111111",
  61725=>"000000001",
  61726=>"000000111",
  61727=>"001000111",
  61728=>"010100000",
  61729=>"111011000",
  61730=>"011011010",
  61731=>"000111111",
  61732=>"000000011",
  61733=>"000000000",
  61734=>"111111000",
  61735=>"111000000",
  61736=>"111111111",
  61737=>"000111100",
  61738=>"111011011",
  61739=>"111000000",
  61740=>"000000000",
  61741=>"100101000",
  61742=>"000000000",
  61743=>"110111010",
  61744=>"000000000",
  61745=>"000110111",
  61746=>"111100000",
  61747=>"000010010",
  61748=>"110111000",
  61749=>"000111111",
  61750=>"000000000",
  61751=>"111111000",
  61752=>"111111010",
  61753=>"001000111",
  61754=>"000000000",
  61755=>"111000000",
  61756=>"111000000",
  61757=>"111111111",
  61758=>"100111111",
  61759=>"000000111",
  61760=>"111111111",
  61761=>"110111111",
  61762=>"001000000",
  61763=>"011001001",
  61764=>"000111111",
  61765=>"111111111",
  61766=>"000011111",
  61767=>"000000000",
  61768=>"000000000",
  61769=>"111000000",
  61770=>"101111110",
  61771=>"100001001",
  61772=>"100110111",
  61773=>"111111000",
  61774=>"000000000",
  61775=>"000000000",
  61776=>"000001001",
  61777=>"111010000",
  61778=>"111111000",
  61779=>"111111110",
  61780=>"100000000",
  61781=>"000011001",
  61782=>"000111011",
  61783=>"000000110",
  61784=>"111101111",
  61785=>"111000000",
  61786=>"011111110",
  61787=>"111111001",
  61788=>"010011000",
  61789=>"100100000",
  61790=>"000100110",
  61791=>"001001010",
  61792=>"000111111",
  61793=>"000111001",
  61794=>"000101111",
  61795=>"111111100",
  61796=>"000001011",
  61797=>"001000000",
  61798=>"000000000",
  61799=>"111110111",
  61800=>"100100010",
  61801=>"111111111",
  61802=>"100000011",
  61803=>"010010111",
  61804=>"001000000",
  61805=>"100111111",
  61806=>"011111111",
  61807=>"001110000",
  61808=>"111111111",
  61809=>"000000000",
  61810=>"010101111",
  61811=>"011111111",
  61812=>"000000010",
  61813=>"111100000",
  61814=>"111000001",
  61815=>"000111000",
  61816=>"010000011",
  61817=>"010000111",
  61818=>"000000110",
  61819=>"100000011",
  61820=>"111111111",
  61821=>"100100111",
  61822=>"010010000",
  61823=>"000000000",
  61824=>"000000110",
  61825=>"000100111",
  61826=>"100110111",
  61827=>"111000000",
  61828=>"111011111",
  61829=>"011011000",
  61830=>"101111101",
  61831=>"011001110",
  61832=>"111000101",
  61833=>"000000000",
  61834=>"111011011",
  61835=>"111111011",
  61836=>"101101111",
  61837=>"000110110",
  61838=>"000000000",
  61839=>"010111110",
  61840=>"000011111",
  61841=>"001000110",
  61842=>"011001111",
  61843=>"000000000",
  61844=>"111111111",
  61845=>"000011011",
  61846=>"111111111",
  61847=>"001011001",
  61848=>"111100000",
  61849=>"000110101",
  61850=>"000000000",
  61851=>"000000110",
  61852=>"100111000",
  61853=>"000000000",
  61854=>"001000000",
  61855=>"000000111",
  61856=>"000011101",
  61857=>"100101001",
  61858=>"000000000",
  61859=>"111111100",
  61860=>"111111111",
  61861=>"111111110",
  61862=>"001000001",
  61863=>"111001001",
  61864=>"110101001",
  61865=>"100000000",
  61866=>"111111100",
  61867=>"000000100",
  61868=>"111000000",
  61869=>"100111110",
  61870=>"010111111",
  61871=>"000000111",
  61872=>"111111100",
  61873=>"110000000",
  61874=>"001111110",
  61875=>"100100000",
  61876=>"000000010",
  61877=>"111111000",
  61878=>"001000001",
  61879=>"100000010",
  61880=>"111000000",
  61881=>"011111000",
  61882=>"000111111",
  61883=>"000000111",
  61884=>"110000000",
  61885=>"111000000",
  61886=>"110000011",
  61887=>"100000111",
  61888=>"111110000",
  61889=>"101000000",
  61890=>"111010000",
  61891=>"000000000",
  61892=>"111111111",
  61893=>"011111000",
  61894=>"000110100",
  61895=>"111111000",
  61896=>"011111000",
  61897=>"000000000",
  61898=>"001000101",
  61899=>"000000111",
  61900=>"000110001",
  61901=>"001000001",
  61902=>"100000111",
  61903=>"000011111",
  61904=>"000000111",
  61905=>"000111111",
  61906=>"111111000",
  61907=>"111111001",
  61908=>"111101111",
  61909=>"000111111",
  61910=>"111111011",
  61911=>"000000000",
  61912=>"111000000",
  61913=>"000000111",
  61914=>"001000000",
  61915=>"000000000",
  61916=>"010000000",
  61917=>"000110111",
  61918=>"001011000",
  61919=>"000000101",
  61920=>"011111000",
  61921=>"111000000",
  61922=>"000000101",
  61923=>"111111110",
  61924=>"100101100",
  61925=>"000000011",
  61926=>"001101110",
  61927=>"000111111",
  61928=>"000000000",
  61929=>"001000111",
  61930=>"000000011",
  61931=>"000000111",
  61932=>"000000000",
  61933=>"001011010",
  61934=>"111000000",
  61935=>"010000000",
  61936=>"000111111",
  61937=>"100111111",
  61938=>"111111111",
  61939=>"111111000",
  61940=>"000000111",
  61941=>"000111111",
  61942=>"000000000",
  61943=>"011000100",
  61944=>"111011000",
  61945=>"000111111",
  61946=>"000000000",
  61947=>"111001000",
  61948=>"111101001",
  61949=>"000000000",
  61950=>"001000110",
  61951=>"000000100",
  61952=>"110000000",
  61953=>"111011011",
  61954=>"000011000",
  61955=>"000000000",
  61956=>"000000000",
  61957=>"000000000",
  61958=>"111111000",
  61959=>"000000000",
  61960=>"111111111",
  61961=>"100111111",
  61962=>"111111101",
  61963=>"111111000",
  61964=>"011000001",
  61965=>"100000000",
  61966=>"001011001",
  61967=>"000000110",
  61968=>"110111111",
  61969=>"001001111",
  61970=>"111111111",
  61971=>"111111111",
  61972=>"111111111",
  61973=>"000000000",
  61974=>"111101100",
  61975=>"111111111",
  61976=>"011011000",
  61977=>"000010000",
  61978=>"111111001",
  61979=>"000000000",
  61980=>"000000000",
  61981=>"111111111",
  61982=>"111101101",
  61983=>"111111110",
  61984=>"111111111",
  61985=>"000000111",
  61986=>"000110110",
  61987=>"111101111",
  61988=>"111000100",
  61989=>"111111111",
  61990=>"000000000",
  61991=>"111111111",
  61992=>"000000000",
  61993=>"000011010",
  61994=>"111111100",
  61995=>"111110110",
  61996=>"111111000",
  61997=>"011100111",
  61998=>"111011011",
  61999=>"111111000",
  62000=>"000000000",
  62001=>"111111111",
  62002=>"000000000",
  62003=>"011001100",
  62004=>"001011011",
  62005=>"110110110",
  62006=>"000100100",
  62007=>"011111101",
  62008=>"000100000",
  62009=>"011011000",
  62010=>"111111111",
  62011=>"111111010",
  62012=>"001100110",
  62013=>"111111110",
  62014=>"000001011",
  62015=>"000000000",
  62016=>"111111111",
  62017=>"101101000",
  62018=>"111111000",
  62019=>"111111111",
  62020=>"001011000",
  62021=>"111111110",
  62022=>"111111111",
  62023=>"111111111",
  62024=>"000000001",
  62025=>"001011111",
  62026=>"111111111",
  62027=>"101111111",
  62028=>"101111111",
  62029=>"000000000",
  62030=>"001001111",
  62031=>"000110111",
  62032=>"111111111",
  62033=>"000000000",
  62034=>"111111111",
  62035=>"111110000",
  62036=>"000000000",
  62037=>"000110000",
  62038=>"000001001",
  62039=>"101101100",
  62040=>"110111111",
  62041=>"111111111",
  62042=>"000000000",
  62043=>"101111111",
  62044=>"000000000",
  62045=>"000000111",
  62046=>"111111111",
  62047=>"110111111",
  62048=>"111101111",
  62049=>"000001011",
  62050=>"111111111",
  62051=>"111111111",
  62052=>"000000000",
  62053=>"101111111",
  62054=>"111111111",
  62055=>"111111101",
  62056=>"000000000",
  62057=>"000011111",
  62058=>"001100000",
  62059=>"100100111",
  62060=>"100100000",
  62061=>"000000000",
  62062=>"000000000",
  62063=>"111111111",
  62064=>"000000011",
  62065=>"011011110",
  62066=>"011011011",
  62067=>"111111111",
  62068=>"011011000",
  62069=>"000000000",
  62070=>"000000000",
  62071=>"000000000",
  62072=>"011001001",
  62073=>"000000000",
  62074=>"000000000",
  62075=>"000000000",
  62076=>"100000000",
  62077=>"011001100",
  62078=>"000000000",
  62079=>"010000110",
  62080=>"111111111",
  62081=>"000111111",
  62082=>"000000000",
  62083=>"011111001",
  62084=>"000000000",
  62085=>"111111011",
  62086=>"000000110",
  62087=>"000111111",
  62088=>"111111000",
  62089=>"111010000",
  62090=>"001111111",
  62091=>"111111111",
  62092=>"000000111",
  62093=>"100000000",
  62094=>"000110110",
  62095=>"000000101",
  62096=>"000000000",
  62097=>"000000000",
  62098=>"000010000",
  62099=>"000000000",
  62100=>"111111111",
  62101=>"000000111",
  62102=>"101110100",
  62103=>"110111110",
  62104=>"000000000",
  62105=>"000000111",
  62106=>"100111111",
  62107=>"000010000",
  62108=>"000000000",
  62109=>"001011111",
  62110=>"111111101",
  62111=>"111111111",
  62112=>"111111111",
  62113=>"000010111",
  62114=>"010010011",
  62115=>"111111110",
  62116=>"000000010",
  62117=>"101111000",
  62118=>"010111111",
  62119=>"000000011",
  62120=>"000100110",
  62121=>"111111011",
  62122=>"100110111",
  62123=>"111111011",
  62124=>"111111100",
  62125=>"111111011",
  62126=>"111111101",
  62127=>"011011111",
  62128=>"111111111",
  62129=>"110000000",
  62130=>"111111011",
  62131=>"111100100",
  62132=>"110010000",
  62133=>"100000000",
  62134=>"000011011",
  62135=>"111111111",
  62136=>"001111111",
  62137=>"000000000",
  62138=>"001000001",
  62139=>"100000000",
  62140=>"000110111",
  62141=>"000000000",
  62142=>"000000000",
  62143=>"111111111",
  62144=>"000000011",
  62145=>"110111110",
  62146=>"111111111",
  62147=>"001000000",
  62148=>"000000000",
  62149=>"000000000",
  62150=>"011000000",
  62151=>"001011110",
  62152=>"001101000",
  62153=>"000111111",
  62154=>"001011111",
  62155=>"111111011",
  62156=>"000000001",
  62157=>"001110110",
  62158=>"111111000",
  62159=>"001001001",
  62160=>"000000000",
  62161=>"000100111",
  62162=>"111111111",
  62163=>"111111111",
  62164=>"110111110",
  62165=>"001001001",
  62166=>"110110000",
  62167=>"000000001",
  62168=>"111111010",
  62169=>"111111111",
  62170=>"111111111",
  62171=>"001001000",
  62172=>"101111111",
  62173=>"111111011",
  62174=>"000110010",
  62175=>"111111101",
  62176=>"000000000",
  62177=>"111110110",
  62178=>"111111111",
  62179=>"100111111",
  62180=>"011000000",
  62181=>"111111111",
  62182=>"000000000",
  62183=>"000000000",
  62184=>"111111111",
  62185=>"000001100",
  62186=>"000100111",
  62187=>"001001111",
  62188=>"000011000",
  62189=>"000000000",
  62190=>"111111111",
  62191=>"111000110",
  62192=>"000000000",
  62193=>"000000000",
  62194=>"111100100",
  62195=>"111111111",
  62196=>"110110111",
  62197=>"111111111",
  62198=>"001000010",
  62199=>"010110111",
  62200=>"111111111",
  62201=>"000000000",
  62202=>"000011000",
  62203=>"000000000",
  62204=>"011001001",
  62205=>"110110111",
  62206=>"000000000",
  62207=>"011111001",
  62208=>"100111001",
  62209=>"111001001",
  62210=>"111111111",
  62211=>"000000000",
  62212=>"111111111",
  62213=>"111111110",
  62214=>"000000101",
  62215=>"111011000",
  62216=>"000001001",
  62217=>"000000000",
  62218=>"000000000",
  62219=>"011011000",
  62220=>"000010110",
  62221=>"000000010",
  62222=>"000111111",
  62223=>"111110000",
  62224=>"111111101",
  62225=>"111111111",
  62226=>"000000000",
  62227=>"111111000",
  62228=>"101000111",
  62229=>"000000111",
  62230=>"111111011",
  62231=>"000000000",
  62232=>"100000000",
  62233=>"111110000",
  62234=>"000011011",
  62235=>"111110111",
  62236=>"110111111",
  62237=>"111111111",
  62238=>"111111111",
  62239=>"000001011",
  62240=>"001000000",
  62241=>"111111111",
  62242=>"111011001",
  62243=>"111111111",
  62244=>"000000000",
  62245=>"101110111",
  62246=>"000100111",
  62247=>"000000000",
  62248=>"111111001",
  62249=>"111111111",
  62250=>"111111011",
  62251=>"101100100",
  62252=>"111111111",
  62253=>"111111111",
  62254=>"000100111",
  62255=>"111111111",
  62256=>"111111111",
  62257=>"000000000",
  62258=>"011011001",
  62259=>"000000000",
  62260=>"111111111",
  62261=>"100010001",
  62262=>"000000000",
  62263=>"000000001",
  62264=>"000000111",
  62265=>"000000000",
  62266=>"000000000",
  62267=>"111110100",
  62268=>"001001001",
  62269=>"010111111",
  62270=>"000000111",
  62271=>"110100110",
  62272=>"111110111",
  62273=>"111111000",
  62274=>"111101001",
  62275=>"010010010",
  62276=>"000011111",
  62277=>"111111111",
  62278=>"111111111",
  62279=>"011111111",
  62280=>"111111111",
  62281=>"000000111",
  62282=>"110000110",
  62283=>"110000001",
  62284=>"111111000",
  62285=>"111111000",
  62286=>"001111111",
  62287=>"011001001",
  62288=>"011011000",
  62289=>"000000000",
  62290=>"000110111",
  62291=>"000000000",
  62292=>"110111111",
  62293=>"011011001",
  62294=>"111111111",
  62295=>"000000000",
  62296=>"000000000",
  62297=>"111111111",
  62298=>"110000000",
  62299=>"000000000",
  62300=>"100000000",
  62301=>"000000000",
  62302=>"011011111",
  62303=>"000000000",
  62304=>"010000000",
  62305=>"111001011",
  62306=>"011011011",
  62307=>"111111111",
  62308=>"111111010",
  62309=>"000001011",
  62310=>"000100110",
  62311=>"111111001",
  62312=>"111010000",
  62313=>"010010011",
  62314=>"000000111",
  62315=>"100000111",
  62316=>"110010011",
  62317=>"111011001",
  62318=>"110000000",
  62319=>"000011001",
  62320=>"000000110",
  62321=>"111111110",
  62322=>"000010000",
  62323=>"011001000",
  62324=>"100111111",
  62325=>"000000000",
  62326=>"111111111",
  62327=>"000000100",
  62328=>"111111111",
  62329=>"110110111",
  62330=>"001111111",
  62331=>"000000000",
  62332=>"000000000",
  62333=>"000010000",
  62334=>"000000000",
  62335=>"000001111",
  62336=>"110010011",
  62337=>"111111111",
  62338=>"101111111",
  62339=>"000110000",
  62340=>"000000111",
  62341=>"111111111",
  62342=>"010000000",
  62343=>"111111111",
  62344=>"001000100",
  62345=>"110110110",
  62346=>"111110110",
  62347=>"111111111",
  62348=>"111111111",
  62349=>"011011011",
  62350=>"100001001",
  62351=>"111111000",
  62352=>"111000000",
  62353=>"000001001",
  62354=>"000000000",
  62355=>"110110000",
  62356=>"000000000",
  62357=>"000000000",
  62358=>"000001011",
  62359=>"000010011",
  62360=>"000000111",
  62361=>"111001011",
  62362=>"000000000",
  62363=>"111111111",
  62364=>"000000001",
  62365=>"000000000",
  62366=>"000000100",
  62367=>"000111111",
  62368=>"000000000",
  62369=>"000000000",
  62370=>"000000000",
  62371=>"111111000",
  62372=>"000000001",
  62373=>"111111111",
  62374=>"000000000",
  62375=>"000111111",
  62376=>"111111110",
  62377=>"000000110",
  62378=>"111111111",
  62379=>"110010110",
  62380=>"000000101",
  62381=>"110000001",
  62382=>"001000000",
  62383=>"001011000",
  62384=>"110110111",
  62385=>"000000000",
  62386=>"000000000",
  62387=>"000000000",
  62388=>"111011111",
  62389=>"001000011",
  62390=>"000011111",
  62391=>"111111111",
  62392=>"110110000",
  62393=>"000001000",
  62394=>"000000101",
  62395=>"000000000",
  62396=>"000000000",
  62397=>"101101111",
  62398=>"000000001",
  62399=>"011111111",
  62400=>"110111111",
  62401=>"000000000",
  62402=>"000000000",
  62403=>"111111111",
  62404=>"111011111",
  62405=>"100000000",
  62406=>"111011010",
  62407=>"000000000",
  62408=>"000000000",
  62409=>"111111011",
  62410=>"111111111",
  62411=>"111111111",
  62412=>"011000000",
  62413=>"111111111",
  62414=>"111111011",
  62415=>"000110111",
  62416=>"000000000",
  62417=>"001000010",
  62418=>"000000000",
  62419=>"000000000",
  62420=>"110110100",
  62421=>"101000000",
  62422=>"000000111",
  62423=>"100110110",
  62424=>"011111111",
  62425=>"111011000",
  62426=>"000000101",
  62427=>"000100100",
  62428=>"111000101",
  62429=>"000011000",
  62430=>"111111111",
  62431=>"111111111",
  62432=>"000000100",
  62433=>"000000000",
  62434=>"111111111",
  62435=>"000000101",
  62436=>"000000000",
  62437=>"111010000",
  62438=>"000000111",
  62439=>"000011111",
  62440=>"000010000",
  62441=>"000000000",
  62442=>"000000000",
  62443=>"001001000",
  62444=>"001000100",
  62445=>"000011111",
  62446=>"100111111",
  62447=>"111111111",
  62448=>"000000011",
  62449=>"000000000",
  62450=>"111011111",
  62451=>"111111111",
  62452=>"110110110",
  62453=>"000000000",
  62454=>"111111111",
  62455=>"000000000",
  62456=>"111111111",
  62457=>"110110111",
  62458=>"000000000",
  62459=>"111111111",
  62460=>"111111000",
  62461=>"000000110",
  62462=>"111011011",
  62463=>"000000000",
  62464=>"000100110",
  62465=>"100100111",
  62466=>"111111111",
  62467=>"101110000",
  62468=>"001001011",
  62469=>"000000000",
  62470=>"000000010",
  62471=>"111111000",
  62472=>"111111110",
  62473=>"000000001",
  62474=>"111111111",
  62475=>"011000000",
  62476=>"000000000",
  62477=>"011000000",
  62478=>"111011111",
  62479=>"000000100",
  62480=>"111111001",
  62481=>"111101000",
  62482=>"011001000",
  62483=>"111111111",
  62484=>"000000101",
  62485=>"000000011",
  62486=>"111111011",
  62487=>"111000000",
  62488=>"110111001",
  62489=>"011011110",
  62490=>"110111111",
  62491=>"000100100",
  62492=>"111000000",
  62493=>"110110100",
  62494=>"001001111",
  62495=>"000100000",
  62496=>"000000000",
  62497=>"101000011",
  62498=>"001111111",
  62499=>"111111111",
  62500=>"111111111",
  62501=>"000000000",
  62502=>"001000000",
  62503=>"100111010",
  62504=>"111101001",
  62505=>"000000101",
  62506=>"111111111",
  62507=>"111111101",
  62508=>"000000111",
  62509=>"110001011",
  62510=>"000000100",
  62511=>"011111111",
  62512=>"000000000",
  62513=>"000000000",
  62514=>"011101100",
  62515=>"000100100",
  62516=>"011111111",
  62517=>"011011100",
  62518=>"000001111",
  62519=>"000111100",
  62520=>"001010000",
  62521=>"111110000",
  62522=>"000000000",
  62523=>"011000000",
  62524=>"000010000",
  62525=>"001001111",
  62526=>"000000111",
  62527=>"111111111",
  62528=>"100100111",
  62529=>"111111010",
  62530=>"000110111",
  62531=>"111111111",
  62532=>"110110001",
  62533=>"001100100",
  62534=>"110000000",
  62535=>"000000000",
  62536=>"010111110",
  62537=>"000000000",
  62538=>"000001000",
  62539=>"111111111",
  62540=>"111001000",
  62541=>"000101101",
  62542=>"000000101",
  62543=>"111111000",
  62544=>"101000000",
  62545=>"111000000",
  62546=>"000000010",
  62547=>"111101000",
  62548=>"011010110",
  62549=>"110111111",
  62550=>"101001011",
  62551=>"000000000",
  62552=>"001001000",
  62553=>"000000000",
  62554=>"111000000",
  62555=>"000111111",
  62556=>"111000000",
  62557=>"010100011",
  62558=>"000101111",
  62559=>"111001000",
  62560=>"100000000",
  62561=>"000000000",
  62562=>"010111001",
  62563=>"111000111",
  62564=>"000000111",
  62565=>"111000011",
  62566=>"111100111",
  62567=>"000001011",
  62568=>"100100000",
  62569=>"010000111",
  62570=>"000000110",
  62571=>"111111010",
  62572=>"100110000",
  62573=>"110000001",
  62574=>"000000000",
  62575=>"000000000",
  62576=>"000111111",
  62577=>"000011111",
  62578=>"010110111",
  62579=>"111001001",
  62580=>"001000000",
  62581=>"111000000",
  62582=>"111111111",
  62583=>"011011000",
  62584=>"111100000",
  62585=>"111000100",
  62586=>"011001000",
  62587=>"000000111",
  62588=>"001000000",
  62589=>"100101001",
  62590=>"011011000",
  62591=>"001001000",
  62592=>"011001111",
  62593=>"011110000",
  62594=>"111001000",
  62595=>"100111000",
  62596=>"011111111",
  62597=>"000000000",
  62598=>"111111111",
  62599=>"011000000",
  62600=>"000000000",
  62601=>"010111111",
  62602=>"000000111",
  62603=>"011000000",
  62604=>"111111000",
  62605=>"111111111",
  62606=>"100100111",
  62607=>"000000000",
  62608=>"111111000",
  62609=>"000000000",
  62610=>"101000000",
  62611=>"111000000",
  62612=>"011000000",
  62613=>"000000111",
  62614=>"110110000",
  62615=>"000111111",
  62616=>"111000110",
  62617=>"000000000",
  62618=>"111010111",
  62619=>"111101000",
  62620=>"000000000",
  62621=>"111101000",
  62622=>"000111111",
  62623=>"111100100",
  62624=>"000000111",
  62625=>"001000000",
  62626=>"111000000",
  62627=>"111111111",
  62628=>"011011011",
  62629=>"000000000",
  62630=>"000000000",
  62631=>"000100001",
  62632=>"000100000",
  62633=>"111111111",
  62634=>"000110100",
  62635=>"111001011",
  62636=>"111110111",
  62637=>"010011111",
  62638=>"111111111",
  62639=>"000000000",
  62640=>"111111000",
  62641=>"000011111",
  62642=>"111111011",
  62643=>"000100000",
  62644=>"111101111",
  62645=>"111010111",
  62646=>"001011100",
  62647=>"111111110",
  62648=>"001111111",
  62649=>"000000111",
  62650=>"000000000",
  62651=>"000110111",
  62652=>"000000011",
  62653=>"001000111",
  62654=>"000100111",
  62655=>"001000001",
  62656=>"000000111",
  62657=>"111111111",
  62658=>"111111110",
  62659=>"000000000",
  62660=>"000110110",
  62661=>"111111111",
  62662=>"000111111",
  62663=>"000000000",
  62664=>"111000000",
  62665=>"111100000",
  62666=>"010111111",
  62667=>"111111000",
  62668=>"010111110",
  62669=>"001000000",
  62670=>"011000000",
  62671=>"111000010",
  62672=>"000000000",
  62673=>"000000111",
  62674=>"100000111",
  62675=>"000000000",
  62676=>"111000000",
  62677=>"111000000",
  62678=>"110011111",
  62679=>"000111111",
  62680=>"111111111",
  62681=>"111110000",
  62682=>"000000111",
  62683=>"000000000",
  62684=>"000000000",
  62685=>"011111000",
  62686=>"011001001",
  62687=>"111110000",
  62688=>"000000000",
  62689=>"000000000",
  62690=>"010111110",
  62691=>"000000111",
  62692=>"000000000",
  62693=>"000000110",
  62694=>"000000000",
  62695=>"000000000",
  62696=>"000000000",
  62697=>"111111111",
  62698=>"111100110",
  62699=>"000001000",
  62700=>"111010000",
  62701=>"000000111",
  62702=>"111000000",
  62703=>"111011000",
  62704=>"111110111",
  62705=>"100000111",
  62706=>"111000000",
  62707=>"111111110",
  62708=>"010001111",
  62709=>"110110000",
  62710=>"100100000",
  62711=>"111111000",
  62712=>"010000000",
  62713=>"000100100",
  62714=>"100110110",
  62715=>"000110000",
  62716=>"010010100",
  62717=>"100000000",
  62718=>"000000001",
  62719=>"001011001",
  62720=>"000000000",
  62721=>"001011111",
  62722=>"001001011",
  62723=>"111001001",
  62724=>"101000000",
  62725=>"000000000",
  62726=>"000000100",
  62727=>"001011111",
  62728=>"101100100",
  62729=>"111111111",
  62730=>"101111111",
  62731=>"111111111",
  62732=>"000000010",
  62733=>"000100111",
  62734=>"000001111",
  62735=>"000000000",
  62736=>"111011011",
  62737=>"011000000",
  62738=>"000000110",
  62739=>"111001111",
  62740=>"110101001",
  62741=>"111000000",
  62742=>"100111111",
  62743=>"110110000",
  62744=>"111111100",
  62745=>"001001000",
  62746=>"000000000",
  62747=>"111101000",
  62748=>"000111110",
  62749=>"111000111",
  62750=>"001000110",
  62751=>"001000000",
  62752=>"000000000",
  62753=>"011111111",
  62754=>"100000001",
  62755=>"110111111",
  62756=>"110101111",
  62757=>"001111101",
  62758=>"000000000",
  62759=>"000000000",
  62760=>"111000000",
  62761=>"000010110",
  62762=>"111011111",
  62763=>"011111111",
  62764=>"000010000",
  62765=>"110111100",
  62766=>"100010011",
  62767=>"000100000",
  62768=>"001001111",
  62769=>"111111000",
  62770=>"111000000",
  62771=>"000000001",
  62772=>"010000111",
  62773=>"000000111",
  62774=>"000000000",
  62775=>"000011010",
  62776=>"000000000",
  62777=>"000011001",
  62778=>"111111000",
  62779=>"000000110",
  62780=>"111111111",
  62781=>"110000000",
  62782=>"000000000",
  62783=>"111110000",
  62784=>"111000000",
  62785=>"000001111",
  62786=>"000000011",
  62787=>"000000101",
  62788=>"111100100",
  62789=>"110100000",
  62790=>"100111011",
  62791=>"111111001",
  62792=>"000011111",
  62793=>"111000111",
  62794=>"100100111",
  62795=>"001111101",
  62796=>"000000001",
  62797=>"001111111",
  62798=>"011010110",
  62799=>"110110110",
  62800=>"111111110",
  62801=>"111111111",
  62802=>"111111111",
  62803=>"001000000",
  62804=>"000000000",
  62805=>"011000000",
  62806=>"111000000",
  62807=>"000000110",
  62808=>"111110111",
  62809=>"110111111",
  62810=>"000000000",
  62811=>"001111111",
  62812=>"101111111",
  62813=>"000111111",
  62814=>"000000100",
  62815=>"111110110",
  62816=>"111111111",
  62817=>"110100000",
  62818=>"000001100",
  62819=>"000010000",
  62820=>"111001110",
  62821=>"111111111",
  62822=>"000111111",
  62823=>"011010000",
  62824=>"101111111",
  62825=>"111000000",
  62826=>"111011000",
  62827=>"100111111",
  62828=>"001110000",
  62829=>"110101001",
  62830=>"100000000",
  62831=>"000000000",
  62832=>"000100111",
  62833=>"111111111",
  62834=>"110110000",
  62835=>"100000001",
  62836=>"100000000",
  62837=>"000000010",
  62838=>"111101000",
  62839=>"000000000",
  62840=>"000111111",
  62841=>"000110110",
  62842=>"000000000",
  62843=>"000011111",
  62844=>"000110111",
  62845=>"010111101",
  62846=>"111001111",
  62847=>"001000000",
  62848=>"010010000",
  62849=>"000001000",
  62850=>"010001001",
  62851=>"000100111",
  62852=>"111111110",
  62853=>"000010000",
  62854=>"110100110",
  62855=>"000111101",
  62856=>"000000100",
  62857=>"101001001",
  62858=>"111111111",
  62859=>"111111000",
  62860=>"000111111",
  62861=>"110111111",
  62862=>"001011111",
  62863=>"000000000",
  62864=>"100100000",
  62865=>"000010000",
  62866=>"111111001",
  62867=>"101111111",
  62868=>"000000000",
  62869=>"000000000",
  62870=>"001111111",
  62871=>"011011000",
  62872=>"000000000",
  62873=>"111000000",
  62874=>"111111111",
  62875=>"000000000",
  62876=>"001001100",
  62877=>"000000111",
  62878=>"000000000",
  62879=>"011111111",
  62880=>"011001011",
  62881=>"011011011",
  62882=>"000111111",
  62883=>"111111000",
  62884=>"000000001",
  62885=>"111011111",
  62886=>"000000000",
  62887=>"100110111",
  62888=>"100111111",
  62889=>"000000000",
  62890=>"100100101",
  62891=>"000111111",
  62892=>"000000000",
  62893=>"110110111",
  62894=>"101000000",
  62895=>"000011111",
  62896=>"111000000",
  62897=>"111111000",
  62898=>"000000000",
  62899=>"111111110",
  62900=>"001111111",
  62901=>"000000100",
  62902=>"000100000",
  62903=>"110111000",
  62904=>"110000111",
  62905=>"111010011",
  62906=>"000000000",
  62907=>"111100111",
  62908=>"000000000",
  62909=>"000110110",
  62910=>"100000000",
  62911=>"000010011",
  62912=>"011100111",
  62913=>"111111110",
  62914=>"000011000",
  62915=>"000000000",
  62916=>"000000111",
  62917=>"111110100",
  62918=>"100100111",
  62919=>"011001000",
  62920=>"011001000",
  62921=>"000010111",
  62922=>"000111111",
  62923=>"010111000",
  62924=>"000000111",
  62925=>"010000000",
  62926=>"111001011",
  62927=>"000011111",
  62928=>"000101101",
  62929=>"110000000",
  62930=>"011011011",
  62931=>"111000110",
  62932=>"100001001",
  62933=>"101111110",
  62934=>"100111111",
  62935=>"001000000",
  62936=>"000100000",
  62937=>"111110100",
  62938=>"000101111",
  62939=>"111111000",
  62940=>"100100111",
  62941=>"101000111",
  62942=>"111001001",
  62943=>"111010000",
  62944=>"000000111",
  62945=>"000111111",
  62946=>"000000000",
  62947=>"000100100",
  62948=>"111001000",
  62949=>"110110000",
  62950=>"000000000",
  62951=>"000000001",
  62952=>"111100101",
  62953=>"100000111",
  62954=>"111000000",
  62955=>"111000000",
  62956=>"111100110",
  62957=>"110110110",
  62958=>"000000000",
  62959=>"111111110",
  62960=>"000000010",
  62961=>"111111100",
  62962=>"001101111",
  62963=>"000000000",
  62964=>"000000000",
  62965=>"000000111",
  62966=>"001001111",
  62967=>"110110111",
  62968=>"000000111",
  62969=>"000110110",
  62970=>"111111111",
  62971=>"000000100",
  62972=>"101000011",
  62973=>"000000111",
  62974=>"000111111",
  62975=>"000011011",
  62976=>"110110100",
  62977=>"000000000",
  62978=>"000000000",
  62979=>"111111111",
  62980=>"000100100",
  62981=>"010000000",
  62982=>"110000000",
  62983=>"000000000",
  62984=>"000000111",
  62985=>"110110011",
  62986=>"011111000",
  62987=>"000010111",
  62988=>"110110111",
  62989=>"000000000",
  62990=>"000000000",
  62991=>"111111010",
  62992=>"110110011",
  62993=>"100111111",
  62994=>"111111111",
  62995=>"000000000",
  62996=>"000000100",
  62997=>"000000000",
  62998=>"010000000",
  62999=>"000000100",
  63000=>"100000001",
  63001=>"000011110",
  63002=>"111110111",
  63003=>"110111001",
  63004=>"111111110",
  63005=>"111111100",
  63006=>"110010110",
  63007=>"000000000",
  63008=>"000001000",
  63009=>"111111111",
  63010=>"011110110",
  63011=>"000000000",
  63012=>"000111100",
  63013=>"000110111",
  63014=>"011000000",
  63015=>"111111111",
  63016=>"011111110",
  63017=>"100000000",
  63018=>"001000111",
  63019=>"111111111",
  63020=>"111011000",
  63021=>"111111110",
  63022=>"111111111",
  63023=>"110110100",
  63024=>"000000111",
  63025=>"010111111",
  63026=>"111111111",
  63027=>"111000000",
  63028=>"011011001",
  63029=>"110000010",
  63030=>"001001000",
  63031=>"000000000",
  63032=>"011111111",
  63033=>"010000000",
  63034=>"000000000",
  63035=>"000000000",
  63036=>"001000001",
  63037=>"011000000",
  63038=>"001011001",
  63039=>"000000000",
  63040=>"001011000",
  63041=>"000000000",
  63042=>"010000000",
  63043=>"000000000",
  63044=>"010011001",
  63045=>"111111000",
  63046=>"100100111",
  63047=>"000100111",
  63048=>"111111111",
  63049=>"000000001",
  63050=>"111110111",
  63051=>"111001101",
  63052=>"000000000",
  63053=>"001000001",
  63054=>"000010100",
  63055=>"000000111",
  63056=>"000000000",
  63057=>"111111000",
  63058=>"110111110",
  63059=>"111100000",
  63060=>"000000111",
  63061=>"000000000",
  63062=>"000001100",
  63063=>"111111111",
  63064=>"000000000",
  63065=>"111100111",
  63066=>"100111111",
  63067=>"111111111",
  63068=>"111110110",
  63069=>"000000000",
  63070=>"000101111",
  63071=>"001001100",
  63072=>"111111111",
  63073=>"100100111",
  63074=>"101000000",
  63075=>"000000000",
  63076=>"101000000",
  63077=>"001111111",
  63078=>"111111111",
  63079=>"000000110",
  63080=>"001111110",
  63081=>"111110000",
  63082=>"110111111",
  63083=>"001111111",
  63084=>"111110000",
  63085=>"000000000",
  63086=>"000000011",
  63087=>"000001011",
  63088=>"000011000",
  63089=>"000000001",
  63090=>"011001000",
  63091=>"011001001",
  63092=>"000000100",
  63093=>"000001001",
  63094=>"100101000",
  63095=>"000000000",
  63096=>"011111110",
  63097=>"001000000",
  63098=>"110111000",
  63099=>"000000000",
  63100=>"101111100",
  63101=>"011111111",
  63102=>"111111111",
  63103=>"000000000",
  63104=>"001001001",
  63105=>"000000111",
  63106=>"111111111",
  63107=>"011111010",
  63108=>"000000000",
  63109=>"000000000",
  63110=>"111111111",
  63111=>"000000000",
  63112=>"111111111",
  63113=>"000000000",
  63114=>"000000000",
  63115=>"100000100",
  63116=>"000000000",
  63117=>"000001000",
  63118=>"001001001",
  63119=>"000000001",
  63120=>"111110111",
  63121=>"000000000",
  63122=>"111111000",
  63123=>"000111000",
  63124=>"100110111",
  63125=>"111111111",
  63126=>"000111110",
  63127=>"111111111",
  63128=>"000000100",
  63129=>"111111111",
  63130=>"100001001",
  63131=>"011000000",
  63132=>"011000100",
  63133=>"001101001",
  63134=>"000000000",
  63135=>"000000111",
  63136=>"101000000",
  63137=>"000000100",
  63138=>"011111111",
  63139=>"001110010",
  63140=>"111111111",
  63141=>"111011101",
  63142=>"110111111",
  63143=>"001001000",
  63144=>"011000000",
  63145=>"000110110",
  63146=>"000000000",
  63147=>"000000000",
  63148=>"111111001",
  63149=>"000000011",
  63150=>"111111111",
  63151=>"001110000",
  63152=>"100100000",
  63153=>"111111111",
  63154=>"110111111",
  63155=>"000111111",
  63156=>"000000000",
  63157=>"000000010",
  63158=>"000000000",
  63159=>"000101111",
  63160=>"111111111",
  63161=>"000000001",
  63162=>"111000000",
  63163=>"001101001",
  63164=>"111100110",
  63165=>"000000000",
  63166=>"000111011",
  63167=>"110111000",
  63168=>"001000000",
  63169=>"111110000",
  63170=>"111111100",
  63171=>"000000001",
  63172=>"000000000",
  63173=>"111111111",
  63174=>"100001000",
  63175=>"101000000",
  63176=>"000100000",
  63177=>"000000000",
  63178=>"000000000",
  63179=>"111010010",
  63180=>"000111111",
  63181=>"111111111",
  63182=>"000000001",
  63183=>"000000000",
  63184=>"011111110",
  63185=>"011111111",
  63186=>"000110011",
  63187=>"000000000",
  63188=>"101111111",
  63189=>"000000000",
  63190=>"111111111",
  63191=>"111111110",
  63192=>"000000000",
  63193=>"000000000",
  63194=>"000000000",
  63195=>"010011001",
  63196=>"000000111",
  63197=>"000000000",
  63198=>"111111011",
  63199=>"111000000",
  63200=>"000000000",
  63201=>"010000111",
  63202=>"111111100",
  63203=>"111011000",
  63204=>"000010010",
  63205=>"111001000",
  63206=>"111001001",
  63207=>"000000000",
  63208=>"000000001",
  63209=>"000100111",
  63210=>"011101001",
  63211=>"000000000",
  63212=>"000000000",
  63213=>"111111111",
  63214=>"000000000",
  63215=>"100100100",
  63216=>"000000001",
  63217=>"000000000",
  63218=>"000000000",
  63219=>"110110000",
  63220=>"100111110",
  63221=>"000110110",
  63222=>"100011001",
  63223=>"111111111",
  63224=>"100111101",
  63225=>"000000000",
  63226=>"001111111",
  63227=>"000010011",
  63228=>"011111011",
  63229=>"001000000",
  63230=>"110000000",
  63231=>"011111111",
  63232=>"011000000",
  63233=>"110111111",
  63234=>"111111111",
  63235=>"001111011",
  63236=>"000000000",
  63237=>"000000000",
  63238=>"100111111",
  63239=>"000000000",
  63240=>"111111111",
  63241=>"000000000",
  63242=>"111111001",
  63243=>"000000000",
  63244=>"111111111",
  63245=>"111000000",
  63246=>"100000100",
  63247=>"000000000",
  63248=>"000000000",
  63249=>"000100000",
  63250=>"111111000",
  63251=>"111110110",
  63252=>"100000000",
  63253=>"000000000",
  63254=>"001001001",
  63255=>"000000000",
  63256=>"000000100",
  63257=>"000111111",
  63258=>"111000000",
  63259=>"000000000",
  63260=>"110111110",
  63261=>"111111000",
  63262=>"000000000",
  63263=>"111110111",
  63264=>"011111001",
  63265=>"111111111",
  63266=>"110000000",
  63267=>"111101000",
  63268=>"111010010",
  63269=>"000000000",
  63270=>"111100000",
  63271=>"110110100",
  63272=>"000000000",
  63273=>"111100000",
  63274=>"010000000",
  63275=>"000000000",
  63276=>"111111100",
  63277=>"111001011",
  63278=>"000000000",
  63279=>"001111111",
  63280=>"101011011",
  63281=>"000000011",
  63282=>"111111111",
  63283=>"000000000",
  63284=>"000000101",
  63285=>"111010110",
  63286=>"000101111",
  63287=>"000100100",
  63288=>"000111111",
  63289=>"111111111",
  63290=>"011000000",
  63291=>"111111111",
  63292=>"000000000",
  63293=>"000000000",
  63294=>"111111110",
  63295=>"100100111",
  63296=>"000100000",
  63297=>"111111100",
  63298=>"000110010",
  63299=>"101000000",
  63300=>"000000000",
  63301=>"000001101",
  63302=>"111001000",
  63303=>"000000001",
  63304=>"000011111",
  63305=>"110111111",
  63306=>"011100100",
  63307=>"000000100",
  63308=>"001000000",
  63309=>"111110110",
  63310=>"111111111",
  63311=>"010111110",
  63312=>"011011000",
  63313=>"111111111",
  63314=>"000000000",
  63315=>"000000000",
  63316=>"000111001",
  63317=>"011001001",
  63318=>"111111100",
  63319=>"000000111",
  63320=>"110100110",
  63321=>"111111111",
  63322=>"100100000",
  63323=>"000000000",
  63324=>"100000100",
  63325=>"000000000",
  63326=>"111111110",
  63327=>"111000000",
  63328=>"000000101",
  63329=>"111000010",
  63330=>"101001111",
  63331=>"000111111",
  63332=>"100100000",
  63333=>"111100000",
  63334=>"111111111",
  63335=>"111111111",
  63336=>"000000000",
  63337=>"111111011",
  63338=>"000000000",
  63339=>"000000101",
  63340=>"110100000",
  63341=>"111110000",
  63342=>"000011111",
  63343=>"000111111",
  63344=>"000000000",
  63345=>"000000000",
  63346=>"110110111",
  63347=>"011010000",
  63348=>"111111011",
  63349=>"100101001",
  63350=>"000000000",
  63351=>"001000000",
  63352=>"000000000",
  63353=>"000000000",
  63354=>"000000000",
  63355=>"111111111",
  63356=>"011011000",
  63357=>"001000001",
  63358=>"110110111",
  63359=>"001001011",
  63360=>"001001111",
  63361=>"001000000",
  63362=>"111111001",
  63363=>"000000000",
  63364=>"111111100",
  63365=>"000000000",
  63366=>"110111111",
  63367=>"111111111",
  63368=>"111111111",
  63369=>"100000000",
  63370=>"111111111",
  63371=>"000000000",
  63372=>"000000010",
  63373=>"000001000",
  63374=>"000000000",
  63375=>"000000011",
  63376=>"000000111",
  63377=>"100000110",
  63378=>"010111000",
  63379=>"000000100",
  63380=>"111111111",
  63381=>"000000000",
  63382=>"111111111",
  63383=>"111111111",
  63384=>"111111111",
  63385=>"000001111",
  63386=>"111111000",
  63387=>"111111100",
  63388=>"111111111",
  63389=>"000000000",
  63390=>"000000000",
  63391=>"000000000",
  63392=>"000000000",
  63393=>"011111110",
  63394=>"111010110",
  63395=>"100000101",
  63396=>"100100000",
  63397=>"000000000",
  63398=>"000000111",
  63399=>"010111111",
  63400=>"001111100",
  63401=>"000000000",
  63402=>"111111111",
  63403=>"111111000",
  63404=>"000000000",
  63405=>"011111111",
  63406=>"000000000",
  63407=>"110111111",
  63408=>"000000000",
  63409=>"111111111",
  63410=>"000000000",
  63411=>"000000001",
  63412=>"001001000",
  63413=>"101100000",
  63414=>"111100000",
  63415=>"111111111",
  63416=>"000000000",
  63417=>"111110000",
  63418=>"111110000",
  63419=>"000111111",
  63420=>"000000000",
  63421=>"000001100",
  63422=>"000000100",
  63423=>"000000000",
  63424=>"111111000",
  63425=>"111111111",
  63426=>"000010111",
  63427=>"100011010",
  63428=>"111100000",
  63429=>"100001001",
  63430=>"111110000",
  63431=>"011011110",
  63432=>"111111111",
  63433=>"111100000",
  63434=>"111111111",
  63435=>"111011000",
  63436=>"000000001",
  63437=>"000100111",
  63438=>"001111100",
  63439=>"011011011",
  63440=>"000000000",
  63441=>"001101111",
  63442=>"000000000",
  63443=>"000000000",
  63444=>"000111111",
  63445=>"111111111",
  63446=>"111111111",
  63447=>"001100111",
  63448=>"000000000",
  63449=>"000000000",
  63450=>"111111111",
  63451=>"111111111",
  63452=>"111111111",
  63453=>"000100000",
  63454=>"000000100",
  63455=>"110111000",
  63456=>"000011011",
  63457=>"000000000",
  63458=>"111111111",
  63459=>"000000000",
  63460=>"011111000",
  63461=>"000000001",
  63462=>"000001000",
  63463=>"011011011",
  63464=>"010110110",
  63465=>"111111000",
  63466=>"000110110",
  63467=>"000000000",
  63468=>"111111111",
  63469=>"111111111",
  63470=>"110100001",
  63471=>"111001000",
  63472=>"111111111",
  63473=>"000101111",
  63474=>"111100101",
  63475=>"111111010",
  63476=>"011111111",
  63477=>"111111101",
  63478=>"111111111",
  63479=>"111111111",
  63480=>"000101111",
  63481=>"000000000",
  63482=>"110110000",
  63483=>"000000111",
  63484=>"101111111",
  63485=>"000110110",
  63486=>"110111100",
  63487=>"011001000",
  63488=>"001010000",
  63489=>"000000000",
  63490=>"101111111",
  63491=>"111111111",
  63492=>"000100100",
  63493=>"001000000",
  63494=>"000000000",
  63495=>"111111111",
  63496=>"000000000",
  63497=>"111111111",
  63498=>"000000111",
  63499=>"000100001",
  63500=>"000000000",
  63501=>"000111111",
  63502=>"000000101",
  63503=>"000100111",
  63504=>"100000000",
  63505=>"001101100",
  63506=>"000101101",
  63507=>"011111111",
  63508=>"111001000",
  63509=>"111101111",
  63510=>"000000000",
  63511=>"000110110",
  63512=>"001001111",
  63513=>"110110111",
  63514=>"000000000",
  63515=>"111110111",
  63516=>"111001000",
  63517=>"000011000",
  63518=>"000000000",
  63519=>"110110110",
  63520=>"001100111",
  63521=>"000000000",
  63522=>"000000110",
  63523=>"000110000",
  63524=>"000000000",
  63525=>"111110111",
  63526=>"000000000",
  63527=>"111110011",
  63528=>"111111111",
  63529=>"110111111",
  63530=>"000000000",
  63531=>"111111111",
  63532=>"000000000",
  63533=>"110111000",
  63534=>"000000010",
  63535=>"000100111",
  63536=>"110000110",
  63537=>"000000000",
  63538=>"100100100",
  63539=>"011011110",
  63540=>"100111110",
  63541=>"111111111",
  63542=>"001000000",
  63543=>"111111111",
  63544=>"000000000",
  63545=>"000000000",
  63546=>"000001111",
  63547=>"111111111",
  63548=>"000000000",
  63549=>"000011111",
  63550=>"110111111",
  63551=>"111111101",
  63552=>"000000000",
  63553=>"000000000",
  63554=>"111111001",
  63555=>"000001111",
  63556=>"100000000",
  63557=>"001111111",
  63558=>"111111110",
  63559=>"000000000",
  63560=>"000100100",
  63561=>"000000000",
  63562=>"100110111",
  63563=>"111110100",
  63564=>"101111101",
  63565=>"001000000",
  63566=>"111111111",
  63567=>"111111111",
  63568=>"011111111",
  63569=>"111111111",
  63570=>"000000000",
  63571=>"111110110",
  63572=>"000000000",
  63573=>"111101001",
  63574=>"001011111",
  63575=>"000000000",
  63576=>"111111111",
  63577=>"111001000",
  63578=>"110110111",
  63579=>"000000000",
  63580=>"101111010",
  63581=>"001001111",
  63582=>"000000000",
  63583=>"111110111",
  63584=>"000111111",
  63585=>"100110000",
  63586=>"111100110",
  63587=>"100100000",
  63588=>"010000001",
  63589=>"001000001",
  63590=>"000000000",
  63591=>"011011111",
  63592=>"111111011",
  63593=>"110010000",
  63594=>"000000111",
  63595=>"000000000",
  63596=>"111110000",
  63597=>"000000000",
  63598=>"000000101",
  63599=>"000000000",
  63600=>"001001001",
  63601=>"111111111",
  63602=>"111111111",
  63603=>"000000000",
  63604=>"111111111",
  63605=>"100111111",
  63606=>"000000000",
  63607=>"001111000",
  63608=>"001000000",
  63609=>"001111111",
  63610=>"000000000",
  63611=>"000001000",
  63612=>"000000100",
  63613=>"101111111",
  63614=>"001111000",
  63615=>"000000000",
  63616=>"000011111",
  63617=>"111111111",
  63618=>"010111111",
  63619=>"000000000",
  63620=>"001101111",
  63621=>"111101000",
  63622=>"101111111",
  63623=>"010110101",
  63624=>"000000111",
  63625=>"000000000",
  63626=>"000000110",
  63627=>"111111111",
  63628=>"000000111",
  63629=>"000000100",
  63630=>"111110111",
  63631=>"000000010",
  63632=>"101111111",
  63633=>"000100010",
  63634=>"111111111",
  63635=>"000000000",
  63636=>"001101110",
  63637=>"010000000",
  63638=>"111111111",
  63639=>"000000111",
  63640=>"000000000",
  63641=>"000000000",
  63642=>"111111111",
  63643=>"000000101",
  63644=>"111111111",
  63645=>"001000000",
  63646=>"111111111",
  63647=>"000000001",
  63648=>"000000000",
  63649=>"000000000",
  63650=>"000000000",
  63651=>"111110111",
  63652=>"000000000",
  63653=>"000001000",
  63654=>"000000000",
  63655=>"111111111",
  63656=>"111111110",
  63657=>"000001001",
  63658=>"111000010",
  63659=>"111111111",
  63660=>"110010000",
  63661=>"000000000",
  63662=>"001010000",
  63663=>"000000000",
  63664=>"000011111",
  63665=>"110100000",
  63666=>"101111111",
  63667=>"000000001",
  63668=>"101101001",
  63669=>"001001000",
  63670=>"100111110",
  63671=>"110100111",
  63672=>"000000010",
  63673=>"001111111",
  63674=>"000110111",
  63675=>"001111100",
  63676=>"000000000",
  63677=>"011111111",
  63678=>"111111111",
  63679=>"000000000",
  63680=>"001101111",
  63681=>"000000100",
  63682=>"000000010",
  63683=>"111111110",
  63684=>"111111111",
  63685=>"000111111",
  63686=>"111000000",
  63687=>"000000111",
  63688=>"111111111",
  63689=>"000000000",
  63690=>"000000000",
  63691=>"000000000",
  63692=>"000000000",
  63693=>"111100101",
  63694=>"000111111",
  63695=>"000010000",
  63696=>"000100111",
  63697=>"111111111",
  63698=>"000000000",
  63699=>"001000000",
  63700=>"000000000",
  63701=>"001000000",
  63702=>"011011111",
  63703=>"111111000",
  63704=>"111111111",
  63705=>"010000000",
  63706=>"000000100",
  63707=>"000000000",
  63708=>"000000111",
  63709=>"000000000",
  63710=>"000000111",
  63711=>"001000000",
  63712=>"111111001",
  63713=>"010000001",
  63714=>"111000111",
  63715=>"000000000",
  63716=>"000000000",
  63717=>"111111111",
  63718=>"000000111",
  63719=>"001111111",
  63720=>"111111111",
  63721=>"111111101",
  63722=>"011111111",
  63723=>"000010010",
  63724=>"000000000",
  63725=>"000000111",
  63726=>"000000111",
  63727=>"011000000",
  63728=>"111111111",
  63729=>"111110111",
  63730=>"000000111",
  63731=>"110110001",
  63732=>"111111011",
  63733=>"111011111",
  63734=>"111111111",
  63735=>"111100000",
  63736=>"000111111",
  63737=>"000000100",
  63738=>"000100111",
  63739=>"111111011",
  63740=>"000100000",
  63741=>"001000100",
  63742=>"000001001",
  63743=>"111111111",
  63744=>"000000111",
  63745=>"111111111",
  63746=>"111111111",
  63747=>"111101111",
  63748=>"110110110",
  63749=>"111111111",
  63750=>"100111001",
  63751=>"111111111",
  63752=>"000000010",
  63753=>"010010111",
  63754=>"000000101",
  63755=>"010011011",
  63756=>"111000001",
  63757=>"111111111",
  63758=>"001000001",
  63759=>"111110000",
  63760=>"001001000",
  63761=>"000000110",
  63762=>"111101111",
  63763=>"001001000",
  63764=>"000111111",
  63765=>"000000000",
  63766=>"011111111",
  63767=>"000000000",
  63768=>"000000100",
  63769=>"000000000",
  63770=>"001111111",
  63771=>"000000110",
  63772=>"111011000",
  63773=>"110111000",
  63774=>"000001000",
  63775=>"001000011",
  63776=>"111000000",
  63777=>"000000001",
  63778=>"111111111",
  63779=>"000000010",
  63780=>"111111111",
  63781=>"000000011",
  63782=>"011011011",
  63783=>"111110010",
  63784=>"111000100",
  63785=>"101001111",
  63786=>"111111011",
  63787=>"111111111",
  63788=>"010111110",
  63789=>"001001001",
  63790=>"111111000",
  63791=>"000000000",
  63792=>"001001111",
  63793=>"111111111",
  63794=>"101101111",
  63795=>"011001111",
  63796=>"110111000",
  63797=>"000000000",
  63798=>"011101100",
  63799=>"010000010",
  63800=>"010011000",
  63801=>"011001001",
  63802=>"000010000",
  63803=>"111111111",
  63804=>"001000001",
  63805=>"001000111",
  63806=>"100100111",
  63807=>"110000000",
  63808=>"000000000",
  63809=>"000000000",
  63810=>"001101100",
  63811=>"111111011",
  63812=>"000000000",
  63813=>"111111111",
  63814=>"000000111",
  63815=>"010111111",
  63816=>"000000000",
  63817=>"111111011",
  63818=>"000000000",
  63819=>"100000001",
  63820=>"000000000",
  63821=>"000110111",
  63822=>"000000000",
  63823=>"001000000",
  63824=>"001100100",
  63825=>"011000111",
  63826=>"011111101",
  63827=>"000000000",
  63828=>"011111000",
  63829=>"000000000",
  63830=>"010000110",
  63831=>"100100100",
  63832=>"111111111",
  63833=>"000000000",
  63834=>"100100101",
  63835=>"000000000",
  63836=>"000000000",
  63837=>"100111111",
  63838=>"001010010",
  63839=>"000000000",
  63840=>"111111000",
  63841=>"011111001",
  63842=>"000000000",
  63843=>"111000000",
  63844=>"000000100",
  63845=>"001000000",
  63846=>"111111111",
  63847=>"111001101",
  63848=>"100000000",
  63849=>"000000111",
  63850=>"100000000",
  63851=>"101111011",
  63852=>"010010110",
  63853=>"011000000",
  63854=>"011111111",
  63855=>"111110100",
  63856=>"100110110",
  63857=>"100000000",
  63858=>"000000111",
  63859=>"111111111",
  63860=>"000000000",
  63861=>"000110000",
  63862=>"101100100",
  63863=>"110000000",
  63864=>"000000000",
  63865=>"111111111",
  63866=>"101001001",
  63867=>"110110110",
  63868=>"110100100",
  63869=>"000000000",
  63870=>"001001001",
  63871=>"000000000",
  63872=>"000000100",
  63873=>"000000101",
  63874=>"000100111",
  63875=>"111000000",
  63876=>"010000000",
  63877=>"000101000",
  63878=>"101101100",
  63879=>"111010010",
  63880=>"001111111",
  63881=>"000000000",
  63882=>"111111000",
  63883=>"000000000",
  63884=>"000010000",
  63885=>"111111111",
  63886=>"000000000",
  63887=>"000000001",
  63888=>"111111111",
  63889=>"111111111",
  63890=>"001000010",
  63891=>"110010000",
  63892=>"111110000",
  63893=>"000001000",
  63894=>"101100000",
  63895=>"000000000",
  63896=>"101100110",
  63897=>"000100000",
  63898=>"111000000",
  63899=>"000000000",
  63900=>"101111111",
  63901=>"111111111",
  63902=>"000000000",
  63903=>"000000000",
  63904=>"000000000",
  63905=>"000100100",
  63906=>"111111011",
  63907=>"111111101",
  63908=>"000000001",
  63909=>"110001001",
  63910=>"111111000",
  63911=>"101111110",
  63912=>"101000111",
  63913=>"010001000",
  63914=>"001111111",
  63915=>"011111110",
  63916=>"000000000",
  63917=>"000100101",
  63918=>"111111000",
  63919=>"011010111",
  63920=>"000000000",
  63921=>"111111111",
  63922=>"000110000",
  63923=>"111111111",
  63924=>"000000000",
  63925=>"110111111",
  63926=>"110110110",
  63927=>"010000001",
  63928=>"111101111",
  63929=>"111111111",
  63930=>"000000110",
  63931=>"000000000",
  63932=>"010000000",
  63933=>"000000000",
  63934=>"111001000",
  63935=>"111011110",
  63936=>"110011111",
  63937=>"000101111",
  63938=>"011111001",
  63939=>"000110110",
  63940=>"110110000",
  63941=>"111111111",
  63942=>"011000000",
  63943=>"111011000",
  63944=>"000000000",
  63945=>"000000000",
  63946=>"000000000",
  63947=>"000000000",
  63948=>"000000000",
  63949=>"000001011",
  63950=>"100000001",
  63951=>"111101001",
  63952=>"000011011",
  63953=>"000000111",
  63954=>"100001111",
  63955=>"111000000",
  63956=>"000000000",
  63957=>"000000110",
  63958=>"000001111",
  63959=>"000000000",
  63960=>"111111111",
  63961=>"001001000",
  63962=>"000010111",
  63963=>"111110110",
  63964=>"100000100",
  63965=>"111111110",
  63966=>"100000000",
  63967=>"111011011",
  63968=>"101101011",
  63969=>"101000000",
  63970=>"111111111",
  63971=>"111111110",
  63972=>"001111011",
  63973=>"111111100",
  63974=>"110110111",
  63975=>"111111111",
  63976=>"111111001",
  63977=>"001000100",
  63978=>"100100111",
  63979=>"010000000",
  63980=>"000011000",
  63981=>"000010001",
  63982=>"000100111",
  63983=>"001001101",
  63984=>"111111111",
  63985=>"111111111",
  63986=>"100111110",
  63987=>"111111000",
  63988=>"111111111",
  63989=>"000000101",
  63990=>"000000000",
  63991=>"000000000",
  63992=>"010000010",
  63993=>"011101111",
  63994=>"101001001",
  63995=>"101111111",
  63996=>"111111111",
  63997=>"000100110",
  63998=>"000110110",
  63999=>"111001000",
  64000=>"000000000",
  64001=>"001000000",
  64002=>"111111111",
  64003=>"111111111",
  64004=>"000001000",
  64005=>"000000000",
  64006=>"001000000",
  64007=>"000000000",
  64008=>"000000111",
  64009=>"000000110",
  64010=>"000000000",
  64011=>"111101101",
  64012=>"110111110",
  64013=>"001000000",
  64014=>"100011011",
  64015=>"000000100",
  64016=>"111000001",
  64017=>"111000000",
  64018=>"111000000",
  64019=>"000001111",
  64020=>"000000101",
  64021=>"111111111",
  64022=>"000010010",
  64023=>"111111111",
  64024=>"000000000",
  64025=>"111111111",
  64026=>"111111111",
  64027=>"111111010",
  64028=>"000000000",
  64029=>"111111111",
  64030=>"111111111",
  64031=>"000000000",
  64032=>"111111111",
  64033=>"110100011",
  64034=>"000000001",
  64035=>"111000000",
  64036=>"101111111",
  64037=>"111111111",
  64038=>"111111111",
  64039=>"111111000",
  64040=>"000111101",
  64041=>"000000000",
  64042=>"010010000",
  64043=>"111001111",
  64044=>"110111011",
  64045=>"101111100",
  64046=>"111101000",
  64047=>"111000000",
  64048=>"000000000",
  64049=>"001000000",
  64050=>"000110111",
  64051=>"111111111",
  64052=>"111000000",
  64053=>"011111110",
  64054=>"111111000",
  64055=>"001000000",
  64056=>"111111000",
  64057=>"000001111",
  64058=>"000000000",
  64059=>"111001111",
  64060=>"101100101",
  64061=>"000000100",
  64062=>"110110100",
  64063=>"000000000",
  64064=>"111001001",
  64065=>"000000000",
  64066=>"000011011",
  64067=>"000000000",
  64068=>"000000000",
  64069=>"111100110",
  64070=>"101101100",
  64071=>"111111111",
  64072=>"000110110",
  64073=>"000000000",
  64074=>"111111111",
  64075=>"101111111",
  64076=>"000110111",
  64077=>"111111110",
  64078=>"100000000",
  64079=>"000000000",
  64080=>"101001111",
  64081=>"111111111",
  64082=>"111000000",
  64083=>"010000000",
  64084=>"000000000",
  64085=>"000000000",
  64086=>"000000000",
  64087=>"111111001",
  64088=>"111000000",
  64089=>"000000101",
  64090=>"000001111",
  64091=>"111111111",
  64092=>"000000000",
  64093=>"111111111",
  64094=>"110010001",
  64095=>"110010000",
  64096=>"000110111",
  64097=>"111011000",
  64098=>"000000000",
  64099=>"111001000",
  64100=>"001001111",
  64101=>"111000111",
  64102=>"111110010",
  64103=>"111101101",
  64104=>"111011000",
  64105=>"111111111",
  64106=>"111111111",
  64107=>"000000111",
  64108=>"111000000",
  64109=>"111101010",
  64110=>"111111111",
  64111=>"110100110",
  64112=>"111111111",
  64113=>"101001000",
  64114=>"000000000",
  64115=>"110110000",
  64116=>"111111111",
  64117=>"100100111",
  64118=>"111111000",
  64119=>"000000000",
  64120=>"111000000",
  64121=>"000000001",
  64122=>"000111111",
  64123=>"111101100",
  64124=>"001101001",
  64125=>"011001001",
  64126=>"000000111",
  64127=>"100111111",
  64128=>"001100101",
  64129=>"100000001",
  64130=>"011010100",
  64131=>"000111000",
  64132=>"111100000",
  64133=>"111101111",
  64134=>"111111111",
  64135=>"110000000",
  64136=>"000111111",
  64137=>"111101111",
  64138=>"000000000",
  64139=>"101111111",
  64140=>"111111111",
  64141=>"000010010",
  64142=>"111111011",
  64143=>"111111111",
  64144=>"010000000",
  64145=>"111111111",
  64146=>"011001000",
  64147=>"000000111",
  64148=>"111111111",
  64149=>"001000000",
  64150=>"011000000",
  64151=>"000000000",
  64152=>"011001000",
  64153=>"100110100",
  64154=>"001000111",
  64155=>"000000011",
  64156=>"000000000",
  64157=>"110100111",
  64158=>"011100001",
  64159=>"000101000",
  64160=>"000000000",
  64161=>"101101001",
  64162=>"000000000",
  64163=>"111111111",
  64164=>"001011000",
  64165=>"011000000",
  64166=>"000011110",
  64167=>"110100000",
  64168=>"000000111",
  64169=>"000000000",
  64170=>"111111111",
  64171=>"111111111",
  64172=>"100111111",
  64173=>"110110100",
  64174=>"111101001",
  64175=>"111110111",
  64176=>"000000000",
  64177=>"111110110",
  64178=>"111111111",
  64179=>"111111000",
  64180=>"111111100",
  64181=>"101000000",
  64182=>"000111111",
  64183=>"000000000",
  64184=>"111111111",
  64185=>"111000000",
  64186=>"000101101",
  64187=>"010111011",
  64188=>"111000000",
  64189=>"111001000",
  64190=>"101000000",
  64191=>"000000111",
  64192=>"000000000",
  64193=>"100111111",
  64194=>"000000000",
  64195=>"000000000",
  64196=>"011000110",
  64197=>"000000000",
  64198=>"000111011",
  64199=>"000000000",
  64200=>"110011011",
  64201=>"000000000",
  64202=>"001001001",
  64203=>"000000101",
  64204=>"000111101",
  64205=>"011011001",
  64206=>"000001000",
  64207=>"000000000",
  64208=>"110010000",
  64209=>"101000000",
  64210=>"000001000",
  64211=>"000000000",
  64212=>"000000000",
  64213=>"100111111",
  64214=>"111111111",
  64215=>"111110000",
  64216=>"101111111",
  64217=>"111111111",
  64218=>"000000000",
  64219=>"111101100",
  64220=>"111011111",
  64221=>"000100111",
  64222=>"111111111",
  64223=>"011111111",
  64224=>"111111111",
  64225=>"000000110",
  64226=>"010111111",
  64227=>"011111001",
  64228=>"111111111",
  64229=>"111111111",
  64230=>"000010000",
  64231=>"000000000",
  64232=>"010111111",
  64233=>"000000000",
  64234=>"101000000",
  64235=>"000101111",
  64236=>"111010000",
  64237=>"101000000",
  64238=>"110101000",
  64239=>"111000000",
  64240=>"011000111",
  64241=>"111101101",
  64242=>"111111111",
  64243=>"101100111",
  64244=>"000010000",
  64245=>"111111000",
  64246=>"010010100",
  64247=>"011111111",
  64248=>"000111111",
  64249=>"111111110",
  64250=>"000000000",
  64251=>"000000011",
  64252=>"000000000",
  64253=>"001011011",
  64254=>"001111111",
  64255=>"000000100",
  64256=>"000001001",
  64257=>"000000000",
  64258=>"111111001",
  64259=>"011010011",
  64260=>"110111110",
  64261=>"000100110",
  64262=>"000000000",
  64263=>"000000100",
  64264=>"000100000",
  64265=>"111111111",
  64266=>"111111111",
  64267=>"000100001",
  64268=>"001001000",
  64269=>"010000000",
  64270=>"111111111",
  64271=>"110111111",
  64272=>"000000000",
  64273=>"000000000",
  64274=>"000000000",
  64275=>"001011111",
  64276=>"000000000",
  64277=>"000000010",
  64278=>"111111110",
  64279=>"111111000",
  64280=>"000011011",
  64281=>"111110111",
  64282=>"111111110",
  64283=>"110110010",
  64284=>"001001001",
  64285=>"000000000",
  64286=>"111111111",
  64287=>"000000010",
  64288=>"100110100",
  64289=>"000000000",
  64290=>"000100100",
  64291=>"000000000",
  64292=>"000000000",
  64293=>"011111111",
  64294=>"000000000",
  64295=>"100111110",
  64296=>"101000110",
  64297=>"111111101",
  64298=>"111111000",
  64299=>"000000000",
  64300=>"001001000",
  64301=>"110111111",
  64302=>"100111111",
  64303=>"000000000",
  64304=>"000010111",
  64305=>"000000000",
  64306=>"111111011",
  64307=>"001101111",
  64308=>"111001001",
  64309=>"000000111",
  64310=>"000000000",
  64311=>"111011000",
  64312=>"111000000",
  64313=>"000000000",
  64314=>"111111101",
  64315=>"000001001",
  64316=>"000000111",
  64317=>"100000010",
  64318=>"110110110",
  64319=>"110010000",
  64320=>"000000000",
  64321=>"110111111",
  64322=>"111111011",
  64323=>"000000000",
  64324=>"011011001",
  64325=>"111111111",
  64326=>"111001000",
  64327=>"000000110",
  64328=>"111111100",
  64329=>"111000000",
  64330=>"101000000",
  64331=>"000000000",
  64332=>"111000000",
  64333=>"000000000",
  64334=>"000111111",
  64335=>"011010000",
  64336=>"111001001",
  64337=>"001101111",
  64338=>"110110100",
  64339=>"111100000",
  64340=>"000111111",
  64341=>"111111111",
  64342=>"111111111",
  64343=>"000000100",
  64344=>"111000001",
  64345=>"000000000",
  64346=>"000000000",
  64347=>"000000110",
  64348=>"111111101",
  64349=>"101000111",
  64350=>"001000000",
  64351=>"111011011",
  64352=>"001011011",
  64353=>"111110010",
  64354=>"111111111",
  64355=>"000000000",
  64356=>"000000000",
  64357=>"100110111",
  64358=>"011011001",
  64359=>"111111111",
  64360=>"011001001",
  64361=>"000000000",
  64362=>"000000000",
  64363=>"000000100",
  64364=>"110010001",
  64365=>"000101100",
  64366=>"111111111",
  64367=>"000000110",
  64368=>"111111100",
  64369=>"000000000",
  64370=>"000000001",
  64371=>"000000000",
  64372=>"000000000",
  64373=>"111000000",
  64374=>"100100000",
  64375=>"110000110",
  64376=>"101000000",
  64377=>"001000000",
  64378=>"110110111",
  64379=>"011101101",
  64380=>"000000000",
  64381=>"010111111",
  64382=>"111111111",
  64383=>"000000000",
  64384=>"000011111",
  64385=>"111100101",
  64386=>"111000111",
  64387=>"000000011",
  64388=>"000000111",
  64389=>"111111111",
  64390=>"111011000",
  64391=>"110111110",
  64392=>"111001001",
  64393=>"111001000",
  64394=>"111111110",
  64395=>"000000111",
  64396=>"000000111",
  64397=>"000100110",
  64398=>"111111100",
  64399=>"111111111",
  64400=>"000000100",
  64401=>"101001000",
  64402=>"111111111",
  64403=>"000000110",
  64404=>"111111111",
  64405=>"000010000",
  64406=>"111111111",
  64407=>"111000100",
  64408=>"001000000",
  64409=>"111111110",
  64410=>"001001111",
  64411=>"111111101",
  64412=>"000000001",
  64413=>"001001010",
  64414=>"001001001",
  64415=>"000000000",
  64416=>"111101111",
  64417=>"111110100",
  64418=>"011011011",
  64419=>"000111111",
  64420=>"111111111",
  64421=>"100111111",
  64422=>"111001111",
  64423=>"000111010",
  64424=>"111000010",
  64425=>"111110110",
  64426=>"111111111",
  64427=>"001000000",
  64428=>"000000000",
  64429=>"000000000",
  64430=>"000111110",
  64431=>"000000000",
  64432=>"000001000",
  64433=>"000000000",
  64434=>"111111111",
  64435=>"000000000",
  64436=>"111101111",
  64437=>"010110111",
  64438=>"111101001",
  64439=>"000000001",
  64440=>"010111001",
  64441=>"110111011",
  64442=>"111111000",
  64443=>"111111111",
  64444=>"000000000",
  64445=>"011000000",
  64446=>"000010010",
  64447=>"111111011",
  64448=>"000000011",
  64449=>"000000111",
  64450=>"010011111",
  64451=>"111001000",
  64452=>"001101001",
  64453=>"000111111",
  64454=>"111000111",
  64455=>"000000000",
  64456=>"001101000",
  64457=>"000000110",
  64458=>"000000000",
  64459=>"110111000",
  64460=>"111001001",
  64461=>"010111111",
  64462=>"111000000",
  64463=>"111111100",
  64464=>"000000000",
  64465=>"001101111",
  64466=>"001001001",
  64467=>"111111001",
  64468=>"000000000",
  64469=>"011001111",
  64470=>"111111110",
  64471=>"101111011",
  64472=>"000000100",
  64473=>"111001001",
  64474=>"000000000",
  64475=>"000100001",
  64476=>"000011011",
  64477=>"111111111",
  64478=>"000000011",
  64479=>"000110111",
  64480=>"111011000",
  64481=>"111111111",
  64482=>"000000111",
  64483=>"001000110",
  64484=>"111111111",
  64485=>"011000111",
  64486=>"111110110",
  64487=>"000101111",
  64488=>"011001111",
  64489=>"000000000",
  64490=>"001001111",
  64491=>"000000000",
  64492=>"111111001",
  64493=>"111111011",
  64494=>"111111111",
  64495=>"101001000",
  64496=>"000000000",
  64497=>"100000000",
  64498=>"001001000",
  64499=>"000000000",
  64500=>"001001011",
  64501=>"111111111",
  64502=>"000000111",
  64503=>"111111100",
  64504=>"000000111",
  64505=>"111001000",
  64506=>"100000000",
  64507=>"011111111",
  64508=>"111111110",
  64509=>"111111111",
  64510=>"111101100",
  64511=>"111000001",
  64512=>"001101100",
  64513=>"100000111",
  64514=>"111111000",
  64515=>"000001001",
  64516=>"001101000",
  64517=>"110001000",
  64518=>"111000000",
  64519=>"000001111",
  64520=>"111111000",
  64521=>"000000111",
  64522=>"111111110",
  64523=>"000111111",
  64524=>"110010000",
  64525=>"001000000",
  64526=>"100100011",
  64527=>"111111111",
  64528=>"001110111",
  64529=>"000111111",
  64530=>"110110010",
  64531=>"110110101",
  64532=>"110000000",
  64533=>"101000000",
  64534=>"010111000",
  64535=>"011111111",
  64536=>"111111111",
  64537=>"000000000",
  64538=>"000000101",
  64539=>"110100000",
  64540=>"001000101",
  64541=>"001000000",
  64542=>"111111111",
  64543=>"111111011",
  64544=>"000111111",
  64545=>"001100111",
  64546=>"010111000",
  64547=>"000111011",
  64548=>"000000000",
  64549=>"000010000",
  64550=>"000000000",
  64551=>"111000000",
  64552=>"101000111",
  64553=>"000100001",
  64554=>"111111111",
  64555=>"001000111",
  64556=>"111111111",
  64557=>"111011000",
  64558=>"111101000",
  64559=>"100000000",
  64560=>"110111111",
  64561=>"111111000",
  64562=>"111111011",
  64563=>"100111111",
  64564=>"000000111",
  64565=>"011011110",
  64566=>"111000110",
  64567=>"000110110",
  64568=>"101000100",
  64569=>"000000000",
  64570=>"111111111",
  64571=>"111011101",
  64572=>"111111001",
  64573=>"111100000",
  64574=>"111111111",
  64575=>"100000111",
  64576=>"111111111",
  64577=>"000000000",
  64578=>"111111111",
  64579=>"000000000",
  64580=>"111101000",
  64581=>"011000001",
  64582=>"111111000",
  64583=>"111111111",
  64584=>"001000000",
  64585=>"000000111",
  64586=>"001111111",
  64587=>"001000111",
  64588=>"001001000",
  64589=>"010010000",
  64590=>"110101111",
  64591=>"000110111",
  64592=>"110000000",
  64593=>"000001001",
  64594=>"111111111",
  64595=>"100100000",
  64596=>"001000000",
  64597=>"000000000",
  64598=>"000001111",
  64599=>"000001111",
  64600=>"000111111",
  64601=>"111111111",
  64602=>"000010000",
  64603=>"101001000",
  64604=>"000000000",
  64605=>"111001111",
  64606=>"011001100",
  64607=>"100111011",
  64608=>"111101001",
  64609=>"000111111",
  64610=>"000000010",
  64611=>"000000111",
  64612=>"000000000",
  64613=>"011001100",
  64614=>"111111111",
  64615=>"000000000",
  64616=>"010010010",
  64617=>"110101111",
  64618=>"111111100",
  64619=>"000010110",
  64620=>"111111111",
  64621=>"111111111",
  64622=>"111001111",
  64623=>"001101111",
  64624=>"000000111",
  64625=>"000000000",
  64626=>"111000000",
  64627=>"111001000",
  64628=>"111111011",
  64629=>"111111111",
  64630=>"111111000",
  64631=>"111111111",
  64632=>"000010000",
  64633=>"011111111",
  64634=>"000000011",
  64635=>"111110000",
  64636=>"100100000",
  64637=>"000000110",
  64638=>"000000111",
  64639=>"000000000",
  64640=>"111111000",
  64641=>"000000000",
  64642=>"111000100",
  64643=>"111111111",
  64644=>"110111111",
  64645=>"111110111",
  64646=>"100110000",
  64647=>"001000110",
  64648=>"111111111",
  64649=>"000110000",
  64650=>"000000011",
  64651=>"111110111",
  64652=>"010000000",
  64653=>"000000011",
  64654=>"000000010",
  64655=>"111110000",
  64656=>"000000000",
  64657=>"110110111",
  64658=>"011111000",
  64659=>"110111000",
  64660=>"000000011",
  64661=>"000000001",
  64662=>"001011011",
  64663=>"111011001",
  64664=>"001000000",
  64665=>"000001100",
  64666=>"111000001",
  64667=>"000000000",
  64668=>"100010111",
  64669=>"000001111",
  64670=>"100000000",
  64671=>"101100100",
  64672=>"011000000",
  64673=>"111001000",
  64674=>"101000100",
  64675=>"000011111",
  64676=>"010111000",
  64677=>"001101101",
  64678=>"001000000",
  64679=>"111111100",
  64680=>"000100000",
  64681=>"111111000",
  64682=>"000000000",
  64683=>"000000110",
  64684=>"000111111",
  64685=>"000000011",
  64686=>"111111000",
  64687=>"000000000",
  64688=>"111001000",
  64689=>"100111011",
  64690=>"000111010",
  64691=>"000000101",
  64692=>"100000000",
  64693=>"000000111",
  64694=>"000000000",
  64695=>"000000111",
  64696=>"001001111",
  64697=>"000000111",
  64698=>"000000000",
  64699=>"011111111",
  64700=>"000001000",
  64701=>"000000000",
  64702=>"000010000",
  64703=>"111101111",
  64704=>"111111001",
  64705=>"111101111",
  64706=>"111111111",
  64707=>"001111111",
  64708=>"000111000",
  64709=>"000000111",
  64710=>"000001100",
  64711=>"110110000",
  64712=>"111111111",
  64713=>"001000000",
  64714=>"000000100",
  64715=>"111111111",
  64716=>"000000111",
  64717=>"011111110",
  64718=>"111111111",
  64719=>"011111111",
  64720=>"000000000",
  64721=>"010011001",
  64722=>"111111011",
  64723=>"111011000",
  64724=>"111000000",
  64725=>"000100100",
  64726=>"000000001",
  64727=>"000011110",
  64728=>"011100111",
  64729=>"111111000",
  64730=>"000100100",
  64731=>"000110111",
  64732=>"001000000",
  64733=>"111111111",
  64734=>"000000001",
  64735=>"001101111",
  64736=>"001111111",
  64737=>"000010000",
  64738=>"111011000",
  64739=>"101111111",
  64740=>"000000111",
  64741=>"101000110",
  64742=>"111001111",
  64743=>"000000011",
  64744=>"111111011",
  64745=>"011011101",
  64746=>"111110000",
  64747=>"000000111",
  64748=>"111111111",
  64749=>"000010000",
  64750=>"000000111",
  64751=>"000000000",
  64752=>"111111111",
  64753=>"000000000",
  64754=>"111011000",
  64755=>"010111111",
  64756=>"000000111",
  64757=>"111111110",
  64758=>"000000001",
  64759=>"111111000",
  64760=>"000000000",
  64761=>"000001101",
  64762=>"001000000",
  64763=>"001001000",
  64764=>"011001001",
  64765=>"110010000",
  64766=>"011000000",
  64767=>"111111100",
  64768=>"101101111",
  64769=>"000000111",
  64770=>"111111111",
  64771=>"001000001",
  64772=>"111111000",
  64773=>"000000000",
  64774=>"111110100",
  64775=>"101000111",
  64776=>"001000000",
  64777=>"001111011",
  64778=>"000000111",
  64779=>"111111000",
  64780=>"101001101",
  64781=>"101000000",
  64782=>"000000011",
  64783=>"111110111",
  64784=>"000011000",
  64785=>"101000111",
  64786=>"111100000",
  64787=>"001111111",
  64788=>"000000111",
  64789=>"001000111",
  64790=>"011111110",
  64791=>"111000111",
  64792=>"001111111",
  64793=>"111111111",
  64794=>"000000000",
  64795=>"000000000",
  64796=>"001001000",
  64797=>"000100111",
  64798=>"010111111",
  64799=>"000000100",
  64800=>"110111100",
  64801=>"100111111",
  64802=>"000000110",
  64803=>"000000111",
  64804=>"111011110",
  64805=>"001000000",
  64806=>"000000000",
  64807=>"101000100",
  64808=>"111111001",
  64809=>"001000000",
  64810=>"010000000",
  64811=>"000000010",
  64812=>"000000111",
  64813=>"111011000",
  64814=>"000000000",
  64815=>"000000000",
  64816=>"000111111",
  64817=>"111000000",
  64818=>"110111110",
  64819=>"111010000",
  64820=>"110110000",
  64821=>"111111110",
  64822=>"111011000",
  64823=>"100111111",
  64824=>"111111010",
  64825=>"001000000",
  64826=>"000001111",
  64827=>"010010000",
  64828=>"011000001",
  64829=>"011000010",
  64830=>"000110111",
  64831=>"101000000",
  64832=>"000000000",
  64833=>"000000000",
  64834=>"111101000",
  64835=>"000010111",
  64836=>"000000000",
  64837=>"001000111",
  64838=>"111111100",
  64839=>"000010000",
  64840=>"000000111",
  64841=>"111000000",
  64842=>"011001111",
  64843=>"000100100",
  64844=>"011000111",
  64845=>"000011111",
  64846=>"111111111",
  64847=>"000001001",
  64848=>"011101111",
  64849=>"110000010",
  64850=>"000000000",
  64851=>"001000000",
  64852=>"000001000",
  64853=>"011011011",
  64854=>"001111111",
  64855=>"111101111",
  64856=>"111111111",
  64857=>"111000000",
  64858=>"000000111",
  64859=>"000111111",
  64860=>"011111111",
  64861=>"110100000",
  64862=>"111100000",
  64863=>"001000111",
  64864=>"111001110",
  64865=>"111111111",
  64866=>"110111001",
  64867=>"001001001",
  64868=>"000000000",
  64869=>"111111001",
  64870=>"111111101",
  64871=>"000000100",
  64872=>"011011011",
  64873=>"111001000",
  64874=>"000000011",
  64875=>"100011111",
  64876=>"111001000",
  64877=>"000111110",
  64878=>"111111111",
  64879=>"001001001",
  64880=>"110010010",
  64881=>"010111111",
  64882=>"110000000",
  64883=>"010111000",
  64884=>"000000000",
  64885=>"111111111",
  64886=>"000000000",
  64887=>"001000000",
  64888=>"111000110",
  64889=>"010000111",
  64890=>"000001111",
  64891=>"100000000",
  64892=>"111001111",
  64893=>"001011111",
  64894=>"101000000",
  64895=>"000000100",
  64896=>"000111111",
  64897=>"000111111",
  64898=>"111100100",
  64899=>"111111111",
  64900=>"111000000",
  64901=>"110100110",
  64902=>"011111111",
  64903=>"100000000",
  64904=>"111011010",
  64905=>"001011111",
  64906=>"000011111",
  64907=>"000010000",
  64908=>"101111111",
  64909=>"000110111",
  64910=>"111111000",
  64911=>"101111111",
  64912=>"000000000",
  64913=>"001000000",
  64914=>"111000111",
  64915=>"101100100",
  64916=>"010111111",
  64917=>"000001011",
  64918=>"000010111",
  64919=>"110111100",
  64920=>"010000111",
  64921=>"000111111",
  64922=>"111111111",
  64923=>"000000111",
  64924=>"111111111",
  64925=>"111101100",
  64926=>"111111000",
  64927=>"000110111",
  64928=>"001001111",
  64929=>"111110111",
  64930=>"010000111",
  64931=>"000111111",
  64932=>"101111111",
  64933=>"000000000",
  64934=>"000000001",
  64935=>"000000000",
  64936=>"100100011",
  64937=>"000111000",
  64938=>"100000111",
  64939=>"001000000",
  64940=>"000000000",
  64941=>"001111111",
  64942=>"000000000",
  64943=>"111001000",
  64944=>"110000000",
  64945=>"110111000",
  64946=>"000000000",
  64947=>"111001011",
  64948=>"111111000",
  64949=>"111111000",
  64950=>"111011111",
  64951=>"100000000",
  64952=>"000000011",
  64953=>"111101111",
  64954=>"011000001",
  64955=>"111000111",
  64956=>"110111111",
  64957=>"000000111",
  64958=>"000000000",
  64959=>"000111111",
  64960=>"000001000",
  64961=>"000000011",
  64962=>"000000000",
  64963=>"000000111",
  64964=>"000000111",
  64965=>"101000010",
  64966=>"010010111",
  64967=>"111111111",
  64968=>"000001011",
  64969=>"111111000",
  64970=>"100100100",
  64971=>"111101100",
  64972=>"000111111",
  64973=>"111001111",
  64974=>"000100100",
  64975=>"110111111",
  64976=>"111011000",
  64977=>"000000001",
  64978=>"001111111",
  64979=>"111111111",
  64980=>"010011111",
  64981=>"000000111",
  64982=>"000011011",
  64983=>"111111011",
  64984=>"000000000",
  64985=>"001100101",
  64986=>"101111100",
  64987=>"111111000",
  64988=>"001010110",
  64989=>"000000111",
  64990=>"111111000",
  64991=>"000000000",
  64992=>"011111000",
  64993=>"111000000",
  64994=>"010000000",
  64995=>"100000111",
  64996=>"001000101",
  64997=>"000000111",
  64998=>"000000110",
  64999=>"001101000",
  65000=>"111000101",
  65001=>"000000111",
  65002=>"000000110",
  65003=>"110000100",
  65004=>"000000000",
  65005=>"110110000",
  65006=>"011111111",
  65007=>"111111110",
  65008=>"001011000",
  65009=>"000000001",
  65010=>"000000110",
  65011=>"001111001",
  65012=>"000000000",
  65013=>"000100100",
  65014=>"000011101",
  65015=>"110111111",
  65016=>"011000000",
  65017=>"001110111",
  65018=>"111000000",
  65019=>"111001111",
  65020=>"101101000",
  65021=>"101000111",
  65022=>"111111000",
  65023=>"101000000",
  65024=>"110111111",
  65025=>"111111111",
  65026=>"000000100",
  65027=>"111111100",
  65028=>"011111111",
  65029=>"111011111",
  65030=>"000000000",
  65031=>"111111111",
  65032=>"000000001",
  65033=>"000001001",
  65034=>"000000001",
  65035=>"111111111",
  65036=>"000000011",
  65037=>"111100111",
  65038=>"101100100",
  65039=>"111111000",
  65040=>"111111111",
  65041=>"111111111",
  65042=>"000000000",
  65043=>"111111111",
  65044=>"110000000",
  65045=>"000000000",
  65046=>"111111011",
  65047=>"000001000",
  65048=>"011001011",
  65049=>"111111011",
  65050=>"000000000",
  65051=>"010110111",
  65052=>"000000000",
  65053=>"100111000",
  65054=>"111110100",
  65055=>"111111111",
  65056=>"011011001",
  65057=>"000110110",
  65058=>"000000010",
  65059=>"000000110",
  65060=>"111001001",
  65061=>"000111111",
  65062=>"000000111",
  65063=>"000100000",
  65064=>"000001101",
  65065=>"000000000",
  65066=>"001111111",
  65067=>"100101101",
  65068=>"111111111",
  65069=>"111010000",
  65070=>"100000000",
  65071=>"000010000",
  65072=>"111010110",
  65073=>"111110000",
  65074=>"100000001",
  65075=>"000000100",
  65076=>"111111000",
  65077=>"000011011",
  65078=>"000101101",
  65079=>"011000000",
  65080=>"000000000",
  65081=>"101111111",
  65082=>"010010000",
  65083=>"101000000",
  65084=>"000001000",
  65085=>"001011111",
  65086=>"011011010",
  65087=>"111111111",
  65088=>"000001000",
  65089=>"111000000",
  65090=>"111000001",
  65091=>"000000000",
  65092=>"111111100",
  65093=>"110110100",
  65094=>"000000001",
  65095=>"000000000",
  65096=>"111111111",
  65097=>"000100110",
  65098=>"111111111",
  65099=>"000000001",
  65100=>"111110000",
  65101=>"111111111",
  65102=>"000000101",
  65103=>"111111100",
  65104=>"010000000",
  65105=>"110110111",
  65106=>"001100111",
  65107=>"000000000",
  65108=>"111111001",
  65109=>"111110100",
  65110=>"000000001",
  65111=>"111011000",
  65112=>"000000111",
  65113=>"110101111",
  65114=>"000000000",
  65115=>"111111110",
  65116=>"000000001",
  65117=>"111111111",
  65118=>"000000000",
  65119=>"111001001",
  65120=>"000000000",
  65121=>"110110110",
  65122=>"111111011",
  65123=>"000000111",
  65124=>"011001000",
  65125=>"000000000",
  65126=>"011011111",
  65127=>"000100100",
  65128=>"111110000",
  65129=>"000010111",
  65130=>"111111111",
  65131=>"000000000",
  65132=>"000000000",
  65133=>"111111111",
  65134=>"000001001",
  65135=>"000000000",
  65136=>"001111111",
  65137=>"111101000",
  65138=>"101001011",
  65139=>"111111111",
  65140=>"000000000",
  65141=>"111100100",
  65142=>"010000000",
  65143=>"111111111",
  65144=>"001000100",
  65145=>"000100101",
  65146=>"000000000",
  65147=>"000000000",
  65148=>"000100110",
  65149=>"111111110",
  65150=>"000000000",
  65151=>"111110111",
  65152=>"111011011",
  65153=>"000110111",
  65154=>"111000000",
  65155=>"111101110",
  65156=>"111111111",
  65157=>"111111011",
  65158=>"100110110",
  65159=>"000010000",
  65160=>"001000000",
  65161=>"101000000",
  65162=>"011011011",
  65163=>"001001000",
  65164=>"000000000",
  65165=>"111110000",
  65166=>"111111111",
  65167=>"000000110",
  65168=>"000000000",
  65169=>"111101001",
  65170=>"011001011",
  65171=>"111111111",
  65172=>"000000000",
  65173=>"000000111",
  65174=>"000000000",
  65175=>"111101100",
  65176=>"001000001",
  65177=>"000000000",
  65178=>"000000000",
  65179=>"111000000",
  65180=>"000000111",
  65181=>"001000001",
  65182=>"111111111",
  65183=>"100000001",
  65184=>"000011000",
  65185=>"000011101",
  65186=>"111100111",
  65187=>"111001111",
  65188=>"000000000",
  65189=>"111111000",
  65190=>"111111000",
  65191=>"111111111",
  65192=>"000000000",
  65193=>"111000000",
  65194=>"010111111",
  65195=>"000010000",
  65196=>"011001001",
  65197=>"001100100",
  65198=>"111111111",
  65199=>"111101101",
  65200=>"000000000",
  65201=>"111001000",
  65202=>"011111011",
  65203=>"111111001",
  65204=>"010011111",
  65205=>"111111111",
  65206=>"111111111",
  65207=>"111111111",
  65208=>"110110111",
  65209=>"111111011",
  65210=>"000011000",
  65211=>"111111110",
  65212=>"111111011",
  65213=>"000000100",
  65214=>"000111111",
  65215=>"000000000",
  65216=>"011111111",
  65217=>"111111111",
  65218=>"000100111",
  65219=>"111111111",
  65220=>"000000000",
  65221=>"000000011",
  65222=>"000000000",
  65223=>"111111111",
  65224=>"111111111",
  65225=>"001001001",
  65226=>"000000000",
  65227=>"000000000",
  65228=>"000101101",
  65229=>"111111111",
  65230=>"110001111",
  65231=>"001101001",
  65232=>"111110110",
  65233=>"000000111",
  65234=>"000001111",
  65235=>"000000000",
  65236=>"000110110",
  65237=>"000000000",
  65238=>"111001000",
  65239=>"100000100",
  65240=>"111111111",
  65241=>"000000001",
  65242=>"000000000",
  65243=>"000011111",
  65244=>"101110110",
  65245=>"000110101",
  65246=>"110111111",
  65247=>"000000001",
  65248=>"000000000",
  65249=>"000010000",
  65250=>"100111111",
  65251=>"111111111",
  65252=>"001001001",
  65253=>"111111101",
  65254=>"111111111",
  65255=>"000001011",
  65256=>"000000111",
  65257=>"111100111",
  65258=>"000000101",
  65259=>"111111111",
  65260=>"111111111",
  65261=>"000000000",
  65262=>"011011000",
  65263=>"000001001",
  65264=>"111101101",
  65265=>"000000000",
  65266=>"111111111",
  65267=>"000101101",
  65268=>"000000000",
  65269=>"100100100",
  65270=>"000000000",
  65271=>"000100110",
  65272=>"000000000",
  65273=>"100101111",
  65274=>"000111110",
  65275=>"001000000",
  65276=>"111110000",
  65277=>"000000110",
  65278=>"000000000",
  65279=>"100000000",
  65280=>"000110000",
  65281=>"011001111",
  65282=>"000000000",
  65283=>"011111111",
  65284=>"111111111",
  65285=>"000001011",
  65286=>"000000000",
  65287=>"001000000",
  65288=>"000000000",
  65289=>"000000000",
  65290=>"111000011",
  65291=>"111101001",
  65292=>"111000000",
  65293=>"011000001",
  65294=>"100101111",
  65295=>"110100111",
  65296=>"000000000",
  65297=>"000000001",
  65298=>"010111111",
  65299=>"000000000",
  65300=>"000000011",
  65301=>"000000000",
  65302=>"111111100",
  65303=>"000000000",
  65304=>"111111111",
  65305=>"001101111",
  65306=>"000000100",
  65307=>"111111111",
  65308=>"010111111",
  65309=>"000001111",
  65310=>"110111111",
  65311=>"000000111",
  65312=>"000000000",
  65313=>"000001011",
  65314=>"000000000",
  65315=>"000000101",
  65316=>"111000010",
  65317=>"111111111",
  65318=>"100100100",
  65319=>"000111111",
  65320=>"111111111",
  65321=>"000000000",
  65322=>"000000000",
  65323=>"000000110",
  65324=>"110111111",
  65325=>"000000100",
  65326=>"111111111",
  65327=>"000001001",
  65328=>"000000111",
  65329=>"111111111",
  65330=>"111111111",
  65331=>"111111111",
  65332=>"111111011",
  65333=>"000000111",
  65334=>"000000010",
  65335=>"000000111",
  65336=>"000000000",
  65337=>"000000000",
  65338=>"111100000",
  65339=>"000000000",
  65340=>"011011011",
  65341=>"000000111",
  65342=>"111111111",
  65343=>"111111001",
  65344=>"000010000",
  65345=>"110111111",
  65346=>"000000111",
  65347=>"000100110",
  65348=>"000000000",
  65349=>"000000011",
  65350=>"111111111",
  65351=>"000000000",
  65352=>"111111001",
  65353=>"111111111",
  65354=>"100001001",
  65355=>"011011011",
  65356=>"110110110",
  65357=>"000101111",
  65358=>"000000001",
  65359=>"100001111",
  65360=>"110111111",
  65361=>"010001001",
  65362=>"111111110",
  65363=>"000000011",
  65364=>"001000000",
  65365=>"000000000",
  65366=>"111111111",
  65367=>"000000111",
  65368=>"111111000",
  65369=>"111011000",
  65370=>"111100000",
  65371=>"110111111",
  65372=>"000000000",
  65373=>"111010000",
  65374=>"111111111",
  65375=>"001001101",
  65376=>"000000000",
  65377=>"111111111",
  65378=>"111011011",
  65379=>"110100000",
  65380=>"111111111",
  65381=>"000001101",
  65382=>"000000000",
  65383=>"000000001",
  65384=>"101100100",
  65385=>"001000001",
  65386=>"100111000",
  65387=>"000000000",
  65388=>"100000001",
  65389=>"000001000",
  65390=>"000011111",
  65391=>"011000000",
  65392=>"111100111",
  65393=>"001111111",
  65394=>"000111111",
  65395=>"011010000",
  65396=>"111111111",
  65397=>"101111111",
  65398=>"000000111",
  65399=>"000000011",
  65400=>"000000000",
  65401=>"101011011",
  65402=>"000110110",
  65403=>"111100000",
  65404=>"111111001",
  65405=>"000111111",
  65406=>"000000000",
  65407=>"000000000",
  65408=>"100111111",
  65409=>"110110100",
  65410=>"000000010",
  65411=>"000000000",
  65412=>"101111001",
  65413=>"000000000",
  65414=>"000000000",
  65415=>"000000110",
  65416=>"000000101",
  65417=>"111111111",
  65418=>"100110000",
  65419=>"000000111",
  65420=>"011011000",
  65421=>"111111111",
  65422=>"011000000",
  65423=>"001000000",
  65424=>"111000000",
  65425=>"111111110",
  65426=>"111111111",
  65427=>"101110111",
  65428=>"000100000",
  65429=>"000010000",
  65430=>"110000011",
  65431=>"000000000",
  65432=>"110110000",
  65433=>"101000100",
  65434=>"010000000",
  65435=>"000001110",
  65436=>"001111111",
  65437=>"111111111",
  65438=>"000000000",
  65439=>"010111111",
  65440=>"001110111",
  65441=>"110111111",
  65442=>"000000000",
  65443=>"000000000",
  65444=>"111101111",
  65445=>"111111111",
  65446=>"110110111",
  65447=>"000010111",
  65448=>"110000100",
  65449=>"111111001",
  65450=>"000000100",
  65451=>"000000000",
  65452=>"000000000",
  65453=>"110110111",
  65454=>"100000001",
  65455=>"000000001",
  65456=>"000000000",
  65457=>"000000000",
  65458=>"011111111",
  65459=>"001111111",
  65460=>"000101111",
  65461=>"000000000",
  65462=>"111111111",
  65463=>"000000001",
  65464=>"000000111",
  65465=>"000100000",
  65466=>"010000000",
  65467=>"000100111",
  65468=>"000110010",
  65469=>"111111101",
  65470=>"001000000",
  65471=>"111111111",
  65472=>"000000110",
  65473=>"111001001",
  65474=>"010011011",
  65475=>"111111111",
  65476=>"110010110",
  65477=>"111001001",
  65478=>"000000000",
  65479=>"000000000",
  65480=>"000000000",
  65481=>"000000000",
  65482=>"000000001",
  65483=>"000100101",
  65484=>"111111110",
  65485=>"000000000",
  65486=>"000000000",
  65487=>"000000100",
  65488=>"111100001",
  65489=>"101111111",
  65490=>"001001101",
  65491=>"010110110",
  65492=>"111111111",
  65493=>"101000101",
  65494=>"000000000",
  65495=>"000000000",
  65496=>"000000001",
  65497=>"111010000",
  65498=>"000000111",
  65499=>"111111101",
  65500=>"000000001",
  65501=>"000001000",
  65502=>"000000111",
  65503=>"001001001",
  65504=>"000000000",
  65505=>"000000000",
  65506=>"000000000",
  65507=>"000110000",
  65508=>"111111111",
  65509=>"000000100",
  65510=>"111110000",
  65511=>"000100111",
  65512=>"000000100",
  65513=>"001000000",
  65514=>"011111111",
  65515=>"110101101",
  65516=>"000000001",
  65517=>"111011001",
  65518=>"011000000",
  65519=>"111111111",
  65520=>"101000000",
  65521=>"111011011",
  65522=>"000000000",
  65523=>"000001001",
  65524=>"000000000",
  65525=>"000000000",
  65526=>"011001000",
  65527=>"001001100",
  65528=>"110111111",
  65529=>"100101001",
  65530=>"111111100",
  65531=>"111010000",
  65532=>"111111011",
  65533=>"110110111",
  65534=>"000001111",
  65535=>"000000000");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;