LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L3_1_WROM IS
    PORT (
        weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
        address : IN unsigned(weightsbitsAddress(3)-1 DOWNTO 0));
END L3_1_WROM;

ARCHITECTURE RTL OF L3_1_WROM IS

    TYPE ROM_mem IS ARRAY (0 TO 1023) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

    CONSTANT ROM_content : ROM_mem := (0=>"100110110",
    1=>"000110110",
    2=>"011011011",
    3=>"100100100",
    4=>"010111111",
    5=>"001001010",
    6=>"110110110",
    7=>"011010010",
    8=>"110010110",
    9=>"011001010",
    10=>"010011011",
    11=>"001001010",
    12=>"000010000",
    13=>"000100101",
    14=>"001001001",
    15=>"010110110",
    16=>"110110110",
    17=>"101101001",
    18=>"100001011",
    19=>"001111010",
    20=>"001001001",
    21=>"110110110",
    22=>"110110100",
    23=>"001101001",
    24=>"001001011",
    25=>"100100101",
    26=>"001001011",
    27=>"100100000",
    28=>"011000011",
    29=>"110110110",
    30=>"001000011",
    31=>"011011011",
    32=>"100100111",
    33=>"000100101",
    34=>"111000000",
    35=>"000000111",
    36=>"000111011",
    37=>"000111100",
    38=>"101111111",
    39=>"000100110",
    40=>"111000000",
    41=>"000000001",
    42=>"010000111",
    43=>"101000000",
    44=>"000001000",
    45=>"100001000",
    46=>"011001111",
    47=>"001011101",
    48=>"110010000",
    49=>"000111111",
    50=>"001101100",
    51=>"111000000",
    52=>"100000111",
    53=>"000111111",
    54=>"101111100",
    55=>"110001000",
    56=>"100001111",
    57=>"111100000",
    58=>"000111111",
    59=>"000010000",
    60=>"001100010",
    61=>"010000010",
    62=>"111010111",
    63=>"101001001",
    64=>"011001001",
    65=>"001011011",
    66=>"100100100",
    67=>"100101101",
    68=>"111001001",
    69=>"011011000",
    70=>"111101111",
    71=>"100100111",
    72=>"011001001",
    73=>"100100100",
    74=>"101111111",
    75=>"000000100",
    76=>"000000000",
    77=>"011000000",
    78=>"100110110",
    79=>"001101011",
    80=>"111111001",
    81=>"010001010",
    82=>"110000100",
    83=>"011011011",
    84=>"001001001",
    85=>"101100100",
    86=>"101111111",
    87=>"000100100",
    88=>"001001011",
    89=>"010010011",
    90=>"011011001",
    91=>"000000000",
    92=>"010011011",
    93=>"011001101",
    94=>"000100110",
    95=>"110101001",
    96=>"000000000",
    97=>"000010000",
    98=>"001101111",
    99=>"010000010",
    100=>"010111111",
    101=>"000000000",
    102=>"100100100",
    103=>"100100000",
    104=>"010101000",
    105=>"000110000",
    106=>"010110011",
    107=>"000111000",
    108=>"001001000",
    109=>"100101011",
    110=>"000111011",
    111=>"011011100",
    112=>"010101110",
    113=>"000010010",
    114=>"010110000",
    115=>"110111000",
    116=>"000100000",
    117=>"000110011",
    118=>"000000000",
    119=>"001100000",
    120=>"110000000",
    121=>"000001101",
    122=>"101111111",
    123=>"011011000",
    124=>"011011110",
    125=>"000000100",
    126=>"111000111",
    127=>"000000000",
    128=>"100101111",
    129=>"100101100",
    130=>"000000001",
    131=>"000000000",
    132=>"111101000",
    133=>"000001001",
    134=>"110111111",
    135=>"000100111",
    136=>"001000000",
    137=>"000100100",
    138=>"001000011",
    139=>"100100110",
    140=>"101001111",
    141=>"100000100",
    142=>"000000000",
    143=>"011111110",
    144=>"001101101",
    145=>"000100100",
    146=>"010000000",
    147=>"111111111",
    148=>"010001000",
    149=>"000000000",
    150=>"100101111",
    151=>"000000100",
    152=>"111110000",
    153=>"110111111",
    154=>"111111111",
    155=>"010111111",
    156=>"000000000",
    157=>"001111111",
    158=>"001001111",
    159=>"111110000",
    160=>"000111111",
    161=>"000000111",
    162=>"001001000",
    163=>"111110111",
    164=>"001001001",
    165=>"110011001",
    166=>"000111111",
    167=>"000110110",
    168=>"010111011",
    169=>"111001000",
    170=>"000000000",
    171=>"011001000",
    172=>"011000000",
    173=>"111110100",
    174=>"000110010",
    175=>"110111111",
    176=>"011011001",
    177=>"111100100",
    178=>"000000100",
    179=>"110111011",
    180=>"011001001",
    181=>"100110111",
    182=>"111111111",
    183=>"011000000",
    184=>"011000100",
    185=>"110110111",
    186=>"000000000",
    187=>"110110111",
    188=>"111011000",
    189=>"000111011",
    190=>"111000000",
    191=>"111001000",
    192=>"011100001",
    193=>"100101000",
    194=>"011100000",
    195=>"100101011",
    196=>"000001110",
    197=>"000111110",
    198=>"111111000",
    199=>"111111100",
    200=>"000111100",
    201=>"100001111",
    202=>"000111100",
    203=>"000110100",
    204=>"000001000",
    205=>"100001111",
    206=>"000001111",
    207=>"011001000",
    208=>"001111100",
    209=>"110000011",
    210=>"000011110",
    211=>"000011110",
    212=>"001110000",
    213=>"011100000",
    214=>"000000011",
    215=>"000000111",
    216=>"001110100",
    217=>"110000011",
    218=>"011110000",
    219=>"000000001",
    220=>"111000111",
    221=>"011110000",
    222=>"000011110",
    223=>"011100110",
    224=>"101001001",
    225=>"101101100",
    226=>"011100011",
    227=>"000000000",
    228=>"110000101",
    229=>"100100110",
    230=>"111000000",
    231=>"111101001",
    232=>"100000000",
    233=>"010110110",
    234=>"111111111",
    235=>"100000001",
    236=>"101000001",
    237=>"000000000",
    238=>"111111111",
    239=>"000001011",
    240=>"101001011",
    241=>"011010110",
    242=>"110101000",
    243=>"000000000",
    244=>"110101101",
    245=>"000000001",
    246=>"100001001",
    247=>"111110110",
    248=>"111111111",
    249=>"000110100",
    250=>"111110100",
    251=>"000000001",
    252=>"010100111",
    253=>"101001001",
    254=>"000111111",
    255=>"110110110",
    256=>"111001000",
    257=>"000101111",
    258=>"100110111",
    259=>"011000100",
    260=>"000000000",
    261=>"100100111",
    262=>"100111011",
    263=>"001001111",
    264=>"110111011",
    265=>"011001100",
    266=>"111111111",
    267=>"001001000",
    268=>"011000000",
    269=>"011111101",
    270=>"011001100",
    271=>"111001001",
    272=>"000000000",
    273=>"000011001",
    274=>"001100110",
    275=>"100110111",
    276=>"001000000",
    277=>"011001100",
    278=>"111101101",
    279=>"111100100",
    280=>"100110111",
    281=>"100110011",
    282=>"000110011",
    283=>"000100110",
    284=>"100110111",
    285=>"001000010",
    286=>"000000111",
    287=>"111001010",
    288=>"000101001",
    289=>"100101100",
    290=>"001000000",
    291=>"000000000",
    292=>"001101111",
    293=>"000101001",
    294=>"100000111",
    295=>"101101101",
    296=>"111111101",
    297=>"001101101",
    298=>"000000100",
    299=>"000000000",
    300=>"101001000",
    301=>"011001011",
    302=>"000000000",
    303=>"000100111",
    304=>"011010111",
    305=>"101000111",
    306=>"000101101",
    307=>"111101101",
    308=>"000001101",
    309=>"011111111",
    310=>"000000000",
    311=>"000000011",
    312=>"100100010",
    313=>"000000100",
    314=>"000100100",
    315=>"101000010",
    316=>"010001110",
    317=>"101100101",
    318=>"000000010",
    319=>"111111111",
    320=>"100001011",
    321=>"100001011",
    322=>"011010001",
    323=>"110111111",
    324=>"110000000",
    325=>"100101111",
    326=>"011111111",
    327=>"001001011",
    328=>"111111000",
    329=>"110100111",
    330=>"100110110",
    331=>"000001001",
    332=>"100100000",
    333=>"011111110",
    334=>"011111111",
    335=>"011001011",
    336=>"000111011",
    337=>"000001001",
    338=>"111100010",
    339=>"111111111",
    340=>"100000000",
    341=>"000000000",
    342=>"001001001",
    343=>"011110110",
    344=>"100001000",
    345=>"000000000",
    346=>"100000001",
    347=>"110111110",
    348=>"000000000",
    349=>"100000100",
    350=>"110111111",
    351=>"111000010",
    352=>"011001001",
    353=>"100100110",
    354=>"000000000",
    355=>"110110110",
    356=>"001000100",
    357=>"000100110",
    358=>"110110001",
    359=>"011011001",
    360=>"100110100",
    361=>"011011001",
    362=>"010011110",
    363=>"011011001",
    364=>"001001101",
    365=>"010000010",
    366=>"101101111",
    367=>"101100101",
    368=>"000110111",
    369=>"011000110",
    370=>"110011000",
    371=>"100000100",
    372=>"100100110",
    373=>"111011000",
    374=>"001000001",
    375=>"011010010",
    376=>"111101111",
    377=>"111001111",
    378=>"000101100",
    379=>"011111001",
    380=>"100110110",
    381=>"001100101",
    382=>"010011010",
    383=>"001101100",
    384=>"000010010",
    385=>"000011000",
    386=>"100100000",
    387=>"001011110",
    388=>"111111011",
    389=>"000010010",
    390=>"001011101",
    391=>"000011000",
    392=>"110000000",
    393=>"010111000",
    394=>"000010000",
    395=>"000110000",
    396=>"010010000",
    397=>"010010010",
    398=>"001011000",
    399=>"010110010",
    400=>"000011000",
    401=>"010010010",
    402=>"000011000",
    403=>"111011010",
    404=>"000011000",
    405=>"000011000",
    406=>"010010010",
    407=>"000110000",
    408=>"000010011",
    409=>"001111000",
    410=>"100110001",
    411=>"000000010",
    412=>"100011001",
    413=>"000101001",
    414=>"111010111",
    415=>"000111010",
    416=>"111010010",
    417=>"010001011",
    418=>"100000010",
    419=>"001001100",
    420=>"111000011",
    421=>"001000011",
    422=>"111000111",
    423=>"010011001",
    424=>"011010000",
    425=>"000111001",
    426=>"110010011",
    427=>"110001000",
    428=>"000000000",
    429=>"011101100",
    430=>"111000111",
    431=>"000000110",
    432=>"010010110",
    433=>"101101101",
    434=>"011011000",
    435=>"101000011",
    436=>"000010010",
    437=>"111000000",
    438=>"101000101",
    439=>"000111000",
    440=>"100111011",
    441=>"011001100",
    442=>"110100001",
    443=>"011000100",
    444=>"000111000",
    445=>"110000111",
    446=>"000111001",
    447=>"000111011",
    448=>"100100110",
    449=>"011001001",
    450=>"010111001",
    451=>"110011011",
    452=>"001000000",
    453=>"011001000",
    454=>"110001101",
    455=>"100110110",
    456=>"111111000",
    457=>"100110110",
    458=>"111111111",
    459=>"001100100",
    460=>"000100100",
    461=>"010000010",
    462=>"101100011",
    463=>"111001101",
    464=>"010001110",
    465=>"010010010",
    466=>"111011001",
    467=>"111110000",
    468=>"011111010",
    469=>"111011010",
    470=>"011000100",
    471=>"001110000",
    472=>"011111110",
    473=>"101101111",
    474=>"000100100",
    475=>"111011011",
    476=>"011011101",
    477=>"100101100",
    478=>"000000110",
    479=>"010010000",
    480=>"100100110",
    481=>"101101000",
    482=>"111111101",
    483=>"111111111",
    484=>"000000001",
    485=>"101111111",
    486=>"111000100",
    487=>"101111001",
    488=>"000000000",
    489=>"111101001",
    490=>"111111111",
    491=>"101001000",
    492=>"110000000",
    493=>"111111111",
    494=>"110101001",
    495=>"011101110",
    496=>"000000000",
    497=>"100000100",
    498=>"111000000",
    499=>"100101011",
    500=>"100001011",
    501=>"100011101",
    502=>"001101101",
    503=>"000000000",
    504=>"111111111",
    505=>"001100110",
    506=>"101011010",
    507=>"011101110",
    508=>"001000000",
    509=>"000000000",
    510=>"000000000",
    511=>"110111001",
    512=>"100001111",
    513=>"000101101",
    514=>"011100100",
    515=>"110001000",
    516=>"100111000",
    517=>"111011000",
    518=>"111000000",
    519=>"110110101",
    520=>"101111000",
    521=>"010000111",
    522=>"111110000",
    523=>"100000000",
    524=>"000001000",
    525=>"001000001",
    526=>"111100110",
    527=>"111001001",
    528=>"111001000",
    529=>"000110111",
    530=>"110111000",
    531=>"010000010",
    532=>"111000010",
    533=>"111000000",
    534=>"000111111",
    535=>"000111111",
    536=>"100110111",
    537=>"111001101",
    538=>"111111010",
    539=>"111001000",
    540=>"000111111",
    541=>"111000000",
    542=>"000111111",
    543=>"000000110",
    544=>"010010010",
    545=>"010000010",
    546=>"100010011",
    547=>"001000101",
    548=>"111010100",
    549=>"011000010",
    550=>"111111000",
    551=>"010010011",
    552=>"111000000",
    553=>"000010010",
    554=>"111111111",
    555=>"000000011",
    556=>"000000001",
    557=>"011011111",
    558=>"000000011",
    559=>"011001000",
    560=>"011011001",
    561=>"001000100",
    562=>"110110011",
    563=>"111111111",
    564=>"000000011",
    565=>"111111110",
    566=>"010000111",
    567=>"000000000",
    568=>"001111111",
    569=>"000010000",
    570=>"100000100",
    571=>"111111111",
    572=>"000000000",
    573=>"101101000",
    574=>"000000000",
    575=>"010101111",
    576=>"100100100",
    577=>"010011001",
    578=>"101100110",
    579=>"011001001",
    580=>"100110110",
    581=>"010001001",
    582=>"101110110",
    583=>"000011001",
    584=>"110010000",
    585=>"010000001",
    586=>"100110111",
    587=>"010010000",
    588=>"001100000",
    589=>"011011000",
    590=>"001001100",
    591=>"110010001",
    592=>"100110110",
    593=>"011001100",
    594=>"011001001",
    595=>"010010010",
    596=>"000001011",
    597=>"001001001",
    598=>"100100110",
    599=>"011101100",
    600=>"100100111",
    601=>"110011001",
    602=>"100110111",
    603=>"110001000",
    604=>"011000001",
    605=>"100110010",
    606=>"010000001",
    607=>"011011011",
    608=>"000100101",
    609=>"001100001",
    610=>"011100000",
    611=>"100001111",
    612=>"001110100",
    613=>"001110100",
    614=>"100011010",
    615=>"000110001",
    616=>"001011100",
    617=>"001110000",
    618=>"111110000",
    619=>"011100000",
    620=>"001000000",
    621=>"101001111",
    622=>"111000001",
    623=>"010010101",
    624=>"000100000",
    625=>"100001111",
    626=>"011110000",
    627=>"110100011",
    628=>"111100000",
    629=>"001011110",
    630=>"110000001",
    631=>"100000110",
    632=>"000100100",
    633=>"100001111",
    634=>"010110100",
    635=>"000001100",
    636=>"000011110",
    637=>"010110010",
    638=>"000001101",
    639=>"011100001",
    640=>"011011010",
    641=>"011001011",
    642=>"000011011",
    643=>"000100100",
    644=>"110011010",
    645=>"100100111",
    646=>"111011001",
    647=>"000100110",
    648=>"101101110",
    649=>"001100011",
    650=>"110111001",
    651=>"000000011",
    652=>"000000000",
    653=>"100110010",
    654=>"100100110",
    655=>"010011000",
    656=>"101101010",
    657=>"111011000",
    658=>"100111111",
    659=>"001010011",
    660=>"100100100",
    661=>"000110110",
    662=>"011011011",
    663=>"100011000",
    664=>"000011001",
    665=>"101110010",
    666=>"010000000",
    667=>"000100110",
    668=>"000111111",
    669=>"010010011",
    670=>"000011000",
    671=>"000100110",
    672=>"000010010",
    673=>"011011111",
    674=>"000000011",
    675=>"111111111",
    676=>"111110111",
    677=>"011101101",
    678=>"001000000",
    679=>"000111111",
    680=>"000000010",
    681=>"010111011",
    682=>"110100011",
    683=>"111111011",
    684=>"111111111",
    685=>"000000010",
    686=>"100110111",
    687=>"100111011",
    688=>"000000000",
    689=>"100010110",
    690=>"111111101",
    691=>"111111001",
    692=>"011001001",
    693=>"111111111",
    694=>"000000100",
    695=>"000111111",
    696=>"101110110",
    697=>"010011101",
    698=>"111111001",
    699=>"000000000",
    700=>"000100001",
    701=>"001011100",
    702=>"110011111",
    703=>"110111011",
    704=>"011111101",
    705=>"101100101",
    706=>"001000001",
    707=>"000000000",
    708=>"101100000",
    709=>"101100100",
    710=>"111111111",
    711=>"100101001",
    712=>"111000110",
    713=>"101101001",
    714=>"001010010",
    715=>"100100000",
    716=>"100000000",
    717=>"000000000",
    718=>"001000000",
    719=>"001001001",
    720=>"001011111",
    721=>"111011011",
    722=>"100100101",
    723=>"000000111",
    724=>"001000001",
    725=>"101111000",
    726=>"001000001",
    727=>"000000100",
    728=>"000000000",
    729=>"100000100",
    730=>"100000000",
    731=>"000110111",
    732=>"001001000",
    733=>"010010111",
    734=>"001000000",
    735=>"110100100",
    736=>"000000111",
    737=>"111100000",
    738=>"110000001",
    739=>"111101001",
    740=>"111111011",
    741=>"111000000",
    742=>"111100000",
    743=>"000000111",
    744=>"101101001",
    745=>"000010111",
    746=>"010110010",
    747=>"000001111",
    748=>"010001011",
    749=>"101011111",
    750=>"011111101",
    751=>"000000111",
    752=>"100000100",
    753=>"111000001",
    754=>"001010100",
    755=>"111101111",
    756=>"001000110",
    757=>"100000001",
    758=>"001000001",
    759=>"100000000",
    760=>"010111111",
    761=>"000011000",
    762=>"111110010",
    763=>"100110101",
    764=>"001000001",
    765=>"100001001",
    766=>"000011101",
    767=>"100000011",
    768=>"001101101",
    769=>"101100100",
    770=>"000000000",
    771=>"100000100",
    772=>"101111101",
    773=>"111010110",
    774=>"101101101",
    775=>"101100111",
    776=>"111111111",
    777=>"000000011",
    778=>"000000000",
    779=>"101100111",
    780=>"000000000",
    781=>"000000000",
    782=>"111100111",
    783=>"000110000",
    784=>"111111111",
    785=>"111000011",
    786=>"001000100",
    787=>"111001100",
    788=>"011111101",
    789=>"100111101",
    790=>"001000101",
    791=>"111000111",
    792=>"000000000",
    793=>"111001111",
    794=>"011011011",
    795=>"000000000",
    796=>"111000111",
    797=>"101101100",
    798=>"110111111",
    799=>"111000111",
    800=>"010010010",
    801=>"010010011",
    802=>"111110001",
    803=>"000000000",
    804=>"000001000",
    805=>"010011011",
    806=>"100100101",
    807=>"000011111",
    808=>"000000000",
    809=>"000011111",
    810=>"001000001",
    811=>"000000001",
    812=>"010000010",
    813=>"101100000",
    814=>"111111111",
    815=>"110111111",
    816=>"110100000",
    817=>"111100000",
    818=>"001001011",
    819=>"100100000",
    820=>"010000100",
    821=>"011001001",
    822=>"111100000",
    823=>"111100001",
    824=>"000000000",
    825=>"011111111",
    826=>"111110101",
    827=>"010001100",
    828=>"111011011",
    829=>"000101000",
    830=>"111100110",
    831=>"011111111",
    832=>"011110011",
    833=>"011110000",
    834=>"111111111",
    835=>"000000000",
    836=>"011111110",
    837=>"000010001",
    838=>"000111111",
    839=>"011010000",
    840=>"011011111",
    841=>"010000011",
    842=>"011111111",
    843=>"111000001",
    844=>"110000000",
    845=>"100000000",
    846=>"000011111",
    847=>"010100000",
    848=>"100101101",
    849=>"111000000",
    850=>"010000001",
    851=>"111111111",
    852=>"010110101",
    853=>"000001011",
    854=>"111110000",
    855=>"111100000",
    856=>"011011111",
    857=>"000000000",
    858=>"001011111",
    859=>"000000000",
    860=>"111000001",
    861=>"000111111",
    862=>"110000001",
    863=>"111000000",
    864=>"001001001",
    865=>"000001011",
    866=>"011011101",
    867=>"100111010",
    868=>"000111000",
    869=>"111100000",
    870=>"011110100",
    871=>"000011011",
    872=>"101100101",
    873=>"111100100",
    874=>"001111100",
    875=>"111010000",
    876=>"001111000",
    877=>"001111100",
    878=>"000100100",
    879=>"000000101",
    880=>"111110000",
    881=>"111100100",
    882=>"000111110",
    883=>"000000111",
    884=>"000001111",
    885=>"000000001",
    886=>"001011011",
    887=>"011100010",
    888=>"110111110",
    889=>"100101001",
    890=>"100100101",
    891=>"010101110",
    892=>"111110000",
    893=>"100101100",
    894=>"010110100",
    895=>"011001011",
    896=>"010000000",
    897=>"000000000",
    898=>"000001001",
    899=>"011111111",
    900=>"000000101",
    901=>"000000000",
    902=>"000010010",
    903=>"010000000",
    904=>"111000000",
    905=>"010111000",
    906=>"100011001",
    907=>"000000000",
    908=>"011111101",
    909=>"111110011",
    910=>"110110011",
    911=>"000110000",
    912=>"010100001",
    913=>"000011010",
    914=>"111111111",
    915=>"000000111",
    916=>"011111111",
    917=>"010110110",
    918=>"001000101",
    919=>"100110011",
    920=>"111011010",
    921=>"000100110",
    922=>"111011110",
    923=>"101000000",
    924=>"010011000",
    925=>"010011111",
    926=>"000101100",
    927=>"111011000",
    928=>"101100101",
    929=>"101000101",
    930=>"000000000",
    931=>"001101100",
    932=>"000000000",
    933=>"111001001",
    934=>"100000111",
    935=>"101000100",
    936=>"111000000",
    937=>"101000100",
    938=>"111111111",
    939=>"001000000",
    940=>"001000000",
    941=>"110010011",
    942=>"001001000",
    943=>"001000001",
    944=>"100111111",
    945=>"001000101",
    946=>"111101101",
    947=>"000000000",
    948=>"000000000",
    949=>"001000000",
    950=>"111111111",
    951=>"100100100",
    952=>"110110110",
    953=>"101101101",
    954=>"100000000",
    955=>"101101011",
    956=>"011001001",
    957=>"010010010",
    958=>"111111111",
    959=>"001000001",
    960=>"010000101",
    961=>"000000110",
    962=>"011100100",
    963=>"000111001",
    964=>"011100010",
    965=>"000110011",
    966=>"000111110",
    967=>"000100111",
    968=>"011110011",
    969=>"011000111",
    970=>"000001000",
    971=>"000000111",
    972=>"000000001",
    973=>"100000000",
    974=>"111111000",
    975=>"000100011",
    976=>"000110011",
    977=>"111001100",
    978=>"111101000",
    979=>"001000111",
    980=>"000011001",
    981=>"100111000",
    982=>"001000111",
    983=>"111001100",
    984=>"111001100",
    985=>"001000111",
    986=>"001000111",
    987=>"000111011",
    988=>"100000111",
    989=>"000111001",
    990=>"000001001",
    991=>"110001111",
    992=>"011001111",
    993=>"000100010",
    994=>"110110001",
    995=>"001100110",
    996=>"000000000",
    997=>"011001110",
    998=>"000000011",
    999=>"000001111",
    1000=>"111011111",
    1001=>"100000000",
    1002=>"111001001",
    1003=>"000000000",
    1004=>"111111010",
    1005=>"011111110",
    1006=>"010001001",
    1007=>"100110110",
    1008=>"010010010",
    1009=>"000001110",
    1010=>"011001011",
    1011=>"000011010",
    1012=>"111111111",
    1013=>"111111000",
    1014=>"100100111",
    1015=>"111111001",
    1016=>"110000001",
    1017=>"101110110",
    1018=>"110100111",
    1019=>"011101011",
    1020=>"001011100",
    1021=>"011000011",
    1022=>"101110011",
    1023=>"111111011");

BEGIN
    weight <= ROM_content(to_integer(address));
END RTL;