LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_1_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    address : IN unsigned(5 DOWNTO 0));
END L8_1_BNROM;

ARCHITECTURE RTL OF L8_1_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 63) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  --Contenido bias || scale
  (0=>"0010000111011100"&"0010000100010011",
  1=>"0000111000100011"&"0010001101010101",
  2=>"0010100000101011"&"0001111101111000",
  3=>"0001001111000001"&"0010000100101000",
  4=>"0001000001011010"&"0010010001101111",
  5=>"0001101101111011"&"0010001101000001",
  6=>"0000101011000110"&"0001110001110011",
  7=>"0001101101010001"&"0010010000100101",
  8=>"0001101010010100"&"0010001101101111",
  9=>"0010100100010100"&"0010100010101101",
  10=>"0000111100011011"&"0010001010011010",
  11=>"0001100001101011"&"0010001001100101",
  12=>"0001011000011011"&"0010010010010101",
  13=>"0000110011101111"&"0001111001011000",
  14=>"0010011111100101"&"0010000111001100",
  15=>"0001100100000001"&"0010010010101101",
  16=>"0010000001000010"&"0010010101101010",
  17=>"0001000010101111"&"0010010101011111",
  18=>"0001111110101100"&"0010010110111101",
  19=>"0010000100110000"&"0010010101100011",
  20=>"0001010100101110"&"0010101000011001",
  21=>"0010000011011010"&"0010001001111110",
  22=>"0001100010010111"&"0010001001011010",
  23=>"0001010111010110"&"0010001010101001",
  24=>"0001110110000010"&"0010001101100111",
  25=>"0000010000111011"&"0010000110110101",
  26=>"0001111111010101"&"0010001100111001",
  27=>"0010001010011100"&"0010000000111101",
  28=>"0000111101010100"&"0001110011001010",
  29=>"0000111100010101"&"0010000101100011",
  30=>"0000111110110000"&"0010001001100101",
  31=>"1111010110001101"&"0010000101110101",
  32=>"0000110011001011"&"0010011100100111",
  33=>"0001000011001011"&"0010000001001110",
  34=>"0000011001000000"&"0010010100101101",
  35=>"0000000110111100"&"0001110111011011",
  36=>"0000010011001111"&"0001111101111100",
  37=>"0010100010110000"&"0010010000110110",
  38=>"0001100011000001"&"0010001101100011",
  39=>"0000100001001010"&"0010000011010011",
  40=>"0001001101101100"&"0010001011011000",
  41=>"0001101111011100"&"0010001111111001",
  42=>"0001000111010001"&"0010010001011011",
  43=>"0001001110001000"&"0010001100001111",
  44=>"0010101100111110"&"0010000011011100",
  45=>"0000101010000100"&"0001011111000010",
  46=>"0010000110011111"&"0001110101100101",
  47=>"0010100001110110"&"0010001000010101",
  48=>"0010101111011011"&"0001111100101011",
  49=>"0001111000010101"&"0010001110001000",
  50=>"0001011010010111"&"0010011100001010",
  51=>"0001111011101111"&"0010001011101010",
  52=>"0001011101101010"&"0001100100110100",
  53=>"0001000111001110"&"0010010101100101",
  54=>"0010001111100010"&"0001100101100111",
  55=>"0001011100011111"&"0010001100000101",
  56=>"0001001011111001"&"0010100010111110",
  57=>"0010000010101100"&"0010001011000111",
  58=>"0001100100010000"&"0010001100100011",
  59=>"0001000111000111"&"0010001100001101",
  60=>"0010010101101111"&"0010001000011010",
  61=>"0000110011111001"&"0001110101110001",
  62=>"0001010100100110"&"0010010001010010",
  63=>"0010001001110110"&"0010000100101001");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;