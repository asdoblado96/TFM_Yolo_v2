LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L7_1_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(7) - 1 DOWNTO 0));
END L7_1_WROM;

ARCHITECTURE RTL OF L7_1_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"000011011",
  1=>"001001101",
  2=>"000000111",
  3=>"000000000",
  4=>"011001000",
  5=>"000111111",
  6=>"000000000",
  7=>"111111111",
  8=>"101101111",
  9=>"111111111",
  10=>"001001000",
  11=>"111111110",
  12=>"000110000",
  13=>"100000000",
  14=>"101001001",
  15=>"000001011",
  16=>"000000011",
  17=>"110101111",
  18=>"111010001",
  19=>"000000000",
  20=>"000000000",
  21=>"110000000",
  22=>"000000011",
  23=>"011001000",
  24=>"111111111",
  25=>"000000110",
  26=>"000011000",
  27=>"000100111",
  28=>"111111001",
  29=>"111110100",
  30=>"011000100",
  31=>"111000000",
  32=>"110110000",
  33=>"000111111",
  34=>"001000000",
  35=>"000100100",
  36=>"000000101",
  37=>"101111110",
  38=>"000000111",
  39=>"111001000",
  40=>"000000011",
  41=>"000000000",
  42=>"000111111",
  43=>"000111001",
  44=>"110000000",
  45=>"110000000",
  46=>"000000000",
  47=>"000000000",
  48=>"000010110",
  49=>"000010110",
  50=>"010000000",
  51=>"000000000",
  52=>"111100000",
  53=>"111011011",
  54=>"000111101",
  55=>"000000000",
  56=>"111001000",
  57=>"000010011",
  58=>"000000000",
  59=>"111111110",
  60=>"001001111",
  61=>"111101111",
  62=>"100110110",
  63=>"000000000",
  64=>"100100100",
  65=>"111111110",
  66=>"000111110",
  67=>"111111111",
  68=>"111110010",
  69=>"011111100",
  70=>"000000000",
  71=>"000000001",
  72=>"100111111",
  73=>"101000000",
  74=>"100100100",
  75=>"110100000",
  76=>"000000001",
  77=>"001101111",
  78=>"000001111",
  79=>"001111111",
  80=>"111011000",
  81=>"111011001",
  82=>"111111111",
  83=>"010110110",
  84=>"111000000",
  85=>"100000000",
  86=>"000111111",
  87=>"111111111",
  88=>"101000000",
  89=>"000101111",
  90=>"100000111",
  91=>"010000100",
  92=>"110010000",
  93=>"111111111",
  94=>"100100111",
  95=>"100100101",
  96=>"000000000",
  97=>"101000100",
  98=>"000000111",
  99=>"000111111",
  100=>"000000000",
  101=>"000000000",
  102=>"101000000",
  103=>"111111101",
  104=>"111100000",
  105=>"111100111",
  106=>"000000011",
  107=>"001001001",
  108=>"010111111",
  109=>"000000000",
  110=>"111111111",
  111=>"111111111",
  112=>"000000000",
  113=>"000000000",
  114=>"111111111",
  115=>"100000000",
  116=>"101000000",
  117=>"000000000",
  118=>"111000000",
  119=>"000000000",
  120=>"100111111",
  121=>"000100000",
  122=>"000000100",
  123=>"001000000",
  124=>"011111111",
  125=>"000100000",
  126=>"100100110",
  127=>"001100111",
  128=>"000000000",
  129=>"110111101",
  130=>"011111111",
  131=>"000111111",
  132=>"111111111",
  133=>"111000111",
  134=>"110110110",
  135=>"011111000",
  136=>"000110111",
  137=>"000000000",
  138=>"111110100",
  139=>"101001000",
  140=>"111100000",
  141=>"111100000",
  142=>"100100000",
  143=>"000000000",
  144=>"011011010",
  145=>"111100101",
  146=>"111110111",
  147=>"000111111",
  148=>"000000010",
  149=>"110111111",
  150=>"101111011",
  151=>"111111111",
  152=>"000000001",
  153=>"111111000",
  154=>"010000111",
  155=>"000111000",
  156=>"000000100",
  157=>"010110111",
  158=>"111111111",
  159=>"000000001",
  160=>"000000111",
  161=>"111111111",
  162=>"110110010",
  163=>"000000000",
  164=>"000110000",
  165=>"010000001",
  166=>"000010110",
  167=>"001111100",
  168=>"011111000",
  169=>"000111111",
  170=>"111101000",
  171=>"111110110",
  172=>"011000001",
  173=>"100110000",
  174=>"011111111",
  175=>"101111110",
  176=>"000000000",
  177=>"111111111",
  178=>"111111111",
  179=>"110000111",
  180=>"000000000",
  181=>"111111011",
  182=>"111111111",
  183=>"000111111",
  184=>"000011111",
  185=>"111111111",
  186=>"000011111",
  187=>"111111111",
  188=>"000000100",
  189=>"000000000",
  190=>"000110111",
  191=>"111111001",
  192=>"000000000",
  193=>"000000101",
  194=>"111111111",
  195=>"111111111",
  196=>"111111110",
  197=>"000111111",
  198=>"000000000",
  199=>"111111111",
  200=>"000000000",
  201=>"000100111",
  202=>"000000110",
  203=>"000000000",
  204=>"011111111",
  205=>"001001000",
  206=>"110000000",
  207=>"000000000",
  208=>"000111111",
  209=>"000000001",
  210=>"000010011",
  211=>"000000100",
  212=>"000000000",
  213=>"010001000",
  214=>"000000111",
  215=>"110111111",
  216=>"000001000",
  217=>"100101111",
  218=>"000100111",
  219=>"000000000",
  220=>"111111111",
  221=>"001000100",
  222=>"111000000",
  223=>"001011111",
  224=>"000000001",
  225=>"101000000",
  226=>"111101000",
  227=>"000000000",
  228=>"100000000",
  229=>"000000011",
  230=>"100110110",
  231=>"110110110",
  232=>"111000000",
  233=>"000100111",
  234=>"111111111",
  235=>"000000110",
  236=>"011000000",
  237=>"111000111",
  238=>"111111001",
  239=>"111001001",
  240=>"011011010",
  241=>"000111001",
  242=>"000000000",
  243=>"111000000",
  244=>"111111000",
  245=>"111001111",
  246=>"001111110",
  247=>"111111111",
  248=>"101111000",
  249=>"100001111",
  250=>"000000111",
  251=>"111111111",
  252=>"101001001",
  253=>"111000000",
  254=>"111111110",
  255=>"111111000",
  256=>"000000000",
  257=>"000110110",
  258=>"110000000",
  259=>"111111000",
  260=>"000110000",
  261=>"011001111",
  262=>"111111111",
  263=>"000000111",
  264=>"000111111",
  265=>"111111111",
  266=>"100000000",
  267=>"000100111",
  268=>"111111111",
  269=>"111000001",
  270=>"111111111",
  271=>"000000000",
  272=>"000000000",
  273=>"000000000",
  274=>"111010010",
  275=>"000000000",
  276=>"000000000",
  277=>"000000111",
  278=>"011111110",
  279=>"110101101",
  280=>"100100100",
  281=>"010111000",
  282=>"111111111",
  283=>"111000010",
  284=>"101111110",
  285=>"000000110",
  286=>"111000000",
  287=>"111011101",
  288=>"000000011",
  289=>"110111011",
  290=>"000010011",
  291=>"111001111",
  292=>"011000001",
  293=>"010000000",
  294=>"100100001",
  295=>"000000111",
  296=>"000000101",
  297=>"000000110",
  298=>"000000101",
  299=>"111100110",
  300=>"110101111",
  301=>"101101111",
  302=>"000110110",
  303=>"000000000",
  304=>"001111101",
  305=>"111101111",
  306=>"100000100",
  307=>"000000110",
  308=>"000110110",
  309=>"000001000",
  310=>"101000000",
  311=>"010000001",
  312=>"000111110",
  313=>"111111111",
  314=>"111000000",
  315=>"000000000",
  316=>"111000000",
  317=>"000111110",
  318=>"111101100",
  319=>"111111111",
  320=>"001111111",
  321=>"110110010",
  322=>"111111111",
  323=>"111101000",
  324=>"111111110",
  325=>"011011000",
  326=>"000010110",
  327=>"111000000",
  328=>"111100101",
  329=>"011000000",
  330=>"110111110",
  331=>"001001001",
  332=>"010000000",
  333=>"010111010",
  334=>"000111111",
  335=>"000000111",
  336=>"110000000",
  337=>"000000000",
  338=>"111111111",
  339=>"111100111",
  340=>"000000110",
  341=>"000111111",
  342=>"111011111",
  343=>"000111111",
  344=>"011111111",
  345=>"010000000",
  346=>"111000101",
  347=>"000001000",
  348=>"000000000",
  349=>"111111101",
  350=>"000000000",
  351=>"001010110",
  352=>"000010010",
  353=>"111110000",
  354=>"010111011",
  355=>"000000001",
  356=>"111110110",
  357=>"000000100",
  358=>"011000111",
  359=>"000000000",
  360=>"110100100",
  361=>"000111111",
  362=>"101101111",
  363=>"110111100",
  364=>"001111011",
  365=>"000010000",
  366=>"000000000",
  367=>"011111000",
  368=>"000000100",
  369=>"001001011",
  370=>"100111111",
  371=>"000000110",
  372=>"000110000",
  373=>"100111000",
  374=>"000011000",
  375=>"111101111",
  376=>"111001001",
  377=>"111110111",
  378=>"000101111",
  379=>"000101111",
  380=>"010111100",
  381=>"111111111",
  382=>"100100111",
  383=>"110000000",
  384=>"010111110",
  385=>"111000111",
  386=>"110111111",
  387=>"111111111",
  388=>"000111111",
  389=>"100100100",
  390=>"000111111",
  391=>"001010110",
  392=>"000000000",
  393=>"011111100",
  394=>"110110000",
  395=>"111001111",
  396=>"000001000",
  397=>"000001001",
  398=>"000000001",
  399=>"000110110",
  400=>"111100000",
  401=>"110010000",
  402=>"111000000",
  403=>"111010000",
  404=>"101001111",
  405=>"000000000",
  406=>"100110111",
  407=>"000001011",
  408=>"000000100",
  409=>"010000000",
  410=>"010110000",
  411=>"000111111",
  412=>"111111101",
  413=>"111101111",
  414=>"111001000",
  415=>"000111111",
  416=>"000000111",
  417=>"001011011",
  418=>"100000100",
  419=>"100000000",
  420=>"000000001",
  421=>"111111101",
  422=>"000000000",
  423=>"111000000",
  424=>"000100111",
  425=>"110111111",
  426=>"000000000",
  427=>"100100101",
  428=>"111100111",
  429=>"111000000",
  430=>"111111000",
  431=>"000101111",
  432=>"001001000",
  433=>"100111111",
  434=>"000000000",
  435=>"001111000",
  436=>"000000000",
  437=>"000000000",
  438=>"110010000",
  439=>"111000000",
  440=>"110110000",
  441=>"111001001",
  442=>"000000100",
  443=>"000000111",
  444=>"000000000",
  445=>"000001001",
  446=>"001001000",
  447=>"011011010",
  448=>"000000000",
  449=>"111111111",
  450=>"111000010",
  451=>"111000001",
  452=>"111110000",
  453=>"000100100",
  454=>"000000000",
  455=>"000101011",
  456=>"000000000",
  457=>"000101111",
  458=>"001000000",
  459=>"111111000",
  460=>"000000100",
  461=>"000000000",
  462=>"000000111",
  463=>"000110000",
  464=>"011111111",
  465=>"000110110",
  466=>"000100000",
  467=>"000110111",
  468=>"100111111",
  469=>"000000000",
  470=>"000100101",
  471=>"001000000",
  472=>"000001111",
  473=>"111101110",
  474=>"000000100",
  475=>"000000000",
  476=>"001011111",
  477=>"111111000",
  478=>"000000000",
  479=>"001000000",
  480=>"000011011",
  481=>"000111101",
  482=>"011000000",
  483=>"000000000",
  484=>"111111111",
  485=>"000000000",
  486=>"001000000",
  487=>"100101101",
  488=>"010000000",
  489=>"111111010",
  490=>"110100111",
  491=>"111111111",
  492=>"111111111",
  493=>"000000100",
  494=>"111111111",
  495=>"110111111",
  496=>"000000000",
  497=>"111111111",
  498=>"000000111",
  499=>"000000000",
  500=>"000000000",
  501=>"110000000",
  502=>"100100100",
  503=>"100110110",
  504=>"110110110",
  505=>"000110000",
  506=>"111111111",
  507=>"110100000",
  508=>"000000000",
  509=>"111111111",
  510=>"000000011",
  511=>"010000000",
  512=>"000000000",
  513=>"111110110",
  514=>"101000101",
  515=>"111111111",
  516=>"101011001",
  517=>"011011000",
  518=>"011111011",
  519=>"111111111",
  520=>"000100000",
  521=>"000000000",
  522=>"010111111",
  523=>"111111001",
  524=>"010111111",
  525=>"000111111",
  526=>"100110111",
  527=>"111111111",
  528=>"110111000",
  529=>"000000000",
  530=>"111111111",
  531=>"000000001",
  532=>"000000100",
  533=>"111111000",
  534=>"000000000",
  535=>"011011011",
  536=>"100101111",
  537=>"111111111",
  538=>"111111110",
  539=>"001100001",
  540=>"000000000",
  541=>"000000111",
  542=>"000000000",
  543=>"000100100",
  544=>"100111000",
  545=>"000000000",
  546=>"111111111",
  547=>"101110101",
  548=>"111101001",
  549=>"011001000",
  550=>"111111111",
  551=>"000100111",
  552=>"000000000",
  553=>"111111111",
  554=>"111111111",
  555=>"000010111",
  556=>"101000000",
  557=>"111111100",
  558=>"111111111",
  559=>"011000000",
  560=>"111111111",
  561=>"101000000",
  562=>"111100000",
  563=>"000001011",
  564=>"110111111",
  565=>"110100100",
  566=>"111100110",
  567=>"000110111",
  568=>"000001111",
  569=>"001000100",
  570=>"110111111",
  571=>"000000111",
  572=>"000000000",
  573=>"111111111",
  574=>"111011000",
  575=>"111100110",
  576=>"111110000",
  577=>"110111000",
  578=>"000000100",
  579=>"000111111",
  580=>"110111111",
  581=>"000000000",
  582=>"000000001",
  583=>"111111110",
  584=>"111111111",
  585=>"000110111",
  586=>"111000000",
  587=>"000011111",
  588=>"001000100",
  589=>"111111111",
  590=>"000000000",
  591=>"000111001",
  592=>"000000100",
  593=>"111011011",
  594=>"111101101",
  595=>"100101100",
  596=>"011001000",
  597=>"111110111",
  598=>"011000100",
  599=>"000000000",
  600=>"000000000",
  601=>"111111111",
  602=>"000000000",
  603=>"011011000",
  604=>"000000000",
  605=>"101100000",
  606=>"001110111",
  607=>"011111000",
  608=>"000101111",
  609=>"000000000",
  610=>"011111111",
  611=>"000101111",
  612=>"000000000",
  613=>"000100110",
  614=>"000000000",
  615=>"000000000",
  616=>"001111011",
  617=>"000000111",
  618=>"111110111",
  619=>"001011011",
  620=>"111011000",
  621=>"111100000",
  622=>"100111111",
  623=>"111111111",
  624=>"111000000",
  625=>"111100100",
  626=>"111100000",
  627=>"000000000",
  628=>"111111001",
  629=>"000000000",
  630=>"010110110",
  631=>"011000000",
  632=>"000000000",
  633=>"111000001",
  634=>"111000000",
  635=>"000000000",
  636=>"100100100",
  637=>"111111111",
  638=>"111001111",
  639=>"111000000",
  640=>"111011011",
  641=>"000000000",
  642=>"000100011",
  643=>"001001001",
  644=>"110100111",
  645=>"000000000",
  646=>"111111111",
  647=>"111101000",
  648=>"001000000",
  649=>"000000100",
  650=>"000100111",
  651=>"000000000",
  652=>"111100100",
  653=>"111100100",
  654=>"000000001",
  655=>"000000000",
  656=>"010000110",
  657=>"111111000",
  658=>"111101000",
  659=>"111111111",
  660=>"111111111",
  661=>"000011111",
  662=>"000000000",
  663=>"111111111",
  664=>"111101100",
  665=>"111111011",
  666=>"000000000",
  667=>"000000111",
  668=>"111111111",
  669=>"110101100",
  670=>"111011111",
  671=>"000000111",
  672=>"000010011",
  673=>"111111111",
  674=>"000000100",
  675=>"000000000",
  676=>"111111111",
  677=>"111011011",
  678=>"111000000",
  679=>"000000000",
  680=>"111111111",
  681=>"011001000",
  682=>"001001000",
  683=>"000000000",
  684=>"111111000",
  685=>"000000000",
  686=>"111111111",
  687=>"000001101",
  688=>"110101111",
  689=>"111111111",
  690=>"111111111",
  691=>"011000000",
  692=>"000000000",
  693=>"000000000",
  694=>"000000000",
  695=>"011111111",
  696=>"000011101",
  697=>"111111111",
  698=>"010111111",
  699=>"000000000",
  700=>"111100000",
  701=>"000000100",
  702=>"111010000",
  703=>"000000000",
  704=>"000000111",
  705=>"001001111",
  706=>"111111111",
  707=>"111111111",
  708=>"101100110",
  709=>"000111111",
  710=>"100000110",
  711=>"000000000",
  712=>"011111111",
  713=>"111111010",
  714=>"000000000",
  715=>"000000000",
  716=>"111011111",
  717=>"101111111",
  718=>"000000000",
  719=>"111010010",
  720=>"111111111",
  721=>"001001000",
  722=>"111111111",
  723=>"000010010",
  724=>"011000111",
  725=>"010010110",
  726=>"111111011",
  727=>"011001000",
  728=>"000001001",
  729=>"111111111",
  730=>"000000111",
  731=>"000000000",
  732=>"000110110",
  733=>"111111111",
  734=>"000001111",
  735=>"111111111",
  736=>"000000000",
  737=>"000000000",
  738=>"000000000",
  739=>"000000000",
  740=>"111111111",
  741=>"100001001",
  742=>"001000000",
  743=>"000000111",
  744=>"111111111",
  745=>"000000011",
  746=>"111111111",
  747=>"111111111",
  748=>"000000000",
  749=>"000000000",
  750=>"111111111",
  751=>"011000000",
  752=>"011011101",
  753=>"000000001",
  754=>"011011011",
  755=>"000000100",
  756=>"111111111",
  757=>"111100000",
  758=>"000000000",
  759=>"111111000",
  760=>"000000100",
  761=>"000100111",
  762=>"000000000",
  763=>"101101001",
  764=>"110110000",
  765=>"000000000",
  766=>"011001001",
  767=>"000000101",
  768=>"111111111",
  769=>"111111011",
  770=>"000000001",
  771=>"111111110",
  772=>"001000000",
  773=>"111000111",
  774=>"111111111",
  775=>"111111110",
  776=>"111111111",
  777=>"000000001",
  778=>"000111111",
  779=>"101111111",
  780=>"100100110",
  781=>"101000001",
  782=>"100111111",
  783=>"111111011",
  784=>"001010000",
  785=>"000101111",
  786=>"000000100",
  787=>"000000000",
  788=>"101101001",
  789=>"001111111",
  790=>"000000000",
  791=>"111111111",
  792=>"110111111",
  793=>"110100111",
  794=>"000000000",
  795=>"000000111",
  796=>"111111111",
  797=>"000110110",
  798=>"111111110",
  799=>"000000111",
  800=>"000000001",
  801=>"110110110",
  802=>"000000000",
  803=>"111111111",
  804=>"011111111",
  805=>"111101111",
  806=>"001111111",
  807=>"000000100",
  808=>"111101000",
  809=>"001101111",
  810=>"001000000",
  811=>"000000000",
  812=>"001011011",
  813=>"000000000",
  814=>"000111000",
  815=>"000100111",
  816=>"011000000",
  817=>"010000000",
  818=>"000000000",
  819=>"000100111",
  820=>"111101100",
  821=>"000000000",
  822=>"000000000",
  823=>"000000000",
  824=>"100000000",
  825=>"100111111",
  826=>"000111111",
  827=>"111111111",
  828=>"001000000",
  829=>"001010010",
  830=>"000000000",
  831=>"011111111",
  832=>"111111111",
  833=>"111111111",
  834=>"111111111",
  835=>"010110100",
  836=>"000000111",
  837=>"111111111",
  838=>"000000111",
  839=>"110111111",
  840=>"000000000",
  841=>"011000001",
  842=>"111111111",
  843=>"111111111",
  844=>"000000010",
  845=>"111111111",
  846=>"001111111",
  847=>"100110110",
  848=>"000101111",
  849=>"000000110",
  850=>"111000000",
  851=>"110001111",
  852=>"000110111",
  853=>"001011011",
  854=>"111111000",
  855=>"001000000",
  856=>"000000100",
  857=>"000000000",
  858=>"001000000",
  859=>"100000000",
  860=>"000000111",
  861=>"111111111",
  862=>"111111111",
  863=>"110111111",
  864=>"001011111",
  865=>"000000000",
  866=>"000000000",
  867=>"100000001",
  868=>"000000000",
  869=>"111111111",
  870=>"100000011",
  871=>"111111001",
  872=>"110010110",
  873=>"111111000",
  874=>"000110000",
  875=>"110000000",
  876=>"100101111",
  877=>"000010000",
  878=>"010111000",
  879=>"000000000",
  880=>"111111111",
  881=>"000000000",
  882=>"111111111",
  883=>"111111111",
  884=>"111111010",
  885=>"111111111",
  886=>"000000000",
  887=>"000100101",
  888=>"111111111",
  889=>"111111111",
  890=>"000000000",
  891=>"000000000",
  892=>"010010001",
  893=>"111000001",
  894=>"001000000",
  895=>"000000000",
  896=>"110000000",
  897=>"000000000",
  898=>"000000000",
  899=>"111011000",
  900=>"111100100",
  901=>"000110110",
  902=>"010110111",
  903=>"111111110",
  904=>"110110111",
  905=>"110011000",
  906=>"111011011",
  907=>"111100110",
  908=>"000000000",
  909=>"110110110",
  910=>"111111111",
  911=>"000000011",
  912=>"001010010",
  913=>"011001000",
  914=>"100001111",
  915=>"011000110",
  916=>"111111111",
  917=>"000000000",
  918=>"011001001",
  919=>"001111000",
  920=>"000000000",
  921=>"010000001",
  922=>"000000000",
  923=>"000000000",
  924=>"001011011",
  925=>"110110111",
  926=>"000000001",
  927=>"110110000",
  928=>"000000000",
  929=>"000010001",
  930=>"001100100",
  931=>"111111000",
  932=>"001000000",
  933=>"001001000",
  934=>"101001001",
  935=>"011000000",
  936=>"111111011",
  937=>"111111111",
  938=>"011000000",
  939=>"000000001",
  940=>"111101101",
  941=>"001001000",
  942=>"000011001",
  943=>"000000001",
  944=>"111110000",
  945=>"000000000",
  946=>"110111111",
  947=>"111111111",
  948=>"000000100",
  949=>"111111111",
  950=>"101111111",
  951=>"100000000",
  952=>"001001000",
  953=>"001000000",
  954=>"111111011",
  955=>"000000000",
  956=>"100100110",
  957=>"011000000",
  958=>"011000000",
  959=>"000111100",
  960=>"000000010",
  961=>"000000110",
  962=>"000000000",
  963=>"000000000",
  964=>"011010111",
  965=>"000000000",
  966=>"100100000",
  967=>"111101111",
  968=>"000100000",
  969=>"110110111",
  970=>"000000000",
  971=>"111111110",
  972=>"000100000",
  973=>"111000000",
  974=>"111011000",
  975=>"010000000",
  976=>"110011111",
  977=>"101111111",
  978=>"111111011",
  979=>"111101111",
  980=>"111101000",
  981=>"111111001",
  982=>"111111111",
  983=>"000000010",
  984=>"000000100",
  985=>"000000000",
  986=>"100100000",
  987=>"011001111",
  988=>"000000000",
  989=>"100100100",
  990=>"000000000",
  991=>"000000000",
  992=>"100000000",
  993=>"000111010",
  994=>"000000000",
  995=>"111101000",
  996=>"111000111",
  997=>"111101111",
  998=>"101000100",
  999=>"010000000",
  1000=>"101000101",
  1001=>"011011011",
  1002=>"111110100",
  1003=>"111110110",
  1004=>"000101111",
  1005=>"011001000",
  1006=>"000100110",
  1007=>"111011110",
  1008=>"000000011",
  1009=>"010111111",
  1010=>"111000000",
  1011=>"111111011",
  1012=>"111111111",
  1013=>"011001001",
  1014=>"111111111",
  1015=>"100000000",
  1016=>"010011011",
  1017=>"011010010",
  1018=>"101011011",
  1019=>"000000000",
  1020=>"111111011",
  1021=>"001000000",
  1022=>"111111111",
  1023=>"111111111",
  1024=>"111111111",
  1025=>"111111101",
  1026=>"000010011",
  1027=>"111111110",
  1028=>"111001111",
  1029=>"000000110",
  1030=>"000000000",
  1031=>"111001001",
  1032=>"000000000",
  1033=>"111011001",
  1034=>"111100101",
  1035=>"100011011",
  1036=>"011001001",
  1037=>"100111111",
  1038=>"000000000",
  1039=>"111101101",
  1040=>"111101001",
  1041=>"000000000",
  1042=>"111111111",
  1043=>"111111111",
  1044=>"000000001",
  1045=>"000111111",
  1046=>"100111111",
  1047=>"111111011",
  1048=>"100100000",
  1049=>"000100100",
  1050=>"101001011",
  1051=>"111111111",
  1052=>"111111111",
  1053=>"111111111",
  1054=>"001111111",
  1055=>"000000001",
  1056=>"001000101",
  1057=>"000000001",
  1058=>"101101101",
  1059=>"000000100",
  1060=>"000100100",
  1061=>"000100111",
  1062=>"111100000",
  1063=>"111001000",
  1064=>"000101101",
  1065=>"000000000",
  1066=>"110111111",
  1067=>"101111101",
  1068=>"111111111",
  1069=>"110010000",
  1070=>"011011000",
  1071=>"100000000",
  1072=>"000000000",
  1073=>"110101100",
  1074=>"111001111",
  1075=>"000000000",
  1076=>"111001001",
  1077=>"101000000",
  1078=>"100100100",
  1079=>"000111111",
  1080=>"111111111",
  1081=>"111011000",
  1082=>"000110111",
  1083=>"010000000",
  1084=>"100000000",
  1085=>"111111111",
  1086=>"111001000",
  1087=>"000000110",
  1088=>"100000000",
  1089=>"011001011",
  1090=>"111110110",
  1091=>"011011111",
  1092=>"000000001",
  1093=>"110110000",
  1094=>"000000000",
  1095=>"111001001",
  1096=>"011011001",
  1097=>"000000000",
  1098=>"111111110",
  1099=>"001001001",
  1100=>"010011110",
  1101=>"100101000",
  1102=>"000011100",
  1103=>"000000000",
  1104=>"101111100",
  1105=>"110111111",
  1106=>"111000000",
  1107=>"111110111",
  1108=>"110110111",
  1109=>"001111111",
  1110=>"111111111",
  1111=>"111111111",
  1112=>"111111000",
  1113=>"111000000",
  1114=>"111111001",
  1115=>"001001000",
  1116=>"000000001",
  1117=>"000000111",
  1118=>"000000000",
  1119=>"000000000",
  1120=>"111000000",
  1121=>"111111111",
  1122=>"100111111",
  1123=>"011000000",
  1124=>"011000000",
  1125=>"101000010",
  1126=>"111111000",
  1127=>"111111111",
  1128=>"000000011",
  1129=>"011001111",
  1130=>"000010010",
  1131=>"000100000",
  1132=>"100100000",
  1133=>"111000100",
  1134=>"000110000",
  1135=>"110111010",
  1136=>"111100110",
  1137=>"001001100",
  1138=>"011011111",
  1139=>"001000000",
  1140=>"111111111",
  1141=>"101101001",
  1142=>"111111011",
  1143=>"000000000",
  1144=>"111111111",
  1145=>"110110110",
  1146=>"100101101",
  1147=>"000000000",
  1148=>"100100100",
  1149=>"000111111",
  1150=>"000000001",
  1151=>"011111111",
  1152=>"000000000",
  1153=>"110000000",
  1154=>"100110110",
  1155=>"001001001",
  1156=>"100100110",
  1157=>"000000000",
  1158=>"000110110",
  1159=>"011010010",
  1160=>"110110110",
  1161=>"111111111",
  1162=>"000000000",
  1163=>"111111110",
  1164=>"111101000",
  1165=>"111111111",
  1166=>"000111111",
  1167=>"001001011",
  1168=>"111111111",
  1169=>"000111111",
  1170=>"000000110",
  1171=>"000000000",
  1172=>"000000000",
  1173=>"100100000",
  1174=>"000000000",
  1175=>"000110110",
  1176=>"111111101",
  1177=>"111111111",
  1178=>"100100000",
  1179=>"000000000",
  1180=>"111111111",
  1181=>"110010000",
  1182=>"000000000",
  1183=>"100000000",
  1184=>"110101001",
  1185=>"111111111",
  1186=>"001001001",
  1187=>"110111110",
  1188=>"101111111",
  1189=>"011011000",
  1190=>"110000000",
  1191=>"011011001",
  1192=>"110010001",
  1193=>"000000000",
  1194=>"000000000",
  1195=>"000000000",
  1196=>"100101001",
  1197=>"101011000",
  1198=>"000001111",
  1199=>"000000000",
  1200=>"111111000",
  1201=>"110110011",
  1202=>"110111110",
  1203=>"010000011",
  1204=>"000000000",
  1205=>"111100000",
  1206=>"000000000",
  1207=>"100000000",
  1208=>"101101111",
  1209=>"111111110",
  1210=>"101100000",
  1211=>"101000110",
  1212=>"010010000",
  1213=>"111111111",
  1214=>"111111111",
  1215=>"000100111",
  1216=>"100101111",
  1217=>"111111111",
  1218=>"000000000",
  1219=>"111111111",
  1220=>"111111110",
  1221=>"011000001",
  1222=>"100101111",
  1223=>"000000101",
  1224=>"000110101",
  1225=>"101111111",
  1226=>"000100101",
  1227=>"110110010",
  1228=>"000000101",
  1229=>"000010010",
  1230=>"000110111",
  1231=>"111111111",
  1232=>"111111011",
  1233=>"000000101",
  1234=>"110000000",
  1235=>"100000000",
  1236=>"000001101",
  1237=>"000000000",
  1238=>"011010010",
  1239=>"000000000",
  1240=>"111111111",
  1241=>"011010100",
  1242=>"000000000",
  1243=>"011000000",
  1244=>"000000100",
  1245=>"111111000",
  1246=>"111111111",
  1247=>"100100000",
  1248=>"000000000",
  1249=>"010011000",
  1250=>"111111111",
  1251=>"101110000",
  1252=>"100000000",
  1253=>"100000111",
  1254=>"110110110",
  1255=>"111111111",
  1256=>"111111011",
  1257=>"111111111",
  1258=>"000000001",
  1259=>"000111011",
  1260=>"010011001",
  1261=>"011000010",
  1262=>"000000001",
  1263=>"110111111",
  1264=>"101111111",
  1265=>"111111111",
  1266=>"100110000",
  1267=>"001011111",
  1268=>"100000000",
  1269=>"001000000",
  1270=>"000000000",
  1271=>"000000010",
  1272=>"111110110",
  1273=>"010110010",
  1274=>"001001000",
  1275=>"001011011",
  1276=>"000100110",
  1277=>"110110100",
  1278=>"000000000",
  1279=>"001111111",
  1280=>"111111111",
  1281=>"000000001",
  1282=>"111111111",
  1283=>"000000000",
  1284=>"100000100",
  1285=>"000101101",
  1286=>"101101101",
  1287=>"000100000",
  1288=>"111111111",
  1289=>"000000001",
  1290=>"100110111",
  1291=>"111111001",
  1292=>"100000000",
  1293=>"111111111",
  1294=>"111111111",
  1295=>"110011000",
  1296=>"100100100",
  1297=>"000000000",
  1298=>"110110111",
  1299=>"110111111",
  1300=>"000100100",
  1301=>"111111100",
  1302=>"100111111",
  1303=>"101101111",
  1304=>"100000001",
  1305=>"000100100",
  1306=>"111111111",
  1307=>"000000100",
  1308=>"000001001",
  1309=>"001000000",
  1310=>"000100110",
  1311=>"100000011",
  1312=>"111111011",
  1313=>"000000000",
  1314=>"101111011",
  1315=>"100111111",
  1316=>"111111111",
  1317=>"111111011",
  1318=>"000000001",
  1319=>"011001101",
  1320=>"111111000",
  1321=>"000000010",
  1322=>"011000000",
  1323=>"000000000",
  1324=>"000000110",
  1325=>"111111110",
  1326=>"111000001",
  1327=>"000000000",
  1328=>"001111000",
  1329=>"000000000",
  1330=>"011111111",
  1331=>"000000000",
  1332=>"000000000",
  1333=>"111111111",
  1334=>"110111111",
  1335=>"000000000",
  1336=>"000000000",
  1337=>"100000100",
  1338=>"000000000",
  1339=>"000000000",
  1340=>"000000110",
  1341=>"000000111",
  1342=>"000101100",
  1343=>"100000100",
  1344=>"000000000",
  1345=>"100111111",
  1346=>"101111101",
  1347=>"111011111",
  1348=>"001001101",
  1349=>"111111111",
  1350=>"100100101",
  1351=>"111111111",
  1352=>"000000101",
  1353=>"000000000",
  1354=>"100000000",
  1355=>"100000000",
  1356=>"101001101",
  1357=>"000000000",
  1358=>"111111111",
  1359=>"000000011",
  1360=>"100110110",
  1361=>"111100000",
  1362=>"000110111",
  1363=>"111100111",
  1364=>"000000000",
  1365=>"001001001",
  1366=>"000100110",
  1367=>"110110111",
  1368=>"111111111",
  1369=>"100100111",
  1370=>"011000000",
  1371=>"000000000",
  1372=>"111111101",
  1373=>"111111111",
  1374=>"011000000",
  1375=>"000001111",
  1376=>"000000110",
  1377=>"000000000",
  1378=>"011011001",
  1379=>"101001111",
  1380=>"101111111",
  1381=>"000000000",
  1382=>"000000000",
  1383=>"000000000",
  1384=>"100110101",
  1385=>"011000011",
  1386=>"000001000",
  1387=>"000001111",
  1388=>"011111111",
  1389=>"101111111",
  1390=>"101000100",
  1391=>"000000000",
  1392=>"000001000",
  1393=>"000000000",
  1394=>"000000000",
  1395=>"001000000",
  1396=>"110010110",
  1397=>"111110001",
  1398=>"000000000",
  1399=>"001000000",
  1400=>"111000000",
  1401=>"000000000",
  1402=>"000000000",
  1403=>"100000000",
  1404=>"100100101",
  1405=>"000000000",
  1406=>"000000000",
  1407=>"100000000",
  1408=>"111111011",
  1409=>"000000111",
  1410=>"111111011",
  1411=>"000000000",
  1412=>"110011000",
  1413=>"000000000",
  1414=>"001001001",
  1415=>"000000100",
  1416=>"000000100",
  1417=>"000001011",
  1418=>"000100101",
  1419=>"000010111",
  1420=>"111111111",
  1421=>"111110100",
  1422=>"111111111",
  1423=>"111111011",
  1424=>"010010000",
  1425=>"000000100",
  1426=>"001001000",
  1427=>"110110110",
  1428=>"001011111",
  1429=>"000000000",
  1430=>"101101101",
  1431=>"001001000",
  1432=>"110110011",
  1433=>"100000000",
  1434=>"111111111",
  1435=>"001001000",
  1436=>"000000000",
  1437=>"010011111",
  1438=>"000000000",
  1439=>"000000000",
  1440=>"111101100",
  1441=>"001001000",
  1442=>"000000011",
  1443=>"111111111",
  1444=>"001101101",
  1445=>"111111011",
  1446=>"111110111",
  1447=>"010011111",
  1448=>"100000010",
  1449=>"001100110",
  1450=>"001111101",
  1451=>"000000000",
  1452=>"100110110",
  1453=>"000111100",
  1454=>"100111001",
  1455=>"000000001",
  1456=>"010000000",
  1457=>"000000000",
  1458=>"111111111",
  1459=>"001111111",
  1460=>"000000100",
  1461=>"000000000",
  1462=>"101101111",
  1463=>"111111111",
  1464=>"001000000",
  1465=>"100000011",
  1466=>"011000000",
  1467=>"100100000",
  1468=>"000000001",
  1469=>"111000001",
  1470=>"110000000",
  1471=>"101111111",
  1472=>"000000010",
  1473=>"111111111",
  1474=>"011000011",
  1475=>"111111110",
  1476=>"011000000",
  1477=>"000000000",
  1478=>"001001000",
  1479=>"111011001",
  1480=>"001000011",
  1481=>"000000110",
  1482=>"000000000",
  1483=>"100001001",
  1484=>"000000000",
  1485=>"001010000",
  1486=>"000000001",
  1487=>"111111111",
  1488=>"001000000",
  1489=>"000000100",
  1490=>"101001000",
  1491=>"000000000",
  1492=>"000000111",
  1493=>"000000000",
  1494=>"000000000",
  1495=>"111100111",
  1496=>"000000000",
  1497=>"100111111",
  1498=>"011010000",
  1499=>"101111111",
  1500=>"100100110",
  1501=>"111110100",
  1502=>"001011111",
  1503=>"100101111",
  1504=>"000000001",
  1505=>"111000000",
  1506=>"111110000",
  1507=>"111011001",
  1508=>"101111000",
  1509=>"000000000",
  1510=>"111110000",
  1511=>"010111111",
  1512=>"101000001",
  1513=>"111101001",
  1514=>"000000011",
  1515=>"000000001",
  1516=>"111000000",
  1517=>"100100100",
  1518=>"011111111",
  1519=>"110110111",
  1520=>"000000000",
  1521=>"000000000",
  1522=>"011111111",
  1523=>"010000000",
  1524=>"000000000",
  1525=>"111010100",
  1526=>"111111111",
  1527=>"000000000",
  1528=>"111111111",
  1529=>"100000100",
  1530=>"101111111",
  1531=>"000000000",
  1532=>"000000000",
  1533=>"000000000",
  1534=>"110111110",
  1535=>"100100110",
  1536=>"111111111",
  1537=>"110110100",
  1538=>"110000000",
  1539=>"011000000",
  1540=>"111111111",
  1541=>"000000000",
  1542=>"111111111",
  1543=>"111000000",
  1544=>"111111111",
  1545=>"111001001",
  1546=>"001000001",
  1547=>"111100000",
  1548=>"111001000",
  1549=>"000100000",
  1550=>"110111111",
  1551=>"111011111",
  1552=>"000000000",
  1553=>"111111111",
  1554=>"000000000",
  1555=>"000000001",
  1556=>"110000000",
  1557=>"110010000",
  1558=>"110010000",
  1559=>"000000000",
  1560=>"111111111",
  1561=>"011001011",
  1562=>"101000000",
  1563=>"111111110",
  1564=>"001001111",
  1565=>"011000011",
  1566=>"000010111",
  1567=>"000000000",
  1568=>"000000011",
  1569=>"000000000",
  1570=>"011001001",
  1571=>"010010111",
  1572=>"001101000",
  1573=>"111001011",
  1574=>"111100110",
  1575=>"000000111",
  1576=>"001000000",
  1577=>"000000000",
  1578=>"111111111",
  1579=>"011011011",
  1580=>"110010011",
  1581=>"110000000",
  1582=>"011011011",
  1583=>"111111111",
  1584=>"001000111",
  1585=>"011001000",
  1586=>"001000101",
  1587=>"011111111",
  1588=>"011011011",
  1589=>"111011011",
  1590=>"001000000",
  1591=>"111000000",
  1592=>"001000000",
  1593=>"111111111",
  1594=>"000000000",
  1595=>"010110010",
  1596=>"000000000",
  1597=>"111100100",
  1598=>"111111111",
  1599=>"111000100",
  1600=>"000000001",
  1601=>"101001101",
  1602=>"001000111",
  1603=>"000000000",
  1604=>"000000000",
  1605=>"000000000",
  1606=>"110110000",
  1607=>"111111111",
  1608=>"001001001",
  1609=>"000000000",
  1610=>"111111111",
  1611=>"110000101",
  1612=>"111111111",
  1613=>"100000111",
  1614=>"000011011",
  1615=>"000000000",
  1616=>"100000001",
  1617=>"000000000",
  1618=>"011011011",
  1619=>"011011111",
  1620=>"000000000",
  1621=>"000000000",
  1622=>"101101111",
  1623=>"011011001",
  1624=>"000010000",
  1625=>"000000000",
  1626=>"111000101",
  1627=>"001000110",
  1628=>"111111111",
  1629=>"111111110",
  1630=>"000000000",
  1631=>"000000000",
  1632=>"111000000",
  1633=>"000000000",
  1634=>"100100000",
  1635=>"011111111",
  1636=>"000111111",
  1637=>"000000000",
  1638=>"111111000",
  1639=>"101100111",
  1640=>"111111111",
  1641=>"111111111",
  1642=>"000100111",
  1643=>"000000001",
  1644=>"111111111",
  1645=>"000000000",
  1646=>"000000000",
  1647=>"000000010",
  1648=>"000000000",
  1649=>"111111101",
  1650=>"000000001",
  1651=>"111011011",
  1652=>"111111111",
  1653=>"100100000",
  1654=>"111111111",
  1655=>"000000000",
  1656=>"000000000",
  1657=>"011011010",
  1658=>"000001111",
  1659=>"011000000",
  1660=>"000000010",
  1661=>"110110000",
  1662=>"000000001",
  1663=>"000000000",
  1664=>"110111010",
  1665=>"000000000",
  1666=>"000000010",
  1667=>"111111111",
  1668=>"100100100",
  1669=>"001001111",
  1670=>"100000000",
  1671=>"001001110",
  1672=>"111111111",
  1673=>"011011001",
  1674=>"000000000",
  1675=>"111111111",
  1676=>"000000000",
  1677=>"111111111",
  1678=>"111111111",
  1679=>"000001001",
  1680=>"111111111",
  1681=>"111111111",
  1682=>"111111111",
  1683=>"000000000",
  1684=>"000000000",
  1685=>"000000000",
  1686=>"000010111",
  1687=>"001001011",
  1688=>"111111111",
  1689=>"001101101",
  1690=>"111111111",
  1691=>"101000000",
  1692=>"110110000",
  1693=>"100001111",
  1694=>"100000000",
  1695=>"000000000",
  1696=>"000000000",
  1697=>"000000000",
  1698=>"000000001",
  1699=>"111111111",
  1700=>"001000100",
  1701=>"111111000",
  1702=>"111111111",
  1703=>"111111110",
  1704=>"111111110",
  1705=>"000000000",
  1706=>"000000000",
  1707=>"000000000",
  1708=>"000000000",
  1709=>"000000000",
  1710=>"111111111",
  1711=>"000011011",
  1712=>"111000111",
  1713=>"011001001",
  1714=>"111111111",
  1715=>"000000000",
  1716=>"111111001",
  1717=>"011000000",
  1718=>"111111011",
  1719=>"110110010",
  1720=>"110110110",
  1721=>"000000000",
  1722=>"111001001",
  1723=>"111101111",
  1724=>"010010010",
  1725=>"000000011",
  1726=>"010111000",
  1727=>"111111111",
  1728=>"011011011",
  1729=>"100000001",
  1730=>"111111111",
  1731=>"000000000",
  1732=>"100111111",
  1733=>"010001000",
  1734=>"000000000",
  1735=>"101111111",
  1736=>"001000000",
  1737=>"100000001",
  1738=>"000001011",
  1739=>"000000000",
  1740=>"001100111",
  1741=>"000000111",
  1742=>"000100111",
  1743=>"001011111",
  1744=>"111111111",
  1745=>"111111011",
  1746=>"110110000",
  1747=>"000000101",
  1748=>"111111111",
  1749=>"000100111",
  1750=>"000000000",
  1751=>"001111100",
  1752=>"000000111",
  1753=>"001000000",
  1754=>"000000000",
  1755=>"111111111",
  1756=>"111111110",
  1757=>"000011011",
  1758=>"111111111",
  1759=>"101000000",
  1760=>"111111111",
  1761=>"111110110",
  1762=>"000000000",
  1763=>"110001111",
  1764=>"000000010",
  1765=>"000000000",
  1766=>"000011111",
  1767=>"000000000",
  1768=>"111001000",
  1769=>"000000111",
  1770=>"000000000",
  1771=>"111111111",
  1772=>"000000000",
  1773=>"111111111",
  1774=>"111100000",
  1775=>"000000000",
  1776=>"000111010",
  1777=>"110111111",
  1778=>"111111111",
  1779=>"000000001",
  1780=>"111111111",
  1781=>"000000000",
  1782=>"100100000",
  1783=>"111111011",
  1784=>"111000000",
  1785=>"000000100",
  1786=>"111111111",
  1787=>"100000111",
  1788=>"000000001",
  1789=>"000000000",
  1790=>"111111011",
  1791=>"100111111",
  1792=>"111000001",
  1793=>"000000100",
  1794=>"001001000",
  1795=>"111001000",
  1796=>"001000011",
  1797=>"111000000",
  1798=>"000000000",
  1799=>"001100100",
  1800=>"000000011",
  1801=>"000000010",
  1802=>"111111111",
  1803=>"101101001",
  1804=>"111111111",
  1805=>"100101111",
  1806=>"111110000",
  1807=>"000000000",
  1808=>"000000000",
  1809=>"011011011",
  1810=>"000000000",
  1811=>"111100100",
  1812=>"000000000",
  1813=>"000000111",
  1814=>"011011001",
  1815=>"000000000",
  1816=>"011011111",
  1817=>"000000000",
  1818=>"000000100",
  1819=>"100000000",
  1820=>"110011111",
  1821=>"000000000",
  1822=>"000000000",
  1823=>"000000000",
  1824=>"111111011",
  1825=>"111111111",
  1826=>"000000000",
  1827=>"001111000",
  1828=>"000000111",
  1829=>"010000000",
  1830=>"110111111",
  1831=>"111000001",
  1832=>"000000000",
  1833=>"111111111",
  1834=>"111111000",
  1835=>"110111111",
  1836=>"000000000",
  1837=>"000000000",
  1838=>"111000000",
  1839=>"000000000",
  1840=>"111111111",
  1841=>"101000101",
  1842=>"111111111",
  1843=>"111111110",
  1844=>"100000111",
  1845=>"111111011",
  1846=>"000100011",
  1847=>"000000000",
  1848=>"000000000",
  1849=>"000000111",
  1850=>"111001000",
  1851=>"100000000",
  1852=>"111111111",
  1853=>"000000000",
  1854=>"001011111",
  1855=>"111111010",
  1856=>"001001000",
  1857=>"000000110",
  1858=>"110000001",
  1859=>"000000000",
  1860=>"000101111",
  1861=>"111000000",
  1862=>"000000000",
  1863=>"000000000",
  1864=>"000000000",
  1865=>"011011000",
  1866=>"111111111",
  1867=>"000100000",
  1868=>"000000000",
  1869=>"111111111",
  1870=>"000000111",
  1871=>"000000000",
  1872=>"000000001",
  1873=>"000001000",
  1874=>"000100100",
  1875=>"110111111",
  1876=>"000000000",
  1877=>"111111011",
  1878=>"010010000",
  1879=>"000000000",
  1880=>"000000001",
  1881=>"111111111",
  1882=>"000000111",
  1883=>"111111111",
  1884=>"111111111",
  1885=>"010000000",
  1886=>"110010110",
  1887=>"100110111",
  1888=>"111111110",
  1889=>"000000000",
  1890=>"100100000",
  1891=>"101001111",
  1892=>"111111111",
  1893=>"000000100",
  1894=>"111000010",
  1895=>"000000001",
  1896=>"000001001",
  1897=>"000000100",
  1898=>"000111010",
  1899=>"000100101",
  1900=>"011010001",
  1901=>"000000111",
  1902=>"100000000",
  1903=>"000000000",
  1904=>"000000010",
  1905=>"111000000",
  1906=>"000010111",
  1907=>"110100111",
  1908=>"000000011",
  1909=>"001001001",
  1910=>"000000000",
  1911=>"111001000",
  1912=>"000000000",
  1913=>"100111111",
  1914=>"111111111",
  1915=>"000000000",
  1916=>"000000011",
  1917=>"000000000",
  1918=>"110111111",
  1919=>"000011111",
  1920=>"011001010",
  1921=>"001000001",
  1922=>"000000000",
  1923=>"000000100",
  1924=>"111110111",
  1925=>"000000000",
  1926=>"110010011",
  1927=>"000000000",
  1928=>"000000000",
  1929=>"111011111",
  1930=>"101001001",
  1931=>"101111111",
  1932=>"111111111",
  1933=>"100100100",
  1934=>"000000111",
  1935=>"000000000",
  1936=>"000000000",
  1937=>"111001000",
  1938=>"000000111",
  1939=>"010000001",
  1940=>"000000000",
  1941=>"000000000",
  1942=>"111111111",
  1943=>"111111111",
  1944=>"110111111",
  1945=>"111111101",
  1946=>"001001001",
  1947=>"000000111",
  1948=>"111110111",
  1949=>"111110000",
  1950=>"111111111",
  1951=>"111111110",
  1952=>"000000000",
  1953=>"111011001",
  1954=>"000000001",
  1955=>"000000000",
  1956=>"010000000",
  1957=>"111111111",
  1958=>"000000000",
  1959=>"111111111",
  1960=>"000000000",
  1961=>"111101000",
  1962=>"111000000",
  1963=>"111111111",
  1964=>"000000000",
  1965=>"000000000",
  1966=>"111111111",
  1967=>"001101111",
  1968=>"111011111",
  1969=>"000000000",
  1970=>"111101001",
  1971=>"000000000",
  1972=>"110010000",
  1973=>"111111111",
  1974=>"011001011",
  1975=>"111111111",
  1976=>"000100100",
  1977=>"111111001",
  1978=>"111110000",
  1979=>"010011000",
  1980=>"110000000",
  1981=>"000111110",
  1982=>"000001011",
  1983=>"111111111",
  1984=>"111101111",
  1985=>"111111111",
  1986=>"000000000",
  1987=>"000000000",
  1988=>"100100111",
  1989=>"111110111",
  1990=>"000000100",
  1991=>"111111101",
  1992=>"011000100",
  1993=>"000000111",
  1994=>"000000000",
  1995=>"111001000",
  1996=>"000000000",
  1997=>"011000011",
  1998=>"001000000",
  1999=>"000001001",
  2000=>"000010110",
  2001=>"111111010",
  2002=>"111111111",
  2003=>"000000000",
  2004=>"100000000",
  2005=>"001101111",
  2006=>"100000000",
  2007=>"011101000",
  2008=>"011011011",
  2009=>"100001001",
  2010=>"111111100",
  2011=>"111111011",
  2012=>"000000000",
  2013=>"010000000",
  2014=>"111111111",
  2015=>"000000110",
  2016=>"111111111",
  2017=>"000100100",
  2018=>"111000111",
  2019=>"010000000",
  2020=>"111000000",
  2021=>"111010000",
  2022=>"110000000",
  2023=>"100111111",
  2024=>"001000000",
  2025=>"110111001",
  2026=>"001000000",
  2027=>"000000000",
  2028=>"000000000",
  2029=>"000100110",
  2030=>"000110110",
  2031=>"111011100",
  2032=>"100101101",
  2033=>"011111000",
  2034=>"011011111",
  2035=>"000000000",
  2036=>"000000011",
  2037=>"111111111",
  2038=>"111111111",
  2039=>"011011001",
  2040=>"000000000",
  2041=>"010111011",
  2042=>"000000101",
  2043=>"111111110",
  2044=>"000111000",
  2045=>"000000001",
  2046=>"000000111",
  2047=>"111111111",
  2048=>"111011111",
  2049=>"111111001",
  2050=>"000000000",
  2051=>"111111000",
  2052=>"000000000",
  2053=>"111001111",
  2054=>"110000000",
  2055=>"111111110",
  2056=>"011011000",
  2057=>"100111111",
  2058=>"111100000",
  2059=>"111111111",
  2060=>"000100000",
  2061=>"111111000",
  2062=>"000000000",
  2063=>"000000000",
  2064=>"000000000",
  2065=>"110110011",
  2066=>"111111111",
  2067=>"111111111",
  2068=>"111111001",
  2069=>"000111111",
  2070=>"000000000",
  2071=>"011011111",
  2072=>"110000010",
  2073=>"100000000",
  2074=>"000000000",
  2075=>"110111111",
  2076=>"111111111",
  2077=>"111001100",
  2078=>"000000000",
  2079=>"100000000",
  2080=>"000001001",
  2081=>"111111111",
  2082=>"110110100",
  2083=>"000001111",
  2084=>"111101111",
  2085=>"010011111",
  2086=>"101101101",
  2087=>"111111010",
  2088=>"000000000",
  2089=>"000000000",
  2090=>"000000000",
  2091=>"111111111",
  2092=>"111011000",
  2093=>"111111110",
  2094=>"111111000",
  2095=>"100000000",
  2096=>"000010010",
  2097=>"111111001",
  2098=>"011011010",
  2099=>"011111110",
  2100=>"000000000",
  2101=>"000000000",
  2102=>"000000000",
  2103=>"000000000",
  2104=>"111110000",
  2105=>"111100010",
  2106=>"011011011",
  2107=>"000000000",
  2108=>"101101111",
  2109=>"111011000",
  2110=>"111100000",
  2111=>"000000000",
  2112=>"111111111",
  2113=>"101011001",
  2114=>"000000100",
  2115=>"111111110",
  2116=>"000000000",
  2117=>"111111111",
  2118=>"111111111",
  2119=>"000100111",
  2120=>"011001111",
  2121=>"111111111",
  2122=>"111111100",
  2123=>"111000000",
  2124=>"110000100",
  2125=>"000000000",
  2126=>"000000000",
  2127=>"111000100",
  2128=>"111011011",
  2129=>"000000000",
  2130=>"111111110",
  2131=>"000000001",
  2132=>"000000000",
  2133=>"000001101",
  2134=>"000000111",
  2135=>"111111111",
  2136=>"000001001",
  2137=>"000000101",
  2138=>"111111111",
  2139=>"100000100",
  2140=>"111111111",
  2141=>"000011111",
  2142=>"111111111",
  2143=>"111111111",
  2144=>"111111111",
  2145=>"111111111",
  2146=>"111111111",
  2147=>"111011001",
  2148=>"000000000",
  2149=>"000000001",
  2150=>"111111111",
  2151=>"111111111",
  2152=>"000000000",
  2153=>"000111100",
  2154=>"011011110",
  2155=>"111111111",
  2156=>"001000000",
  2157=>"000000000",
  2158=>"000000000",
  2159=>"000100000",
  2160=>"000000000",
  2161=>"000000111",
  2162=>"000000000",
  2163=>"111111111",
  2164=>"111111111",
  2165=>"000000000",
  2166=>"000000000",
  2167=>"111000010",
  2168=>"000000000",
  2169=>"000000000",
  2170=>"110000100",
  2171=>"000000000",
  2172=>"110111110",
  2173=>"000000000",
  2174=>"111101000",
  2175=>"100000000",
  2176=>"111111111",
  2177=>"000000000",
  2178=>"000000000",
  2179=>"000101111",
  2180=>"111111111",
  2181=>"111111100",
  2182=>"000000000",
  2183=>"000010010",
  2184=>"111111011",
  2185=>"000111111",
  2186=>"000000000",
  2187=>"111111011",
  2188=>"101111111",
  2189=>"111111111",
  2190=>"110111111",
  2191=>"111111111",
  2192=>"110000000",
  2193=>"000001001",
  2194=>"011111110",
  2195=>"011111111",
  2196=>"001000000",
  2197=>"111111111",
  2198=>"111110010",
  2199=>"001000000",
  2200=>"111110110",
  2201=>"000000010",
  2202=>"000000000",
  2203=>"011011000",
  2204=>"111101110",
  2205=>"000000000",
  2206=>"111111111",
  2207=>"000000000",
  2208=>"100000000",
  2209=>"000000000",
  2210=>"111111111",
  2211=>"001001001",
  2212=>"100001000",
  2213=>"000000000",
  2214=>"000000000",
  2215=>"000000000",
  2216=>"000111011",
  2217=>"101001111",
  2218=>"000000110",
  2219=>"111111111",
  2220=>"001001111",
  2221=>"110110100",
  2222=>"000000000",
  2223=>"000000000",
  2224=>"111001011",
  2225=>"000000000",
  2226=>"110111110",
  2227=>"110111101",
  2228=>"111111111",
  2229=>"000000110",
  2230=>"000101010",
  2231=>"111111111",
  2232=>"111111111",
  2233=>"000000000",
  2234=>"000000000",
  2235=>"000000111",
  2236=>"000111111",
  2237=>"111011000",
  2238=>"111100111",
  2239=>"110111111",
  2240=>"000000000",
  2241=>"001111111",
  2242=>"000000000",
  2243=>"000000000",
  2244=>"100111000",
  2245=>"110110111",
  2246=>"010000000",
  2247=>"101001000",
  2248=>"111111111",
  2249=>"001111111",
  2250=>"000000000",
  2251=>"100111111",
  2252=>"111111111",
  2253=>"001111111",
  2254=>"000000000",
  2255=>"011011011",
  2256=>"000001001",
  2257=>"111111111",
  2258=>"111111111",
  2259=>"000000000",
  2260=>"000000000",
  2261=>"011010110",
  2262=>"000000000",
  2263=>"001101111",
  2264=>"111111111",
  2265=>"011011010",
  2266=>"000000000",
  2267=>"000111110",
  2268=>"011001000",
  2269=>"111111111",
  2270=>"011111111",
  2271=>"111010010",
  2272=>"011111111",
  2273=>"000000000",
  2274=>"110110110",
  2275=>"010011011",
  2276=>"100110110",
  2277=>"000001001",
  2278=>"111001000",
  2279=>"111111011",
  2280=>"000000000",
  2281=>"111111111",
  2282=>"111111111",
  2283=>"101001111",
  2284=>"111111000",
  2285=>"000001001",
  2286=>"000000000",
  2287=>"000000001",
  2288=>"001011111",
  2289=>"111111111",
  2290=>"100100100",
  2291=>"111101110",
  2292=>"110010000",
  2293=>"110110111",
  2294=>"111111100",
  2295=>"111111111",
  2296=>"100100101",
  2297=>"111111111",
  2298=>"011011111",
  2299=>"000110100",
  2300=>"000000011",
  2301=>"111111111",
  2302=>"110000111",
  2303=>"111111111",
  2304=>"111111110",
  2305=>"111111111",
  2306=>"111111111",
  2307=>"111000000",
  2308=>"111111111",
  2309=>"000000000",
  2310=>"000000000",
  2311=>"111111111",
  2312=>"111000000",
  2313=>"000000000",
  2314=>"000000000",
  2315=>"010011011",
  2316=>"111101111",
  2317=>"000000000",
  2318=>"011111111",
  2319=>"110000000",
  2320=>"110000000",
  2321=>"000001001",
  2322=>"000000001",
  2323=>"111001001",
  2324=>"111111011",
  2325=>"111001000",
  2326=>"111111111",
  2327=>"000100000",
  2328=>"011001000",
  2329=>"000110001",
  2330=>"001001001",
  2331=>"000100111",
  2332=>"000000111",
  2333=>"111111111",
  2334=>"000000000",
  2335=>"000000000",
  2336=>"000000011",
  2337=>"000000000",
  2338=>"111100100",
  2339=>"000000000",
  2340=>"001001111",
  2341=>"111011011",
  2342=>"111111111",
  2343=>"000000000",
  2344=>"001001000",
  2345=>"000000000",
  2346=>"111100111",
  2347=>"111111111",
  2348=>"000010111",
  2349=>"000000000",
  2350=>"111010011",
  2351=>"000001100",
  2352=>"001111111",
  2353=>"000000000",
  2354=>"111011000",
  2355=>"000100100",
  2356=>"111111111",
  2357=>"110100100",
  2358=>"100000000",
  2359=>"111000001",
  2360=>"101001000",
  2361=>"111111111",
  2362=>"000111111",
  2363=>"000000000",
  2364=>"000000001",
  2365=>"111111111",
  2366=>"000000001",
  2367=>"111111111",
  2368=>"000000000",
  2369=>"111111111",
  2370=>"111111111",
  2371=>"111111111",
  2372=>"000000000",
  2373=>"111111101",
  2374=>"111111111",
  2375=>"000000000",
  2376=>"111111111",
  2377=>"001001000",
  2378=>"101000000",
  2379=>"000011011",
  2380=>"000000000",
  2381=>"111111110",
  2382=>"000000000",
  2383=>"011011111",
  2384=>"000011000",
  2385=>"000000100",
  2386=>"000000111",
  2387=>"111001001",
  2388=>"000000100",
  2389=>"000000001",
  2390=>"111111111",
  2391=>"111111111",
  2392=>"111111111",
  2393=>"111111111",
  2394=>"000000000",
  2395=>"110000100",
  2396=>"000000000",
  2397=>"111111111",
  2398=>"011001000",
  2399=>"000100110",
  2400=>"000000101",
  2401=>"000000000",
  2402=>"000000110",
  2403=>"101101111",
  2404=>"110110010",
  2405=>"000000000",
  2406=>"000000000",
  2407=>"110100000",
  2408=>"000110110",
  2409=>"111111111",
  2410=>"111000111",
  2411=>"111111111",
  2412=>"000000100",
  2413=>"111111111",
  2414=>"000000000",
  2415=>"000110110",
  2416=>"000000000",
  2417=>"010111111",
  2418=>"111111111",
  2419=>"000000000",
  2420=>"000000000",
  2421=>"000000000",
  2422=>"111111110",
  2423=>"000000000",
  2424=>"111111111",
  2425=>"000100000",
  2426=>"111111011",
  2427=>"100110110",
  2428=>"000000100",
  2429=>"111111111",
  2430=>"000000000",
  2431=>"000000000",
  2432=>"010001011",
  2433=>"000000111",
  2434=>"111111101",
  2435=>"000111111",
  2436=>"111111011",
  2437=>"111111000",
  2438=>"000000111",
  2439=>"111111111",
  2440=>"000000000",
  2441=>"000000100",
  2442=>"111111111",
  2443=>"111111111",
  2444=>"000101111",
  2445=>"111111111",
  2446=>"000001000",
  2447=>"000000000",
  2448=>"000000000",
  2449=>"111111111",
  2450=>"000000000",
  2451=>"000000000",
  2452=>"100111111",
  2453=>"000000000",
  2454=>"111111111",
  2455=>"100100000",
  2456=>"000000000",
  2457=>"111111111",
  2458=>"100100000",
  2459=>"111111111",
  2460=>"101111111",
  2461=>"110110111",
  2462=>"000000000",
  2463=>"001111110",
  2464=>"000000000",
  2465=>"010000000",
  2466=>"111111111",
  2467=>"011110110",
  2468=>"000000000",
  2469=>"111111111",
  2470=>"111111111",
  2471=>"010011111",
  2472=>"000000000",
  2473=>"000000100",
  2474=>"110110110",
  2475=>"000000000",
  2476=>"000101101",
  2477=>"001000000",
  2478=>"010000110",
  2479=>"011011111",
  2480=>"111111111",
  2481=>"111110000",
  2482=>"101001011",
  2483=>"000000000",
  2484=>"111111111",
  2485=>"100000000",
  2486=>"100000000",
  2487=>"111111111",
  2488=>"001001000",
  2489=>"000011010",
  2490=>"111011001",
  2491=>"111010011",
  2492=>"111111111",
  2493=>"000000000",
  2494=>"000000100",
  2495=>"100100111",
  2496=>"000000000",
  2497=>"001001000",
  2498=>"111111111",
  2499=>"110111011",
  2500=>"111000100",
  2501=>"111000100",
  2502=>"000000000",
  2503=>"001000001",
  2504=>"000000000",
  2505=>"111111111",
  2506=>"000000000",
  2507=>"000111000",
  2508=>"000000000",
  2509=>"111111110",
  2510=>"111111111",
  2511=>"000000000",
  2512=>"000000000",
  2513=>"101001111",
  2514=>"111111111",
  2515=>"111111111",
  2516=>"000001011",
  2517=>"111110111",
  2518=>"000000000",
  2519=>"000001011",
  2520=>"111001111",
  2521=>"111111010",
  2522=>"000000000",
  2523=>"110010000",
  2524=>"011011001",
  2525=>"111111111",
  2526=>"000000000",
  2527=>"100100100",
  2528=>"111111110",
  2529=>"000001111",
  2530=>"111111111",
  2531=>"000000000",
  2532=>"111011000",
  2533=>"000000000",
  2534=>"111111111",
  2535=>"111111111",
  2536=>"111101111",
  2537=>"000000000",
  2538=>"000001001",
  2539=>"100000001",
  2540=>"000000000",
  2541=>"001001001",
  2542=>"000000000",
  2543=>"010000000",
  2544=>"111111111",
  2545=>"110111111",
  2546=>"111111111",
  2547=>"000000000",
  2548=>"000000000",
  2549=>"000000000",
  2550=>"111111111",
  2551=>"000000000",
  2552=>"000111000",
  2553=>"011110110",
  2554=>"111110010",
  2555=>"111111000",
  2556=>"110110010",
  2557=>"000000000",
  2558=>"100100111",
  2559=>"111110100",
  2560=>"000000000",
  2561=>"111111111",
  2562=>"111111000",
  2563=>"000001011",
  2564=>"000000101",
  2565=>"011010000",
  2566=>"111001001",
  2567=>"000001111",
  2568=>"110110010",
  2569=>"110111111",
  2570=>"111110111",
  2571=>"110111111",
  2572=>"100100100",
  2573=>"100111010",
  2574=>"000001111",
  2575=>"000000000",
  2576=>"000000000",
  2577=>"000000011",
  2578=>"000010000",
  2579=>"011111111",
  2580=>"000000000",
  2581=>"000111111",
  2582=>"101110111",
  2583=>"110111111",
  2584=>"111111111",
  2585=>"010010111",
  2586=>"000111111",
  2587=>"111111011",
  2588=>"111111111",
  2589=>"000101011",
  2590=>"011011011",
  2591=>"100100110",
  2592=>"011001000",
  2593=>"000000000",
  2594=>"111111110",
  2595=>"111111111",
  2596=>"111100100",
  2597=>"000000001",
  2598=>"111111011",
  2599=>"000100000",
  2600=>"001000000",
  2601=>"000000100",
  2602=>"000000100",
  2603=>"011001001",
  2604=>"111111110",
  2605=>"101100111",
  2606=>"000000000",
  2607=>"111110000",
  2608=>"111011111",
  2609=>"000000000",
  2610=>"111111111",
  2611=>"010111111",
  2612=>"000000100",
  2613=>"100110111",
  2614=>"000111111",
  2615=>"001001100",
  2616=>"011111000",
  2617=>"000000000",
  2618=>"111111111",
  2619=>"010111111",
  2620=>"000000000",
  2621=>"000010100",
  2622=>"111111111",
  2623=>"111111111",
  2624=>"111111001",
  2625=>"111111000",
  2626=>"111111111",
  2627=>"111110110",
  2628=>"110100001",
  2629=>"000000100",
  2630=>"100000100",
  2631=>"111111001",
  2632=>"111111010",
  2633=>"001000000",
  2634=>"011000000",
  2635=>"100000000",
  2636=>"000000111",
  2637=>"101100111",
  2638=>"011010100",
  2639=>"000111111",
  2640=>"001000111",
  2641=>"111111100",
  2642=>"110111111",
  2643=>"111001000",
  2644=>"000000000",
  2645=>"110110110",
  2646=>"111111100",
  2647=>"111110000",
  2648=>"010010100",
  2649=>"000001111",
  2650=>"111101000",
  2651=>"110110100",
  2652=>"001000011",
  2653=>"111101000",
  2654=>"000001100",
  2655=>"111111111",
  2656=>"000000000",
  2657=>"111011001",
  2658=>"111000101",
  2659=>"000000000",
  2660=>"000000000",
  2661=>"001001111",
  2662=>"011111111",
  2663=>"111100001",
  2664=>"000000000",
  2665=>"000000000",
  2666=>"110111001",
  2667=>"111111111",
  2668=>"000000000",
  2669=>"000000000",
  2670=>"000000101",
  2671=>"101001100",
  2672=>"011011000",
  2673=>"000000001",
  2674=>"001001111",
  2675=>"001001000",
  2676=>"000000100",
  2677=>"011001000",
  2678=>"111111111",
  2679=>"111111000",
  2680=>"111111111",
  2681=>"000101101",
  2682=>"000000000",
  2683=>"000011111",
  2684=>"001011011",
  2685=>"000000000",
  2686=>"111011010",
  2687=>"001001000",
  2688=>"000000000",
  2689=>"101000000",
  2690=>"000000111",
  2691=>"011100110",
  2692=>"110111011",
  2693=>"111111111",
  2694=>"000001110",
  2695=>"000000000",
  2696=>"111011000",
  2697=>"111111111",
  2698=>"111111111",
  2699=>"010111001",
  2700=>"000001111",
  2701=>"011011100",
  2702=>"011011000",
  2703=>"111111011",
  2704=>"111111111",
  2705=>"111111111",
  2706=>"011000100",
  2707=>"000001101",
  2708=>"111111110",
  2709=>"100000000",
  2710=>"111111111",
  2711=>"111101000",
  2712=>"110100111",
  2713=>"110110110",
  2714=>"111100000",
  2715=>"111111100",
  2716=>"000100000",
  2717=>"011111011",
  2718=>"000110000",
  2719=>"000000000",
  2720=>"000100010",
  2721=>"000000000",
  2722=>"000100110",
  2723=>"011000000",
  2724=>"000000000",
  2725=>"011111111",
  2726=>"111101111",
  2727=>"110010110",
  2728=>"000000110",
  2729=>"111000000",
  2730=>"111101101",
  2731=>"000111111",
  2732=>"100110111",
  2733=>"101001001",
  2734=>"011111111",
  2735=>"111110111",
  2736=>"000001011",
  2737=>"011111111",
  2738=>"000000000",
  2739=>"111000000",
  2740=>"101111111",
  2741=>"110000000",
  2742=>"000000001",
  2743=>"111111111",
  2744=>"100100100",
  2745=>"111111111",
  2746=>"000000000",
  2747=>"000001011",
  2748=>"000100100",
  2749=>"111111111",
  2750=>"100000000",
  2751=>"001000111",
  2752=>"101100100",
  2753=>"111000000",
  2754=>"101111111",
  2755=>"110111111",
  2756=>"111111000",
  2757=>"000000010",
  2758=>"000000000",
  2759=>"000000110",
  2760=>"000100000",
  2761=>"111101100",
  2762=>"000000011",
  2763=>"000000000",
  2764=>"000000000",
  2765=>"110111011",
  2766=>"000010110",
  2767=>"100111111",
  2768=>"100000000",
  2769=>"110111111",
  2770=>"100000000",
  2771=>"001001101",
  2772=>"111000100",
  2773=>"010110100",
  2774=>"000000111",
  2775=>"001000001",
  2776=>"000001111",
  2777=>"000000000",
  2778=>"011111111",
  2779=>"011111111",
  2780=>"001000000",
  2781=>"000000000",
  2782=>"111100100",
  2783=>"000000100",
  2784=>"111111111",
  2785=>"001000001",
  2786=>"111111111",
  2787=>"000000000",
  2788=>"111111001",
  2789=>"011111011",
  2790=>"010000000",
  2791=>"111111100",
  2792=>"000000000",
  2793=>"000000010",
  2794=>"011010110",
  2795=>"101011001",
  2796=>"010110010",
  2797=>"111111110",
  2798=>"000100111",
  2799=>"100000000",
  2800=>"111000000",
  2801=>"000000000",
  2802=>"111111111",
  2803=>"111111110",
  2804=>"000000001",
  2805=>"111111111",
  2806=>"000110110",
  2807=>"000111000",
  2808=>"000000000",
  2809=>"000000100",
  2810=>"000111111",
  2811=>"000111110",
  2812=>"111001111",
  2813=>"100000100",
  2814=>"111111110",
  2815=>"111111100",
  2816=>"000000111",
  2817=>"010011011",
  2818=>"011101000",
  2819=>"000000000",
  2820=>"111100100",
  2821=>"111111111",
  2822=>"111111111",
  2823=>"000000001",
  2824=>"011111110",
  2825=>"011011111",
  2826=>"000000000",
  2827=>"111111111",
  2828=>"100110110",
  2829=>"000000000",
  2830=>"000001101",
  2831=>"111111111",
  2832=>"111001000",
  2833=>"000111000",
  2834=>"000000000",
  2835=>"000000111",
  2836=>"011011001",
  2837=>"100111111",
  2838=>"011001001",
  2839=>"000101110",
  2840=>"111111111",
  2841=>"110111000",
  2842=>"111111111",
  2843=>"000100111",
  2844=>"010110110",
  2845=>"011000000",
  2846=>"111101111",
  2847=>"111111111",
  2848=>"000000111",
  2849=>"001111111",
  2850=>"000000000",
  2851=>"111111000",
  2852=>"000101111",
  2853=>"111000000",
  2854=>"000000000",
  2855=>"000100101",
  2856=>"010000100",
  2857=>"000000000",
  2858=>"111111101",
  2859=>"111101111",
  2860=>"111111001",
  2861=>"000001101",
  2862=>"111111001",
  2863=>"000100110",
  2864=>"000000000",
  2865=>"101100111",
  2866=>"111111111",
  2867=>"111100111",
  2868=>"000000000",
  2869=>"000000000",
  2870=>"000100111",
  2871=>"000011000",
  2872=>"000000000",
  2873=>"111111001",
  2874=>"000000000",
  2875=>"000010011",
  2876=>"101100101",
  2877=>"000000010",
  2878=>"010100000",
  2879=>"001101101",
  2880=>"000100111",
  2881=>"111111001",
  2882=>"000110000",
  2883=>"000000000",
  2884=>"011111111",
  2885=>"111000000",
  2886=>"000000000",
  2887=>"111111111",
  2888=>"110111111",
  2889=>"111000000",
  2890=>"111000000",
  2891=>"111110100",
  2892=>"111111111",
  2893=>"100101000",
  2894=>"111111111",
  2895=>"110111110",
  2896=>"100110110",
  2897=>"111110110",
  2898=>"111110111",
  2899=>"001001001",
  2900=>"110111111",
  2901=>"001001111",
  2902=>"111111100",
  2903=>"111111111",
  2904=>"000000000",
  2905=>"000111111",
  2906=>"000000000",
  2907=>"000111111",
  2908=>"000100110",
  2909=>"000000000",
  2910=>"111000000",
  2911=>"111111111",
  2912=>"001000000",
  2913=>"111101111",
  2914=>"000000000",
  2915=>"111111111",
  2916=>"011111110",
  2917=>"000000011",
  2918=>"111100111",
  2919=>"000000000",
  2920=>"001001011",
  2921=>"010110111",
  2922=>"000000000",
  2923=>"111111111",
  2924=>"100001001",
  2925=>"111001000",
  2926=>"111111111",
  2927=>"000000000",
  2928=>"111111111",
  2929=>"000001111",
  2930=>"111111000",
  2931=>"000000111",
  2932=>"000000000",
  2933=>"000000001",
  2934=>"000000010",
  2935=>"000100110",
  2936=>"011000111",
  2937=>"000000000",
  2938=>"111111111",
  2939=>"111101111",
  2940=>"111001111",
  2941=>"111001111",
  2942=>"100000000",
  2943=>"000100100",
  2944=>"111111011",
  2945=>"001000000",
  2946=>"001001001",
  2947=>"000000000",
  2948=>"111111111",
  2949=>"011001000",
  2950=>"111111110",
  2951=>"111111111",
  2952=>"000000101",
  2953=>"111111110",
  2954=>"111110111",
  2955=>"111111111",
  2956=>"000000000",
  2957=>"001001000",
  2958=>"000000110",
  2959=>"000000111",
  2960=>"111111111",
  2961=>"111111111",
  2962=>"000000000",
  2963=>"001001001",
  2964=>"000000111",
  2965=>"111011101",
  2966=>"000000111",
  2967=>"010010000",
  2968=>"110100111",
  2969=>"101001000",
  2970=>"111101111",
  2971=>"000000010",
  2972=>"000000000",
  2973=>"000000000",
  2974=>"000011000",
  2975=>"100100110",
  2976=>"111111111",
  2977=>"111111111",
  2978=>"011011000",
  2979=>"000100101",
  2980=>"011011011",
  2981=>"111111010",
  2982=>"110000000",
  2983=>"110011011",
  2984=>"000000000",
  2985=>"011111111",
  2986=>"000000000",
  2987=>"000000000",
  2988=>"111111111",
  2989=>"001000010",
  2990=>"101100000",
  2991=>"111101100",
  2992=>"110111011",
  2993=>"100111100",
  2994=>"111000100",
  2995=>"111000100",
  2996=>"000000000",
  2997=>"000000100",
  2998=>"000000000",
  2999=>"111111111",
  3000=>"000000000",
  3001=>"111111100",
  3002=>"101111111",
  3003=>"101101001",
  3004=>"000011111",
  3005=>"110000000",
  3006=>"001000000",
  3007=>"011011010",
  3008=>"111111110",
  3009=>"111111111",
  3010=>"000011011",
  3011=>"111111111",
  3012=>"000000010",
  3013=>"100110110",
  3014=>"000000000",
  3015=>"001011010",
  3016=>"000000000",
  3017=>"111111010",
  3018=>"001111111",
  3019=>"011111000",
  3020=>"000000000",
  3021=>"011111111",
  3022=>"000000000",
  3023=>"111111000",
  3024=>"100110110",
  3025=>"010111111",
  3026=>"101001000",
  3027=>"000000100",
  3028=>"101100111",
  3029=>"100101111",
  3030=>"000000000",
  3031=>"010010000",
  3032=>"000010011",
  3033=>"111010000",
  3034=>"010000000",
  3035=>"111111111",
  3036=>"001111111",
  3037=>"000111000",
  3038=>"100000000",
  3039=>"011011111",
  3040=>"000000000",
  3041=>"101110110",
  3042=>"111111111",
  3043=>"000001111",
  3044=>"010010110",
  3045=>"110110100",
  3046=>"000000000",
  3047=>"000100100",
  3048=>"111111111",
  3049=>"111111111",
  3050=>"000010000",
  3051=>"000000000",
  3052=>"000000000",
  3053=>"000000100",
  3054=>"010111111",
  3055=>"000110110",
  3056=>"000000000",
  3057=>"110111110",
  3058=>"011001000",
  3059=>"000000000",
  3060=>"001001111",
  3061=>"111111100",
  3062=>"111111111",
  3063=>"000000001",
  3064=>"010010011",
  3065=>"100100100",
  3066=>"010000000",
  3067=>"000000100",
  3068=>"111111111",
  3069=>"001011111",
  3070=>"000001001",
  3071=>"000000000",
  3072=>"001011001",
  3073=>"000000000",
  3074=>"000001111",
  3075=>"110111101",
  3076=>"100000000",
  3077=>"110111110",
  3078=>"100111011",
  3079=>"111001101",
  3080=>"111001111",
  3081=>"101000000",
  3082=>"000000000",
  3083=>"000000110",
  3084=>"000000000",
  3085=>"000000111",
  3086=>"110001000",
  3087=>"111111111",
  3088=>"000000000",
  3089=>"100110111",
  3090=>"111111000",
  3091=>"111110000",
  3092=>"001001101",
  3093=>"000000000",
  3094=>"111111000",
  3095=>"000001001",
  3096=>"100000100",
  3097=>"111101111",
  3098=>"000001001",
  3099=>"100110100",
  3100=>"000000000",
  3101=>"111111000",
  3102=>"100101111",
  3103=>"000000111",
  3104=>"001001000",
  3105=>"110111111",
  3106=>"100001111",
  3107=>"111111111",
  3108=>"000000000",
  3109=>"000000111",
  3110=>"110110111",
  3111=>"000000101",
  3112=>"000000000",
  3113=>"111111111",
  3114=>"000001000",
  3115=>"000111110",
  3116=>"001000000",
  3117=>"111111000",
  3118=>"000000110",
  3119=>"001000000",
  3120=>"101001001",
  3121=>"000000111",
  3122=>"000001100",
  3123=>"100000000",
  3124=>"000001000",
  3125=>"000011110",
  3126=>"001101111",
  3127=>"111111111",
  3128=>"001111111",
  3129=>"111111111",
  3130=>"110011111",
  3131=>"000000000",
  3132=>"001000000",
  3133=>"100111011",
  3134=>"100110100",
  3135=>"101001001",
  3136=>"000000100",
  3137=>"110100111",
  3138=>"000000010",
  3139=>"111100100",
  3140=>"000000000",
  3141=>"111111111",
  3142=>"111111111",
  3143=>"000000000",
  3144=>"000111111",
  3145=>"101111111",
  3146=>"000000000",
  3147=>"111110010",
  3148=>"000001001",
  3149=>"000000001",
  3150=>"000000010",
  3151=>"101111111",
  3152=>"000000000",
  3153=>"110110000",
  3154=>"001111111",
  3155=>"000000100",
  3156=>"000010010",
  3157=>"000001101",
  3158=>"000000100",
  3159=>"111111011",
  3160=>"111111101",
  3161=>"111101111",
  3162=>"111111111",
  3163=>"000010111",
  3164=>"111000111",
  3165=>"111111111",
  3166=>"101111111",
  3167=>"000111111",
  3168=>"111000011",
  3169=>"110111101",
  3170=>"111111101",
  3171=>"011111111",
  3172=>"111111101",
  3173=>"111100100",
  3174=>"000000111",
  3175=>"111111111",
  3176=>"111000011",
  3177=>"011000101",
  3178=>"111111111",
  3179=>"000101100",
  3180=>"001011111",
  3181=>"000111010",
  3182=>"000000111",
  3183=>"001001101",
  3184=>"111101101",
  3185=>"000111111",
  3186=>"000000000",
  3187=>"010110001",
  3188=>"111011000",
  3189=>"000000100",
  3190=>"111111111",
  3191=>"111111111",
  3192=>"111011011",
  3193=>"100101001",
  3194=>"111100000",
  3195=>"111011011",
  3196=>"100110111",
  3197=>"001011111",
  3198=>"000000000",
  3199=>"000000000",
  3200=>"000000000",
  3201=>"111111001",
  3202=>"000101111",
  3203=>"111001001",
  3204=>"000000000",
  3205=>"110101001",
  3206=>"000000001",
  3207=>"111111101",
  3208=>"000000000",
  3209=>"000100100",
  3210=>"110111111",
  3211=>"000000000",
  3212=>"100011111",
  3213=>"000000000",
  3214=>"111111111",
  3215=>"110111000",
  3216=>"000001111",
  3217=>"000000001",
  3218=>"000010111",
  3219=>"001001000",
  3220=>"000010100",
  3221=>"000000011",
  3222=>"111011010",
  3223=>"100000000",
  3224=>"111011111",
  3225=>"000000000",
  3226=>"000000000",
  3227=>"111111111",
  3228=>"011001001",
  3229=>"011001001",
  3230=>"001001001",
  3231=>"000100000",
  3232=>"000000100",
  3233=>"110000110",
  3234=>"110111111",
  3235=>"111111111",
  3236=>"000101011",
  3237=>"111111110",
  3238=>"111110000",
  3239=>"011111111",
  3240=>"000000000",
  3241=>"010010000",
  3242=>"000000000",
  3243=>"000010111",
  3244=>"111111111",
  3245=>"000000110",
  3246=>"111111101",
  3247=>"000000000",
  3248=>"000111111",
  3249=>"100100100",
  3250=>"110111010",
  3251=>"000000000",
  3252=>"000001001",
  3253=>"010000000",
  3254=>"000000010",
  3255=>"011111111",
  3256=>"111110000",
  3257=>"111111111",
  3258=>"101000000",
  3259=>"001001111",
  3260=>"000001000",
  3261=>"001001111",
  3262=>"000000000",
  3263=>"111111111",
  3264=>"111111111",
  3265=>"111111111",
  3266=>"111111111",
  3267=>"111111111",
  3268=>"111111111",
  3269=>"000000000",
  3270=>"011111011",
  3271=>"000111111",
  3272=>"111010110",
  3273=>"000000001",
  3274=>"000000000",
  3275=>"001100111",
  3276=>"111101101",
  3277=>"000010010",
  3278=>"000000111",
  3279=>"000000000",
  3280=>"000000000",
  3281=>"000000010",
  3282=>"011011111",
  3283=>"000000000",
  3284=>"000000000",
  3285=>"111000001",
  3286=>"011000000",
  3287=>"000000001",
  3288=>"100001111",
  3289=>"111011000",
  3290=>"111111111",
  3291=>"000111011",
  3292=>"000000111",
  3293=>"101101111",
  3294=>"111111000",
  3295=>"001011110",
  3296=>"000000000",
  3297=>"111111111",
  3298=>"111001000",
  3299=>"000000000",
  3300=>"111111010",
  3301=>"110000000",
  3302=>"111111111",
  3303=>"001000000",
  3304=>"000000000",
  3305=>"111000001",
  3306=>"001000001",
  3307=>"010000000",
  3308=>"111101000",
  3309=>"011111111",
  3310=>"111000000",
  3311=>"000000000",
  3312=>"100000000",
  3313=>"001011001",
  3314=>"001111111",
  3315=>"000011011",
  3316=>"000111111",
  3317=>"000100110",
  3318=>"011111110",
  3319=>"001000100",
  3320=>"001111111",
  3321=>"000110100",
  3322=>"101111111",
  3323=>"111111110",
  3324=>"000010000",
  3325=>"001001101",
  3326=>"100110000",
  3327=>"100111011",
  3328=>"111111000",
  3329=>"000100111",
  3330=>"110111111",
  3331=>"111111101",
  3332=>"101111111",
  3333=>"010001010",
  3334=>"111011001",
  3335=>"101101101",
  3336=>"111111111",
  3337=>"100100100",
  3338=>"111111110",
  3339=>"111111000",
  3340=>"000000100",
  3341=>"111110000",
  3342=>"100000000",
  3343=>"000110110",
  3344=>"000111111",
  3345=>"000000111",
  3346=>"011111111",
  3347=>"111111111",
  3348=>"000000111",
  3349=>"000000000",
  3350=>"100100111",
  3351=>"111111111",
  3352=>"011001000",
  3353=>"001000011",
  3354=>"101111111",
  3355=>"000000000",
  3356=>"111111111",
  3357=>"111111111",
  3358=>"011001000",
  3359=>"111011111",
  3360=>"001011111",
  3361=>"111111010",
  3362=>"110111111",
  3363=>"000000001",
  3364=>"000010000",
  3365=>"100100101",
  3366=>"000000000",
  3367=>"000111111",
  3368=>"100110010",
  3369=>"111011000",
  3370=>"111111111",
  3371=>"011011111",
  3372=>"000111100",
  3373=>"111111111",
  3374=>"000000111",
  3375=>"000100000",
  3376=>"000000111",
  3377=>"000000000",
  3378=>"000000000",
  3379=>"000000111",
  3380=>"010110010",
  3381=>"000100110",
  3382=>"000000110",
  3383=>"011000000",
  3384=>"000111111",
  3385=>"111000111",
  3386=>"000100100",
  3387=>"000000000",
  3388=>"001001111",
  3389=>"100000111",
  3390=>"000000100",
  3391=>"000000001",
  3392=>"000000000",
  3393=>"100011011",
  3394=>"111111111",
  3395=>"111111111",
  3396=>"000000000",
  3397=>"111111100",
  3398=>"111111111",
  3399=>"000000100",
  3400=>"000110111",
  3401=>"000000000",
  3402=>"000000001",
  3403=>"011001001",
  3404=>"000011000",
  3405=>"000000010",
  3406=>"000000000",
  3407=>"100110110",
  3408=>"001001100",
  3409=>"000110111",
  3410=>"111111111",
  3411=>"101101111",
  3412=>"000001001",
  3413=>"011011011",
  3414=>"000001110",
  3415=>"000000011",
  3416=>"111111111",
  3417=>"111001111",
  3418=>"000000101",
  3419=>"111111100",
  3420=>"111111111",
  3421=>"000000011",
  3422=>"000110111",
  3423=>"111111111",
  3424=>"000000100",
  3425=>"111111011",
  3426=>"000110111",
  3427=>"111101101",
  3428=>"000110110",
  3429=>"001101111",
  3430=>"000000010",
  3431=>"111111011",
  3432=>"100100110",
  3433=>"111111111",
  3434=>"000001001",
  3435=>"000000000",
  3436=>"111111111",
  3437=>"001111111",
  3438=>"000001100",
  3439=>"000000000",
  3440=>"000000000",
  3441=>"000011010",
  3442=>"110110111",
  3443=>"100111111",
  3444=>"000000000",
  3445=>"000000000",
  3446=>"111001101",
  3447=>"000000000",
  3448=>"111111111",
  3449=>"000000000",
  3450=>"000000001",
  3451=>"101111001",
  3452=>"111111101",
  3453=>"001101001",
  3454=>"101101101",
  3455=>"101000000",
  3456=>"001001111",
  3457=>"000010101",
  3458=>"111111111",
  3459=>"000110111",
  3460=>"011111000",
  3461=>"110111110",
  3462=>"011111111",
  3463=>"000000010",
  3464=>"000001111",
  3465=>"000000110",
  3466=>"110110110",
  3467=>"110110000",
  3468=>"000000100",
  3469=>"110110110",
  3470=>"100111111",
  3471=>"011011000",
  3472=>"100111111",
  3473=>"000000000",
  3474=>"111111111",
  3475=>"000000011",
  3476=>"101001000",
  3477=>"000000000",
  3478=>"111110000",
  3479=>"100100010",
  3480=>"111000100",
  3481=>"111111110",
  3482=>"110110000",
  3483=>"111011111",
  3484=>"111111111",
  3485=>"100110111",
  3486=>"001000000",
  3487=>"111111000",
  3488=>"000000000",
  3489=>"001011011",
  3490=>"111101101",
  3491=>"000000011",
  3492=>"111111111",
  3493=>"111111111",
  3494=>"000000011",
  3495=>"000000011",
  3496=>"111111111",
  3497=>"000010000",
  3498=>"111111111",
  3499=>"100100111",
  3500=>"000000000",
  3501=>"111111111",
  3502=>"111111111",
  3503=>"111111010",
  3504=>"000100011",
  3505=>"000001000",
  3506=>"000000000",
  3507=>"000110010",
  3508=>"000001111",
  3509=>"000000001",
  3510=>"111111111",
  3511=>"000000000",
  3512=>"111111111",
  3513=>"111110000",
  3514=>"111110000",
  3515=>"001001111",
  3516=>"111111011",
  3517=>"111111111",
  3518=>"010000000",
  3519=>"100100111",
  3520=>"000000000",
  3521=>"111111111",
  3522=>"000000000",
  3523=>"111101000",
  3524=>"000000101",
  3525=>"101111111",
  3526=>"111011000",
  3527=>"001111111",
  3528=>"100000000",
  3529=>"100100000",
  3530=>"100110100",
  3531=>"010111111",
  3532=>"010111111",
  3533=>"000100000",
  3534=>"111111101",
  3535=>"010000100",
  3536=>"001000001",
  3537=>"100110111",
  3538=>"000101001",
  3539=>"111001000",
  3540=>"000000000",
  3541=>"011111000",
  3542=>"111111001",
  3543=>"101101001",
  3544=>"111111100",
  3545=>"110111000",
  3546=>"001000001",
  3547=>"100100111",
  3548=>"111111111",
  3549=>"100000000",
  3550=>"000000101",
  3551=>"001101100",
  3552=>"100101101",
  3553=>"110110111",
  3554=>"101000000",
  3555=>"111111111",
  3556=>"001011111",
  3557=>"100100100",
  3558=>"000000000",
  3559=>"000001001",
  3560=>"110010001",
  3561=>"101001111",
  3562=>"111000001",
  3563=>"100000110",
  3564=>"001001000",
  3565=>"010001001",
  3566=>"111111111",
  3567=>"100000000",
  3568=>"100100100",
  3569=>"111101111",
  3570=>"110000000",
  3571=>"001001001",
  3572=>"001001000",
  3573=>"000000000",
  3574=>"000000000",
  3575=>"000001101",
  3576=>"111000000",
  3577=>"001001001",
  3578=>"000000000",
  3579=>"001000000",
  3580=>"000000101",
  3581=>"101011011",
  3582=>"000000000",
  3583=>"100000000",
  3584=>"111111111",
  3585=>"100000001",
  3586=>"101001000",
  3587=>"111111111",
  3588=>"110111111",
  3589=>"100100110",
  3590=>"000010010",
  3591=>"111111111",
  3592=>"111001000",
  3593=>"000001001",
  3594=>"111001000",
  3595=>"111100001",
  3596=>"000000000",
  3597=>"111111010",
  3598=>"011011011",
  3599=>"000000000",
  3600=>"001001001",
  3601=>"011111111",
  3602=>"100001111",
  3603=>"001000000",
  3604=>"000000011",
  3605=>"000000001",
  3606=>"000001000",
  3607=>"001000100",
  3608=>"011001001",
  3609=>"110010010",
  3610=>"011011000",
  3611=>"111011010",
  3612=>"011000000",
  3613=>"000000000",
  3614=>"011011011",
  3615=>"010011000",
  3616=>"110110000",
  3617=>"111011000",
  3618=>"000000100",
  3619=>"111111111",
  3620=>"011011011",
  3621=>"110011011",
  3622=>"000000001",
  3623=>"000000000",
  3624=>"111011010",
  3625=>"000000000",
  3626=>"000000000",
  3627=>"000000100",
  3628=>"111111111",
  3629=>"011111111",
  3630=>"100101001",
  3631=>"000000111",
  3632=>"000000000",
  3633=>"010010010",
  3634=>"110110110",
  3635=>"111111011",
  3636=>"110110111",
  3637=>"011011010",
  3638=>"001000000",
  3639=>"001111011",
  3640=>"011000100",
  3641=>"000000011",
  3642=>"000000111",
  3643=>"101101100",
  3644=>"110110111",
  3645=>"110010011",
  3646=>"111110010",
  3647=>"000000001",
  3648=>"000000000",
  3649=>"001000000",
  3650=>"001111111",
  3651=>"000000100",
  3652=>"011011000",
  3653=>"000000010",
  3654=>"010000000",
  3655=>"000000011",
  3656=>"000110100",
  3657=>"001001111",
  3658=>"001001101",
  3659=>"001000000",
  3660=>"000000000",
  3661=>"111111111",
  3662=>"111100101",
  3663=>"000000000",
  3664=>"110010111",
  3665=>"001001101",
  3666=>"101000010",
  3667=>"110110110",
  3668=>"110000110",
  3669=>"000000000",
  3670=>"100101101",
  3671=>"010000000",
  3672=>"000011000",
  3673=>"000000000",
  3674=>"100100000",
  3675=>"011000000",
  3676=>"001101000",
  3677=>"001000100",
  3678=>"100000110",
  3679=>"110000000",
  3680=>"000110010",
  3681=>"111101001",
  3682=>"100100100",
  3683=>"111011000",
  3684=>"000001011",
  3685=>"101001000",
  3686=>"111000000",
  3687=>"000000101",
  3688=>"011010000",
  3689=>"001000001",
  3690=>"010111010",
  3691=>"110111111",
  3692=>"111011000",
  3693=>"110110011",
  3694=>"001001101",
  3695=>"101001000",
  3696=>"000001001",
  3697=>"000000101",
  3698=>"101000000",
  3699=>"111000000",
  3700=>"111001000",
  3701=>"001011010",
  3702=>"111111111",
  3703=>"111111111",
  3704=>"111101000",
  3705=>"111111011",
  3706=>"001101111",
  3707=>"101101001",
  3708=>"100101101",
  3709=>"010000000",
  3710=>"111111111",
  3711=>"110110111",
  3712=>"111111111",
  3713=>"000000101",
  3714=>"111111111",
  3715=>"011011011",
  3716=>"010000000",
  3717=>"000100111",
  3718=>"011011111",
  3719=>"000110110",
  3720=>"110110110",
  3721=>"101101101",
  3722=>"001000000",
  3723=>"010110100",
  3724=>"100100110",
  3725=>"000001111",
  3726=>"000000001",
  3727=>"110110000",
  3728=>"100000000",
  3729=>"110110000",
  3730=>"111010010",
  3731=>"111110010",
  3732=>"100100000",
  3733=>"101100111",
  3734=>"101101100",
  3735=>"001000000",
  3736=>"000000000",
  3737=>"000000000",
  3738=>"111001000",
  3739=>"101100000",
  3740=>"001000000",
  3741=>"101101111",
  3742=>"101000111",
  3743=>"000000000",
  3744=>"000000010",
  3745=>"110110110",
  3746=>"111110000",
  3747=>"000101111",
  3748=>"110110000",
  3749=>"111111111",
  3750=>"110110110",
  3751=>"010010100",
  3752=>"100100101",
  3753=>"000001001",
  3754=>"110000000",
  3755=>"111111111",
  3756=>"011001101",
  3757=>"001000100",
  3758=>"111111110",
  3759=>"000000000",
  3760=>"111111010",
  3761=>"001000000",
  3762=>"111111011",
  3763=>"010010000",
  3764=>"010000111",
  3765=>"000001000",
  3766=>"110000000",
  3767=>"111111111",
  3768=>"001000001",
  3769=>"001111000",
  3770=>"001001001",
  3771=>"110010000",
  3772=>"100101100",
  3773=>"001000000",
  3774=>"100101001",
  3775=>"001001001",
  3776=>"000000000",
  3777=>"001001001",
  3778=>"111111111",
  3779=>"000100100",
  3780=>"111100111",
  3781=>"000000011",
  3782=>"001000011",
  3783=>"111101111",
  3784=>"110111111",
  3785=>"000000110",
  3786=>"000000001",
  3787=>"110111011",
  3788=>"000010000",
  3789=>"100110100",
  3790=>"111011010",
  3791=>"101101111",
  3792=>"100000000",
  3793=>"101101111",
  3794=>"000000100",
  3795=>"000000111",
  3796=>"000110111",
  3797=>"111001001",
  3798=>"001001101",
  3799=>"000010000",
  3800=>"111111100",
  3801=>"000000000",
  3802=>"111100000",
  3803=>"000000100",
  3804=>"111111111",
  3805=>"101001001",
  3806=>"111111111",
  3807=>"101001011",
  3808=>"111000000",
  3809=>"111111111",
  3810=>"101100100",
  3811=>"000000000",
  3812=>"000001101",
  3813=>"110010110",
  3814=>"000000000",
  3815=>"110111000",
  3816=>"101111000",
  3817=>"111111011",
  3818=>"111111010",
  3819=>"110010000",
  3820=>"001000000",
  3821=>"101111111",
  3822=>"111110110",
  3823=>"110111111",
  3824=>"000111011",
  3825=>"001001111",
  3826=>"000010000",
  3827=>"110110110",
  3828=>"000000000",
  3829=>"000000000",
  3830=>"100110111",
  3831=>"101111111",
  3832=>"000110111",
  3833=>"000000100",
  3834=>"110110110",
  3835=>"000000100",
  3836=>"110110110",
  3837=>"100000001",
  3838=>"111101001",
  3839=>"000011001",
  3840=>"000000000",
  3841=>"011011011",
  3842=>"000010001",
  3843=>"000000011",
  3844=>"010010000",
  3845=>"001001011",
  3846=>"000001111",
  3847=>"000001100",
  3848=>"111110111",
  3849=>"000000000",
  3850=>"101101001",
  3851=>"111111010",
  3852=>"100000100",
  3853=>"110110111",
  3854=>"000000000",
  3855=>"000000000",
  3856=>"000110111",
  3857=>"110011011",
  3858=>"101001111",
  3859=>"000110110",
  3860=>"001101000",
  3861=>"000101001",
  3862=>"110110110",
  3863=>"000000000",
  3864=>"111111111",
  3865=>"101010010",
  3866=>"100000011",
  3867=>"000111011",
  3868=>"111111011",
  3869=>"101000000",
  3870=>"000000000",
  3871=>"111110111",
  3872=>"110110011",
  3873=>"011000000",
  3874=>"011011000",
  3875=>"000000110",
  3876=>"111100000",
  3877=>"000000110",
  3878=>"011011011",
  3879=>"111001001",
  3880=>"111101101",
  3881=>"000000001",
  3882=>"110010011",
  3883=>"011000000",
  3884=>"000000000",
  3885=>"111111010",
  3886=>"101000001",
  3887=>"100000000",
  3888=>"000100100",
  3889=>"111111001",
  3890=>"111111111",
  3891=>"110000000",
  3892=>"000000000",
  3893=>"111111111",
  3894=>"111101101",
  3895=>"111111111",
  3896=>"000000000",
  3897=>"111111111",
  3898=>"000000100",
  3899=>"001001001",
  3900=>"110000000",
  3901=>"000010011",
  3902=>"000000000",
  3903=>"111011011",
  3904=>"101100000",
  3905=>"111000000",
  3906=>"101000000",
  3907=>"000000101",
  3908=>"000001001",
  3909=>"000001000",
  3910=>"000001000",
  3911=>"000000101",
  3912=>"110110000",
  3913=>"111101100",
  3914=>"110110010",
  3915=>"100100100",
  3916=>"111111000",
  3917=>"111011111",
  3918=>"111111011",
  3919=>"100100110",
  3920=>"000011010",
  3921=>"000000101",
  3922=>"110111010",
  3923=>"000000000",
  3924=>"111111110",
  3925=>"001011011",
  3926=>"111111010",
  3927=>"000001000",
  3928=>"001001001",
  3929=>"111111100",
  3930=>"000001011",
  3931=>"110110100",
  3932=>"001001001",
  3933=>"000000000",
  3934=>"110110000",
  3935=>"001001000",
  3936=>"101100101",
  3937=>"100000000",
  3938=>"110000000",
  3939=>"110110110",
  3940=>"011011011",
  3941=>"110110010",
  3942=>"001011111",
  3943=>"011011111",
  3944=>"110001011",
  3945=>"001001000",
  3946=>"111111111",
  3947=>"001111111",
  3948=>"110110100",
  3949=>"010010011",
  3950=>"000011111",
  3951=>"111000000",
  3952=>"110000000",
  3953=>"111111000",
  3954=>"110111110",
  3955=>"000011011",
  3956=>"000010000",
  3957=>"100110111",
  3958=>"111011011",
  3959=>"000000000",
  3960=>"000000001",
  3961=>"111010100",
  3962=>"111111010",
  3963=>"000000000",
  3964=>"001110110",
  3965=>"000000111",
  3966=>"100000000",
  3967=>"000000100",
  3968=>"001111110",
  3969=>"111111111",
  3970=>"100000001",
  3971=>"101001001",
  3972=>"111100100",
  3973=>"000001001",
  3974=>"101101111",
  3975=>"111100110",
  3976=>"101001001",
  3977=>"111001000",
  3978=>"101000100",
  3979=>"000111111",
  3980=>"100100101",
  3981=>"011000000",
  3982=>"000000111",
  3983=>"111110010",
  3984=>"111111011",
  3985=>"000011111",
  3986=>"000110111",
  3987=>"001000000",
  3988=>"100111101",
  3989=>"000000000",
  3990=>"111111111",
  3991=>"011000000",
  3992=>"000000111",
  3993=>"101100000",
  3994=>"111101011",
  3995=>"010010000",
  3996=>"000101101",
  3997=>"011011011",
  3998=>"000000000",
  3999=>"111111000",
  4000=>"000000000",
  4001=>"011011001",
  4002=>"100000101",
  4003=>"101001000",
  4004=>"100000101",
  4005=>"010111110",
  4006=>"111111000",
  4007=>"111111111",
  4008=>"000000000",
  4009=>"101000110",
  4010=>"011000000",
  4011=>"100000000",
  4012=>"101101101",
  4013=>"101001000",
  4014=>"111000000",
  4015=>"111100101",
  4016=>"001111111",
  4017=>"000000000",
  4018=>"010110010",
  4019=>"111001111",
  4020=>"101001001",
  4021=>"111111010",
  4022=>"111111100",
  4023=>"000000000",
  4024=>"111101111",
  4025=>"000100111",
  4026=>"111010000",
  4027=>"100000000",
  4028=>"000100000",
  4029=>"011001001",
  4030=>"111010110",
  4031=>"111110001",
  4032=>"001001111",
  4033=>"011111000",
  4034=>"111101100",
  4035=>"001010000",
  4036=>"111011111",
  4037=>"100000100",
  4038=>"111111111",
  4039=>"101101111",
  4040=>"000000101",
  4041=>"111011011",
  4042=>"000000000",
  4043=>"000000111",
  4044=>"010010000",
  4045=>"000001111",
  4046=>"001000001",
  4047=>"101101101",
  4048=>"111110010",
  4049=>"000000000",
  4050=>"101101100",
  4051=>"000011111",
  4052=>"100100000",
  4053=>"111110001",
  4054=>"110011110",
  4055=>"000000110",
  4056=>"111111011",
  4057=>"110110110",
  4058=>"000000000",
  4059=>"111000001",
  4060=>"000000000",
  4061=>"111111111",
  4062=>"000000000",
  4063=>"011011011",
  4064=>"000000000",
  4065=>"111101000",
  4066=>"011000000",
  4067=>"111111101",
  4068=>"110110110",
  4069=>"101101101",
  4070=>"011011111",
  4071=>"111101111",
  4072=>"110110011",
  4073=>"111111111",
  4074=>"110000000",
  4075=>"000111111",
  4076=>"011000000",
  4077=>"000110111",
  4078=>"111111011",
  4079=>"000000000",
  4080=>"010011010",
  4081=>"000000001",
  4082=>"000000000",
  4083=>"001001000",
  4084=>"111101111",
  4085=>"111111111",
  4086=>"111111111",
  4087=>"100110110",
  4088=>"000000000",
  4089=>"100000011",
  4090=>"001000000",
  4091=>"001101001",
  4092=>"100101001",
  4093=>"101001000",
  4094=>"100000110",
  4095=>"000000100",
  4096=>"000000000",
  4097=>"101000001",
  4098=>"101101100",
  4099=>"111111101",
  4100=>"110111011",
  4101=>"111111000",
  4102=>"100000000",
  4103=>"000101101",
  4104=>"111111110",
  4105=>"000000000",
  4106=>"000000001",
  4107=>"011001111",
  4108=>"000000001",
  4109=>"000111111",
  4110=>"010010011",
  4111=>"000000000",
  4112=>"110111101",
  4113=>"000110011",
  4114=>"000100111",
  4115=>"000000000",
  4116=>"000000001",
  4117=>"000001001",
  4118=>"000000000",
  4119=>"001001101",
  4120=>"000010000",
  4121=>"001001001",
  4122=>"001000000",
  4123=>"011111111",
  4124=>"010011000",
  4125=>"101001000",
  4126=>"110100100",
  4127=>"000000000",
  4128=>"000000001",
  4129=>"111111111",
  4130=>"101111111",
  4131=>"111111111",
  4132=>"111110110",
  4133=>"000000000",
  4134=>"111111110",
  4135=>"000000011",
  4136=>"111110100",
  4137=>"000000000",
  4138=>"011111111",
  4139=>"100000001",
  4140=>"011001111",
  4141=>"111111111",
  4142=>"111110111",
  4143=>"000000000",
  4144=>"110000001",
  4145=>"011111010",
  4146=>"000000000",
  4147=>"111011010",
  4148=>"101101111",
  4149=>"000000000",
  4150=>"000000000",
  4151=>"000000100",
  4152=>"000000010",
  4153=>"001001001",
  4154=>"101001001",
  4155=>"000000000",
  4156=>"000100100",
  4157=>"100100000",
  4158=>"001000100",
  4159=>"111001111",
  4160=>"111110111",
  4161=>"001001000",
  4162=>"000000000",
  4163=>"111110000",
  4164=>"000011011",
  4165=>"001000000",
  4166=>"111111101",
  4167=>"111101000",
  4168=>"111101111",
  4169=>"001001000",
  4170=>"111111111",
  4171=>"000000000",
  4172=>"000000111",
  4173=>"000000000",
  4174=>"100000000",
  4175=>"111111111",
  4176=>"000000000",
  4177=>"000000000",
  4178=>"000100111",
  4179=>"000111100",
  4180=>"000000000",
  4181=>"110111111",
  4182=>"000011001",
  4183=>"000000001",
  4184=>"000000000",
  4185=>"000000000",
  4186=>"101111101",
  4187=>"011110110",
  4188=>"000000000",
  4189=>"000000000",
  4190=>"000000000",
  4191=>"111110100",
  4192=>"111111011",
  4193=>"001001001",
  4194=>"001000000",
  4195=>"111110111",
  4196=>"000000000",
  4197=>"011111111",
  4198=>"010110110",
  4199=>"000000000",
  4200=>"111111111",
  4201=>"111101001",
  4202=>"000000111",
  4203=>"011000000",
  4204=>"000011110",
  4205=>"000000111",
  4206=>"111111111",
  4207=>"001001000",
  4208=>"000111110",
  4209=>"111111110",
  4210=>"101100100",
  4211=>"000000110",
  4212=>"001000000",
  4213=>"100100111",
  4214=>"110101101",
  4215=>"000000100",
  4216=>"011111111",
  4217=>"101101111",
  4218=>"000000110",
  4219=>"000000000",
  4220=>"110110110",
  4221=>"111111011",
  4222=>"000000100",
  4223=>"100000000",
  4224=>"111011111",
  4225=>"100111100",
  4226=>"001000000",
  4227=>"111111111",
  4228=>"111111110",
  4229=>"101001101",
  4230=>"000000000",
  4231=>"000001000",
  4232=>"000001000",
  4233=>"000000101",
  4234=>"000000000",
  4235=>"111011011",
  4236=>"001000000",
  4237=>"000000000",
  4238=>"111110111",
  4239=>"101001001",
  4240=>"000010111",
  4241=>"111010000",
  4242=>"010110111",
  4243=>"111100100",
  4244=>"111111110",
  4245=>"111000101",
  4246=>"000000001",
  4247=>"100000000",
  4248=>"000000000",
  4249=>"000000001",
  4250=>"000000001",
  4251=>"000010110",
  4252=>"001111111",
  4253=>"000000111",
  4254=>"001101111",
  4255=>"101001101",
  4256=>"011011000",
  4257=>"100001001",
  4258=>"100111011",
  4259=>"000011001",
  4260=>"000000011",
  4261=>"110111111",
  4262=>"010110010",
  4263=>"110111111",
  4264=>"111111101",
  4265=>"110111110",
  4266=>"111000000",
  4267=>"100000111",
  4268=>"000111111",
  4269=>"100110011",
  4270=>"001111111",
  4271=>"011111010",
  4272=>"010110000",
  4273=>"100111100",
  4274=>"111111111",
  4275=>"111111111",
  4276=>"000000010",
  4277=>"111111111",
  4278=>"001001011",
  4279=>"000011111",
  4280=>"000110101",
  4281=>"001001101",
  4282=>"000000000",
  4283=>"000000000",
  4284=>"000000000",
  4285=>"110110110",
  4286=>"101111101",
  4287=>"010101000",
  4288=>"000010111",
  4289=>"000000000",
  4290=>"100110000",
  4291=>"111000000",
  4292=>"011111111",
  4293=>"011111000",
  4294=>"000010111",
  4295=>"011010000",
  4296=>"000000100",
  4297=>"100000000",
  4298=>"111001000",
  4299=>"111111111",
  4300=>"111101011",
  4301=>"111111111",
  4302=>"111111111",
  4303=>"100001011",
  4304=>"000100111",
  4305=>"010010000",
  4306=>"011000000",
  4307=>"000000000",
  4308=>"111001111",
  4309=>"001011111",
  4310=>"000000000",
  4311=>"100000110",
  4312=>"100001111",
  4313=>"111101101",
  4314=>"000101000",
  4315=>"000100111",
  4316=>"111111111",
  4317=>"111011111",
  4318=>"111110111",
  4319=>"000111111",
  4320=>"111111111",
  4321=>"011111010",
  4322=>"001000000",
  4323=>"111111001",
  4324=>"110111111",
  4325=>"010011011",
  4326=>"001000000",
  4327=>"000000000",
  4328=>"111101111",
  4329=>"001001001",
  4330=>"110111111",
  4331=>"000101111",
  4332=>"000000111",
  4333=>"000000000",
  4334=>"100111111",
  4335=>"111001000",
  4336=>"001000111",
  4337=>"111111001",
  4338=>"111111001",
  4339=>"000000000",
  4340=>"100111111",
  4341=>"111000110",
  4342=>"011011110",
  4343=>"111000000",
  4344=>"001011001",
  4345=>"000000000",
  4346=>"100111111",
  4347=>"100110111",
  4348=>"111011011",
  4349=>"101001111",
  4350=>"000000000",
  4351=>"111111101",
  4352=>"000000000",
  4353=>"111110000",
  4354=>"000000000",
  4355=>"000000000",
  4356=>"000011010",
  4357=>"000000000",
  4358=>"111111111",
  4359=>"101101101",
  4360=>"111111111",
  4361=>"101101101",
  4362=>"000000000",
  4363=>"111111111",
  4364=>"000000010",
  4365=>"010110011",
  4366=>"000000011",
  4367=>"000000110",
  4368=>"111111101",
  4369=>"000111111",
  4370=>"001000000",
  4371=>"111100000",
  4372=>"000100000",
  4373=>"111101111",
  4374=>"111111111",
  4375=>"111111000",
  4376=>"110111111",
  4377=>"000000000",
  4378=>"111111111",
  4379=>"001001001",
  4380=>"011011111",
  4381=>"001000000",
  4382=>"111011000",
  4383=>"011111010",
  4384=>"111110111",
  4385=>"110111000",
  4386=>"010010111",
  4387=>"001000001",
  4388=>"111101111",
  4389=>"100000001",
  4390=>"000010000",
  4391=>"000000001",
  4392=>"000111111",
  4393=>"000000000",
  4394=>"111100000",
  4395=>"000000000",
  4396=>"000010111",
  4397=>"000111111",
  4398=>"000000001",
  4399=>"111111110",
  4400=>"111111111",
  4401=>"111110111",
  4402=>"000000111",
  4403=>"000000111",
  4404=>"000001011",
  4405=>"100000000",
  4406=>"111101000",
  4407=>"011000000",
  4408=>"010011110",
  4409=>"111101111",
  4410=>"000000111",
  4411=>"010000000",
  4412=>"101111100",
  4413=>"000010110",
  4414=>"000000000",
  4415=>"100100011",
  4416=>"000000000",
  4417=>"110111111",
  4418=>"000000000",
  4419=>"000110110",
  4420=>"111101001",
  4421=>"001001111",
  4422=>"011011010",
  4423=>"101000001",
  4424=>"111111111",
  4425=>"111001000",
  4426=>"001000000",
  4427=>"111110011",
  4428=>"000011111",
  4429=>"000000110",
  4430=>"000000111",
  4431=>"010010010",
  4432=>"110010000",
  4433=>"111111100",
  4434=>"010000000",
  4435=>"111111111",
  4436=>"000000001",
  4437=>"011011011",
  4438=>"001111111",
  4439=>"101111111",
  4440=>"000000000",
  4441=>"111111011",
  4442=>"110110110",
  4443=>"000111000",
  4444=>"000001000",
  4445=>"001000011",
  4446=>"000001000",
  4447=>"100100110",
  4448=>"110111000",
  4449=>"110010111",
  4450=>"011111111",
  4451=>"111111000",
  4452=>"111101111",
  4453=>"111010110",
  4454=>"111111000",
  4455=>"110111110",
  4456=>"110111101",
  4457=>"111111000",
  4458=>"111001001",
  4459=>"010000001",
  4460=>"110110100",
  4461=>"000111011",
  4462=>"000000000",
  4463=>"000110100",
  4464=>"111101100",
  4465=>"000110110",
  4466=>"011111111",
  4467=>"111011011",
  4468=>"000001000",
  4469=>"000111111",
  4470=>"000010010",
  4471=>"110100000",
  4472=>"000100111",
  4473=>"110111111",
  4474=>"011000111",
  4475=>"110111111",
  4476=>"001000000",
  4477=>"010111111",
  4478=>"000000000",
  4479=>"111000111",
  4480=>"110110110",
  4481=>"000011001",
  4482=>"100000100",
  4483=>"000000111",
  4484=>"100001001",
  4485=>"111111110",
  4486=>"000001111",
  4487=>"100100000",
  4488=>"001000001",
  4489=>"100110000",
  4490=>"111111111",
  4491=>"000000000",
  4492=>"111111101",
  4493=>"111001001",
  4494=>"000000110",
  4495=>"000000000",
  4496=>"011111010",
  4497=>"100000011",
  4498=>"101000000",
  4499=>"111111011",
  4500=>"110111111",
  4501=>"000000000",
  4502=>"111011001",
  4503=>"110110111",
  4504=>"111111111",
  4505=>"011010011",
  4506=>"111111111",
  4507=>"111111111",
  4508=>"110111111",
  4509=>"100111111",
  4510=>"110111111",
  4511=>"010111000",
  4512=>"110111111",
  4513=>"000100111",
  4514=>"000111101",
  4515=>"111101111",
  4516=>"000110110",
  4517=>"000110111",
  4518=>"110110111",
  4519=>"010010111",
  4520=>"100000000",
  4521=>"101100000",
  4522=>"000000001",
  4523=>"000000000",
  4524=>"000000000",
  4525=>"001000000",
  4526=>"111111111",
  4527=>"001000000",
  4528=>"111101101",
  4529=>"000000111",
  4530=>"000000000",
  4531=>"111110111",
  4532=>"111111111",
  4533=>"111001101",
  4534=>"110111111",
  4535=>"000000000",
  4536=>"110010000",
  4537=>"010000000",
  4538=>"101000000",
  4539=>"010011111",
  4540=>"001001000",
  4541=>"111101001",
  4542=>"000000000",
  4543=>"100110111",
  4544=>"111001001",
  4545=>"111111111",
  4546=>"000000000",
  4547=>"001001000",
  4548=>"111111001",
  4549=>"000001000",
  4550=>"110110000",
  4551=>"111101000",
  4552=>"000000000",
  4553=>"000000000",
  4554=>"001000100",
  4555=>"111111111",
  4556=>"111111010",
  4557=>"000000111",
  4558=>"110111000",
  4559=>"000110111",
  4560=>"000000000",
  4561=>"000000110",
  4562=>"100110111",
  4563=>"101011111",
  4564=>"101101001",
  4565=>"111001111",
  4566=>"111111111",
  4567=>"100100100",
  4568=>"111111111",
  4569=>"000111111",
  4570=>"000000000",
  4571=>"010011111",
  4572=>"111011011",
  4573=>"001111110",
  4574=>"100100111",
  4575=>"100000000",
  4576=>"001111111",
  4577=>"110010111",
  4578=>"110010000",
  4579=>"111111111",
  4580=>"000111011",
  4581=>"111111101",
  4582=>"001000101",
  4583=>"111111111",
  4584=>"000000000",
  4585=>"111001000",
  4586=>"111111000",
  4587=>"000000000",
  4588=>"111111111",
  4589=>"011111111",
  4590=>"000000101",
  4591=>"000000001",
  4592=>"000000111",
  4593=>"000000000",
  4594=>"000110100",
  4595=>"111111010",
  4596=>"110110010",
  4597=>"111111111",
  4598=>"010111110",
  4599=>"000000001",
  4600=>"111101101",
  4601=>"011011110",
  4602=>"111111000",
  4603=>"001001001",
  4604=>"000001001",
  4605=>"111111111",
  4606=>"000000000",
  4607=>"111110010",
  4608=>"000101111",
  4609=>"001111111",
  4610=>"000000000",
  4611=>"000000010",
  4612=>"100100000",
  4613=>"010000001",
  4614=>"111000000",
  4615=>"111111110",
  4616=>"110000000",
  4617=>"111111111",
  4618=>"001011111",
  4619=>"000000000",
  4620=>"011010111",
  4621=>"111101111",
  4622=>"000000110",
  4623=>"000011001",
  4624=>"111111001",
  4625=>"001000000",
  4626=>"001111111",
  4627=>"000000000",
  4628=>"000000011",
  4629=>"000000000",
  4630=>"011111100",
  4631=>"001101001",
  4632=>"110110100",
  4633=>"000000000",
  4634=>"111100111",
  4635=>"111111000",
  4636=>"111110000",
  4637=>"101111111",
  4638=>"000001011",
  4639=>"000000000",
  4640=>"001011000",
  4641=>"000001000",
  4642=>"111111110",
  4643=>"111111000",
  4644=>"111111111",
  4645=>"111001101",
  4646=>"000000111",
  4647=>"111111111",
  4648=>"111111111",
  4649=>"000000000",
  4650=>"000000000",
  4651=>"111111111",
  4652=>"111111001",
  4653=>"001000000",
  4654=>"011111111",
  4655=>"000000001",
  4656=>"001011000",
  4657=>"001011101",
  4658=>"000010000",
  4659=>"100100111",
  4660=>"000111111",
  4661=>"000000110",
  4662=>"011111111",
  4663=>"111111111",
  4664=>"111111000",
  4665=>"110000000",
  4666=>"111000000",
  4667=>"111111111",
  4668=>"111001001",
  4669=>"111111011",
  4670=>"001010011",
  4671=>"100000000",
  4672=>"000000000",
  4673=>"111000000",
  4674=>"111111111",
  4675=>"111110000",
  4676=>"111000000",
  4677=>"000000000",
  4678=>"111001100",
  4679=>"110100000",
  4680=>"011000000",
  4681=>"001000011",
  4682=>"110110111",
  4683=>"100000000",
  4684=>"111111111",
  4685=>"111111111",
  4686=>"011000000",
  4687=>"001001110",
  4688=>"000111000",
  4689=>"001011111",
  4690=>"000010010",
  4691=>"000110111",
  4692=>"001111111",
  4693=>"100100110",
  4694=>"110100000",
  4695=>"011111010",
  4696=>"111111111",
  4697=>"000000111",
  4698=>"111111000",
  4699=>"000000000",
  4700=>"110111111",
  4701=>"111111011",
  4702=>"000000011",
  4703=>"011001000",
  4704=>"111111111",
  4705=>"111111111",
  4706=>"111111111",
  4707=>"000000001",
  4708=>"111111111",
  4709=>"000000000",
  4710=>"101111000",
  4711=>"000110111",
  4712=>"110110110",
  4713=>"111111111",
  4714=>"000000000",
  4715=>"010100000",
  4716=>"000000011",
  4717=>"111111111",
  4718=>"000000000",
  4719=>"000111110",
  4720=>"000000000",
  4721=>"001000000",
  4722=>"001001111",
  4723=>"000000000",
  4724=>"000000000",
  4725=>"001101111",
  4726=>"000000000",
  4727=>"000000101",
  4728=>"000000000",
  4729=>"111000100",
  4730=>"101100100",
  4731=>"011111111",
  4732=>"110110110",
  4733=>"000000000",
  4734=>"111100101",
  4735=>"000000000",
  4736=>"000000001",
  4737=>"111111011",
  4738=>"000000001",
  4739=>"011111111",
  4740=>"000000000",
  4741=>"000000110",
  4742=>"011000000",
  4743=>"111111111",
  4744=>"000000000",
  4745=>"111111000",
  4746=>"111111111",
  4747=>"100100000",
  4748=>"001011111",
  4749=>"000000111",
  4750=>"010000010",
  4751=>"100000000",
  4752=>"111111111",
  4753=>"000000000",
  4754=>"111111101",
  4755=>"000000100",
  4756=>"000011011",
  4757=>"011000111",
  4758=>"000000000",
  4759=>"111101101",
  4760=>"111011011",
  4761=>"111111111",
  4762=>"100101101",
  4763=>"000000000",
  4764=>"110100000",
  4765=>"100011001",
  4766=>"000000000",
  4767=>"011000000",
  4768=>"000000000",
  4769=>"111011001",
  4770=>"111110111",
  4771=>"000000000",
  4772=>"111011111",
  4773=>"110000111",
  4774=>"000101000",
  4775=>"001011011",
  4776=>"111111111",
  4777=>"000000101",
  4778=>"000000111",
  4779=>"111111011",
  4780=>"010100000",
  4781=>"110010000",
  4782=>"001000100",
  4783=>"101000000",
  4784=>"111111111",
  4785=>"001001000",
  4786=>"111111110",
  4787=>"111111111",
  4788=>"000000000",
  4789=>"111111101",
  4790=>"000000000",
  4791=>"110000110",
  4792=>"000001111",
  4793=>"111111101",
  4794=>"001000000",
  4795=>"000000111",
  4796=>"000110011",
  4797=>"000001011",
  4798=>"110100100",
  4799=>"000000101",
  4800=>"111111111",
  4801=>"110100000",
  4802=>"001000001",
  4803=>"000001111",
  4804=>"000110111",
  4805=>"000100111",
  4806=>"110000000",
  4807=>"101000000",
  4808=>"000111111",
  4809=>"001000000",
  4810=>"111111111",
  4811=>"111010111",
  4812=>"111110111",
  4813=>"111111111",
  4814=>"111111111",
  4815=>"111111111",
  4816=>"110110100",
  4817=>"011111110",
  4818=>"111111111",
  4819=>"111111111",
  4820=>"100101111",
  4821=>"110110111",
  4822=>"000010111",
  4823=>"111000101",
  4824=>"111110111",
  4825=>"111100000",
  4826=>"011000000",
  4827=>"111111111",
  4828=>"111111101",
  4829=>"111111111",
  4830=>"111011011",
  4831=>"000000000",
  4832=>"000000110",
  4833=>"000000010",
  4834=>"000110110",
  4835=>"110000001",
  4836=>"100000000",
  4837=>"011001000",
  4838=>"111111111",
  4839=>"000000000",
  4840=>"000000000",
  4841=>"100110011",
  4842=>"011001110",
  4843=>"111111100",
  4844=>"111111000",
  4845=>"000000111",
  4846=>"000000000",
  4847=>"011001110",
  4848=>"111111110",
  4849=>"000000000",
  4850=>"011000000",
  4851=>"001000000",
  4852=>"111111001",
  4853=>"000000000",
  4854=>"011000111",
  4855=>"000010110",
  4856=>"110111111",
  4857=>"111111000",
  4858=>"000000000",
  4859=>"100110011",
  4860=>"000110110",
  4861=>"100111111",
  4862=>"010110011",
  4863=>"000000000",
  4864=>"111001001",
  4865=>"000000000",
  4866=>"111110000",
  4867=>"110000000",
  4868=>"000000000",
  4869=>"010000000",
  4870=>"101000000",
  4871=>"101000000",
  4872=>"100100000",
  4873=>"000000100",
  4874=>"000111111",
  4875=>"000000011",
  4876=>"111111111",
  4877=>"011001111",
  4878=>"100100100",
  4879=>"011011000",
  4880=>"000000001",
  4881=>"001001000",
  4882=>"110000000",
  4883=>"111111100",
  4884=>"111100000",
  4885=>"111011000",
  4886=>"110110000",
  4887=>"111011001",
  4888=>"000110110",
  4889=>"100000000",
  4890=>"110110110",
  4891=>"110111111",
  4892=>"000000000",
  4893=>"111111001",
  4894=>"000000000",
  4895=>"111000000",
  4896=>"111111110",
  4897=>"111111111",
  4898=>"000000000",
  4899=>"111111111",
  4900=>"000001000",
  4901=>"011111110",
  4902=>"001001100",
  4903=>"000001111",
  4904=>"000000110",
  4905=>"011011011",
  4906=>"011010000",
  4907=>"111110110",
  4908=>"011000100",
  4909=>"101111110",
  4910=>"111111110",
  4911=>"000000111",
  4912=>"000000100",
  4913=>"001101111",
  4914=>"111111111",
  4915=>"000110111",
  4916=>"111111111",
  4917=>"011110110",
  4918=>"000111111",
  4919=>"111111111",
  4920=>"000000000",
  4921=>"000110111",
  4922=>"000011001",
  4923=>"000010011",
  4924=>"001000000",
  4925=>"111110110",
  4926=>"111111111",
  4927=>"000111110",
  4928=>"000000110",
  4929=>"000000101",
  4930=>"101111111",
  4931=>"110111111",
  4932=>"111011000",
  4933=>"000011111",
  4934=>"110111111",
  4935=>"000000000",
  4936=>"000000011",
  4937=>"000000000",
  4938=>"100111100",
  4939=>"000110110",
  4940=>"000100111",
  4941=>"011110111",
  4942=>"111111111",
  4943=>"100100110",
  4944=>"000010000",
  4945=>"011001000",
  4946=>"101111111",
  4947=>"111111111",
  4948=>"000000000",
  4949=>"011011111",
  4950=>"010111111",
  4951=>"111111111",
  4952=>"111111111",
  4953=>"000000100",
  4954=>"001111110",
  4955=>"001011001",
  4956=>"000000000",
  4957=>"001001001",
  4958=>"111111101",
  4959=>"111111111",
  4960=>"111101111",
  4961=>"111111111",
  4962=>"001000100",
  4963=>"011111111",
  4964=>"110111110",
  4965=>"111000100",
  4966=>"000000000",
  4967=>"111110011",
  4968=>"000000011",
  4969=>"010110000",
  4970=>"111111111",
  4971=>"001001111",
  4972=>"000100100",
  4973=>"001000000",
  4974=>"000000000",
  4975=>"000111111",
  4976=>"101001011",
  4977=>"001001000",
  4978=>"000101111",
  4979=>"111111111",
  4980=>"111110100",
  4981=>"111011111",
  4982=>"000000000",
  4983=>"010010100",
  4984=>"111000000",
  4985=>"101000000",
  4986=>"000000000",
  4987=>"000000000",
  4988=>"000000100",
  4989=>"000000000",
  4990=>"010111111",
  4991=>"000000000",
  4992=>"000000000",
  4993=>"100110110",
  4994=>"000000111",
  4995=>"000000000",
  4996=>"000000110",
  4997=>"111111000",
  4998=>"000000101",
  4999=>"000000000",
  5000=>"000010000",
  5001=>"001000100",
  5002=>"000000001",
  5003=>"010000000",
  5004=>"111101111",
  5005=>"100100111",
  5006=>"001101111",
  5007=>"000000001",
  5008=>"011011000",
  5009=>"111111101",
  5010=>"111111000",
  5011=>"000010010",
  5012=>"011111111",
  5013=>"000000000",
  5014=>"001111111",
  5015=>"000000000",
  5016=>"000000100",
  5017=>"000000100",
  5018=>"000000000",
  5019=>"100100110",
  5020=>"000000000",
  5021=>"100000000",
  5022=>"001001111",
  5023=>"000000000",
  5024=>"111111000",
  5025=>"011000000",
  5026=>"111111111",
  5027=>"111111111",
  5028=>"000000110",
  5029=>"000101111",
  5030=>"111000000",
  5031=>"111111111",
  5032=>"111111111",
  5033=>"000000110",
  5034=>"110111001",
  5035=>"101001000",
  5036=>"000000000",
  5037=>"000001111",
  5038=>"000100001",
  5039=>"110000110",
  5040=>"111111111",
  5041=>"111111000",
  5042=>"110111111",
  5043=>"101111111",
  5044=>"111111111",
  5045=>"111111011",
  5046=>"000000000",
  5047=>"000000110",
  5048=>"110000000",
  5049=>"000000000",
  5050=>"111111111",
  5051=>"110000000",
  5052=>"000000111",
  5053=>"000000111",
  5054=>"011111111",
  5055=>"110110110",
  5056=>"010000000",
  5057=>"000011111",
  5058=>"111111111",
  5059=>"111111000",
  5060=>"001001001",
  5061=>"100100100",
  5062=>"000100110",
  5063=>"000000010",
  5064=>"000000001",
  5065=>"000000000",
  5066=>"000000000",
  5067=>"111111100",
  5068=>"001000000",
  5069=>"001111111",
  5070=>"000111111",
  5071=>"000000000",
  5072=>"000000100",
  5073=>"000010110",
  5074=>"000101111",
  5075=>"000000101",
  5076=>"101000000",
  5077=>"100000000",
  5078=>"000000000",
  5079=>"111111111",
  5080=>"110111000",
  5081=>"000011011",
  5082=>"001000000",
  5083=>"000000000",
  5084=>"000000000",
  5085=>"100110101",
  5086=>"011010010",
  5087=>"001001001",
  5088=>"111001000",
  5089=>"000000111",
  5090=>"000000111",
  5091=>"001000111",
  5092=>"111001101",
  5093=>"001111111",
  5094=>"111000100",
  5095=>"111111000",
  5096=>"111000000",
  5097=>"000000000",
  5098=>"000000000",
  5099=>"000000100",
  5100=>"101101000",
  5101=>"001000000",
  5102=>"000001000",
  5103=>"000011111",
  5104=>"111101111",
  5105=>"111111111",
  5106=>"111111111",
  5107=>"000000000",
  5108=>"001000010",
  5109=>"010100111",
  5110=>"000000111",
  5111=>"100011111",
  5112=>"000000000",
  5113=>"000011011",
  5114=>"000100100",
  5115=>"111111101",
  5116=>"000000000",
  5117=>"000111011",
  5118=>"111111111",
  5119=>"111111111",
  5120=>"110100100",
  5121=>"000000000",
  5122=>"001000000",
  5123=>"000011001",
  5124=>"101111111",
  5125=>"111010110",
  5126=>"100000001",
  5127=>"000000000",
  5128=>"001001000",
  5129=>"110111011",
  5130=>"100110110",
  5131=>"000011111",
  5132=>"000000111",
  5133=>"000000110",
  5134=>"111001011",
  5135=>"111111011",
  5136=>"111111111",
  5137=>"011000001",
  5138=>"111111111",
  5139=>"111001001",
  5140=>"000000000",
  5141=>"011110111",
  5142=>"000000001",
  5143=>"110010100",
  5144=>"001001101",
  5145=>"000001000",
  5146=>"000010110",
  5147=>"100000010",
  5148=>"111110110",
  5149=>"000010010",
  5150=>"000000001",
  5151=>"000101111",
  5152=>"110000000",
  5153=>"100111111",
  5154=>"100000001",
  5155=>"000000011",
  5156=>"000000001",
  5157=>"110100111",
  5158=>"110110100",
  5159=>"111101111",
  5160=>"111100000",
  5161=>"000000110",
  5162=>"100000000",
  5163=>"111111110",
  5164=>"111000000",
  5165=>"100101000",
  5166=>"111111111",
  5167=>"111111111",
  5168=>"111110111",
  5169=>"000001001",
  5170=>"000000011",
  5171=>"111111010",
  5172=>"111111111",
  5173=>"000001110",
  5174=>"100100000",
  5175=>"001000001",
  5176=>"000000010",
  5177=>"100000011",
  5178=>"101111111",
  5179=>"001001001",
  5180=>"000111111",
  5181=>"110111101",
  5182=>"000000001",
  5183=>"111111111",
  5184=>"110111111",
  5185=>"011111100",
  5186=>"111111111",
  5187=>"110110111",
  5188=>"001011111",
  5189=>"001000001",
  5190=>"110101111",
  5191=>"111111111",
  5192=>"011011001",
  5193=>"111111111",
  5194=>"000000000",
  5195=>"100111111",
  5196=>"000000000",
  5197=>"111100001",
  5198=>"001000100",
  5199=>"000000000",
  5200=>"111111101",
  5201=>"000111110",
  5202=>"000000000",
  5203=>"001111000",
  5204=>"001000000",
  5205=>"111111000",
  5206=>"000000000",
  5207=>"000110110",
  5208=>"000011000",
  5209=>"010010000",
  5210=>"000000011",
  5211=>"111111111",
  5212=>"000000000",
  5213=>"111111111",
  5214=>"111111001",
  5215=>"110111111",
  5216=>"000000000",
  5217=>"001111111",
  5218=>"000000000",
  5219=>"000000010",
  5220=>"011111100",
  5221=>"000000011",
  5222=>"101101001",
  5223=>"001011010",
  5224=>"111111111",
  5225=>"111111111",
  5226=>"010000000",
  5227=>"001011001",
  5228=>"000000110",
  5229=>"111111000",
  5230=>"101000000",
  5231=>"111111111",
  5232=>"000000111",
  5233=>"000111111",
  5234=>"111111111",
  5235=>"000111111",
  5236=>"100000001",
  5237=>"001001101",
  5238=>"011010010",
  5239=>"000000001",
  5240=>"111010110",
  5241=>"000110110",
  5242=>"000000001",
  5243=>"111111111",
  5244=>"111111110",
  5245=>"111111111",
  5246=>"000000000",
  5247=>"111000110",
  5248=>"111111111",
  5249=>"111111111",
  5250=>"111000100",
  5251=>"111111111",
  5252=>"111111111",
  5253=>"000000000",
  5254=>"110110111",
  5255=>"111010101",
  5256=>"111111001",
  5257=>"111110111",
  5258=>"111111111",
  5259=>"111111111",
  5260=>"000000000",
  5261=>"100001001",
  5262=>"111111001",
  5263=>"001001001",
  5264=>"010000000",
  5265=>"111111111",
  5266=>"001111110",
  5267=>"111111111",
  5268=>"000110110",
  5269=>"001001111",
  5270=>"111111000",
  5271=>"000000100",
  5272=>"000000000",
  5273=>"100000000",
  5274=>"000000000",
  5275=>"111100100",
  5276=>"111111111",
  5277=>"001100111",
  5278=>"110100000",
  5279=>"110110110",
  5280=>"110100100",
  5281=>"111000000",
  5282=>"111111111",
  5283=>"111111111",
  5284=>"000000000",
  5285=>"100001000",
  5286=>"100000101",
  5287=>"100000010",
  5288=>"111111111",
  5289=>"000011110",
  5290=>"111111101",
  5291=>"001011111",
  5292=>"100110011",
  5293=>"001110111",
  5294=>"111111111",
  5295=>"000000110",
  5296=>"111111100",
  5297=>"101001111",
  5298=>"100000100",
  5299=>"011101111",
  5300=>"100100100",
  5301=>"011111111",
  5302=>"000000000",
  5303=>"110111000",
  5304=>"111110110",
  5305=>"001000000",
  5306=>"000000000",
  5307=>"101001001",
  5308=>"111111111",
  5309=>"111011011",
  5310=>"111111110",
  5311=>"001001111",
  5312=>"111111111",
  5313=>"000000110",
  5314=>"101111111",
  5315=>"000000000",
  5316=>"111111010",
  5317=>"000000000",
  5318=>"010001011",
  5319=>"000000110",
  5320=>"010000000",
  5321=>"100111111",
  5322=>"000000100",
  5323=>"000000100",
  5324=>"110010111",
  5325=>"000000000",
  5326=>"000000000",
  5327=>"000000111",
  5328=>"111001111",
  5329=>"111011100",
  5330=>"000000100",
  5331=>"000000000",
  5332=>"000110000",
  5333=>"000011001",
  5334=>"111111110",
  5335=>"111111111",
  5336=>"000000000",
  5337=>"111111100",
  5338=>"111111100",
  5339=>"100000000",
  5340=>"110111000",
  5341=>"111111110",
  5342=>"111111111",
  5343=>"111111111",
  5344=>"000000000",
  5345=>"011011011",
  5346=>"000000100",
  5347=>"111111001",
  5348=>"111101111",
  5349=>"111111110",
  5350=>"111111111",
  5351=>"000000000",
  5352=>"111000100",
  5353=>"000011111",
  5354=>"000000111",
  5355=>"000000011",
  5356=>"000110111",
  5357=>"001011001",
  5358=>"000000000",
  5359=>"000010000",
  5360=>"111100000",
  5361=>"111111111",
  5362=>"111111111",
  5363=>"010110111",
  5364=>"111111011",
  5365=>"111111111",
  5366=>"100000010",
  5367=>"010000000",
  5368=>"000001011",
  5369=>"111111111",
  5370=>"000000000",
  5371=>"000111011",
  5372=>"111111111",
  5373=>"110111111",
  5374=>"000000111",
  5375=>"110110000",
  5376=>"100000000",
  5377=>"000000001",
  5378=>"000000111",
  5379=>"111111111",
  5380=>"110110001",
  5381=>"111101000",
  5382=>"010110110",
  5383=>"000100110",
  5384=>"000000010",
  5385=>"000001000",
  5386=>"110110110",
  5387=>"100111100",
  5388=>"000000000",
  5389=>"000000000",
  5390=>"001000000",
  5391=>"001001111",
  5392=>"000000000",
  5393=>"101111111",
  5394=>"111101100",
  5395=>"111111011",
  5396=>"111111011",
  5397=>"100111111",
  5398=>"001111111",
  5399=>"111111111",
  5400=>"100101000",
  5401=>"001111111",
  5402=>"111111110",
  5403=>"111011011",
  5404=>"011111111",
  5405=>"000000000",
  5406=>"101001001",
  5407=>"000000100",
  5408=>"110000111",
  5409=>"111111111",
  5410=>"111111111",
  5411=>"110111000",
  5412=>"000000000",
  5413=>"110100000",
  5414=>"000100100",
  5415=>"010110100",
  5416=>"100110111",
  5417=>"110000001",
  5418=>"111111111",
  5419=>"000010011",
  5420=>"111011001",
  5421=>"001101111",
  5422=>"110111000",
  5423=>"110110100",
  5424=>"001001101",
  5425=>"111101000",
  5426=>"000000000",
  5427=>"001011000",
  5428=>"000000000",
  5429=>"110110110",
  5430=>"000000110",
  5431=>"000000001",
  5432=>"000001111",
  5433=>"010011000",
  5434=>"100001001",
  5435=>"110000000",
  5436=>"111101101",
  5437=>"001010111",
  5438=>"111111110",
  5439=>"111010000",
  5440=>"000111111",
  5441=>"111001100",
  5442=>"001011011",
  5443=>"000000000",
  5444=>"011011111",
  5445=>"000000011",
  5446=>"111100000",
  5447=>"000000001",
  5448=>"101000000",
  5449=>"111111011",
  5450=>"111011000",
  5451=>"111111111",
  5452=>"111111111",
  5453=>"001000000",
  5454=>"100001000",
  5455=>"100110100",
  5456=>"011111111",
  5457=>"000000101",
  5458=>"000000000",
  5459=>"111111111",
  5460=>"000000000",
  5461=>"010110000",
  5462=>"000001001",
  5463=>"100000100",
  5464=>"101001100",
  5465=>"100111000",
  5466=>"100110111",
  5467=>"110100100",
  5468=>"011010111",
  5469=>"000000000",
  5470=>"001001101",
  5471=>"110111111",
  5472=>"000001111",
  5473=>"000000000",
  5474=>"100011011",
  5475=>"100000000",
  5476=>"101101111",
  5477=>"100101111",
  5478=>"000000100",
  5479=>"111111110",
  5480=>"111111111",
  5481=>"111011111",
  5482=>"101111111",
  5483=>"000111111",
  5484=>"000000000",
  5485=>"000000000",
  5486=>"000010111",
  5487=>"111111111",
  5488=>"111111111",
  5489=>"001000001",
  5490=>"111111111",
  5491=>"000000000",
  5492=>"000000000",
  5493=>"100000000",
  5494=>"000000111",
  5495=>"011001001",
  5496=>"000000000",
  5497=>"001001000",
  5498=>"100010111",
  5499=>"111110010",
  5500=>"111011111",
  5501=>"000000000",
  5502=>"111111000",
  5503=>"111100100",
  5504=>"100000000",
  5505=>"000000000",
  5506=>"000000100",
  5507=>"111011000",
  5508=>"111111111",
  5509=>"100100100",
  5510=>"001100000",
  5511=>"111001001",
  5512=>"000000000",
  5513=>"111111111",
  5514=>"100100100",
  5515=>"000101111",
  5516=>"111111111",
  5517=>"111111111",
  5518=>"000000000",
  5519=>"111111111",
  5520=>"011000101",
  5521=>"111101100",
  5522=>"101001110",
  5523=>"110000000",
  5524=>"001001000",
  5525=>"111111111",
  5526=>"100100111",
  5527=>"001001111",
  5528=>"011011111",
  5529=>"111111011",
  5530=>"100000000",
  5531=>"111111111",
  5532=>"111011111",
  5533=>"000000111",
  5534=>"000000000",
  5535=>"111111011",
  5536=>"000000000",
  5537=>"011011001",
  5538=>"100100100",
  5539=>"011111111",
  5540=>"110111111",
  5541=>"001101010",
  5542=>"000011010",
  5543=>"001000000",
  5544=>"111111111",
  5545=>"000000000",
  5546=>"101000000",
  5547=>"000101101",
  5548=>"111100110",
  5549=>"111111111",
  5550=>"111011001",
  5551=>"100111111",
  5552=>"111111011",
  5553=>"001000000",
  5554=>"000000000",
  5555=>"111111111",
  5556=>"000000011",
  5557=>"000000001",
  5558=>"011111111",
  5559=>"111111111",
  5560=>"000011111",
  5561=>"111111111",
  5562=>"011110110",
  5563=>"100011110",
  5564=>"100000010",
  5565=>"000000000",
  5566=>"111111000",
  5567=>"100001111",
  5568=>"110110011",
  5569=>"111100000",
  5570=>"000000010",
  5571=>"111111111",
  5572=>"000001011",
  5573=>"100000000",
  5574=>"100111111",
  5575=>"111100000",
  5576=>"000010010",
  5577=>"111011111",
  5578=>"110010110",
  5579=>"100110110",
  5580=>"000110111",
  5581=>"101000010",
  5582=>"001011010",
  5583=>"011011000",
  5584=>"101111111",
  5585=>"010110100",
  5586=>"011111110",
  5587=>"111011011",
  5588=>"000110001",
  5589=>"111110111",
  5590=>"100100100",
  5591=>"000001001",
  5592=>"000000000",
  5593=>"110100100",
  5594=>"000000000",
  5595=>"000000101",
  5596=>"000001011",
  5597=>"000111111",
  5598=>"001001100",
  5599=>"000000001",
  5600=>"000011011",
  5601=>"111111111",
  5602=>"000000000",
  5603=>"100111000",
  5604=>"111111100",
  5605=>"111101111",
  5606=>"000101111",
  5607=>"111011101",
  5608=>"111110110",
  5609=>"100100001",
  5610=>"111000000",
  5611=>"111111100",
  5612=>"000000100",
  5613=>"100100110",
  5614=>"000000000",
  5615=>"000000000",
  5616=>"000000000",
  5617=>"111111011",
  5618=>"000000000",
  5619=>"100100110",
  5620=>"000000000",
  5621=>"111111111",
  5622=>"000000000",
  5623=>"110011110",
  5624=>"000000111",
  5625=>"000110100",
  5626=>"000111111",
  5627=>"000000000",
  5628=>"111111111",
  5629=>"111111111",
  5630=>"000011111",
  5631=>"000000000",
  5632=>"111111111",
  5633=>"010000000",
  5634=>"000000000",
  5635=>"001000000",
  5636=>"111011011",
  5637=>"000100100",
  5638=>"000000000",
  5639=>"101100100",
  5640=>"000000001",
  5641=>"001101111",
  5642=>"001001001",
  5643=>"000000101",
  5644=>"010111111",
  5645=>"000000100",
  5646=>"000000111",
  5647=>"000110110",
  5648=>"110111111",
  5649=>"000100111",
  5650=>"001011111",
  5651=>"001001111",
  5652=>"000000000",
  5653=>"000000000",
  5654=>"100110110",
  5655=>"011011011",
  5656=>"111111110",
  5657=>"111111111",
  5658=>"101101111",
  5659=>"111111111",
  5660=>"111111111",
  5661=>"111001111",
  5662=>"110110000",
  5663=>"000000100",
  5664=>"110100000",
  5665=>"000000000",
  5666=>"000000000",
  5667=>"111001001",
  5668=>"111111110",
  5669=>"111011011",
  5670=>"001000000",
  5671=>"101100000",
  5672=>"110110011",
  5673=>"111101100",
  5674=>"000111111",
  5675=>"011011000",
  5676=>"000000000",
  5677=>"000001111",
  5678=>"111110110",
  5679=>"111110111",
  5680=>"000000000",
  5681=>"000000000",
  5682=>"001011011",
  5683=>"111111111",
  5684=>"111100111",
  5685=>"101011011",
  5686=>"000001011",
  5687=>"100100111",
  5688=>"111101111",
  5689=>"111000111",
  5690=>"011111111",
  5691=>"001000000",
  5692=>"000000100",
  5693=>"001000000",
  5694=>"110111111",
  5695=>"000000110",
  5696=>"111100100",
  5697=>"011111111",
  5698=>"111110110",
  5699=>"000000000",
  5700=>"000110110",
  5701=>"110110000",
  5702=>"000010000",
  5703=>"111111111",
  5704=>"001000000",
  5705=>"101101001",
  5706=>"000000000",
  5707=>"000000000",
  5708=>"000000000",
  5709=>"100111111",
  5710=>"000000000",
  5711=>"001101111",
  5712=>"100110000",
  5713=>"111111111",
  5714=>"000001010",
  5715=>"011001000",
  5716=>"000000001",
  5717=>"111100101",
  5718=>"001000000",
  5719=>"000000000",
  5720=>"000111111",
  5721=>"011011011",
  5722=>"111000000",
  5723=>"001111001",
  5724=>"000000000",
  5725=>"111000000",
  5726=>"001011111",
  5727=>"111111000",
  5728=>"111001111",
  5729=>"000000000",
  5730=>"100000101",
  5731=>"000000000",
  5732=>"000000110",
  5733=>"000100100",
  5734=>"111111111",
  5735=>"000000000",
  5736=>"001000000",
  5737=>"111000100",
  5738=>"000000000",
  5739=>"000010110",
  5740=>"111111111",
  5741=>"111111111",
  5742=>"111111111",
  5743=>"000100000",
  5744=>"111110110",
  5745=>"011001011",
  5746=>"001001011",
  5747=>"000011011",
  5748=>"111111010",
  5749=>"111110000",
  5750=>"011001001",
  5751=>"001111111",
  5752=>"000010111",
  5753=>"000111111",
  5754=>"000000000",
  5755=>"111111110",
  5756=>"000000000",
  5757=>"100110111",
  5758=>"110100000",
  5759=>"111111111",
  5760=>"010000000",
  5761=>"110010000",
  5762=>"000000000",
  5763=>"000010111",
  5764=>"111111111",
  5765=>"111111111",
  5766=>"000000000",
  5767=>"011011011",
  5768=>"000000100",
  5769=>"000110111",
  5770=>"111111111",
  5771=>"111111111",
  5772=>"100000101",
  5773=>"101111111",
  5774=>"111111111",
  5775=>"000000000",
  5776=>"111101100",
  5777=>"100100101",
  5778=>"111111111",
  5779=>"100000000",
  5780=>"000000100",
  5781=>"100100100",
  5782=>"000000000",
  5783=>"001000000",
  5784=>"111111111",
  5785=>"000000000",
  5786=>"000000000",
  5787=>"000000111",
  5788=>"000000000",
  5789=>"010011111",
  5790=>"111111111",
  5791=>"010111100",
  5792=>"110100111",
  5793=>"111000000",
  5794=>"111111111",
  5795=>"000011111",
  5796=>"000001001",
  5797=>"110111111",
  5798=>"101111111",
  5799=>"111111111",
  5800=>"111000000",
  5801=>"000000000",
  5802=>"000000000",
  5803=>"000000000",
  5804=>"111110001",
  5805=>"000000000",
  5806=>"011111111",
  5807=>"001000000",
  5808=>"000000000",
  5809=>"110111111",
  5810=>"111111000",
  5811=>"000000000",
  5812=>"110111100",
  5813=>"111111101",
  5814=>"110110000",
  5815=>"000111111",
  5816=>"111111111",
  5817=>"000000000",
  5818=>"100001000",
  5819=>"000000000",
  5820=>"011111111",
  5821=>"111111111",
  5822=>"010000000",
  5823=>"111011001",
  5824=>"111001111",
  5825=>"111111011",
  5826=>"011000101",
  5827=>"000000000",
  5828=>"000000000",
  5829=>"000000001",
  5830=>"111111011",
  5831=>"011111011",
  5832=>"010011001",
  5833=>"000000000",
  5834=>"100100000",
  5835=>"110110000",
  5836=>"000000010",
  5837=>"000110111",
  5838=>"111110111",
  5839=>"000000111",
  5840=>"001000100",
  5841=>"111111111",
  5842=>"000000100",
  5843=>"110100000",
  5844=>"100000100",
  5845=>"111111111",
  5846=>"000000001",
  5847=>"001100111",
  5848=>"000000110",
  5849=>"111111111",
  5850=>"011111111",
  5851=>"001000000",
  5852=>"100100010",
  5853=>"011000100",
  5854=>"010000000",
  5855=>"111111111",
  5856=>"111001111",
  5857=>"001001011",
  5858=>"111111000",
  5859=>"111011011",
  5860=>"000000000",
  5861=>"100101001",
  5862=>"000000000",
  5863=>"111110100",
  5864=>"111011111",
  5865=>"000000000",
  5866=>"111111111",
  5867=>"111010000",
  5868=>"000000000",
  5869=>"010000000",
  5870=>"000010111",
  5871=>"000000000",
  5872=>"011000110",
  5873=>"000000011",
  5874=>"110100000",
  5875=>"000000001",
  5876=>"000000000",
  5877=>"111111010",
  5878=>"001101111",
  5879=>"111111111",
  5880=>"000000000",
  5881=>"110111011",
  5882=>"111111000",
  5883=>"111111000",
  5884=>"100100111",
  5885=>"100100000",
  5886=>"000000001",
  5887=>"111111111",
  5888=>"111111111",
  5889=>"011111011",
  5890=>"101000111",
  5891=>"111011011",
  5892=>"111101111",
  5893=>"100000000",
  5894=>"100000000",
  5895=>"111111110",
  5896=>"111001111",
  5897=>"000000000",
  5898=>"110111111",
  5899=>"000000000",
  5900=>"111111111",
  5901=>"011111111",
  5902=>"010111111",
  5903=>"000000000",
  5904=>"000100110",
  5905=>"110000000",
  5906=>"000000100",
  5907=>"000000000",
  5908=>"000000000",
  5909=>"000000000",
  5910=>"000100000",
  5911=>"000000011",
  5912=>"111111111",
  5913=>"000010000",
  5914=>"111110110",
  5915=>"000000001",
  5916=>"100000010",
  5917=>"000001001",
  5918=>"000111111",
  5919=>"111001000",
  5920=>"001000010",
  5921=>"000000000",
  5922=>"100111111",
  5923=>"111111111",
  5924=>"111111101",
  5925=>"111100000",
  5926=>"000000011",
  5927=>"011111100",
  5928=>"000000000",
  5929=>"000000000",
  5930=>"011000000",
  5931=>"001000000",
  5932=>"000100000",
  5933=>"111111110",
  5934=>"000000000",
  5935=>"000000000",
  5936=>"111111111",
  5937=>"111111111",
  5938=>"000000110",
  5939=>"111111111",
  5940=>"011111111",
  5941=>"111111111",
  5942=>"000000000",
  5943=>"000001111",
  5944=>"000000000",
  5945=>"100101111",
  5946=>"000000000",
  5947=>"000000000",
  5948=>"000000000",
  5949=>"001001101",
  5950=>"000110111",
  5951=>"000000000",
  5952=>"111101100",
  5953=>"101001011",
  5954=>"111111111",
  5955=>"000000000",
  5956=>"000111100",
  5957=>"000000000",
  5958=>"010111111",
  5959=>"111111111",
  5960=>"110111111",
  5961=>"000000001",
  5962=>"111111010",
  5963=>"000000000",
  5964=>"000000100",
  5965=>"100111111",
  5966=>"010000000",
  5967=>"000000000",
  5968=>"100100100",
  5969=>"011011111",
  5970=>"111110000",
  5971=>"000000000",
  5972=>"000011011",
  5973=>"011000000",
  5974=>"111111111",
  5975=>"111110111",
  5976=>"001101111",
  5977=>"111000000",
  5978=>"111111000",
  5979=>"000000001",
  5980=>"111111111",
  5981=>"000000000",
  5982=>"111111111",
  5983=>"111111111",
  5984=>"000100111",
  5985=>"111111111",
  5986=>"001000000",
  5987=>"111111111",
  5988=>"100101000",
  5989=>"010000000",
  5990=>"000000000",
  5991=>"001001011",
  5992=>"000000000",
  5993=>"111111111",
  5994=>"111111111",
  5995=>"000101101",
  5996=>"100001001",
  5997=>"000000001",
  5998=>"000111011",
  5999=>"000100000",
  6000=>"000000000",
  6001=>"000000000",
  6002=>"111111010",
  6003=>"111100100",
  6004=>"000111110",
  6005=>"111000000",
  6006=>"000010000",
  6007=>"111111111",
  6008=>"000000000",
  6009=>"000000000",
  6010=>"000000000",
  6011=>"110111011",
  6012=>"000000111",
  6013=>"111111111",
  6014=>"000000000",
  6015=>"111011111",
  6016=>"100000000",
  6017=>"000000000",
  6018=>"100001001",
  6019=>"111111000",
  6020=>"110110111",
  6021=>"000000000",
  6022=>"011011100",
  6023=>"001001110",
  6024=>"111110000",
  6025=>"000000000",
  6026=>"000011001",
  6027=>"000011010",
  6028=>"111111111",
  6029=>"000000110",
  6030=>"111111111",
  6031=>"000000000",
  6032=>"000000001",
  6033=>"111001101",
  6034=>"000100111",
  6035=>"000000001",
  6036=>"111111010",
  6037=>"010110000",
  6038=>"110000000",
  6039=>"001011001",
  6040=>"111111111",
  6041=>"010011011",
  6042=>"000000000",
  6043=>"011111100",
  6044=>"111111011",
  6045=>"111111110",
  6046=>"111000000",
  6047=>"111011011",
  6048=>"111111111",
  6049=>"001000000",
  6050=>"101101111",
  6051=>"110111111",
  6052=>"000000110",
  6053=>"111111111",
  6054=>"000000111",
  6055=>"000000111",
  6056=>"110110110",
  6057=>"001000000",
  6058=>"000011111",
  6059=>"111101111",
  6060=>"000000000",
  6061=>"000000001",
  6062=>"100111111",
  6063=>"111000000",
  6064=>"111111000",
  6065=>"000000011",
  6066=>"111111111",
  6067=>"000000000",
  6068=>"000000000",
  6069=>"111111000",
  6070=>"111111111",
  6071=>"100110100",
  6072=>"000000110",
  6073=>"001000010",
  6074=>"111111111",
  6075=>"100101111",
  6076=>"001001111",
  6077=>"110111000",
  6078=>"011000111",
  6079=>"000000000",
  6080=>"000001011",
  6081=>"011111111",
  6082=>"111111000",
  6083=>"000000000",
  6084=>"011000000",
  6085=>"110011000",
  6086=>"011010100",
  6087=>"000000100",
  6088=>"000011111",
  6089=>"000000111",
  6090=>"011000110",
  6091=>"110110110",
  6092=>"000000000",
  6093=>"000000000",
  6094=>"000000100",
  6095=>"000011100",
  6096=>"011110000",
  6097=>"111100011",
  6098=>"111010010",
  6099=>"111111111",
  6100=>"010110100",
  6101=>"000000111",
  6102=>"101110100",
  6103=>"111111111",
  6104=>"000000000",
  6105=>"110111111",
  6106=>"100110110",
  6107=>"010011011",
  6108=>"000000001",
  6109=>"110110100",
  6110=>"111111111",
  6111=>"001011111",
  6112=>"001001101",
  6113=>"000110000",
  6114=>"011111111",
  6115=>"111111111",
  6116=>"001100111",
  6117=>"000000000",
  6118=>"001000111",
  6119=>"000000000",
  6120=>"111110100",
  6121=>"111111111",
  6122=>"111111110",
  6123=>"000000000",
  6124=>"010000000",
  6125=>"000000000",
  6126=>"000000101",
  6127=>"000000000",
  6128=>"100100000",
  6129=>"111111111",
  6130=>"111111111",
  6131=>"011011111",
  6132=>"001111111",
  6133=>"111100000",
  6134=>"111111111",
  6135=>"110110110",
  6136=>"000000100",
  6137=>"011001101",
  6138=>"000011001",
  6139=>"001001000",
  6140=>"111001111",
  6141=>"000000000",
  6142=>"101001111",
  6143=>"000000000",
  6144=>"000000000",
  6145=>"111000001",
  6146=>"111111000",
  6147=>"100000000",
  6148=>"001111111",
  6149=>"111111001",
  6150=>"110111110",
  6151=>"000000000",
  6152=>"111111111",
  6153=>"111111111",
  6154=>"000000000",
  6155=>"001000000",
  6156=>"000010111",
  6157=>"111000110",
  6158=>"100001001",
  6159=>"111111111",
  6160=>"011111000",
  6161=>"111100111",
  6162=>"111100000",
  6163=>"000000000",
  6164=>"010000111",
  6165=>"000001000",
  6166=>"100010000",
  6167=>"111111111",
  6168=>"111110100",
  6169=>"000000000",
  6170=>"111110000",
  6171=>"111111100",
  6172=>"000110010",
  6173=>"011100100",
  6174=>"110110100",
  6175=>"100100110",
  6176=>"111111111",
  6177=>"100000000",
  6178=>"001000000",
  6179=>"000110100",
  6180=>"011011011",
  6181=>"111111111",
  6182=>"000000001",
  6183=>"000010110",
  6184=>"011111011",
  6185=>"000000000",
  6186=>"110100100",
  6187=>"110000000",
  6188=>"011011111",
  6189=>"111011101",
  6190=>"111111111",
  6191=>"000000000",
  6192=>"001000000",
  6193=>"000000000",
  6194=>"000000000",
  6195=>"111011011",
  6196=>"000000000",
  6197=>"111111111",
  6198=>"111111111",
  6199=>"111101101",
  6200=>"000000000",
  6201=>"111000001",
  6202=>"100100101",
  6203=>"000000000",
  6204=>"111111111",
  6205=>"000000000",
  6206=>"000001001",
  6207=>"000000000",
  6208=>"011000111",
  6209=>"000000000",
  6210=>"000000000",
  6211=>"000110100",
  6212=>"000000100",
  6213=>"111110110",
  6214=>"111000111",
  6215=>"111111111",
  6216=>"001011001",
  6217=>"111101110",
  6218=>"111111010",
  6219=>"001110000",
  6220=>"000000000",
  6221=>"100100101",
  6222=>"000000101",
  6223=>"111100111",
  6224=>"000010000",
  6225=>"101001000",
  6226=>"011000101",
  6227=>"000100101",
  6228=>"111111111",
  6229=>"000000111",
  6230=>"111000000",
  6231=>"000000000",
  6232=>"000001001",
  6233=>"000000000",
  6234=>"000000110",
  6235=>"101101001",
  6236=>"111111011",
  6237=>"111111100",
  6238=>"000101111",
  6239=>"011111000",
  6240=>"111111111",
  6241=>"001000000",
  6242=>"000000000",
  6243=>"011111111",
  6244=>"111101001",
  6245=>"111010000",
  6246=>"110111111",
  6247=>"111101100",
  6248=>"000000000",
  6249=>"000000000",
  6250=>"011011011",
  6251=>"000000100",
  6252=>"000000010",
  6253=>"010000100",
  6254=>"101111111",
  6255=>"000001111",
  6256=>"000000011",
  6257=>"011011110",
  6258=>"000110011",
  6259=>"000000000",
  6260=>"111111111",
  6261=>"000000001",
  6262=>"111111110",
  6263=>"000000001",
  6264=>"100110100",
  6265=>"000000000",
  6266=>"000100100",
  6267=>"111100100",
  6268=>"000100110",
  6269=>"111011001",
  6270=>"000000000",
  6271=>"001011011",
  6272=>"000010000",
  6273=>"010010000",
  6274=>"111111111",
  6275=>"111111111",
  6276=>"000000011",
  6277=>"000000000",
  6278=>"100000000",
  6279=>"110000000",
  6280=>"111001000",
  6281=>"000000111",
  6282=>"000111111",
  6283=>"111001011",
  6284=>"100010010",
  6285=>"111111111",
  6286=>"000001111",
  6287=>"111111011",
  6288=>"000000000",
  6289=>"111111111",
  6290=>"000011000",
  6291=>"000011111",
  6292=>"001000000",
  6293=>"111111110",
  6294=>"010100110",
  6295=>"011011011",
  6296=>"001000000",
  6297=>"111110010",
  6298=>"000000000",
  6299=>"010111111",
  6300=>"111110111",
  6301=>"111000000",
  6302=>"000000000",
  6303=>"000001001",
  6304=>"000000000",
  6305=>"111110111",
  6306=>"111111101",
  6307=>"011111111",
  6308=>"000100110",
  6309=>"111111111",
  6310=>"001111111",
  6311=>"110110111",
  6312=>"111000111",
  6313=>"000000001",
  6314=>"111111111",
  6315=>"111111011",
  6316=>"001011011",
  6317=>"100110100",
  6318=>"001001011",
  6319=>"101000001",
  6320=>"111111000",
  6321=>"100100011",
  6322=>"001001011",
  6323=>"110111111",
  6324=>"001111111",
  6325=>"100000000",
  6326=>"000001111",
  6327=>"011111111",
  6328=>"010000000",
  6329=>"111111111",
  6330=>"000110110",
  6331=>"010010000",
  6332=>"000000111",
  6333=>"000101111",
  6334=>"110010010",
  6335=>"100111000",
  6336=>"101100111",
  6337=>"000000000",
  6338=>"000000000",
  6339=>"000011000",
  6340=>"111111001",
  6341=>"000000000",
  6342=>"111111111",
  6343=>"000001000",
  6344=>"000000000",
  6345=>"000111011",
  6346=>"001111111",
  6347=>"000001010",
  6348=>"111101101",
  6349=>"011011101",
  6350=>"000000111",
  6351=>"000000000",
  6352=>"111111111",
  6353=>"000000001",
  6354=>"101101111",
  6355=>"111101000",
  6356=>"000000110",
  6357=>"111111111",
  6358=>"000000000",
  6359=>"000001011",
  6360=>"000000000",
  6361=>"000000000",
  6362=>"000010000",
  6363=>"111101111",
  6364=>"100100110",
  6365=>"000000111",
  6366=>"000000000",
  6367=>"000000110",
  6368=>"000000001",
  6369=>"000000000",
  6370=>"111111111",
  6371=>"111000111",
  6372=>"101101111",
  6373=>"100100111",
  6374=>"111111111",
  6375=>"001000000",
  6376=>"100000100",
  6377=>"111111111",
  6378=>"111011111",
  6379=>"000000100",
  6380=>"110000000",
  6381=>"000000000",
  6382=>"000000111",
  6383=>"000000111",
  6384=>"011011010",
  6385=>"001000000",
  6386=>"100000100",
  6387=>"000110111",
  6388=>"010110110",
  6389=>"111100000",
  6390=>"111111110",
  6391=>"001000100",
  6392=>"010110000",
  6393=>"010010011",
  6394=>"111111111",
  6395=>"000000000",
  6396=>"001001001",
  6397=>"111110111",
  6398=>"000010011",
  6399=>"000000000",
  6400=>"100110100",
  6401=>"001001000",
  6402=>"110111100",
  6403=>"111110000",
  6404=>"011000000",
  6405=>"111111111",
  6406=>"111111110",
  6407=>"011011000",
  6408=>"110110011",
  6409=>"000000000",
  6410=>"100100100",
  6411=>"000000000",
  6412=>"000000000",
  6413=>"000000111",
  6414=>"011011000",
  6415=>"010111110",
  6416=>"000000000",
  6417=>"100110111",
  6418=>"100100110",
  6419=>"000000000",
  6420=>"000000100",
  6421=>"011111111",
  6422=>"100100100",
  6423=>"000000001",
  6424=>"111111111",
  6425=>"000011111",
  6426=>"101101000",
  6427=>"111101111",
  6428=>"000000000",
  6429=>"110110111",
  6430=>"111111111",
  6431=>"000000001",
  6432=>"100111111",
  6433=>"100110111",
  6434=>"000011111",
  6435=>"000000111",
  6436=>"001000001",
  6437=>"000000000",
  6438=>"000000001",
  6439=>"000000111",
  6440=>"001101101",
  6441=>"000000000",
  6442=>"000000000",
  6443=>"000000000",
  6444=>"000000101",
  6445=>"001100111",
  6446=>"000111111",
  6447=>"111111111",
  6448=>"011011011",
  6449=>"100000000",
  6450=>"011000000",
  6451=>"001001000",
  6452=>"000000000",
  6453=>"001101001",
  6454=>"111110000",
  6455=>"000000111",
  6456=>"010111001",
  6457=>"000000000",
  6458=>"000100100",
  6459=>"011000010",
  6460=>"000000000",
  6461=>"001000001",
  6462=>"000000000",
  6463=>"000000011",
  6464=>"111001111",
  6465=>"000000000",
  6466=>"000000000",
  6467=>"000111011",
  6468=>"010111000",
  6469=>"110111111",
  6470=>"000000000",
  6471=>"111111111",
  6472=>"000000000",
  6473=>"010000111",
  6474=>"000000111",
  6475=>"001001000",
  6476=>"111111111",
  6477=>"111111111",
  6478=>"111111111",
  6479=>"001011111",
  6480=>"010001111",
  6481=>"111111111",
  6482=>"000000010",
  6483=>"001011111",
  6484=>"000111111",
  6485=>"110110111",
  6486=>"000000000",
  6487=>"111110100",
  6488=>"000000000",
  6489=>"111111111",
  6490=>"111100100",
  6491=>"100000111",
  6492=>"010000111",
  6493=>"111100111",
  6494=>"111111111",
  6495=>"111111110",
  6496=>"000110011",
  6497=>"111111111",
  6498=>"001001011",
  6499=>"000000000",
  6500=>"011011011",
  6501=>"110110111",
  6502=>"000000000",
  6503=>"110000000",
  6504=>"010000000",
  6505=>"111111111",
  6506=>"111111111",
  6507=>"111011000",
  6508=>"111111011",
  6509=>"111110010",
  6510=>"111111111",
  6511=>"000000000",
  6512=>"000000101",
  6513=>"001111111",
  6514=>"111000000",
  6515=>"000000101",
  6516=>"000000000",
  6517=>"011010111",
  6518=>"011111011",
  6519=>"000000011",
  6520=>"000000000",
  6521=>"000000000",
  6522=>"111111111",
  6523=>"000000000",
  6524=>"111111111",
  6525=>"000000011",
  6526=>"101000000",
  6527=>"111000000",
  6528=>"111111111",
  6529=>"000000000",
  6530=>"110110111",
  6531=>"000000000",
  6532=>"110111111",
  6533=>"111011000",
  6534=>"011001001",
  6535=>"001000001",
  6536=>"111111111",
  6537=>"010000000",
  6538=>"001101101",
  6539=>"000000011",
  6540=>"111111111",
  6541=>"111100100",
  6542=>"000000001",
  6543=>"000010000",
  6544=>"011011011",
  6545=>"111110111",
  6546=>"111111111",
  6547=>"000000000",
  6548=>"010000000",
  6549=>"000000100",
  6550=>"000000100",
  6551=>"000000000",
  6552=>"111111111",
  6553=>"001000111",
  6554=>"100000000",
  6555=>"111111111",
  6556=>"110110110",
  6557=>"111111111",
  6558=>"000010010",
  6559=>"111101110",
  6560=>"100000000",
  6561=>"000000000",
  6562=>"000000000",
  6563=>"000000110",
  6564=>"001000000",
  6565=>"111111111",
  6566=>"111111111",
  6567=>"110111111",
  6568=>"111111111",
  6569=>"000000000",
  6570=>"000000101",
  6571=>"000000110",
  6572=>"011000000",
  6573=>"100000000",
  6574=>"000000000",
  6575=>"111111011",
  6576=>"111111111",
  6577=>"011000000",
  6578=>"111011000",
  6579=>"101000101",
  6580=>"000001011",
  6581=>"011010111",
  6582=>"000011111",
  6583=>"101000001",
  6584=>"000000000",
  6585=>"000111111",
  6586=>"111111100",
  6587=>"111111111",
  6588=>"000110110",
  6589=>"011011011",
  6590=>"001001011",
  6591=>"000100000",
  6592=>"000000011",
  6593=>"000000000",
  6594=>"000000000",
  6595=>"111111111",
  6596=>"100010011",
  6597=>"100110011",
  6598=>"010011111",
  6599=>"000111111",
  6600=>"110000000",
  6601=>"000000000",
  6602=>"111101111",
  6603=>"111111111",
  6604=>"111111111",
  6605=>"000111111",
  6606=>"110111011",
  6607=>"111100100",
  6608=>"001001001",
  6609=>"000000000",
  6610=>"000010100",
  6611=>"001001000",
  6612=>"000000001",
  6613=>"111111111",
  6614=>"101101111",
  6615=>"111111111",
  6616=>"111111111",
  6617=>"101001101",
  6618=>"011111010",
  6619=>"111111111",
  6620=>"000011111",
  6621=>"000000000",
  6622=>"110110111",
  6623=>"001111011",
  6624=>"000000000",
  6625=>"000011001",
  6626=>"001000000",
  6627=>"001011111",
  6628=>"111000111",
  6629=>"111111111",
  6630=>"110110111",
  6631=>"011001000",
  6632=>"000010011",
  6633=>"111001111",
  6634=>"011001000",
  6635=>"111011000",
  6636=>"111000000",
  6637=>"100001011",
  6638=>"001000000",
  6639=>"111111111",
  6640=>"000010000",
  6641=>"111111111",
  6642=>"000000000",
  6643=>"000010011",
  6644=>"000000001",
  6645=>"111010000",
  6646=>"000000000",
  6647=>"110110110",
  6648=>"001001000",
  6649=>"000011001",
  6650=>"000000000",
  6651=>"001001011",
  6652=>"111111111",
  6653=>"011111100",
  6654=>"101111111",
  6655=>"000000000",
  6656=>"110100000",
  6657=>"111000000",
  6658=>"101101111",
  6659=>"010111111",
  6660=>"000000000",
  6661=>"010000000",
  6662=>"000000000",
  6663=>"111000111",
  6664=>"100100000",
  6665=>"000111100",
  6666=>"111010111",
  6667=>"000001100",
  6668=>"000000110",
  6669=>"001111111",
  6670=>"110110000",
  6671=>"000000100",
  6672=>"011111000",
  6673=>"101111111",
  6674=>"000010000",
  6675=>"000000000",
  6676=>"000000111",
  6677=>"111101000",
  6678=>"111100000",
  6679=>"111111000",
  6680=>"111111101",
  6681=>"101100000",
  6682=>"111111111",
  6683=>"111111001",
  6684=>"000111111",
  6685=>"111011000",
  6686=>"011110110",
  6687=>"111111101",
  6688=>"110000001",
  6689=>"011111111",
  6690=>"111111111",
  6691=>"100110000",
  6692=>"111111111",
  6693=>"111111111",
  6694=>"000000000",
  6695=>"000001111",
  6696=>"111100000",
  6697=>"000000000",
  6698=>"000000111",
  6699=>"000111111",
  6700=>"110100100",
  6701=>"111111111",
  6702=>"111000000",
  6703=>"111110110",
  6704=>"111100000",
  6705=>"000000000",
  6706=>"111100000",
  6707=>"110110000",
  6708=>"000000000",
  6709=>"000001001",
  6710=>"000000111",
  6711=>"001000100",
  6712=>"000011000",
  6713=>"000101101",
  6714=>"000000000",
  6715=>"100011011",
  6716=>"111111000",
  6717=>"000000000",
  6718=>"001001000",
  6719=>"111110000",
  6720=>"111111111",
  6721=>"000000111",
  6722=>"100111111",
  6723=>"100100110",
  6724=>"111110000",
  6725=>"000000000",
  6726=>"111011011",
  6727=>"111111111",
  6728=>"111011001",
  6729=>"000000000",
  6730=>"111111111",
  6731=>"011111111",
  6732=>"111111111",
  6733=>"001101111",
  6734=>"110110111",
  6735=>"111111000",
  6736=>"000000000",
  6737=>"000000000",
  6738=>"000010100",
  6739=>"101111000",
  6740=>"000001111",
  6741=>"100000000",
  6742=>"001011001",
  6743=>"000000000",
  6744=>"000000000",
  6745=>"101000000",
  6746=>"111111010",
  6747=>"000000000",
  6748=>"000111111",
  6749=>"000000000",
  6750=>"101111111",
  6751=>"011111111",
  6752=>"000100000",
  6753=>"111111100",
  6754=>"001000000",
  6755=>"000001111",
  6756=>"000000000",
  6757=>"000000001",
  6758=>"001111111",
  6759=>"001111111",
  6760=>"000011000",
  6761=>"000011111",
  6762=>"111100000",
  6763=>"110111110",
  6764=>"110000000",
  6765=>"111111000",
  6766=>"111111111",
  6767=>"000111000",
  6768=>"010111111",
  6769=>"111111111",
  6770=>"000111111",
  6771=>"000001000",
  6772=>"111110111",
  6773=>"000100110",
  6774=>"011001001",
  6775=>"001000001",
  6776=>"001001000",
  6777=>"000000111",
  6778=>"000000000",
  6779=>"111111000",
  6780=>"011001111",
  6781=>"111010000",
  6782=>"100000000",
  6783=>"000001101",
  6784=>"111111111",
  6785=>"111111000",
  6786=>"000111111",
  6787=>"000110000",
  6788=>"111111000",
  6789=>"000000111",
  6790=>"101110111",
  6791=>"000000001",
  6792=>"111010111",
  6793=>"000000011",
  6794=>"000010000",
  6795=>"000000000",
  6796=>"111111000",
  6797=>"110111111",
  6798=>"100100111",
  6799=>"000100111",
  6800=>"000000110",
  6801=>"011111111",
  6802=>"000000000",
  6803=>"111100000",
  6804=>"000000000",
  6805=>"111111111",
  6806=>"001000000",
  6807=>"111010000",
  6808=>"100111000",
  6809=>"011011111",
  6810=>"011001000",
  6811=>"100110111",
  6812=>"111101111",
  6813=>"000000011",
  6814=>"100100110",
  6815=>"100000010",
  6816=>"000000000",
  6817=>"111111111",
  6818=>"111000001",
  6819=>"111111111",
  6820=>"001000000",
  6821=>"101101000",
  6822=>"000110111",
  6823=>"000110100",
  6824=>"111111111",
  6825=>"111100110",
  6826=>"111001000",
  6827=>"101000000",
  6828=>"101111100",
  6829=>"100101111",
  6830=>"000000000",
  6831=>"000011111",
  6832=>"010000000",
  6833=>"111110110",
  6834=>"011111111",
  6835=>"111101110",
  6836=>"111111000",
  6837=>"111111111",
  6838=>"000000000",
  6839=>"100100000",
  6840=>"111000000",
  6841=>"111111000",
  6842=>"001000000",
  6843=>"101100000",
  6844=>"111000000",
  6845=>"000100000",
  6846=>"110111111",
  6847=>"011011010",
  6848=>"000000011",
  6849=>"011000000",
  6850=>"000000111",
  6851=>"111110000",
  6852=>"111111010",
  6853=>"000111111",
  6854=>"111000000",
  6855=>"001111111",
  6856=>"111111000",
  6857=>"011111111",
  6858=>"111110000",
  6859=>"011111001",
  6860=>"111110111",
  6861=>"011111111",
  6862=>"001111110",
  6863=>"111001000",
  6864=>"011000000",
  6865=>"111000000",
  6866=>"111111111",
  6867=>"111111000",
  6868=>"111000000",
  6869=>"001101000",
  6870=>"001000000",
  6871=>"000000000",
  6872=>"000000000",
  6873=>"001011000",
  6874=>"000001111",
  6875=>"100000111",
  6876=>"000000000",
  6877=>"000000100",
  6878=>"011000000",
  6879=>"100100110",
  6880=>"000000001",
  6881=>"000000000",
  6882=>"000111011",
  6883=>"111000011",
  6884=>"111110000",
  6885=>"000100111",
  6886=>"011111001",
  6887=>"111000000",
  6888=>"011011111",
  6889=>"011000001",
  6890=>"101001001",
  6891=>"111111000",
  6892=>"000000111",
  6893=>"000000111",
  6894=>"111111111",
  6895=>"111111001",
  6896=>"111100000",
  6897=>"000100111",
  6898=>"111001000",
  6899=>"111111101",
  6900=>"000000000",
  6901=>"111110100",
  6902=>"000100111",
  6903=>"000000000",
  6904=>"000000111",
  6905=>"000000000",
  6906=>"000000000",
  6907=>"000011001",
  6908=>"011111000",
  6909=>"001001111",
  6910=>"100100000",
  6911=>"000010111",
  6912=>"111100000",
  6913=>"010111111",
  6914=>"100001000",
  6915=>"000000100",
  6916=>"110000110",
  6917=>"000000111",
  6918=>"111111000",
  6919=>"111111100",
  6920=>"111110000",
  6921=>"000110111",
  6922=>"111100000",
  6923=>"000000100",
  6924=>"000000110",
  6925=>"000001001",
  6926=>"000101000",
  6927=>"000011010",
  6928=>"110111111",
  6929=>"111111011",
  6930=>"111000000",
  6931=>"111000001",
  6932=>"001111000",
  6933=>"111111111",
  6934=>"111100000",
  6935=>"000000111",
  6936=>"000101111",
  6937=>"000000000",
  6938=>"000111101",
  6939=>"000000111",
  6940=>"001001000",
  6941=>"000001011",
  6942=>"111111111",
  6943=>"011010111",
  6944=>"000000001",
  6945=>"010100110",
  6946=>"000110000",
  6947=>"111101101",
  6948=>"000011111",
  6949=>"111111111",
  6950=>"011111100",
  6951=>"111111010",
  6952=>"111111110",
  6953=>"000000000",
  6954=>"000000000",
  6955=>"000000000",
  6956=>"001010000",
  6957=>"001000000",
  6958=>"000011111",
  6959=>"011111111",
  6960=>"001101111",
  6961=>"001111111",
  6962=>"000010000",
  6963=>"000000000",
  6964=>"000000000",
  6965=>"000000010",
  6966=>"000000000",
  6967=>"111111001",
  6968=>"000010111",
  6969=>"110000111",
  6970=>"100000000",
  6971=>"000010000",
  6972=>"000100000",
  6973=>"001111111",
  6974=>"001111111",
  6975=>"110111111",
  6976=>"111111000",
  6977=>"000000000",
  6978=>"000110111",
  6979=>"001001010",
  6980=>"111010111",
  6981=>"000000110",
  6982=>"011110110",
  6983=>"111100100",
  6984=>"000000000",
  6985=>"000000001",
  6986=>"100000111",
  6987=>"111101000",
  6988=>"000000100",
  6989=>"000000001",
  6990=>"111111101",
  6991=>"000011111",
  6992=>"000001001",
  6993=>"111000000",
  6994=>"000110000",
  6995=>"000100000",
  6996=>"000010010",
  6997=>"111111111",
  6998=>"000000001",
  6999=>"000000111",
  7000=>"111111111",
  7001=>"000000001",
  7002=>"111110110",
  7003=>"111001000",
  7004=>"100110101",
  7005=>"111111111",
  7006=>"000000111",
  7007=>"011110100",
  7008=>"000111111",
  7009=>"000000000",
  7010=>"101101001",
  7011=>"111000000",
  7012=>"011000000",
  7013=>"000000011",
  7014=>"111011111",
  7015=>"000000111",
  7016=>"111110110",
  7017=>"111101111",
  7018=>"000000111",
  7019=>"111001001",
  7020=>"110111011",
  7021=>"000000001",
  7022=>"000101111",
  7023=>"000111111",
  7024=>"000000000",
  7025=>"000111111",
  7026=>"100100111",
  7027=>"011111100",
  7028=>"111000000",
  7029=>"010000010",
  7030=>"000101111",
  7031=>"000000101",
  7032=>"000100111",
  7033=>"111001111",
  7034=>"000101111",
  7035=>"111001001",
  7036=>"000001000",
  7037=>"111111101",
  7038=>"010111010",
  7039=>"000111111",
  7040=>"110111111",
  7041=>"101101001",
  7042=>"000000000",
  7043=>"000000000",
  7044=>"000000000",
  7045=>"000000111",
  7046=>"110001111",
  7047=>"111000111",
  7048=>"000000111",
  7049=>"101111000",
  7050=>"111100000",
  7051=>"001111111",
  7052=>"111111111",
  7053=>"000110110",
  7054=>"111111001",
  7055=>"111000111",
  7056=>"111111010",
  7057=>"111100100",
  7058=>"011011000",
  7059=>"011011000",
  7060=>"111101000",
  7061=>"000000001",
  7062=>"111111111",
  7063=>"000101111",
  7064=>"000000111",
  7065=>"111011001",
  7066=>"111001001",
  7067=>"000000111",
  7068=>"110111111",
  7069=>"111110000",
  7070=>"000000000",
  7071=>"000000111",
  7072=>"000000000",
  7073=>"110111111",
  7074=>"000100111",
  7075=>"111111111",
  7076=>"100100111",
  7077=>"111000000",
  7078=>"111100000",
  7079=>"001111111",
  7080=>"111011111",
  7081=>"000000100",
  7082=>"000011111",
  7083=>"001111111",
  7084=>"000000000",
  7085=>"111111100",
  7086=>"000100000",
  7087=>"000100110",
  7088=>"111000000",
  7089=>"110000111",
  7090=>"000000000",
  7091=>"111000000",
  7092=>"000111111",
  7093=>"000100000",
  7094=>"111111111",
  7095=>"111111100",
  7096=>"000001111",
  7097=>"110000111",
  7098=>"001111111",
  7099=>"011011110",
  7100=>"111001000",
  7101=>"111000000",
  7102=>"111111000",
  7103=>"000010011",
  7104=>"100100000",
  7105=>"111100000",
  7106=>"000000111",
  7107=>"111111000",
  7108=>"001001000",
  7109=>"000000101",
  7110=>"000000011",
  7111=>"111011001",
  7112=>"000000000",
  7113=>"011111111",
  7114=>"000100111",
  7115=>"000000111",
  7116=>"001011000",
  7117=>"000001111",
  7118=>"011111111",
  7119=>"111111111",
  7120=>"100111111",
  7121=>"000010110",
  7122=>"000000000",
  7123=>"000000000",
  7124=>"111111001",
  7125=>"000000111",
  7126=>"111100000",
  7127=>"000001001",
  7128=>"000100111",
  7129=>"110000000",
  7130=>"000000111",
  7131=>"111011111",
  7132=>"011011101",
  7133=>"001101100",
  7134=>"100011011",
  7135=>"111100001",
  7136=>"011000000",
  7137=>"111111011",
  7138=>"110110111",
  7139=>"111011111",
  7140=>"111111001",
  7141=>"000000011",
  7142=>"001000000",
  7143=>"000011111",
  7144=>"111001101",
  7145=>"000000000",
  7146=>"011010010",
  7147=>"000111001",
  7148=>"000000111",
  7149=>"000000111",
  7150=>"111000000",
  7151=>"001000000",
  7152=>"111111111",
  7153=>"100110000",
  7154=>"100000000",
  7155=>"111101000",
  7156=>"111101000",
  7157=>"111010000",
  7158=>"000000100",
  7159=>"111001000",
  7160=>"111011000",
  7161=>"111001111",
  7162=>"110100001",
  7163=>"111000000",
  7164=>"000000000",
  7165=>"011111110",
  7166=>"110000001",
  7167=>"000000000",
  7168=>"011010011",
  7169=>"011111110",
  7170=>"000000000",
  7171=>"000000000",
  7172=>"100100101",
  7173=>"001000100",
  7174=>"000000000",
  7175=>"000000000",
  7176=>"111100000",
  7177=>"011111101",
  7178=>"111111111",
  7179=>"000000110",
  7180=>"111111100",
  7181=>"000111000",
  7182=>"100100000",
  7183=>"000000000",
  7184=>"001000001",
  7185=>"100111111",
  7186=>"000000000",
  7187=>"111111111",
  7188=>"111111101",
  7189=>"000000101",
  7190=>"111000000",
  7191=>"000000000",
  7192=>"001001001",
  7193=>"010010010",
  7194=>"001100100",
  7195=>"111111000",
  7196=>"000100110",
  7197=>"000000000",
  7198=>"111111001",
  7199=>"001111001",
  7200=>"000100100",
  7201=>"111000100",
  7202=>"000000000",
  7203=>"010110110",
  7204=>"000000001",
  7205=>"000000111",
  7206=>"001000000",
  7207=>"000000001",
  7208=>"000000000",
  7209=>"011001111",
  7210=>"000000000",
  7211=>"000111111",
  7212=>"001001001",
  7213=>"111001001",
  7214=>"100000000",
  7215=>"100111110",
  7216=>"001011011",
  7217=>"000000111",
  7218=>"000111111",
  7219=>"000000000",
  7220=>"100000011",
  7221=>"100110010",
  7222=>"001001001",
  7223=>"111000000",
  7224=>"000000000",
  7225=>"000000111",
  7226=>"000000000",
  7227=>"110111111",
  7228=>"111001111",
  7229=>"101111100",
  7230=>"101001001",
  7231=>"001000000",
  7232=>"011000001",
  7233=>"110000000",
  7234=>"111111111",
  7235=>"110000000",
  7236=>"000000010",
  7237=>"111111111",
  7238=>"000000100",
  7239=>"111111111",
  7240=>"111111111",
  7241=>"111110110",
  7242=>"001000000",
  7243=>"000000000",
  7244=>"001000000",
  7245=>"001001111",
  7246=>"001010010",
  7247=>"000000000",
  7248=>"111110110",
  7249=>"111111111",
  7250=>"000000111",
  7251=>"111111011",
  7252=>"000000000",
  7253=>"001001000",
  7254=>"000100110",
  7255=>"111111100",
  7256=>"000000100",
  7257=>"111111110",
  7258=>"011111111",
  7259=>"100000100",
  7260=>"011000000",
  7261=>"111100100",
  7262=>"000000000",
  7263=>"011011111",
  7264=>"000000111",
  7265=>"101100100",
  7266=>"000111111",
  7267=>"000001111",
  7268=>"000011011",
  7269=>"000000000",
  7270=>"111110001",
  7271=>"010000000",
  7272=>"000100100",
  7273=>"000000000",
  7274=>"111010000",
  7275=>"111111111",
  7276=>"110110100",
  7277=>"111000100",
  7278=>"000001000",
  7279=>"000000001",
  7280=>"000101111",
  7281=>"111110100",
  7282=>"111000001",
  7283=>"001001010",
  7284=>"111111000",
  7285=>"000001000",
  7286=>"000000000",
  7287=>"000000000",
  7288=>"000000001",
  7289=>"000000100",
  7290=>"001011111",
  7291=>"000000000",
  7292=>"110000000",
  7293=>"111111111",
  7294=>"111111111",
  7295=>"000000000",
  7296=>"111100000",
  7297=>"000000000",
  7298=>"111111010",
  7299=>"111100110",
  7300=>"110110110",
  7301=>"000000000",
  7302=>"110111001",
  7303=>"001000100",
  7304=>"111111100",
  7305=>"101111111",
  7306=>"000000000",
  7307=>"000000000",
  7308=>"000001011",
  7309=>"001111111",
  7310=>"000110101",
  7311=>"000010000",
  7312=>"000000111",
  7313=>"011011000",
  7314=>"011000111",
  7315=>"111111111",
  7316=>"001111011",
  7317=>"010100100",
  7318=>"000000000",
  7319=>"111100000",
  7320=>"111100100",
  7321=>"111111100",
  7322=>"111111111",
  7323=>"111111011",
  7324=>"111111101",
  7325=>"010001011",
  7326=>"000100101",
  7327=>"000000000",
  7328=>"111111111",
  7329=>"000110000",
  7330=>"001001111",
  7331=>"000000000",
  7332=>"011011111",
  7333=>"000000111",
  7334=>"000000100",
  7335=>"011001001",
  7336=>"111111111",
  7337=>"111111011",
  7338=>"000111000",
  7339=>"111111111",
  7340=>"001111111",
  7341=>"110110000",
  7342=>"001000100",
  7343=>"011100010",
  7344=>"110000000",
  7345=>"100100001",
  7346=>"000100100",
  7347=>"000000000",
  7348=>"100101111",
  7349=>"011011111",
  7350=>"000000000",
  7351=>"111000000",
  7352=>"001000000",
  7353=>"111111000",
  7354=>"000000000",
  7355=>"011001001",
  7356=>"111100101",
  7357=>"111111111",
  7358=>"111111111",
  7359=>"000000000",
  7360=>"000000000",
  7361=>"011101111",
  7362=>"001001000",
  7363=>"001001000",
  7364=>"000110110",
  7365=>"111111110",
  7366=>"001011000",
  7367=>"001000100",
  7368=>"000111111",
  7369=>"000000000",
  7370=>"111111111",
  7371=>"011111111",
  7372=>"100100000",
  7373=>"001001100",
  7374=>"100100100",
  7375=>"000000011",
  7376=>"110100000",
  7377=>"111000000",
  7378=>"111100000",
  7379=>"111111110",
  7380=>"011001101",
  7381=>"000001000",
  7382=>"111111111",
  7383=>"001100000",
  7384=>"000000000",
  7385=>"011011111",
  7386=>"000000000",
  7387=>"001011111",
  7388=>"000000000",
  7389=>"000000100",
  7390=>"111001101",
  7391=>"110110110",
  7392=>"000000000",
  7393=>"000000000",
  7394=>"110111111",
  7395=>"011001111",
  7396=>"111111001",
  7397=>"001100100",
  7398=>"111111111",
  7399=>"111001111",
  7400=>"111111110",
  7401=>"000101111",
  7402=>"011011010",
  7403=>"111111111",
  7404=>"111111111",
  7405=>"100011011",
  7406=>"000111101",
  7407=>"000110111",
  7408=>"000000000",
  7409=>"011000000",
  7410=>"000001011",
  7411=>"011000001",
  7412=>"000000000",
  7413=>"000110111",
  7414=>"111111111",
  7415=>"000000000",
  7416=>"100000000",
  7417=>"000000000",
  7418=>"000000101",
  7419=>"000001001",
  7420=>"000000000",
  7421=>"000000000",
  7422=>"111000100",
  7423=>"000000100",
  7424=>"000001100",
  7425=>"000000000",
  7426=>"111111110",
  7427=>"000000100",
  7428=>"000100100",
  7429=>"110110000",
  7430=>"111111111",
  7431=>"110110000",
  7432=>"111111000",
  7433=>"000000000",
  7434=>"100100111",
  7435=>"011011100",
  7436=>"100100000",
  7437=>"011111111",
  7438=>"001100111",
  7439=>"000100100",
  7440=>"111110110",
  7441=>"101000000",
  7442=>"111111101",
  7443=>"000000111",
  7444=>"000000001",
  7445=>"000110111",
  7446=>"111111011",
  7447=>"000100000",
  7448=>"111011011",
  7449=>"111111111",
  7450=>"000000000",
  7451=>"000001111",
  7452=>"111111111",
  7453=>"001111111",
  7454=>"111110000",
  7455=>"111110110",
  7456=>"000100111",
  7457=>"000000101",
  7458=>"000100111",
  7459=>"111111001",
  7460=>"000000110",
  7461=>"011000000",
  7462=>"111111111",
  7463=>"111111001",
  7464=>"111110000",
  7465=>"000000000",
  7466=>"011000000",
  7467=>"000000001",
  7468=>"111111001",
  7469=>"111001101",
  7470=>"100111010",
  7471=>"000000111",
  7472=>"000111111",
  7473=>"000000000",
  7474=>"111111111",
  7475=>"111111100",
  7476=>"100000110",
  7477=>"001000000",
  7478=>"111111111",
  7479=>"000011111",
  7480=>"111100101",
  7481=>"100100101",
  7482=>"000000101",
  7483=>"111111111",
  7484=>"001101100",
  7485=>"111101001",
  7486=>"000000111",
  7487=>"111000000",
  7488=>"111111111",
  7489=>"111111110",
  7490=>"011001000",
  7491=>"111010110",
  7492=>"011101001",
  7493=>"111111111",
  7494=>"100100011",
  7495=>"110110010",
  7496=>"000110110",
  7497=>"111111110",
  7498=>"011111110",
  7499=>"111110111",
  7500=>"111111111",
  7501=>"111100000",
  7502=>"001001001",
  7503=>"100100110",
  7504=>"110110111",
  7505=>"000100101",
  7506=>"111111111",
  7507=>"111110111",
  7508=>"100100111",
  7509=>"000001011",
  7510=>"010000000",
  7511=>"111111111",
  7512=>"111111000",
  7513=>"000000110",
  7514=>"000001011",
  7515=>"011001000",
  7516=>"100111011",
  7517=>"000000000",
  7518=>"111010010",
  7519=>"000000001",
  7520=>"111111111",
  7521=>"111100111",
  7522=>"100000000",
  7523=>"000000000",
  7524=>"110100100",
  7525=>"111111111",
  7526=>"001000000",
  7527=>"111100100",
  7528=>"110110110",
  7529=>"000000010",
  7530=>"100111000",
  7531=>"110110111",
  7532=>"011011011",
  7533=>"100000001",
  7534=>"100000000",
  7535=>"000001000",
  7536=>"111011000",
  7537=>"000000111",
  7538=>"000000000",
  7539=>"111111100",
  7540=>"110101111",
  7541=>"011111110",
  7542=>"000000011",
  7543=>"111100000",
  7544=>"111111111",
  7545=>"011001000",
  7546=>"111111100",
  7547=>"100100111",
  7548=>"000010111",
  7549=>"011001001",
  7550=>"011011000",
  7551=>"111111111",
  7552=>"111111101",
  7553=>"000000001",
  7554=>"100100100",
  7555=>"001000000",
  7556=>"101111000",
  7557=>"000110110",
  7558=>"010000000",
  7559=>"001011111",
  7560=>"111001001",
  7561=>"011011000",
  7562=>"100100100",
  7563=>"000000010",
  7564=>"000000000",
  7565=>"100110000",
  7566=>"011000111",
  7567=>"111111111",
  7568=>"111111111",
  7569=>"111000000",
  7570=>"111111111",
  7571=>"111111111",
  7572=>"000111111",
  7573=>"000010000",
  7574=>"111001111",
  7575=>"111001011",
  7576=>"110100100",
  7577=>"000111110",
  7578=>"110000000",
  7579=>"000110111",
  7580=>"000000100",
  7581=>"111111010",
  7582=>"111111111",
  7583=>"000000000",
  7584=>"111001111",
  7585=>"101001000",
  7586=>"000000001",
  7587=>"000000001",
  7588=>"001000001",
  7589=>"111111111",
  7590=>"111111111",
  7591=>"100111111",
  7592=>"000000010",
  7593=>"110110101",
  7594=>"000000000",
  7595=>"111110001",
  7596=>"000000000",
  7597=>"001000001",
  7598=>"000000011",
  7599=>"101111011",
  7600=>"000010010",
  7601=>"000000000",
  7602=>"111111010",
  7603=>"111101100",
  7604=>"000000000",
  7605=>"000000000",
  7606=>"000110000",
  7607=>"000000111",
  7608=>"011111111",
  7609=>"111110101",
  7610=>"111111111",
  7611=>"111111100",
  7612=>"101001000",
  7613=>"111111111",
  7614=>"100000111",
  7615=>"111111000",
  7616=>"100110110",
  7617=>"110111111",
  7618=>"110111111",
  7619=>"001001001",
  7620=>"011111000",
  7621=>"000100111",
  7622=>"000000111",
  7623=>"001001001",
  7624=>"001111111",
  7625=>"001000000",
  7626=>"100100100",
  7627=>"100100100",
  7628=>"111001101",
  7629=>"100101101",
  7630=>"011111100",
  7631=>"000001001",
  7632=>"111111001",
  7633=>"111110100",
  7634=>"111100101",
  7635=>"000000100",
  7636=>"000000000",
  7637=>"111111110",
  7638=>"100100111",
  7639=>"000100111",
  7640=>"000000100",
  7641=>"011010100",
  7642=>"000100111",
  7643=>"000000000",
  7644=>"000110010",
  7645=>"010000000",
  7646=>"000000000",
  7647=>"011101001",
  7648=>"011011111",
  7649=>"110110000",
  7650=>"011000100",
  7651=>"001001000",
  7652=>"011011111",
  7653=>"111101111",
  7654=>"001011000",
  7655=>"111000000",
  7656=>"001000110",
  7657=>"000001001",
  7658=>"111111000",
  7659=>"000000000",
  7660=>"110110110",
  7661=>"111111111",
  7662=>"110000000",
  7663=>"111111111",
  7664=>"000100111",
  7665=>"011001000",
  7666=>"011011000",
  7667=>"000000011",
  7668=>"011010000",
  7669=>"011001001",
  7670=>"011001110",
  7671=>"110111111",
  7672=>"001011011",
  7673=>"000000000",
  7674=>"111111001",
  7675=>"111101111",
  7676=>"001000001",
  7677=>"011000000",
  7678=>"000000001",
  7679=>"111111111",
  7680=>"110110110",
  7681=>"111000000",
  7682=>"111111000",
  7683=>"000111110",
  7684=>"000111111",
  7685=>"001101001",
  7686=>"000001111",
  7687=>"111000111",
  7688=>"000000000",
  7689=>"111111010",
  7690=>"111111111",
  7691=>"110000000",
  7692=>"000000001",
  7693=>"011100100",
  7694=>"001101000",
  7695=>"011000111",
  7696=>"000010011",
  7697=>"010111111",
  7698=>"000000000",
  7699=>"000000000",
  7700=>"100000000",
  7701=>"000110000",
  7702=>"111010000",
  7703=>"000000000",
  7704=>"010110000",
  7705=>"001111111",
  7706=>"000001111",
  7707=>"111000000",
  7708=>"100000111",
  7709=>"111000101",
  7710=>"000000001",
  7711=>"000000001",
  7712=>"010111111",
  7713=>"111100110",
  7714=>"000001001",
  7715=>"111111111",
  7716=>"110100000",
  7717=>"000000000",
  7718=>"000000000",
  7719=>"000000000",
  7720=>"000000011",
  7721=>"000000111",
  7722=>"100110000",
  7723=>"111111111",
  7724=>"111000001",
  7725=>"100111101",
  7726=>"111111100",
  7727=>"000000000",
  7728=>"011000111",
  7729=>"000000100",
  7730=>"000000001",
  7731=>"100011001",
  7732=>"000111100",
  7733=>"000000000",
  7734=>"100000000",
  7735=>"000000000",
  7736=>"010111111",
  7737=>"111111011",
  7738=>"001000001",
  7739=>"000000000",
  7740=>"111111100",
  7741=>"111101000",
  7742=>"001011111",
  7743=>"111001000",
  7744=>"111110001",
  7745=>"000000100",
  7746=>"100000111",
  7747=>"111000000",
  7748=>"010011010",
  7749=>"000000000",
  7750=>"111111010",
  7751=>"100101001",
  7752=>"000000000",
  7753=>"010000001",
  7754=>"111111111",
  7755=>"111000001",
  7756=>"111011001",
  7757=>"000000100",
  7758=>"000000000",
  7759=>"000000110",
  7760=>"111001001",
  7761=>"000000000",
  7762=>"000000000",
  7763=>"111111111",
  7764=>"000111111",
  7765=>"000000111",
  7766=>"111101111",
  7767=>"000000000",
  7768=>"000001001",
  7769=>"000000111",
  7770=>"111111100",
  7771=>"000000110",
  7772=>"000000110",
  7773=>"000000001",
  7774=>"111111001",
  7775=>"100001000",
  7776=>"000000000",
  7777=>"110000000",
  7778=>"110000000",
  7779=>"000101111",
  7780=>"000000111",
  7781=>"000110010",
  7782=>"111111111",
  7783=>"000000111",
  7784=>"111111110",
  7785=>"100100100",
  7786=>"111111000",
  7787=>"000011000",
  7788=>"110111011",
  7789=>"001000000",
  7790=>"110111011",
  7791=>"110111111",
  7792=>"000000000",
  7793=>"111011111",
  7794=>"100110111",
  7795=>"110000000",
  7796=>"111111111",
  7797=>"010000111",
  7798=>"000000110",
  7799=>"111001000",
  7800=>"000000000",
  7801=>"011111111",
  7802=>"000000100",
  7803=>"111000000",
  7804=>"111011000",
  7805=>"011010000",
  7806=>"000000000",
  7807=>"111111111",
  7808=>"111111111",
  7809=>"011000000",
  7810=>"111111111",
  7811=>"000100111",
  7812=>"000000111",
  7813=>"000000000",
  7814=>"110100111",
  7815=>"111011011",
  7816=>"001000000",
  7817=>"000001001",
  7818=>"111111111",
  7819=>"111000111",
  7820=>"000000111",
  7821=>"000111111",
  7822=>"011111000",
  7823=>"110000000",
  7824=>"111100110",
  7825=>"100111111",
  7826=>"000111111",
  7827=>"100010111",
  7828=>"000111111",
  7829=>"011011011",
  7830=>"000000000",
  7831=>"111111000",
  7832=>"001001111",
  7833=>"000000111",
  7834=>"000000001",
  7835=>"000111111",
  7836=>"111111111",
  7837=>"111111000",
  7838=>"111000111",
  7839=>"111111111",
  7840=>"000000011",
  7841=>"111011000",
  7842=>"000111111",
  7843=>"110111111",
  7844=>"000010000",
  7845=>"111111000",
  7846=>"100000000",
  7847=>"001001000",
  7848=>"111100000",
  7849=>"000000000",
  7850=>"111111100",
  7851=>"111111111",
  7852=>"111000110",
  7853=>"100111111",
  7854=>"111111111",
  7855=>"100111000",
  7856=>"011000001",
  7857=>"000100100",
  7858=>"111111111",
  7859=>"111111111",
  7860=>"111111111",
  7861=>"111111001",
  7862=>"000000011",
  7863=>"110000000",
  7864=>"011100011",
  7865=>"111111111",
  7866=>"110111100",
  7867=>"111000001",
  7868=>"000000000",
  7869=>"011011001",
  7870=>"000110000",
  7871=>"111111010",
  7872=>"000011010",
  7873=>"110000000",
  7874=>"000000000",
  7875=>"001110000",
  7876=>"000111000",
  7877=>"001111111",
  7878=>"000010011",
  7879=>"011011011",
  7880=>"000000111",
  7881=>"111001001",
  7882=>"100000001",
  7883=>"000000001",
  7884=>"111001000",
  7885=>"110101111",
  7886=>"100100000",
  7887=>"111000000",
  7888=>"111000000",
  7889=>"000000100",
  7890=>"001000011",
  7891=>"000011001",
  7892=>"101111100",
  7893=>"000001001",
  7894=>"110110000",
  7895=>"000000111",
  7896=>"000000111",
  7897=>"011111111",
  7898=>"000011001",
  7899=>"011111111",
  7900=>"010000000",
  7901=>"111000100",
  7902=>"000000000",
  7903=>"111111000",
  7904=>"111101110",
  7905=>"101000000",
  7906=>"111111111",
  7907=>"111111111",
  7908=>"000000111",
  7909=>"000000111",
  7910=>"111111111",
  7911=>"111111111",
  7912=>"010000000",
  7913=>"110100000",
  7914=>"111111011",
  7915=>"000000111",
  7916=>"000000000",
  7917=>"101110111",
  7918=>"111111111",
  7919=>"111000000",
  7920=>"111011000",
  7921=>"111000000",
  7922=>"000101111",
  7923=>"110100000",
  7924=>"000111111",
  7925=>"011001000",
  7926=>"000011000",
  7927=>"000000000",
  7928=>"101111111",
  7929=>"000000111",
  7930=>"111001111",
  7931=>"101101000",
  7932=>"110111111",
  7933=>"111011110",
  7934=>"111010000",
  7935=>"010110111",
  7936=>"101101111",
  7937=>"000000000",
  7938=>"111111001",
  7939=>"000001000",
  7940=>"000000000",
  7941=>"111101110",
  7942=>"111111111",
  7943=>"000000111",
  7944=>"001000000",
  7945=>"000110111",
  7946=>"111011000",
  7947=>"111111011",
  7948=>"100000100",
  7949=>"001000000",
  7950=>"111010000",
  7951=>"111111000",
  7952=>"110111000",
  7953=>"011111111",
  7954=>"111001011",
  7955=>"111111011",
  7956=>"000000000",
  7957=>"111000010",
  7958=>"000110000",
  7959=>"111111111",
  7960=>"000000000",
  7961=>"000000000",
  7962=>"011000000",
  7963=>"000000000",
  7964=>"000000100",
  7965=>"111111000",
  7966=>"111001111",
  7967=>"000000000",
  7968=>"110100000",
  7969=>"111011001",
  7970=>"111111111",
  7971=>"000110110",
  7972=>"000010111",
  7973=>"001100111",
  7974=>"011100100",
  7975=>"111000011",
  7976=>"111011000",
  7977=>"000000000",
  7978=>"000000000",
  7979=>"101000000",
  7980=>"000000000",
  7981=>"111111000",
  7982=>"111000111",
  7983=>"000000001",
  7984=>"111001111",
  7985=>"111111111",
  7986=>"010101100",
  7987=>"101000000",
  7988=>"100101111",
  7989=>"000000001",
  7990=>"000000000",
  7991=>"101000000",
  7992=>"111000000",
  7993=>"000100100",
  7994=>"100011000",
  7995=>"111000000",
  7996=>"111000001",
  7997=>"100000101",
  7998=>"110111111",
  7999=>"000011111",
  8000=>"101111000",
  8001=>"001000110",
  8002=>"001001111",
  8003=>"000000000",
  8004=>"111111111",
  8005=>"000000111",
  8006=>"010000111",
  8007=>"000000000",
  8008=>"000000100",
  8009=>"000000010",
  8010=>"000000100",
  8011=>"000001011",
  8012=>"111011111",
  8013=>"111110111",
  8014=>"001001000",
  8015=>"000000111",
  8016=>"000000011",
  8017=>"111001001",
  8018=>"000111111",
  8019=>"000111111",
  8020=>"100011000",
  8021=>"011011001",
  8022=>"000000000",
  8023=>"111100110",
  8024=>"000111111",
  8025=>"111110110",
  8026=>"111101111",
  8027=>"001000111",
  8028=>"000000001",
  8029=>"001000000",
  8030=>"011000111",
  8031=>"000000111",
  8032=>"000000000",
  8033=>"000000111",
  8034=>"001001111",
  8035=>"000000111",
  8036=>"111111011",
  8037=>"011111000",
  8038=>"111100000",
  8039=>"000000011",
  8040=>"000000100",
  8041=>"111001000",
  8042=>"000000101",
  8043=>"111000000",
  8044=>"000011001",
  8045=>"000000001",
  8046=>"011011111",
  8047=>"101111111",
  8048=>"010000111",
  8049=>"111111111",
  8050=>"111010000",
  8051=>"101100000",
  8052=>"111110111",
  8053=>"111011001",
  8054=>"000101111",
  8055=>"110000000",
  8056=>"000000000",
  8057=>"010010110",
  8058=>"000000111",
  8059=>"000000111",
  8060=>"111110100",
  8061=>"111010000",
  8062=>"111111111",
  8063=>"111111111",
  8064=>"000001011",
  8065=>"000000000",
  8066=>"000000000",
  8067=>"010100111",
  8068=>"100110000",
  8069=>"000000000",
  8070=>"000000110",
  8071=>"001000000",
  8072=>"111000000",
  8073=>"000000001",
  8074=>"111000000",
  8075=>"000111000",
  8076=>"111111111",
  8077=>"000000100",
  8078=>"001000000",
  8079=>"111000000",
  8080=>"000110111",
  8081=>"000111111",
  8082=>"000011111",
  8083=>"011100110",
  8084=>"011111111",
  8085=>"000010011",
  8086=>"000110111",
  8087=>"111111011",
  8088=>"000000000",
  8089=>"111110111",
  8090=>"111000000",
  8091=>"110111111",
  8092=>"000011111",
  8093=>"111111000",
  8094=>"100111000",
  8095=>"000000000",
  8096=>"110000000",
  8097=>"110111001",
  8098=>"110110011",
  8099=>"111000111",
  8100=>"000000000",
  8101=>"111111111",
  8102=>"000110111",
  8103=>"010000000",
  8104=>"010000001",
  8105=>"001000110",
  8106=>"000111101",
  8107=>"000000101",
  8108=>"010000000",
  8109=>"111100100",
  8110=>"111000000",
  8111=>"111111111",
  8112=>"111111110",
  8113=>"000000000",
  8114=>"000000010",
  8115=>"111111111",
  8116=>"111111000",
  8117=>"001001000",
  8118=>"000000010",
  8119=>"100000000",
  8120=>"001000000",
  8121=>"111000000",
  8122=>"111111111",
  8123=>"011111011",
  8124=>"000000000",
  8125=>"000000111",
  8126=>"000011000",
  8127=>"000000000",
  8128=>"101000000",
  8129=>"111111111",
  8130=>"111000111",
  8131=>"111110111",
  8132=>"101101000",
  8133=>"000000100",
  8134=>"111000000",
  8135=>"111101000",
  8136=>"100000001",
  8137=>"001000100",
  8138=>"111111000",
  8139=>"000001000",
  8140=>"111111111",
  8141=>"001011111",
  8142=>"110111000",
  8143=>"110000110",
  8144=>"000001111",
  8145=>"001111101",
  8146=>"000010110",
  8147=>"000000000",
  8148=>"000000000",
  8149=>"111001101",
  8150=>"111000000",
  8151=>"001000000",
  8152=>"111111011",
  8153=>"111100111",
  8154=>"111110110",
  8155=>"111111111",
  8156=>"000011111",
  8157=>"011111111",
  8158=>"111100111",
  8159=>"100110011",
  8160=>"111111000",
  8161=>"111001000",
  8162=>"111111000",
  8163=>"001010010",
  8164=>"111101111",
  8165=>"000000110",
  8166=>"001011110",
  8167=>"111000100",
  8168=>"011011011",
  8169=>"111000000",
  8170=>"111000010",
  8171=>"101101111",
  8172=>"011001000",
  8173=>"111111111",
  8174=>"111111000",
  8175=>"000000000",
  8176=>"111111001",
  8177=>"011011011",
  8178=>"111111000",
  8179=>"110000000",
  8180=>"100000000",
  8181=>"011111111",
  8182=>"111111000",
  8183=>"001111110",
  8184=>"000000000",
  8185=>"001000111",
  8186=>"011001000",
  8187=>"111111000",
  8188=>"010111111",
  8189=>"001111110",
  8190=>"001000010",
  8191=>"000000000",
  8192=>"000000110",
  8193=>"110000000",
  8194=>"111110000",
  8195=>"001000000",
  8196=>"100000111",
  8197=>"011111001",
  8198=>"001001111",
  8199=>"000011100",
  8200=>"000000000",
  8201=>"000000000",
  8202=>"111000000",
  8203=>"001000001",
  8204=>"000111111",
  8205=>"000000000",
  8206=>"000100011",
  8207=>"000000000",
  8208=>"111011000",
  8209=>"000000000",
  8210=>"111111101",
  8211=>"110111111",
  8212=>"111111111",
  8213=>"110110110",
  8214=>"111111111",
  8215=>"001001111",
  8216=>"110110110",
  8217=>"111100100",
  8218=>"101000000",
  8219=>"111110110",
  8220=>"100101000",
  8221=>"000000000",
  8222=>"111111111",
  8223=>"111110100",
  8224=>"110111111",
  8225=>"000000000",
  8226=>"111111111",
  8227=>"001001001",
  8228=>"000000000",
  8229=>"001011111",
  8230=>"000010000",
  8231=>"001110010",
  8232=>"000000100",
  8233=>"000000000",
  8234=>"001111111",
  8235=>"000000000",
  8236=>"000000000",
  8237=>"000000000",
  8238=>"111111111",
  8239=>"000000100",
  8240=>"111111111",
  8241=>"111111111",
  8242=>"001000000",
  8243=>"111111111",
  8244=>"111111111",
  8245=>"000100100",
  8246=>"000000101",
  8247=>"000000000",
  8248=>"000000000",
  8249=>"011011000",
  8250=>"000011011",
  8251=>"000000000",
  8252=>"000011111",
  8253=>"011011110",
  8254=>"001000000",
  8255=>"000000000",
  8256=>"111110100",
  8257=>"111111000",
  8258=>"000100001",
  8259=>"111100100",
  8260=>"000000101",
  8261=>"000000000",
  8262=>"111111111",
  8263=>"000000000",
  8264=>"111111111",
  8265=>"000000000",
  8266=>"001000000",
  8267=>"100000111",
  8268=>"000000000",
  8269=>"111001001",
  8270=>"000000000",
  8271=>"100001010",
  8272=>"011011000",
  8273=>"111111111",
  8274=>"000101111",
  8275=>"100100000",
  8276=>"011011000",
  8277=>"000000001",
  8278=>"001101101",
  8279=>"101111111",
  8280=>"111111111",
  8281=>"111111111",
  8282=>"111111000",
  8283=>"000000000",
  8284=>"111111111",
  8285=>"000000000",
  8286=>"000000000",
  8287=>"001001000",
  8288=>"111111111",
  8289=>"000000000",
  8290=>"111001001",
  8291=>"110000111",
  8292=>"100100000",
  8293=>"111111111",
  8294=>"000000010",
  8295=>"100000000",
  8296=>"000000000",
  8297=>"111111111",
  8298=>"011011000",
  8299=>"111001000",
  8300=>"111000000",
  8301=>"011011001",
  8302=>"111111111",
  8303=>"111111000",
  8304=>"000001001",
  8305=>"000000000",
  8306=>"011010000",
  8307=>"111111111",
  8308=>"111111111",
  8309=>"000010000",
  8310=>"000110111",
  8311=>"000000100",
  8312=>"000000000",
  8313=>"111101000",
  8314=>"111111111",
  8315=>"110111000",
  8316=>"110100000",
  8317=>"011011010",
  8318=>"111111000",
  8319=>"010110111",
  8320=>"111111111",
  8321=>"000000110",
  8322=>"111110000",
  8323=>"000000000",
  8324=>"000000001",
  8325=>"111111111",
  8326=>"110000100",
  8327=>"000000000",
  8328=>"000110000",
  8329=>"000000011",
  8330=>"001011111",
  8331=>"011001000",
  8332=>"000000000",
  8333=>"110111111",
  8334=>"001000100",
  8335=>"111011111",
  8336=>"111111111",
  8337=>"000010011",
  8338=>"111011010",
  8339=>"011001001",
  8340=>"000000000",
  8341=>"111111111",
  8342=>"111111111",
  8343=>"111111111",
  8344=>"001000101",
  8345=>"000100111",
  8346=>"110000100",
  8347=>"111111111",
  8348=>"111111111",
  8349=>"110111111",
  8350=>"111001000",
  8351=>"000111111",
  8352=>"000010111",
  8353=>"011000000",
  8354=>"111111111",
  8355=>"111111011",
  8356=>"100000001",
  8357=>"000100100",
  8358=>"111111111",
  8359=>"001001000",
  8360=>"111110111",
  8361=>"111111111",
  8362=>"111111111",
  8363=>"000000100",
  8364=>"111111111",
  8365=>"000000100",
  8366=>"001000101",
  8367=>"011011111",
  8368=>"100111000",
  8369=>"111011011",
  8370=>"000000000",
  8371=>"000000000",
  8372=>"111111111",
  8373=>"011111011",
  8374=>"000000000",
  8375=>"011111111",
  8376=>"111111111",
  8377=>"111111000",
  8378=>"110100100",
  8379=>"001001000",
  8380=>"000011011",
  8381=>"001110110",
  8382=>"111111111",
  8383=>"000011010",
  8384=>"000000010",
  8385=>"111111110",
  8386=>"000000000",
  8387=>"111111000",
  8388=>"000000000",
  8389=>"000000000",
  8390=>"111111111",
  8391=>"000000000",
  8392=>"000000000",
  8393=>"001001111",
  8394=>"000000000",
  8395=>"001011010",
  8396=>"111111111",
  8397=>"001111111",
  8398=>"111111111",
  8399=>"011000000",
  8400=>"000010000",
  8401=>"000001111",
  8402=>"111111000",
  8403=>"001000000",
  8404=>"111111111",
  8405=>"001001001",
  8406=>"000010000",
  8407=>"101001101",
  8408=>"111000000",
  8409=>"110110010",
  8410=>"000000000",
  8411=>"000000000",
  8412=>"111110111",
  8413=>"100100000",
  8414=>"000000000",
  8415=>"000000000",
  8416=>"000000111",
  8417=>"000000000",
  8418=>"000000111",
  8419=>"001011010",
  8420=>"111111111",
  8421=>"111000000",
  8422=>"000000000",
  8423=>"000001111",
  8424=>"000111111",
  8425=>"110101101",
  8426=>"000001111",
  8427=>"000000110",
  8428=>"001000001",
  8429=>"010110010",
  8430=>"000000110",
  8431=>"110111111",
  8432=>"111000000",
  8433=>"111111000",
  8434=>"010111011",
  8435=>"000000000",
  8436=>"000000001",
  8437=>"001011000",
  8438=>"000000000",
  8439=>"000000000",
  8440=>"111111011",
  8441=>"101111111",
  8442=>"001011111",
  8443=>"011011011",
  8444=>"110110111",
  8445=>"001001110",
  8446=>"001000110",
  8447=>"000000000",
  8448=>"000000000",
  8449=>"011111111",
  8450=>"111111111",
  8451=>"111111111",
  8452=>"000000000",
  8453=>"100000000",
  8454=>"000000000",
  8455=>"000000111",
  8456=>"111111111",
  8457=>"000011111",
  8458=>"000000000",
  8459=>"111111111",
  8460=>"111110110",
  8461=>"000000000",
  8462=>"101111101",
  8463=>"010000000",
  8464=>"111101001",
  8465=>"011011111",
  8466=>"111011001",
  8467=>"000000000",
  8468=>"111111001",
  8469=>"100000000",
  8470=>"111111111",
  8471=>"111111000",
  8472=>"000000000",
  8473=>"000000000",
  8474=>"111010000",
  8475=>"000010100",
  8476=>"111111110",
  8477=>"000000000",
  8478=>"111111111",
  8479=>"000000111",
  8480=>"000000000",
  8481=>"101111111",
  8482=>"101000000",
  8483=>"000000111",
  8484=>"000000010",
  8485=>"000000001",
  8486=>"111110111",
  8487=>"000000000",
  8488=>"011000000",
  8489=>"001001111",
  8490=>"011111111",
  8491=>"000110111",
  8492=>"110110110",
  8493=>"100100000",
  8494=>"111111000",
  8495=>"111111111",
  8496=>"000000000",
  8497=>"000111111",
  8498=>"111111111",
  8499=>"011011000",
  8500=>"000000000",
  8501=>"000000000",
  8502=>"000000010",
  8503=>"101111011",
  8504=>"100000000",
  8505=>"100100000",
  8506=>"111111110",
  8507=>"000000000",
  8508=>"000100110",
  8509=>"000111111",
  8510=>"001101111",
  8511=>"100111000",
  8512=>"000010110",
  8513=>"111111111",
  8514=>"011111110",
  8515=>"101100100",
  8516=>"000010111",
  8517=>"111111111",
  8518=>"000000000",
  8519=>"000000111",
  8520=>"111111111",
  8521=>"111111000",
  8522=>"110110111",
  8523=>"000000000",
  8524=>"110010000",
  8525=>"111111111",
  8526=>"111000000",
  8527=>"000011111",
  8528=>"001001000",
  8529=>"110110110",
  8530=>"011010111",
  8531=>"000000000",
  8532=>"000111111",
  8533=>"011011001",
  8534=>"111111111",
  8535=>"101000000",
  8536=>"000110110",
  8537=>"000111111",
  8538=>"000000001",
  8539=>"000100111",
  8540=>"110110110",
  8541=>"101001111",
  8542=>"011000110",
  8543=>"000000000",
  8544=>"000000000",
  8545=>"111111011",
  8546=>"100110111",
  8547=>"111111111",
  8548=>"100101110",
  8549=>"000000000",
  8550=>"000000000",
  8551=>"011111111",
  8552=>"011011011",
  8553=>"001001000",
  8554=>"000100110",
  8555=>"000000000",
  8556=>"000000000",
  8557=>"110111111",
  8558=>"000101111",
  8559=>"001111111",
  8560=>"000000000",
  8561=>"000000000",
  8562=>"001101111",
  8563=>"000100111",
  8564=>"111110111",
  8565=>"000100000",
  8566=>"000000111",
  8567=>"000100111",
  8568=>"111111111",
  8569=>"000000100",
  8570=>"100100000",
  8571=>"000011111",
  8572=>"000000011",
  8573=>"110100110",
  8574=>"000011111",
  8575=>"111111111",
  8576=>"001001011",
  8577=>"011111111",
  8578=>"000000000",
  8579=>"111111111",
  8580=>"000000111",
  8581=>"000000000",
  8582=>"111111111",
  8583=>"010000000",
  8584=>"000000000",
  8585=>"111110110",
  8586=>"111111111",
  8587=>"111111000",
  8588=>"111111111",
  8589=>"001011111",
  8590=>"000000001",
  8591=>"001111011",
  8592=>"111111111",
  8593=>"111111111",
  8594=>"000000000",
  8595=>"000000000",
  8596=>"000111111",
  8597=>"000000000",
  8598=>"001000000",
  8599=>"001001100",
  8600=>"000110111",
  8601=>"110000000",
  8602=>"111111111",
  8603=>"111101101",
  8604=>"111111111",
  8605=>"000000001",
  8606=>"111011011",
  8607=>"000000111",
  8608=>"000000000",
  8609=>"000011011",
  8610=>"001001000",
  8611=>"111111111",
  8612=>"111100111",
  8613=>"000010011",
  8614=>"000000000",
  8615=>"000110110",
  8616=>"001001001",
  8617=>"000111111",
  8618=>"000000111",
  8619=>"000000000",
  8620=>"000001001",
  8621=>"110110110",
  8622=>"111111111",
  8623=>"111111111",
  8624=>"000000000",
  8625=>"111111111",
  8626=>"010110111",
  8627=>"000000000",
  8628=>"111111111",
  8629=>"010110110",
  8630=>"111111111",
  8631=>"000001111",
  8632=>"000000000",
  8633=>"010001000",
  8634=>"000000111",
  8635=>"111111111",
  8636=>"110000000",
  8637=>"000000101",
  8638=>"000000000",
  8639=>"011111111",
  8640=>"011001001",
  8641=>"000000000",
  8642=>"011111111",
  8643=>"111111101",
  8644=>"011111111",
  8645=>"000000001",
  8646=>"001000000",
  8647=>"111101101",
  8648=>"110110000",
  8649=>"000100110",
  8650=>"111101101",
  8651=>"000000000",
  8652=>"000100000",
  8653=>"100111111",
  8654=>"000000000",
  8655=>"111111000",
  8656=>"111100110",
  8657=>"111111111",
  8658=>"000000000",
  8659=>"111111001",
  8660=>"110110111",
  8661=>"001001001",
  8662=>"111111000",
  8663=>"011011111",
  8664=>"011011111",
  8665=>"000000101",
  8666=>"000001001",
  8667=>"111111101",
  8668=>"100111111",
  8669=>"111111111",
  8670=>"000000000",
  8671=>"101001000",
  8672=>"111111111",
  8673=>"000000000",
  8674=>"010111111",
  8675=>"101101111",
  8676=>"111111111",
  8677=>"001000000",
  8678=>"000000100",
  8679=>"111111000",
  8680=>"000001111",
  8681=>"000110110",
  8682=>"011010000",
  8683=>"111111111",
  8684=>"000000001",
  8685=>"000000111",
  8686=>"000000111",
  8687=>"111110000",
  8688=>"000000000",
  8689=>"111011000",
  8690=>"000000000",
  8691=>"111111111",
  8692=>"111100100",
  8693=>"000000000",
  8694=>"111111011",
  8695=>"000000000",
  8696=>"111000000",
  8697=>"111111111",
  8698=>"000000000",
  8699=>"000000000",
  8700=>"000000000",
  8701=>"000000000",
  8702=>"000000000",
  8703=>"000000000",
  8704=>"001001110",
  8705=>"111101111",
  8706=>"111111111",
  8707=>"111101000",
  8708=>"000010111",
  8709=>"111111111",
  8710=>"011111000",
  8711=>"111111111",
  8712=>"001000111",
  8713=>"001111001",
  8714=>"111111111",
  8715=>"000100000",
  8716=>"111111110",
  8717=>"111111011",
  8718=>"010111111",
  8719=>"000011111",
  8720=>"111011111",
  8721=>"111111000",
  8722=>"000000000",
  8723=>"000000000",
  8724=>"111111100",
  8725=>"111111111",
  8726=>"001000111",
  8727=>"111111111",
  8728=>"111111000",
  8729=>"001000000",
  8730=>"000010111",
  8731=>"100100000",
  8732=>"110011001",
  8733=>"110011000",
  8734=>"000001001",
  8735=>"000000011",
  8736=>"000000110",
  8737=>"110111111",
  8738=>"100100000",
  8739=>"110000000",
  8740=>"001000110",
  8741=>"111100000",
  8742=>"111111111",
  8743=>"111101101",
  8744=>"000111111",
  8745=>"111100111",
  8746=>"000000110",
  8747=>"111111111",
  8748=>"000001100",
  8749=>"111001110",
  8750=>"111100110",
  8751=>"000000000",
  8752=>"100100101",
  8753=>"111111111",
  8754=>"111111110",
  8755=>"011111010",
  8756=>"000000000",
  8757=>"100111110",
  8758=>"000000101",
  8759=>"000000111",
  8760=>"111111111",
  8761=>"000000100",
  8762=>"111111111",
  8763=>"111111111",
  8764=>"111111111",
  8765=>"000000000",
  8766=>"111011111",
  8767=>"111101111",
  8768=>"100110111",
  8769=>"111001000",
  8770=>"111110100",
  8771=>"000000101",
  8772=>"000000000",
  8773=>"000000000",
  8774=>"111111111",
  8775=>"111111111",
  8776=>"011001111",
  8777=>"000001111",
  8778=>"111111000",
  8779=>"101001001",
  8780=>"010010111",
  8781=>"110100100",
  8782=>"000000000",
  8783=>"000110010",
  8784=>"111001000",
  8785=>"111011000",
  8786=>"000000000",
  8787=>"100110000",
  8788=>"110110000",
  8789=>"001000000",
  8790=>"111111111",
  8791=>"000000100",
  8792=>"111111000",
  8793=>"000000011",
  8794=>"000000000",
  8795=>"111111101",
  8796=>"111111010",
  8797=>"111111111",
  8798=>"011111111",
  8799=>"000000100",
  8800=>"111001000",
  8801=>"000010000",
  8802=>"110111001",
  8803=>"000000000",
  8804=>"100111110",
  8805=>"111110111",
  8806=>"111010000",
  8807=>"111111111",
  8808=>"000100000",
  8809=>"111111111",
  8810=>"011011011",
  8811=>"111100100",
  8812=>"000000000",
  8813=>"000000000",
  8814=>"100110000",
  8815=>"111111111",
  8816=>"111111111",
  8817=>"111111111",
  8818=>"110100100",
  8819=>"000000000",
  8820=>"110111111",
  8821=>"111111110",
  8822=>"010100110",
  8823=>"111111010",
  8824=>"110110100",
  8825=>"011000000",
  8826=>"111110100",
  8827=>"000000001",
  8828=>"100000000",
  8829=>"000000100",
  8830=>"100100101",
  8831=>"001000000",
  8832=>"110111110",
  8833=>"111111111",
  8834=>"000000000",
  8835=>"011111000",
  8836=>"111111000",
  8837=>"101001111",
  8838=>"001111000",
  8839=>"111000000",
  8840=>"110110111",
  8841=>"111111111",
  8842=>"000000001",
  8843=>"111111111",
  8844=>"100100000",
  8845=>"011111000",
  8846=>"111000111",
  8847=>"001000101",
  8848=>"000100000",
  8849=>"111000000",
  8850=>"000111111",
  8851=>"000000110",
  8852=>"000000000",
  8853=>"110110000",
  8854=>"000000000",
  8855=>"000001000",
  8856=>"011001001",
  8857=>"000000000",
  8858=>"011111110",
  8859=>"111111000",
  8860=>"011011111",
  8861=>"100000000",
  8862=>"100000000",
  8863=>"111101111",
  8864=>"101000111",
  8865=>"111100000",
  8866=>"111111000",
  8867=>"000000100",
  8868=>"010000000",
  8869=>"111001011",
  8870=>"000000010",
  8871=>"000000000",
  8872=>"000000100",
  8873=>"100111111",
  8874=>"111111111",
  8875=>"111110111",
  8876=>"000000011",
  8877=>"100111001",
  8878=>"100100101",
  8879=>"011111111",
  8880=>"000001011",
  8881=>"000000000",
  8882=>"110010010",
  8883=>"111100001",
  8884=>"001000111",
  8885=>"111111111",
  8886=>"011011011",
  8887=>"000000011",
  8888=>"000010110",
  8889=>"011011010",
  8890=>"111111111",
  8891=>"011111111",
  8892=>"111000000",
  8893=>"110111111",
  8894=>"111000011",
  8895=>"000000111",
  8896=>"000000000",
  8897=>"000000011",
  8898=>"000111111",
  8899=>"111001001",
  8900=>"011111111",
  8901=>"111111111",
  8902=>"111111111",
  8903=>"110111111",
  8904=>"000111111",
  8905=>"111111111",
  8906=>"100110111",
  8907=>"111111101",
  8908=>"111111000",
  8909=>"111111111",
  8910=>"111111110",
  8911=>"111111001",
  8912=>"111111111",
  8913=>"001100111",
  8914=>"100111111",
  8915=>"100000000",
  8916=>"000000000",
  8917=>"011110110",
  8918=>"111111010",
  8919=>"001101110",
  8920=>"001001001",
  8921=>"101101001",
  8922=>"111111100",
  8923=>"111001000",
  8924=>"001101101",
  8925=>"000000000",
  8926=>"111111100",
  8927=>"111111001",
  8928=>"001000000",
  8929=>"111111111",
  8930=>"100111111",
  8931=>"011000000",
  8932=>"000000000",
  8933=>"110111111",
  8934=>"011110000",
  8935=>"000000000",
  8936=>"111111000",
  8937=>"000000000",
  8938=>"000011111",
  8939=>"000000111",
  8940=>"110110110",
  8941=>"000000000",
  8942=>"000000000",
  8943=>"000000000",
  8944=>"000000000",
  8945=>"001000111",
  8946=>"000100111",
  8947=>"111011000",
  8948=>"000000000",
  8949=>"001001000",
  8950=>"010010010",
  8951=>"111111011",
  8952=>"000011000",
  8953=>"000100111",
  8954=>"011001000",
  8955=>"111111000",
  8956=>"000000100",
  8957=>"000000110",
  8958=>"111111111",
  8959=>"000000000",
  8960=>"000000101",
  8961=>"111111111",
  8962=>"011011011",
  8963=>"111111111",
  8964=>"110000100",
  8965=>"111111111",
  8966=>"001011000",
  8967=>"111111111",
  8968=>"001000101",
  8969=>"000000000",
  8970=>"011000000",
  8971=>"001101000",
  8972=>"000000000",
  8973=>"111111111",
  8974=>"000000000",
  8975=>"111111111",
  8976=>"000000000",
  8977=>"001111111",
  8978=>"000001000",
  8979=>"110110110",
  8980=>"100100100",
  8981=>"000000000",
  8982=>"111101001",
  8983=>"011001111",
  8984=>"000001011",
  8985=>"111111111",
  8986=>"111111111",
  8987=>"011000000",
  8988=>"101111111",
  8989=>"111000000",
  8990=>"000000001",
  8991=>"111111111",
  8992=>"100100111",
  8993=>"111110111",
  8994=>"100100000",
  8995=>"000000001",
  8996=>"000000001",
  8997=>"000000000",
  8998=>"000001011",
  8999=>"101101111",
  9000=>"111011000",
  9001=>"000000010",
  9002=>"110100111",
  9003=>"011001000",
  9004=>"111111101",
  9005=>"000000011",
  9006=>"000001000",
  9007=>"000011000",
  9008=>"100110011",
  9009=>"111100100",
  9010=>"000100110",
  9011=>"100111111",
  9012=>"111111011",
  9013=>"000100110",
  9014=>"000000000",
  9015=>"100101111",
  9016=>"000000000",
  9017=>"000000000",
  9018=>"000000000",
  9019=>"000001000",
  9020=>"000000000",
  9021=>"110010110",
  9022=>"100000000",
  9023=>"000000100",
  9024=>"000100101",
  9025=>"100111000",
  9026=>"111111111",
  9027=>"000000000",
  9028=>"000000000",
  9029=>"000111110",
  9030=>"000111111",
  9031=>"000000000",
  9032=>"111011011",
  9033=>"100000000",
  9034=>"111111111",
  9035=>"000000000",
  9036=>"000111001",
  9037=>"110111101",
  9038=>"001001101",
  9039=>"111111111",
  9040=>"000110000",
  9041=>"001000000",
  9042=>"100111111",
  9043=>"111111001",
  9044=>"100110000",
  9045=>"111111111",
  9046=>"111111111",
  9047=>"011111111",
  9048=>"100111111",
  9049=>"111101000",
  9050=>"110111101",
  9051=>"000111111",
  9052=>"111111110",
  9053=>"000000000",
  9054=>"101111001",
  9055=>"000011111",
  9056=>"111101111",
  9057=>"011010111",
  9058=>"010111110",
  9059=>"111111111",
  9060=>"000000000",
  9061=>"000001000",
  9062=>"111111111",
  9063=>"001101001",
  9064=>"001000000",
  9065=>"000000111",
  9066=>"000000111",
  9067=>"000000000",
  9068=>"001011011",
  9069=>"111111011",
  9070=>"000010000",
  9071=>"000000111",
  9072=>"111111101",
  9073=>"000000000",
  9074=>"100100111",
  9075=>"110011111",
  9076=>"000000011",
  9077=>"000000000",
  9078=>"011111111",
  9079=>"111101111",
  9080=>"111111111",
  9081=>"000000000",
  9082=>"011000111",
  9083=>"111111100",
  9084=>"111011111",
  9085=>"000000000",
  9086=>"000000000",
  9087=>"000000000",
  9088=>"100100000",
  9089=>"111011001",
  9090=>"000000000",
  9091=>"111101101",
  9092=>"111111111",
  9093=>"110000000",
  9094=>"001000101",
  9095=>"000100111",
  9096=>"000000000",
  9097=>"001001001",
  9098=>"111111111",
  9099=>"101001001",
  9100=>"000000010",
  9101=>"110110110",
  9102=>"000000100",
  9103=>"000000000",
  9104=>"000000000",
  9105=>"000000000",
  9106=>"111011000",
  9107=>"000000000",
  9108=>"001000000",
  9109=>"001000000",
  9110=>"101100111",
  9111=>"101101000",
  9112=>"111111111",
  9113=>"011011111",
  9114=>"111111110",
  9115=>"100111100",
  9116=>"111111111",
  9117=>"000000000",
  9118=>"000000001",
  9119=>"010010000",
  9120=>"111111111",
  9121=>"100100110",
  9122=>"101101101",
  9123=>"000000010",
  9124=>"111111111",
  9125=>"011001000",
  9126=>"011011111",
  9127=>"000000000",
  9128=>"001101111",
  9129=>"000000000",
  9130=>"001011111",
  9131=>"100000000",
  9132=>"000000000",
  9133=>"111111111",
  9134=>"101100000",
  9135=>"111111111",
  9136=>"111111111",
  9137=>"111111111",
  9138=>"111111111",
  9139=>"000000011",
  9140=>"010111111",
  9141=>"101101000",
  9142=>"010100110",
  9143=>"000000000",
  9144=>"111111111",
  9145=>"000000110",
  9146=>"000011011",
  9147=>"001111111",
  9148=>"001111001",
  9149=>"111111111",
  9150=>"100111000",
  9151=>"011011011",
  9152=>"000111010",
  9153=>"110011001",
  9154=>"000000000",
  9155=>"000010110",
  9156=>"111111111",
  9157=>"001011011",
  9158=>"000000000",
  9159=>"000000000",
  9160=>"111011100",
  9161=>"000111111",
  9162=>"111111001",
  9163=>"000000000",
  9164=>"000001000",
  9165=>"111111111",
  9166=>"111111110",
  9167=>"111001000",
  9168=>"000000000",
  9169=>"000001010",
  9170=>"111001001",
  9171=>"111111111",
  9172=>"000110111",
  9173=>"001101111",
  9174=>"111111111",
  9175=>"011001011",
  9176=>"000111111",
  9177=>"001111111",
  9178=>"111110111",
  9179=>"000000111",
  9180=>"001100111",
  9181=>"111101100",
  9182=>"000000000",
  9183=>"001001111",
  9184=>"111111111",
  9185=>"111111111",
  9186=>"000000101",
  9187=>"000011111",
  9188=>"000000111",
  9189=>"000000000",
  9190=>"000010011",
  9191=>"001000000",
  9192=>"111111111",
  9193=>"000000000",
  9194=>"111000000",
  9195=>"001011001",
  9196=>"000000000",
  9197=>"011011000",
  9198=>"111111111",
  9199=>"111011000",
  9200=>"000000100",
  9201=>"111001111",
  9202=>"011001000",
  9203=>"111100100",
  9204=>"100000000",
  9205=>"000000000",
  9206=>"000001100",
  9207=>"001001001",
  9208=>"111111111",
  9209=>"100110110",
  9210=>"000000000",
  9211=>"000000000",
  9212=>"111111111",
  9213=>"111100110",
  9214=>"111111111",
  9215=>"111111111",
  9216=>"111001001",
  9217=>"000000000",
  9218=>"111111100",
  9219=>"000000000",
  9220=>"111000000",
  9221=>"000000000",
  9222=>"000001111",
  9223=>"111111111",
  9224=>"111110000",
  9225=>"110111111",
  9226=>"000000000",
  9227=>"000111111",
  9228=>"000000110",
  9229=>"000000000",
  9230=>"100111111",
  9231=>"111001011",
  9232=>"100010011",
  9233=>"000000101",
  9234=>"000000010",
  9235=>"000111111",
  9236=>"111111001",
  9237=>"101000000",
  9238=>"000000000",
  9239=>"101101111",
  9240=>"111101111",
  9241=>"000001001",
  9242=>"001000111",
  9243=>"111111110",
  9244=>"100000000",
  9245=>"000000100",
  9246=>"000100100",
  9247=>"100000010",
  9248=>"100100111",
  9249=>"001001000",
  9250=>"111111111",
  9251=>"000000000",
  9252=>"000000000",
  9253=>"111000000",
  9254=>"100000000",
  9255=>"111111000",
  9256=>"111111111",
  9257=>"111010000",
  9258=>"101101111",
  9259=>"110111111",
  9260=>"111111111",
  9261=>"000000101",
  9262=>"011101111",
  9263=>"000000111",
  9264=>"111111101",
  9265=>"000000000",
  9266=>"001100100",
  9267=>"111111111",
  9268=>"100101101",
  9269=>"010011111",
  9270=>"000000000",
  9271=>"000000000",
  9272=>"001111111",
  9273=>"111111110",
  9274=>"111111111",
  9275=>"111111111",
  9276=>"000000000",
  9277=>"000000001",
  9278=>"000000000",
  9279=>"001111111",
  9280=>"000001000",
  9281=>"000111000",
  9282=>"111111111",
  9283=>"000000111",
  9284=>"000000000",
  9285=>"111111111",
  9286=>"000000000",
  9287=>"000000000",
  9288=>"001000000",
  9289=>"111000111",
  9290=>"111111111",
  9291=>"111111111",
  9292=>"011111000",
  9293=>"111111001",
  9294=>"000000000",
  9295=>"000000000",
  9296=>"000110110",
  9297=>"000000000",
  9298=>"111110110",
  9299=>"000011111",
  9300=>"001011001",
  9301=>"001111011",
  9302=>"111001011",
  9303=>"111111110",
  9304=>"101000001",
  9305=>"100000111",
  9306=>"000000000",
  9307=>"000000000",
  9308=>"101111110",
  9309=>"000000000",
  9310=>"000000100",
  9311=>"001011001",
  9312=>"001000111",
  9313=>"011111111",
  9314=>"000000111",
  9315=>"000010000",
  9316=>"111111110",
  9317=>"000000000",
  9318=>"000000000",
  9319=>"100101001",
  9320=>"111111000",
  9321=>"111111111",
  9322=>"110011000",
  9323=>"010011111",
  9324=>"000000000",
  9325=>"111111111",
  9326=>"000000000",
  9327=>"000111111",
  9328=>"101100000",
  9329=>"000000000",
  9330=>"011111001",
  9331=>"000101111",
  9332=>"001000000",
  9333=>"110111011",
  9334=>"000000001",
  9335=>"110010000",
  9336=>"111111100",
  9337=>"111111111",
  9338=>"111011000",
  9339=>"111111111",
  9340=>"000000000",
  9341=>"000000000",
  9342=>"110100000",
  9343=>"110100000",
  9344=>"111111111",
  9345=>"111110110",
  9346=>"000000000",
  9347=>"101001001",
  9348=>"111111000",
  9349=>"101111111",
  9350=>"111011000",
  9351=>"000000000",
  9352=>"111111111",
  9353=>"111111111",
  9354=>"000000000",
  9355=>"000000000",
  9356=>"111011011",
  9357=>"111111111",
  9358=>"111101111",
  9359=>"111100110",
  9360=>"100000000",
  9361=>"111111111",
  9362=>"000100100",
  9363=>"111011000",
  9364=>"101111100",
  9365=>"000000111",
  9366=>"111111111",
  9367=>"000000100",
  9368=>"100000001",
  9369=>"111111111",
  9370=>"110000011",
  9371=>"000000000",
  9372=>"111001000",
  9373=>"000000100",
  9374=>"000000000",
  9375=>"111111111",
  9376=>"111110100",
  9377=>"011000000",
  9378=>"111111111",
  9379=>"111100000",
  9380=>"000000110",
  9381=>"111101111",
  9382=>"100110100",
  9383=>"001000000",
  9384=>"111111110",
  9385=>"000000111",
  9386=>"000000101",
  9387=>"111000000",
  9388=>"111110110",
  9389=>"000110110",
  9390=>"010000000",
  9391=>"000000001",
  9392=>"000111011",
  9393=>"111111101",
  9394=>"111111000",
  9395=>"000000000",
  9396=>"010111111",
  9397=>"111111111",
  9398=>"011111000",
  9399=>"111110000",
  9400=>"000000111",
  9401=>"100000000",
  9402=>"100001001",
  9403=>"000001000",
  9404=>"000000000",
  9405=>"111111111",
  9406=>"000000000",
  9407=>"011011111",
  9408=>"000000000",
  9409=>"000000000",
  9410=>"001001001",
  9411=>"001000000",
  9412=>"111111111",
  9413=>"000000000",
  9414=>"101101111",
  9415=>"100000000",
  9416=>"000110111",
  9417=>"111111111",
  9418=>"000000000",
  9419=>"000000111",
  9420=>"111111111",
  9421=>"000000111",
  9422=>"111111111",
  9423=>"111111111",
  9424=>"111101111",
  9425=>"100111111",
  9426=>"011000001",
  9427=>"111111111",
  9428=>"001000110",
  9429=>"111111111",
  9430=>"000000000",
  9431=>"000001111",
  9432=>"000110100",
  9433=>"000000000",
  9434=>"111110000",
  9435=>"111101100",
  9436=>"000000001",
  9437=>"000000000",
  9438=>"100000000",
  9439=>"000001001",
  9440=>"000000000",
  9441=>"000000000",
  9442=>"110011000",
  9443=>"111000000",
  9444=>"000001000",
  9445=>"100000100",
  9446=>"010000111",
  9447=>"000000000",
  9448=>"000000111",
  9449=>"111000111",
  9450=>"110000111",
  9451=>"111111111",
  9452=>"001001011",
  9453=>"000000000",
  9454=>"000000100",
  9455=>"111110000",
  9456=>"000000000",
  9457=>"000000000",
  9458=>"001111111",
  9459=>"111111011",
  9460=>"000010111",
  9461=>"110100000",
  9462=>"111110111",
  9463=>"111111111",
  9464=>"000000000",
  9465=>"111011000",
  9466=>"111111111",
  9467=>"000100000",
  9468=>"100111111",
  9469=>"000000000",
  9470=>"111110000",
  9471=>"000100111",
  9472=>"001001001",
  9473=>"011111111",
  9474=>"101000000",
  9475=>"111111111",
  9476=>"100011011",
  9477=>"111111111",
  9478=>"100100000",
  9479=>"111111111",
  9480=>"000000000",
  9481=>"000100100",
  9482=>"000000000",
  9483=>"111111111",
  9484=>"100100100",
  9485=>"000000000",
  9486=>"111111111",
  9487=>"000000000",
  9488=>"000000000",
  9489=>"111111011",
  9490=>"000000000",
  9491=>"000101001",
  9492=>"000000000",
  9493=>"011000000",
  9494=>"011111111",
  9495=>"000000000",
  9496=>"111111110",
  9497=>"000111011",
  9498=>"110100101",
  9499=>"000111111",
  9500=>"011001000",
  9501=>"011100000",
  9502=>"000000000",
  9503=>"011011111",
  9504=>"000000000",
  9505=>"000000000",
  9506=>"000011011",
  9507=>"111111111",
  9508=>"000000000",
  9509=>"000000000",
  9510=>"000000001",
  9511=>"000000000",
  9512=>"000000000",
  9513=>"001000011",
  9514=>"000000000",
  9515=>"000000000",
  9516=>"000000111",
  9517=>"000001000",
  9518=>"111100000",
  9519=>"000000000",
  9520=>"000111111",
  9521=>"111111000",
  9522=>"111111111",
  9523=>"111101001",
  9524=>"111101000",
  9525=>"000000000",
  9526=>"101001000",
  9527=>"001000000",
  9528=>"000000000",
  9529=>"111110111",
  9530=>"000000000",
  9531=>"111000100",
  9532=>"001000000",
  9533=>"001001111",
  9534=>"111111110",
  9535=>"000000000",
  9536=>"111111111",
  9537=>"111111111",
  9538=>"000000110",
  9539=>"100000000",
  9540=>"111111111",
  9541=>"000100101",
  9542=>"110000000",
  9543=>"000001111",
  9544=>"010000100",
  9545=>"000100000",
  9546=>"111111111",
  9547=>"110000100",
  9548=>"111111111",
  9549=>"111111111",
  9550=>"000000000",
  9551=>"110111111",
  9552=>"111001000",
  9553=>"100011010",
  9554=>"000011100",
  9555=>"000000000",
  9556=>"111111000",
  9557=>"001001011",
  9558=>"110000000",
  9559=>"101001001",
  9560=>"111111111",
  9561=>"000000000",
  9562=>"000000000",
  9563=>"000000000",
  9564=>"000000000",
  9565=>"000000001",
  9566=>"000000000",
  9567=>"001001001",
  9568=>"001000000",
  9569=>"111101001",
  9570=>"000111011",
  9571=>"011111111",
  9572=>"000000110",
  9573=>"001000001",
  9574=>"111000000",
  9575=>"111111111",
  9576=>"111110101",
  9577=>"110100000",
  9578=>"000000111",
  9579=>"100000000",
  9580=>"100000111",
  9581=>"101100000",
  9582=>"000010000",
  9583=>"111111110",
  9584=>"011111111",
  9585=>"000000011",
  9586=>"000000000",
  9587=>"111111111",
  9588=>"111111111",
  9589=>"000000000",
  9590=>"111111111",
  9591=>"110111000",
  9592=>"000000000",
  9593=>"000000000",
  9594=>"101000000",
  9595=>"001000000",
  9596=>"110000000",
  9597=>"110110000",
  9598=>"011111000",
  9599=>"000111111",
  9600=>"000000000",
  9601=>"111111111",
  9602=>"111111111",
  9603=>"000000000",
  9604=>"100111111",
  9605=>"000000000",
  9606=>"111011011",
  9607=>"000101001",
  9608=>"000000000",
  9609=>"111111000",
  9610=>"101111111",
  9611=>"000000000",
  9612=>"100000110",
  9613=>"000000000",
  9614=>"100110111",
  9615=>"000000000",
  9616=>"100000000",
  9617=>"000011111",
  9618=>"000000000",
  9619=>"110000000",
  9620=>"111111000",
  9621=>"000000111",
  9622=>"000010000",
  9623=>"000000000",
  9624=>"000000000",
  9625=>"010110100",
  9626=>"111111111",
  9627=>"000000100",
  9628=>"001000000",
  9629=>"111111110",
  9630=>"111110100",
  9631=>"111111111",
  9632=>"111111111",
  9633=>"011010000",
  9634=>"001001010",
  9635=>"000000000",
  9636=>"001001111",
  9637=>"001000000",
  9638=>"111001000",
  9639=>"000000000",
  9640=>"000000100",
  9641=>"111010000",
  9642=>"111111111",
  9643=>"011111111",
  9644=>"000000000",
  9645=>"100000000",
  9646=>"111110111",
  9647=>"100100110",
  9648=>"000000110",
  9649=>"100000000",
  9650=>"011000000",
  9651=>"101001111",
  9652=>"111111000",
  9653=>"111011111",
  9654=>"100110110",
  9655=>"111111111",
  9656=>"111111110",
  9657=>"011111111",
  9658=>"001000001",
  9659=>"111101111",
  9660=>"111101111",
  9661=>"111111111",
  9662=>"000000111",
  9663=>"000000000",
  9664=>"000000000",
  9665=>"111111111",
  9666=>"000000000",
  9667=>"000000000",
  9668=>"000000111",
  9669=>"111110100",
  9670=>"101001111",
  9671=>"000000000",
  9672=>"010000000",
  9673=>"000101110",
  9674=>"000000000",
  9675=>"000000011",
  9676=>"111110001",
  9677=>"111111100",
  9678=>"000000000",
  9679=>"111011011",
  9680=>"000000000",
  9681=>"100100100",
  9682=>"111111111",
  9683=>"111111111",
  9684=>"111111000",
  9685=>"000000100",
  9686=>"000000110",
  9687=>"001001001",
  9688=>"000101001",
  9689=>"000000000",
  9690=>"010111011",
  9691=>"000000000",
  9692=>"011000000",
  9693=>"001000000",
  9694=>"111111111",
  9695=>"011001000",
  9696=>"100101000",
  9697=>"001001000",
  9698=>"100101111",
  9699=>"000000000",
  9700=>"100110110",
  9701=>"000000001",
  9702=>"000000011",
  9703=>"111111011",
  9704=>"111111111",
  9705=>"111111000",
  9706=>"000000000",
  9707=>"111111111",
  9708=>"000000000",
  9709=>"000000000",
  9710=>"000000000",
  9711=>"111111111",
  9712=>"000000100",
  9713=>"000001111",
  9714=>"011000101",
  9715=>"000000000",
  9716=>"000000000",
  9717=>"111111111",
  9718=>"001111110",
  9719=>"000000000",
  9720=>"000000000",
  9721=>"101000000",
  9722=>"000000000",
  9723=>"000000000",
  9724=>"000000111",
  9725=>"000000000",
  9726=>"000000000",
  9727=>"001000000",
  9728=>"000000000",
  9729=>"011110010",
  9730=>"111101111",
  9731=>"111111111",
  9732=>"111111111",
  9733=>"001000000",
  9734=>"110110000",
  9735=>"111111111",
  9736=>"000000100",
  9737=>"000111011",
  9738=>"110000100",
  9739=>"110111111",
  9740=>"100110110",
  9741=>"000100000",
  9742=>"000000000",
  9743=>"111111101",
  9744=>"111110110",
  9745=>"000110100",
  9746=>"000000000",
  9747=>"010111111",
  9748=>"111111111",
  9749=>"011111001",
  9750=>"011000000",
  9751=>"011111111",
  9752=>"110100100",
  9753=>"000111111",
  9754=>"111111101",
  9755=>"000000000",
  9756=>"111111100",
  9757=>"111001000",
  9758=>"011011000",
  9759=>"110111110",
  9760=>"000000000",
  9761=>"000000000",
  9762=>"000000000",
  9763=>"001000010",
  9764=>"111111111",
  9765=>"000100000",
  9766=>"001011000",
  9767=>"111111111",
  9768=>"111111111",
  9769=>"111000000",
  9770=>"100100000",
  9771=>"111111111",
  9772=>"111100111",
  9773=>"000000000",
  9774=>"010110111",
  9775=>"000000000",
  9776=>"000000000",
  9777=>"011111111",
  9778=>"000000001",
  9779=>"111111111",
  9780=>"000111111",
  9781=>"011111001",
  9782=>"111111111",
  9783=>"000000100",
  9784=>"111011000",
  9785=>"011110110",
  9786=>"111111111",
  9787=>"110000000",
  9788=>"111000000",
  9789=>"000000110",
  9790=>"000000000",
  9791=>"111000000",
  9792=>"110100000",
  9793=>"110100111",
  9794=>"000001000",
  9795=>"001000110",
  9796=>"000001001",
  9797=>"000000110",
  9798=>"111110000",
  9799=>"000000000",
  9800=>"011011111",
  9801=>"110110111",
  9802=>"111000000",
  9803=>"111111111",
  9804=>"000000000",
  9805=>"000000000",
  9806=>"000010000",
  9807=>"001000100",
  9808=>"000000000",
  9809=>"011000000",
  9810=>"000000000",
  9811=>"001001001",
  9812=>"011111111",
  9813=>"000000000",
  9814=>"101000100",
  9815=>"111111111",
  9816=>"011001000",
  9817=>"101000001",
  9818=>"001000000",
  9819=>"001001001",
  9820=>"000000000",
  9821=>"111111111",
  9822=>"000011111",
  9823=>"100010111",
  9824=>"100111011",
  9825=>"000000001",
  9826=>"111111110",
  9827=>"101101101",
  9828=>"111100000",
  9829=>"111101111",
  9830=>"111111111",
  9831=>"000111110",
  9832=>"100000000",
  9833=>"110100100",
  9834=>"000000000",
  9835=>"000100110",
  9836=>"001000000",
  9837=>"111111111",
  9838=>"000000000",
  9839=>"110110110",
  9840=>"100100111",
  9841=>"000000000",
  9842=>"001000010",
  9843=>"111111111",
  9844=>"000000000",
  9845=>"010111110",
  9846=>"000010000",
  9847=>"000000000",
  9848=>"000000001",
  9849=>"100100000",
  9850=>"111111110",
  9851=>"000100100",
  9852=>"111001111",
  9853=>"000000111",
  9854=>"000000000",
  9855=>"000000000",
  9856=>"000000100",
  9857=>"111111111",
  9858=>"000111111",
  9859=>"111111111",
  9860=>"111111000",
  9861=>"100100111",
  9862=>"111111111",
  9863=>"110111100",
  9864=>"000001011",
  9865=>"111111111",
  9866=>"110111110",
  9867=>"111111111",
  9868=>"110101111",
  9869=>"111100100",
  9870=>"111000000",
  9871=>"000000100",
  9872=>"001000000",
  9873=>"011111111",
  9874=>"111111111",
  9875=>"111111111",
  9876=>"100101000",
  9877=>"011111111",
  9878=>"001000000",
  9879=>"111100000",
  9880=>"000000001",
  9881=>"111111111",
  9882=>"000000000",
  9883=>"000000000",
  9884=>"110111111",
  9885=>"010010010",
  9886=>"001100110",
  9887=>"111110010",
  9888=>"000001111",
  9889=>"001000000",
  9890=>"100001101",
  9891=>"110110110",
  9892=>"000000000",
  9893=>"111111100",
  9894=>"100000000",
  9895=>"000100000",
  9896=>"000100111",
  9897=>"000000000",
  9898=>"111111111",
  9899=>"011001000",
  9900=>"110111111",
  9901=>"000000001",
  9902=>"001001001",
  9903=>"111111111",
  9904=>"111111111",
  9905=>"110100100",
  9906=>"111111011",
  9907=>"000000000",
  9908=>"110110000",
  9909=>"111100111",
  9910=>"000000000",
  9911=>"011111111",
  9912=>"001111111",
  9913=>"111111001",
  9914=>"001011000",
  9915=>"001111111",
  9916=>"011111111",
  9917=>"001111111",
  9918=>"111111111",
  9919=>"111001001",
  9920=>"000000000",
  9921=>"000001001",
  9922=>"111111111",
  9923=>"000000111",
  9924=>"000001111",
  9925=>"000000100",
  9926=>"010010010",
  9927=>"000001101",
  9928=>"111111111",
  9929=>"111111111",
  9930=>"100101000",
  9931=>"011000000",
  9932=>"001000000",
  9933=>"000001001",
  9934=>"001111011",
  9935=>"000000100",
  9936=>"110111011",
  9937=>"110000000",
  9938=>"000100000",
  9939=>"010000000",
  9940=>"111000000",
  9941=>"110110110",
  9942=>"000000000",
  9943=>"100110100",
  9944=>"000000000",
  9945=>"011111000",
  9946=>"111001000",
  9947=>"011111111",
  9948=>"000000000",
  9949=>"000010000",
  9950=>"000111001",
  9951=>"000100100",
  9952=>"111111111",
  9953=>"000010010",
  9954=>"110110110",
  9955=>"001000000",
  9956=>"111111111",
  9957=>"011001100",
  9958=>"111111111",
  9959=>"000000000",
  9960=>"111111111",
  9961=>"000100110",
  9962=>"000000111",
  9963=>"001000000",
  9964=>"111111111",
  9965=>"000100000",
  9966=>"111111111",
  9967=>"000011001",
  9968=>"111111111",
  9969=>"110000111",
  9970=>"111111111",
  9971=>"011011011",
  9972=>"111000000",
  9973=>"000101100",
  9974=>"000100111",
  9975=>"001111001",
  9976=>"110111111",
  9977=>"000100111",
  9978=>"001100101",
  9979=>"111111111",
  9980=>"110111111",
  9981=>"111110110",
  9982=>"111110000",
  9983=>"001111000",
  9984=>"000000000",
  9985=>"100100100",
  9986=>"111111111",
  9987=>"000000000",
  9988=>"001101000",
  9989=>"000000000",
  9990=>"011000000",
  9991=>"111010100",
  9992=>"111111000",
  9993=>"000000100",
  9994=>"000000101",
  9995=>"110111011",
  9996=>"111111111",
  9997=>"111011000",
  9998=>"000001010",
  9999=>"100111111",
  10000=>"111111111",
  10001=>"001001101",
  10002=>"001001001",
  10003=>"000000001",
  10004=>"010110010",
  10005=>"111111111",
  10006=>"100100100",
  10007=>"111111111",
  10008=>"001000001",
  10009=>"111111111",
  10010=>"000000011",
  10011=>"110000100",
  10012=>"000110100",
  10013=>"100100010",
  10014=>"000000000",
  10015=>"111111111",
  10016=>"000100100",
  10017=>"111111111",
  10018=>"001000000",
  10019=>"111111011",
  10020=>"111111000",
  10021=>"111111111",
  10022=>"000000000",
  10023=>"000010111",
  10024=>"110100111",
  10025=>"000000000",
  10026=>"111111111",
  10027=>"111111111",
  10028=>"001000000",
  10029=>"000111111",
  10030=>"000000000",
  10031=>"111111011",
  10032=>"001001111",
  10033=>"111111100",
  10034=>"000000000",
  10035=>"111000000",
  10036=>"000111111",
  10037=>"000000000",
  10038=>"000101111",
  10039=>"000000000",
  10040=>"000000000",
  10041=>"111111000",
  10042=>"011011111",
  10043=>"111111000",
  10044=>"110000110",
  10045=>"101011011",
  10046=>"110110100",
  10047=>"000000000",
  10048=>"100110111",
  10049=>"001001011",
  10050=>"000000000",
  10051=>"111110110",
  10052=>"000000000",
  10053=>"000100100",
  10054=>"000000000",
  10055=>"111111110",
  10056=>"111111000",
  10057=>"000000000",
  10058=>"010111111",
  10059=>"110000100",
  10060=>"100000111",
  10061=>"000000011",
  10062=>"000000100",
  10063=>"010111111",
  10064=>"011000000",
  10065=>"110000000",
  10066=>"000001111",
  10067=>"001001000",
  10068=>"001000011",
  10069=>"011010000",
  10070=>"000001001",
  10071=>"111111111",
  10072=>"001111111",
  10073=>"111111111",
  10074=>"111111111",
  10075=>"111000000",
  10076=>"000000001",
  10077=>"000111111",
  10078=>"001011000",
  10079=>"001111111",
  10080=>"000010000",
  10081=>"000001111",
  10082=>"010110100",
  10083=>"000000000",
  10084=>"000000011",
  10085=>"011011011",
  10086=>"000110100",
  10087=>"110000001",
  10088=>"100001101",
  10089=>"000000000",
  10090=>"111111100",
  10091=>"110000010",
  10092=>"000000000",
  10093=>"000011000",
  10094=>"000000000",
  10095=>"111111111",
  10096=>"000100000",
  10097=>"000000000",
  10098=>"011000000",
  10099=>"111000000",
  10100=>"000010000",
  10101=>"011001001",
  10102=>"111111100",
  10103=>"111111111",
  10104=>"111111000",
  10105=>"000000000",
  10106=>"000001101",
  10107=>"000001111",
  10108=>"110111111",
  10109=>"111100000",
  10110=>"000100110",
  10111=>"000001000",
  10112=>"111111011",
  10113=>"001000000",
  10114=>"100001001",
  10115=>"110100000",
  10116=>"000000000",
  10117=>"010110111",
  10118=>"111000000",
  10119=>"111111000",
  10120=>"001111011",
  10121=>"111111111",
  10122=>"111100000",
  10123=>"000000000",
  10124=>"101101111",
  10125=>"111111110",
  10126=>"011011000",
  10127=>"000000000",
  10128=>"000100000",
  10129=>"111111111",
  10130=>"000000010",
  10131=>"001001000",
  10132=>"000000000",
  10133=>"000000111",
  10134=>"110111110",
  10135=>"011111111",
  10136=>"000011000",
  10137=>"000000000",
  10138=>"000000000",
  10139=>"111111111",
  10140=>"110111111",
  10141=>"111111010",
  10142=>"111111111",
  10143=>"011111000",
  10144=>"000000101",
  10145=>"000000110",
  10146=>"011111101",
  10147=>"000000000",
  10148=>"100001001",
  10149=>"011000011",
  10150=>"111001101",
  10151=>"000000000",
  10152=>"000000000",
  10153=>"111000000",
  10154=>"111111111",
  10155=>"000000111",
  10156=>"100000011",
  10157=>"000001101",
  10158=>"000000111",
  10159=>"011000111",
  10160=>"111111111",
  10161=>"000011111",
  10162=>"010111110",
  10163=>"111111111",
  10164=>"000000001",
  10165=>"011000000",
  10166=>"000000000",
  10167=>"111111111",
  10168=>"111000111",
  10169=>"111111001",
  10170=>"010000001",
  10171=>"010111111",
  10172=>"000000000",
  10173=>"001001000",
  10174=>"100000001",
  10175=>"100100000",
  10176=>"000000000",
  10177=>"000000000",
  10178=>"000000001",
  10179=>"111111000",
  10180=>"111001111",
  10181=>"001001101",
  10182=>"000000001",
  10183=>"101101111",
  10184=>"111000001",
  10185=>"110000000",
  10186=>"000000001",
  10187=>"000000110",
  10188=>"111011000",
  10189=>"000000011",
  10190=>"100100101",
  10191=>"001111110",
  10192=>"111111111",
  10193=>"111111111",
  10194=>"001001000",
  10195=>"101100100",
  10196=>"100000000",
  10197=>"111111000",
  10198=>"001001000",
  10199=>"001000000",
  10200=>"111111011",
  10201=>"001011111",
  10202=>"111111111",
  10203=>"000000000",
  10204=>"111111111",
  10205=>"000000000",
  10206=>"100111101",
  10207=>"000000000",
  10208=>"001001000",
  10209=>"111111111",
  10210=>"111111111",
  10211=>"011000000",
  10212=>"101111111",
  10213=>"111111000",
  10214=>"111111111",
  10215=>"000010110",
  10216=>"000000001",
  10217=>"111111111",
  10218=>"100001111",
  10219=>"111111111",
  10220=>"110111111",
  10221=>"001110111",
  10222=>"111111111",
  10223=>"111111111",
  10224=>"000111111",
  10225=>"000000000",
  10226=>"000000000",
  10227=>"111111111",
  10228=>"111111111",
  10229=>"000000000",
  10230=>"111111111",
  10231=>"010000000",
  10232=>"110110111",
  10233=>"111001001",
  10234=>"100011111",
  10235=>"000100101",
  10236=>"000010000",
  10237=>"000001101",
  10238=>"111110000",
  10239=>"110111111",
  10240=>"000100110",
  10241=>"111000000",
  10242=>"100101111",
  10243=>"000000000",
  10244=>"000000000",
  10245=>"000000000",
  10246=>"000000000",
  10247=>"111100111",
  10248=>"111111000",
  10249=>"110111111",
  10250=>"001000100",
  10251=>"100000000",
  10252=>"000000000",
  10253=>"000000001",
  10254=>"011111111",
  10255=>"000000100",
  10256=>"000001001",
  10257=>"110111000",
  10258=>"000110100",
  10259=>"111111111",
  10260=>"000000111",
  10261=>"000001000",
  10262=>"101111111",
  10263=>"100100100",
  10264=>"111111000",
  10265=>"111101001",
  10266=>"111110111",
  10267=>"011001001",
  10268=>"100111111",
  10269=>"010011111",
  10270=>"011011011",
  10271=>"111001000",
  10272=>"000000000",
  10273=>"111000000",
  10274=>"111111111",
  10275=>"000000000",
  10276=>"111111111",
  10277=>"111110111",
  10278=>"000000111",
  10279=>"111111111",
  10280=>"111000000",
  10281=>"000000010",
  10282=>"010111111",
  10283=>"011111110",
  10284=>"010011001",
  10285=>"010110000",
  10286=>"111111000",
  10287=>"111111111",
  10288=>"111111111",
  10289=>"000000010",
  10290=>"100100110",
  10291=>"111010000",
  10292=>"000100000",
  10293=>"000011011",
  10294=>"000000011",
  10295=>"000000001",
  10296=>"111111000",
  10297=>"111111001",
  10298=>"000000000",
  10299=>"000001111",
  10300=>"111000000",
  10301=>"001000111",
  10302=>"000001000",
  10303=>"111111111",
  10304=>"111111011",
  10305=>"000000111",
  10306=>"110111111",
  10307=>"000000001",
  10308=>"000001011",
  10309=>"000100110",
  10310=>"011101000",
  10311=>"111000000",
  10312=>"000011111",
  10313=>"000001000",
  10314=>"001000000",
  10315=>"010010111",
  10316=>"001001111",
  10317=>"111101111",
  10318=>"010000111",
  10319=>"111111111",
  10320=>"000000111",
  10321=>"110000100",
  10322=>"111000000",
  10323=>"101000000",
  10324=>"000000110",
  10325=>"111111110",
  10326=>"111000100",
  10327=>"111111111",
  10328=>"100000000",
  10329=>"000011111",
  10330=>"001001000",
  10331=>"000111111",
  10332=>"111011000",
  10333=>"000111111",
  10334=>"000000000",
  10335=>"000000111",
  10336=>"000000000",
  10337=>"110000000",
  10338=>"111111111",
  10339=>"000011111",
  10340=>"000000111",
  10341=>"010010111",
  10342=>"000000111",
  10343=>"000000000",
  10344=>"111010000",
  10345=>"010000111",
  10346=>"000000000",
  10347=>"000000110",
  10348=>"000111001",
  10349=>"000000000",
  10350=>"111000000",
  10351=>"111111011",
  10352=>"000000111",
  10353=>"011111111",
  10354=>"111111000",
  10355=>"000000000",
  10356=>"110100100",
  10357=>"111000000",
  10358=>"111111111",
  10359=>"000111111",
  10360=>"000000001",
  10361=>"001000001",
  10362=>"000000100",
  10363=>"111000100",
  10364=>"011011111",
  10365=>"000010111",
  10366=>"011000000",
  10367=>"101111111",
  10368=>"111111001",
  10369=>"000010000",
  10370=>"000010000",
  10371=>"001001011",
  10372=>"111111111",
  10373=>"111000111",
  10374=>"111111111",
  10375=>"111111010",
  10376=>"111111000",
  10377=>"111111111",
  10378=>"000000000",
  10379=>"100000000",
  10380=>"111110011",
  10381=>"100000000",
  10382=>"111111111",
  10383=>"110000000",
  10384=>"010010000",
  10385=>"010000000",
  10386=>"111000000",
  10387=>"101001000",
  10388=>"000011000",
  10389=>"100000000",
  10390=>"111011010",
  10391=>"000000000",
  10392=>"111111000",
  10393=>"111111111",
  10394=>"000000000",
  10395=>"000000000",
  10396=>"110000000",
  10397=>"000001101",
  10398=>"111111111",
  10399=>"111111010",
  10400=>"000100100",
  10401=>"111001001",
  10402=>"000000000",
  10403=>"111111101",
  10404=>"000000000",
  10405=>"111010100",
  10406=>"000111111",
  10407=>"001110100",
  10408=>"000000111",
  10409=>"000000110",
  10410=>"000000000",
  10411=>"111000000",
  10412=>"111001011",
  10413=>"110111001",
  10414=>"101000111",
  10415=>"111111000",
  10416=>"000000111",
  10417=>"111101111",
  10418=>"111111111",
  10419=>"011111010",
  10420=>"111100111",
  10421=>"111111101",
  10422=>"011000111",
  10423=>"101101001",
  10424=>"111100100",
  10425=>"111101000",
  10426=>"000000101",
  10427=>"100111011",
  10428=>"000000000",
  10429=>"111111001",
  10430=>"111000100",
  10431=>"010010001",
  10432=>"000111111",
  10433=>"110100010",
  10434=>"111111111",
  10435=>"000110111",
  10436=>"111111111",
  10437=>"100111011",
  10438=>"100000000",
  10439=>"010000111",
  10440=>"000000000",
  10441=>"001001001",
  10442=>"100000011",
  10443=>"000111111",
  10444=>"101100111",
  10445=>"101100000",
  10446=>"111000000",
  10447=>"000000000",
  10448=>"000000100",
  10449=>"111000000",
  10450=>"111111111",
  10451=>"000001000",
  10452=>"111000000",
  10453=>"011011000",
  10454=>"111100111",
  10455=>"111111001",
  10456=>"111111110",
  10457=>"000000011",
  10458=>"000000111",
  10459=>"000111110",
  10460=>"000000000",
  10461=>"000001001",
  10462=>"111111110",
  10463=>"111000000",
  10464=>"000000000",
  10465=>"000000011",
  10466=>"000001100",
  10467=>"000000000",
  10468=>"111100000",
  10469=>"000110110",
  10470=>"000000000",
  10471=>"111010100",
  10472=>"000000000",
  10473=>"011111111",
  10474=>"111111110",
  10475=>"111000000",
  10476=>"000000011",
  10477=>"000000111",
  10478=>"111011000",
  10479=>"001000010",
  10480=>"000000011",
  10481=>"000011111",
  10482=>"011101101",
  10483=>"000000111",
  10484=>"000011011",
  10485=>"001001001",
  10486=>"000100101",
  10487=>"000000000",
  10488=>"000000111",
  10489=>"111000000",
  10490=>"000000001",
  10491=>"000010000",
  10492=>"001000110",
  10493=>"111000111",
  10494=>"000000111",
  10495=>"011110110",
  10496=>"000000000",
  10497=>"000001001",
  10498=>"111111000",
  10499=>"011010000",
  10500=>"111000000",
  10501=>"000111111",
  10502=>"111101000",
  10503=>"000111111",
  10504=>"111111010",
  10505=>"100000111",
  10506=>"000000000",
  10507=>"010110111",
  10508=>"101011001",
  10509=>"000000000",
  10510=>"000000000",
  10511=>"110110111",
  10512=>"010110000",
  10513=>"111111000",
  10514=>"111100100",
  10515=>"000000000",
  10516=>"000101101",
  10517=>"100000000",
  10518=>"111001111",
  10519=>"000000110",
  10520=>"000000000",
  10521=>"000000111",
  10522=>"000111000",
  10523=>"111001000",
  10524=>"001100110",
  10525=>"100110111",
  10526=>"111000000",
  10527=>"111111000",
  10528=>"110010111",
  10529=>"001111111",
  10530=>"000000000",
  10531=>"111000000",
  10532=>"000111111",
  10533=>"000000000",
  10534=>"000000111",
  10535=>"000000111",
  10536=>"111000000",
  10537=>"000000111",
  10538=>"000110000",
  10539=>"000000111",
  10540=>"000111111",
  10541=>"001001000",
  10542=>"000000111",
  10543=>"011000000",
  10544=>"000011111",
  10545=>"011111111",
  10546=>"000001001",
  10547=>"000000000",
  10548=>"000000000",
  10549=>"000011111",
  10550=>"111010111",
  10551=>"111111000",
  10552=>"000000000",
  10553=>"111111111",
  10554=>"111000000",
  10555=>"000000000",
  10556=>"110100111",
  10557=>"111111000",
  10558=>"111111010",
  10559=>"000000000",
  10560=>"111111000",
  10561=>"110000000",
  10562=>"110111111",
  10563=>"000000000",
  10564=>"111111111",
  10565=>"110111111",
  10566=>"100000000",
  10567=>"000000111",
  10568=>"111111111",
  10569=>"101101111",
  10570=>"000000000",
  10571=>"000000001",
  10572=>"011000000",
  10573=>"111001000",
  10574=>"111100111",
  10575=>"100101101",
  10576=>"100111111",
  10577=>"001000000",
  10578=>"001000111",
  10579=>"111010000",
  10580=>"000000110",
  10581=>"001000000",
  10582=>"100000111",
  10583=>"100110111",
  10584=>"111100000",
  10585=>"000000010",
  10586=>"111000000",
  10587=>"000111100",
  10588=>"111011000",
  10589=>"111111111",
  10590=>"111000000",
  10591=>"000000001",
  10592=>"011011000",
  10593=>"111111000",
  10594=>"111111100",
  10595=>"111101001",
  10596=>"100000000",
  10597=>"000000000",
  10598=>"000000111",
  10599=>"111110000",
  10600=>"000100110",
  10601=>"110111000",
  10602=>"111111111",
  10603=>"111100000",
  10604=>"010111000",
  10605=>"000000000",
  10606=>"111111111",
  10607=>"111111000",
  10608=>"011110000",
  10609=>"100100000",
  10610=>"000100000",
  10611=>"100110100",
  10612=>"100000000",
  10613=>"111111111",
  10614=>"000000111",
  10615=>"000000100",
  10616=>"000111111",
  10617=>"000000101",
  10618=>"111001000",
  10619=>"000000110",
  10620=>"011000000",
  10621=>"000100000",
  10622=>"000111111",
  10623=>"111111111",
  10624=>"100110110",
  10625=>"000000011",
  10626=>"000011011",
  10627=>"000000000",
  10628=>"000011000",
  10629=>"000000111",
  10630=>"000000000",
  10631=>"000010111",
  10632=>"000000001",
  10633=>"111000000",
  10634=>"111000000",
  10635=>"001001011",
  10636=>"111111111",
  10637=>"011101101",
  10638=>"100000000",
  10639=>"010111111",
  10640=>"000000100",
  10641=>"000001111",
  10642=>"001011000",
  10643=>"111111111",
  10644=>"000001111",
  10645=>"000000000",
  10646=>"000000111",
  10647=>"000001111",
  10648=>"111111111",
  10649=>"111111000",
  10650=>"111111111",
  10651=>"100111011",
  10652=>"000000111",
  10653=>"000110000",
  10654=>"110100111",
  10655=>"000000111",
  10656=>"000000000",
  10657=>"110111001",
  10658=>"000000111",
  10659=>"111111111",
  10660=>"110110111",
  10661=>"000111111",
  10662=>"100000001",
  10663=>"110110010",
  10664=>"111110000",
  10665=>"000010000",
  10666=>"000000000",
  10667=>"111100111",
  10668=>"001111111",
  10669=>"000011111",
  10670=>"111111111",
  10671=>"011000111",
  10672=>"000000000",
  10673=>"000000010",
  10674=>"000000000",
  10675=>"111111010",
  10676=>"000111111",
  10677=>"000111111",
  10678=>"111001111",
  10679=>"110000110",
  10680=>"000000110",
  10681=>"011000001",
  10682=>"010111000",
  10683=>"111111100",
  10684=>"111010110",
  10685=>"111111001",
  10686=>"001011000",
  10687=>"110111000",
  10688=>"000111111",
  10689=>"111111111",
  10690=>"111100111",
  10691=>"111111000",
  10692=>"000000101",
  10693=>"111001100",
  10694=>"000011010",
  10695=>"000000011",
  10696=>"111111111",
  10697=>"000111111",
  10698=>"000000111",
  10699=>"000111111",
  10700=>"111000011",
  10701=>"111111000",
  10702=>"000111000",
  10703=>"000011111",
  10704=>"101111111",
  10705=>"011110100",
  10706=>"000000000",
  10707=>"111111000",
  10708=>"110111100",
  10709=>"110000000",
  10710=>"111111111",
  10711=>"001001000",
  10712=>"000100111",
  10713=>"010100000",
  10714=>"000000111",
  10715=>"111111111",
  10716=>"111100000",
  10717=>"111111111",
  10718=>"000000010",
  10719=>"001011011",
  10720=>"000000001",
  10721=>"111000000",
  10722=>"000011011",
  10723=>"111101000",
  10724=>"111111001",
  10725=>"000110100",
  10726=>"000000000",
  10727=>"111111111",
  10728=>"111011000",
  10729=>"111000000",
  10730=>"000001000",
  10731=>"111111111",
  10732=>"111111111",
  10733=>"001111110",
  10734=>"101000111",
  10735=>"111111010",
  10736=>"111010011",
  10737=>"000000000",
  10738=>"000000000",
  10739=>"000101000",
  10740=>"000000000",
  10741=>"110111111",
  10742=>"001000000",
  10743=>"011001000",
  10744=>"111010000",
  10745=>"011011000",
  10746=>"010000110",
  10747=>"001010000",
  10748=>"110101000",
  10749=>"000000000",
  10750=>"100110100",
  10751=>"000000000",
  10752=>"000000000",
  10753=>"001000000",
  10754=>"111000000",
  10755=>"011111111",
  10756=>"100000000",
  10757=>"111111111",
  10758=>"000011011",
  10759=>"111101111",
  10760=>"110000000",
  10761=>"111111111",
  10762=>"000000000",
  10763=>"111111110",
  10764=>"101111111",
  10765=>"000000000",
  10766=>"110111111",
  10767=>"000000000",
  10768=>"000001110",
  10769=>"111111011",
  10770=>"000000111",
  10771=>"111111111",
  10772=>"000000000",
  10773=>"011011111",
  10774=>"000000000",
  10775=>"000000110",
  10776=>"111111001",
  10777=>"111111011",
  10778=>"111001000",
  10779=>"011101101",
  10780=>"100110111",
  10781=>"001001001",
  10782=>"110001001",
  10783=>"000100110",
  10784=>"000000101",
  10785=>"110111111",
  10786=>"000000000",
  10787=>"000110111",
  10788=>"011011111",
  10789=>"111111111",
  10790=>"000000000",
  10791=>"111111111",
  10792=>"000000000",
  10793=>"000000111",
  10794=>"111111100",
  10795=>"101000000",
  10796=>"111111000",
  10797=>"001001011",
  10798=>"000000000",
  10799=>"111011011",
  10800=>"011110000",
  10801=>"111111111",
  10802=>"111101111",
  10803=>"111111111",
  10804=>"000000000",
  10805=>"110111111",
  10806=>"000000000",
  10807=>"000000000",
  10808=>"111111111",
  10809=>"111010000",
  10810=>"000000000",
  10811=>"000000000",
  10812=>"111111111",
  10813=>"000011011",
  10814=>"111011000",
  10815=>"000000000",
  10816=>"001000000",
  10817=>"111011111",
  10818=>"000100000",
  10819=>"000000000",
  10820=>"100000000",
  10821=>"101101111",
  10822=>"000000000",
  10823=>"110100100",
  10824=>"111111011",
  10825=>"000000011",
  10826=>"110010000",
  10827=>"100100100",
  10828=>"111111111",
  10829=>"001101111",
  10830=>"000111111",
  10831=>"111111111",
  10832=>"000010111",
  10833=>"000010111",
  10834=>"000000100",
  10835=>"001001001",
  10836=>"000000000",
  10837=>"110110110",
  10838=>"000111111",
  10839=>"000000000",
  10840=>"111111111",
  10841=>"111000000",
  10842=>"000000000",
  10843=>"001000000",
  10844=>"000000100",
  10845=>"000000010",
  10846=>"101111011",
  10847=>"000000000",
  10848=>"000000011",
  10849=>"000111111",
  10850=>"000000000",
  10851=>"000000111",
  10852=>"100110000",
  10853=>"111011111",
  10854=>"111000010",
  10855=>"111011000",
  10856=>"111111111",
  10857=>"111111111",
  10858=>"111111111",
  10859=>"000000000",
  10860=>"111001000",
  10861=>"100000100",
  10862=>"000000000",
  10863=>"000000000",
  10864=>"100100000",
  10865=>"110111000",
  10866=>"111111000",
  10867=>"001001000",
  10868=>"100000000",
  10869=>"000000000",
  10870=>"000000001",
  10871=>"000000000",
  10872=>"111111111",
  10873=>"111111111",
  10874=>"000000011",
  10875=>"000000000",
  10876=>"010111111",
  10877=>"011111111",
  10878=>"000101111",
  10879=>"111011000",
  10880=>"000000000",
  10881=>"111111001",
  10882=>"111011001",
  10883=>"111111111",
  10884=>"000000000",
  10885=>"000000001",
  10886=>"101000110",
  10887=>"000000000",
  10888=>"000000000",
  10889=>"111011011",
  10890=>"111111001",
  10891=>"111000000",
  10892=>"101001111",
  10893=>"110111111",
  10894=>"111111110",
  10895=>"000111111",
  10896=>"101111110",
  10897=>"111111111",
  10898=>"000000100",
  10899=>"111000000",
  10900=>"011000100",
  10901=>"000011111",
  10902=>"111001000",
  10903=>"010011111",
  10904=>"000000000",
  10905=>"000000100",
  10906=>"011011110",
  10907=>"001001111",
  10908=>"000000001",
  10909=>"001110100",
  10910=>"000100000",
  10911=>"000010111",
  10912=>"011011010",
  10913=>"000000000",
  10914=>"000000000",
  10915=>"010010010",
  10916=>"000100101",
  10917=>"000111001",
  10918=>"000111110",
  10919=>"111111111",
  10920=>"111111000",
  10921=>"000000000",
  10922=>"001000000",
  10923=>"000011110",
  10924=>"111111111",
  10925=>"000000000",
  10926=>"100110111",
  10927=>"000000000",
  10928=>"111100100",
  10929=>"110100100",
  10930=>"110111111",
  10931=>"111110000",
  10932=>"111111111",
  10933=>"001000000",
  10934=>"001111100",
  10935=>"011111111",
  10936=>"000010110",
  10937=>"111011000",
  10938=>"000000000",
  10939=>"111111111",
  10940=>"111111110",
  10941=>"111111000",
  10942=>"000000000",
  10943=>"011011010",
  10944=>"101100000",
  10945=>"000000000",
  10946=>"110010000",
  10947=>"111111111",
  10948=>"111111000",
  10949=>"000000000",
  10950=>"101111111",
  10951=>"011001100",
  10952=>"110000000",
  10953=>"111111111",
  10954=>"100000101",
  10955=>"000000000",
  10956=>"110100000",
  10957=>"100000000",
  10958=>"001011111",
  10959=>"111000000",
  10960=>"000111111",
  10961=>"111000000",
  10962=>"111011000",
  10963=>"111111001",
  10964=>"110111111",
  10965=>"000000000",
  10966=>"111111111",
  10967=>"111000000",
  10968=>"010110000",
  10969=>"000000000",
  10970=>"101000001",
  10971=>"000011101",
  10972=>"110111010",
  10973=>"101100000",
  10974=>"001001000",
  10975=>"111111111",
  10976=>"000000000",
  10977=>"010011111",
  10978=>"111111100",
  10979=>"111111111",
  10980=>"000000011",
  10981=>"000000000",
  10982=>"011000011",
  10983=>"111111111",
  10984=>"011001000",
  10985=>"100101100",
  10986=>"110111110",
  10987=>"111111111",
  10988=>"000000000",
  10989=>"111010000",
  10990=>"000000000",
  10991=>"000110110",
  10992=>"000000001",
  10993=>"110010011",
  10994=>"000001001",
  10995=>"111111010",
  10996=>"001000000",
  10997=>"000000100",
  10998=>"000000000",
  10999=>"111111110",
  11000=>"111111111",
  11001=>"111111111",
  11002=>"000000100",
  11003=>"000000000",
  11004=>"000010011",
  11005=>"001000110",
  11006=>"000000000",
  11007=>"000000000",
  11008=>"000000111",
  11009=>"101000100",
  11010=>"001000000",
  11011=>"000100000",
  11012=>"111111111",
  11013=>"000000000",
  11014=>"111111001",
  11015=>"001100101",
  11016=>"000000000",
  11017=>"100000000",
  11018=>"111111111",
  11019=>"000000000",
  11020=>"111110110",
  11021=>"111110101",
  11022=>"110100000",
  11023=>"000000000",
  11024=>"011111000",
  11025=>"100011000",
  11026=>"011000111",
  11027=>"000000000",
  11028=>"100110111",
  11029=>"000011110",
  11030=>"000000111",
  11031=>"000000011",
  11032=>"111111111",
  11033=>"001000000",
  11034=>"000111111",
  11035=>"000000011",
  11036=>"111111111",
  11037=>"110110110",
  11038=>"110111010",
  11039=>"110111111",
  11040=>"100000011",
  11041=>"111111000",
  11042=>"010000000",
  11043=>"111110111",
  11044=>"111011100",
  11045=>"000000000",
  11046=>"100100100",
  11047=>"100000001",
  11048=>"111111110",
  11049=>"110111000",
  11050=>"000000000",
  11051=>"111111011",
  11052=>"011111111",
  11053=>"000000000",
  11054=>"100000111",
  11055=>"010000000",
  11056=>"001001101",
  11057=>"010011001",
  11058=>"001000000",
  11059=>"111111011",
  11060=>"000000000",
  11061=>"000000111",
  11062=>"001000000",
  11063=>"000010010",
  11064=>"000110000",
  11065=>"101000000",
  11066=>"011111000",
  11067=>"000000000",
  11068=>"001100100",
  11069=>"110000110",
  11070=>"100000000",
  11071=>"000000001",
  11072=>"000000001",
  11073=>"111111111",
  11074=>"001001000",
  11075=>"000000000",
  11076=>"111100100",
  11077=>"011111111",
  11078=>"111111101",
  11079=>"000011011",
  11080=>"000111111",
  11081=>"000000000",
  11082=>"001001000",
  11083=>"100000100",
  11084=>"101011001",
  11085=>"011001001",
  11086=>"000000111",
  11087=>"010000000",
  11088=>"111111111",
  11089=>"000000000",
  11090=>"011010111",
  11091=>"111001000",
  11092=>"010111110",
  11093=>"001101111",
  11094=>"011011001",
  11095=>"001111111",
  11096=>"000000000",
  11097=>"000000100",
  11098=>"111111000",
  11099=>"111111110",
  11100=>"111000000",
  11101=>"111111110",
  11102=>"001000000",
  11103=>"001001110",
  11104=>"111100000",
  11105=>"000000000",
  11106=>"111100000",
  11107=>"001001100",
  11108=>"000000000",
  11109=>"101101101",
  11110=>"000000000",
  11111=>"000000000",
  11112=>"000000000",
  11113=>"111100000",
  11114=>"000000000",
  11115=>"111111111",
  11116=>"010011101",
  11117=>"000100000",
  11118=>"001001011",
  11119=>"001000000",
  11120=>"100101111",
  11121=>"000000011",
  11122=>"111110110",
  11123=>"000100000",
  11124=>"111111111",
  11125=>"111110111",
  11126=>"011000000",
  11127=>"000000111",
  11128=>"000000000",
  11129=>"011001000",
  11130=>"000101111",
  11131=>"010011000",
  11132=>"111111110",
  11133=>"001000000",
  11134=>"110111111",
  11135=>"000000000",
  11136=>"001001011",
  11137=>"000001100",
  11138=>"000011111",
  11139=>"000000011",
  11140=>"110000111",
  11141=>"000001111",
  11142=>"101001101",
  11143=>"011001000",
  11144=>"111111111",
  11145=>"111111111",
  11146=>"110010010",
  11147=>"111111000",
  11148=>"100000001",
  11149=>"010110111",
  11150=>"101111111",
  11151=>"111010000",
  11152=>"000111111",
  11153=>"000000000",
  11154=>"111100100",
  11155=>"100000000",
  11156=>"111111111",
  11157=>"000000000",
  11158=>"000000011",
  11159=>"001001001",
  11160=>"110000011",
  11161=>"111111101",
  11162=>"010000111",
  11163=>"111111111",
  11164=>"010010000",
  11165=>"000000000",
  11166=>"000000000",
  11167=>"000000000",
  11168=>"110001001",
  11169=>"111111011",
  11170=>"100100000",
  11171=>"000000000",
  11172=>"000100000",
  11173=>"111111111",
  11174=>"101100111",
  11175=>"111111111",
  11176=>"011011011",
  11177=>"011011001",
  11178=>"000001011",
  11179=>"000100000",
  11180=>"111111111",
  11181=>"000000000",
  11182=>"011000000",
  11183=>"111111111",
  11184=>"000000001",
  11185=>"011111000",
  11186=>"111011011",
  11187=>"000000000",
  11188=>"111111011",
  11189=>"001000000",
  11190=>"111100111",
  11191=>"011000000",
  11192=>"000000000",
  11193=>"111111111",
  11194=>"011000000",
  11195=>"100100000",
  11196=>"111111011",
  11197=>"101110110",
  11198=>"010111110",
  11199=>"110110110",
  11200=>"111000011",
  11201=>"000100000",
  11202=>"110000010",
  11203=>"110100110",
  11204=>"011011000",
  11205=>"110000000",
  11206=>"011000000",
  11207=>"111000000",
  11208=>"000000000",
  11209=>"111111111",
  11210=>"100000000",
  11211=>"000000011",
  11212=>"110010000",
  11213=>"111111111",
  11214=>"000000000",
  11215=>"111001011",
  11216=>"010111111",
  11217=>"111111111",
  11218=>"111011011",
  11219=>"111111000",
  11220=>"111111001",
  11221=>"001011111",
  11222=>"000011111",
  11223=>"000001000",
  11224=>"000100100",
  11225=>"011111111",
  11226=>"111110000",
  11227=>"101111111",
  11228=>"000000000",
  11229=>"000000000",
  11230=>"111111111",
  11231=>"000000111",
  11232=>"001010000",
  11233=>"011001000",
  11234=>"000000000",
  11235=>"000000000",
  11236=>"101111000",
  11237=>"111000000",
  11238=>"011111000",
  11239=>"000000000",
  11240=>"111010000",
  11241=>"111111011",
  11242=>"101000000",
  11243=>"111111100",
  11244=>"000000000",
  11245=>"100100100",
  11246=>"111111100",
  11247=>"100000000",
  11248=>"110111110",
  11249=>"111111111",
  11250=>"100110111",
  11251=>"111000000",
  11252=>"000010011",
  11253=>"111011111",
  11254=>"111011000",
  11255=>"111110100",
  11256=>"111111111",
  11257=>"100000000",
  11258=>"000000000",
  11259=>"000100111",
  11260=>"000010111",
  11261=>"011110000",
  11262=>"000000111",
  11263=>"111000000",
  11264=>"000000000",
  11265=>"000000000",
  11266=>"001101011",
  11267=>"111100100",
  11268=>"010110111",
  11269=>"001001001",
  11270=>"000000000",
  11271=>"111101101",
  11272=>"110000000",
  11273=>"111110111",
  11274=>"001000000",
  11275=>"110010011",
  11276=>"110111111",
  11277=>"000000000",
  11278=>"000100101",
  11279=>"111111111",
  11280=>"111111111",
  11281=>"000111111",
  11282=>"000001101",
  11283=>"110111111",
  11284=>"000000110",
  11285=>"111111111",
  11286=>"101000111",
  11287=>"110110111",
  11288=>"000001101",
  11289=>"110110110",
  11290=>"000000000",
  11291=>"111100100",
  11292=>"111111111",
  11293=>"111111111",
  11294=>"111100100",
  11295=>"111000111",
  11296=>"101100111",
  11297=>"000000000",
  11298=>"111011111",
  11299=>"111111101",
  11300=>"000111111",
  11301=>"000000000",
  11302=>"101000100",
  11303=>"111000000",
  11304=>"000000110",
  11305=>"011111111",
  11306=>"111111111",
  11307=>"111111111",
  11308=>"000001000",
  11309=>"111111111",
  11310=>"111101111",
  11311=>"011101111",
  11312=>"111011111",
  11313=>"000000000",
  11314=>"111100000",
  11315=>"000000100",
  11316=>"101101000",
  11317=>"001001000",
  11318=>"000100101",
  11319=>"001000000",
  11320=>"000000000",
  11321=>"001001111",
  11322=>"110111111",
  11323=>"111111100",
  11324=>"001000000",
  11325=>"001100000",
  11326=>"000000000",
  11327=>"100111111",
  11328=>"101001000",
  11329=>"010000111",
  11330=>"011011001",
  11331=>"000000000",
  11332=>"000000000",
  11333=>"111111110",
  11334=>"000000000",
  11335=>"000000000",
  11336=>"010110110",
  11337=>"111111111",
  11338=>"100000000",
  11339=>"111010111",
  11340=>"000000001",
  11341=>"100000000",
  11342=>"011001000",
  11343=>"100000001",
  11344=>"111011011",
  11345=>"111010110",
  11346=>"100111110",
  11347=>"000000110",
  11348=>"000111111",
  11349=>"010011000",
  11350=>"000000000",
  11351=>"111111111",
  11352=>"011011001",
  11353=>"000000000",
  11354=>"010110110",
  11355=>"100100000",
  11356=>"000000010",
  11357=>"111111111",
  11358=>"100000111",
  11359=>"011100100",
  11360=>"000000000",
  11361=>"111001000",
  11362=>"000000000",
  11363=>"101000000",
  11364=>"110110000",
  11365=>"111110000",
  11366=>"111111111",
  11367=>"000000000",
  11368=>"010000000",
  11369=>"000111111",
  11370=>"000000000",
  11371=>"100000000",
  11372=>"000000000",
  11373=>"000000101",
  11374=>"000000000",
  11375=>"100100100",
  11376=>"000000100",
  11377=>"000010000",
  11378=>"111111111",
  11379=>"111001111",
  11380=>"111111101",
  11381=>"001111111",
  11382=>"000000001",
  11383=>"000000100",
  11384=>"000000000",
  11385=>"100000000",
  11386=>"101100110",
  11387=>"111100111",
  11388=>"100110110",
  11389=>"001000000",
  11390=>"100100100",
  11391=>"111111111",
  11392=>"000000000",
  11393=>"011011111",
  11394=>"000000001",
  11395=>"000101111",
  11396=>"000000011",
  11397=>"000000000",
  11398=>"001000110",
  11399=>"000001111",
  11400=>"111111111",
  11401=>"000000000",
  11402=>"111000010",
  11403=>"111111111",
  11404=>"001000000",
  11405=>"100000000",
  11406=>"001000110",
  11407=>"111111111",
  11408=>"101001001",
  11409=>"000000000",
  11410=>"000110100",
  11411=>"111000000",
  11412=>"000000010",
  11413=>"000100111",
  11414=>"111111111",
  11415=>"111000100",
  11416=>"000000000",
  11417=>"111111110",
  11418=>"111111111",
  11419=>"010010110",
  11420=>"000000000",
  11421=>"100110111",
  11422=>"111111011",
  11423=>"000000000",
  11424=>"000000000",
  11425=>"101000110",
  11426=>"111111111",
  11427=>"000000111",
  11428=>"001001111",
  11429=>"000000111",
  11430=>"111100000",
  11431=>"111110111",
  11432=>"101000000",
  11433=>"000000000",
  11434=>"011111001",
  11435=>"100100100",
  11436=>"001111111",
  11437=>"110110000",
  11438=>"111111111",
  11439=>"000100110",
  11440=>"000000000",
  11441=>"001000000",
  11442=>"111111111",
  11443=>"111000000",
  11444=>"000001000",
  11445=>"100000000",
  11446=>"111111111",
  11447=>"000000000",
  11448=>"001001001",
  11449=>"000000000",
  11450=>"101100101",
  11451=>"111000000",
  11452=>"000000000",
  11453=>"000000000",
  11454=>"000100100",
  11455=>"010000000",
  11456=>"000000000",
  11457=>"000000000",
  11458=>"000000000",
  11459=>"111111111",
  11460=>"000110111",
  11461=>"000000000",
  11462=>"111111111",
  11463=>"000000000",
  11464=>"000000000",
  11465=>"101001101",
  11466=>"111111111",
  11467=>"000000000",
  11468=>"100110100",
  11469=>"000000101",
  11470=>"000010100",
  11471=>"000000110",
  11472=>"000000000",
  11473=>"101111111",
  11474=>"000000000",
  11475=>"011011010",
  11476=>"100110110",
  11477=>"111111111",
  11478=>"111110111",
  11479=>"001000110",
  11480=>"010010110",
  11481=>"000000000",
  11482=>"111111011",
  11483=>"010000111",
  11484=>"000000000",
  11485=>"111111111",
  11486=>"000000100",
  11487=>"011011000",
  11488=>"011000100",
  11489=>"000000000",
  11490=>"000000110",
  11491=>"111111100",
  11492=>"111011001",
  11493=>"001001110",
  11494=>"111111111",
  11495=>"111001011",
  11496=>"111111111",
  11497=>"010010100",
  11498=>"001001000",
  11499=>"000000110",
  11500=>"100100100",
  11501=>"100110111",
  11502=>"111001111",
  11503=>"100000000",
  11504=>"111010000",
  11505=>"001001000",
  11506=>"001111111",
  11507=>"001000000",
  11508=>"111111111",
  11509=>"101110010",
  11510=>"001001001",
  11511=>"000000000",
  11512=>"000011111",
  11513=>"111111111",
  11514=>"000000000",
  11515=>"111111111",
  11516=>"111111111",
  11517=>"101000000",
  11518=>"110101100",
  11519=>"010111111",
  11520=>"101101001",
  11521=>"111100100",
  11522=>"001111111",
  11523=>"000111111",
  11524=>"111111111",
  11525=>"000111111",
  11526=>"101001100",
  11527=>"110011010",
  11528=>"111111111",
  11529=>"111000000",
  11530=>"000000000",
  11531=>"011010000",
  11532=>"001000000",
  11533=>"110000000",
  11534=>"000000000",
  11535=>"111111111",
  11536=>"011000000",
  11537=>"000000101",
  11538=>"110111111",
  11539=>"000000001",
  11540=>"111111000",
  11541=>"000000000",
  11542=>"100100001",
  11543=>"000000000",
  11544=>"111111111",
  11545=>"000000000",
  11546=>"000000000",
  11547=>"000011011",
  11548=>"111111111",
  11549=>"100110110",
  11550=>"000000000",
  11551=>"001001111",
  11552=>"000001000",
  11553=>"000000111",
  11554=>"011001000",
  11555=>"000000001",
  11556=>"000000110",
  11557=>"111011111",
  11558=>"111111111",
  11559=>"000000000",
  11560=>"111111110",
  11561=>"000000000",
  11562=>"111111011",
  11563=>"001111011",
  11564=>"000101111",
  11565=>"111011111",
  11566=>"000000000",
  11567=>"000000000",
  11568=>"001111111",
  11569=>"100111110",
  11570=>"111000000",
  11571=>"111010111",
  11572=>"000000011",
  11573=>"000000000",
  11574=>"011011111",
  11575=>"000000000",
  11576=>"010111000",
  11577=>"000000000",
  11578=>"000000000",
  11579=>"111111111",
  11580=>"000000100",
  11581=>"000000110",
  11582=>"011111111",
  11583=>"111011011",
  11584=>"000001001",
  11585=>"101001111",
  11586=>"111111111",
  11587=>"010100110",
  11588=>"001001000",
  11589=>"111011011",
  11590=>"010111111",
  11591=>"101001000",
  11592=>"100000000",
  11593=>"000000000",
  11594=>"111111111",
  11595=>"110000000",
  11596=>"000000000",
  11597=>"111110000",
  11598=>"101000000",
  11599=>"011001011",
  11600=>"000100111",
  11601=>"000000000",
  11602=>"110010011",
  11603=>"000000111",
  11604=>"111111111",
  11605=>"011011011",
  11606=>"000000000",
  11607=>"111111000",
  11608=>"111011011",
  11609=>"000100111",
  11610=>"000000000",
  11611=>"111101111",
  11612=>"110111111",
  11613=>"111111111",
  11614=>"110000000",
  11615=>"000000110",
  11616=>"000000000",
  11617=>"110111111",
  11618=>"101000000",
  11619=>"111111111",
  11620=>"000111111",
  11621=>"000000000",
  11622=>"111111011",
  11623=>"100000000",
  11624=>"011000000",
  11625=>"000111111",
  11626=>"010111111",
  11627=>"111101111",
  11628=>"000010111",
  11629=>"101100100",
  11630=>"010000000",
  11631=>"000000001",
  11632=>"000000001",
  11633=>"000000000",
  11634=>"001111100",
  11635=>"000000000",
  11636=>"111111111",
  11637=>"001000000",
  11638=>"110111111",
  11639=>"111111111",
  11640=>"011010000",
  11641=>"000000000",
  11642=>"000000000",
  11643=>"111111111",
  11644=>"000000111",
  11645=>"100000000",
  11646=>"111110110",
  11647=>"000000100",
  11648=>"000011111",
  11649=>"111111111",
  11650=>"100111011",
  11651=>"000000000",
  11652=>"000000111",
  11653=>"000000111",
  11654=>"100000000",
  11655=>"000000000",
  11656=>"111111111",
  11657=>"100100111",
  11658=>"111011111",
  11659=>"010011011",
  11660=>"000000110",
  11661=>"111111111",
  11662=>"110110111",
  11663=>"000000000",
  11664=>"000000000",
  11665=>"000000000",
  11666=>"111111111",
  11667=>"100000000",
  11668=>"111111000",
  11669=>"000000000",
  11670=>"011001000",
  11671=>"000000000",
  11672=>"111111111",
  11673=>"000000000",
  11674=>"000000000",
  11675=>"111111111",
  11676=>"001000000",
  11677=>"000101000",
  11678=>"100101111",
  11679=>"000000000",
  11680=>"111100000",
  11681=>"110000000",
  11682=>"110110110",
  11683=>"110100000",
  11684=>"011111111",
  11685=>"000000001",
  11686=>"100100000",
  11687=>"111111111",
  11688=>"000000001",
  11689=>"000000000",
  11690=>"011000000",
  11691=>"001001101",
  11692=>"000000000",
  11693=>"100100100",
  11694=>"110100111",
  11695=>"100111111",
  11696=>"111111111",
  11697=>"000000000",
  11698=>"100010000",
  11699=>"000110110",
  11700=>"001000000",
  11701=>"111011001",
  11702=>"111001000",
  11703=>"100100110",
  11704=>"000000101",
  11705=>"001000000",
  11706=>"000000000",
  11707=>"011001100",
  11708=>"000110110",
  11709=>"110111111",
  11710=>"000000000",
  11711=>"001000000",
  11712=>"111101100",
  11713=>"100000111",
  11714=>"111111111",
  11715=>"000000000",
  11716=>"110110110",
  11717=>"101110111",
  11718=>"010000000",
  11719=>"001000000",
  11720=>"111111000",
  11721=>"111111011",
  11722=>"100000000",
  11723=>"111111111",
  11724=>"000000000",
  11725=>"100000000",
  11726=>"000011110",
  11727=>"111111111",
  11728=>"000000000",
  11729=>"100100110",
  11730=>"000000000",
  11731=>"000000000",
  11732=>"000000000",
  11733=>"111111111",
  11734=>"111000101",
  11735=>"011001011",
  11736=>"111111111",
  11737=>"000000110",
  11738=>"000000000",
  11739=>"111001101",
  11740=>"000000000",
  11741=>"111111110",
  11742=>"111110111",
  11743=>"100001101",
  11744=>"110111000",
  11745=>"010000000",
  11746=>"110111110",
  11747=>"000000000",
  11748=>"111000000",
  11749=>"111111111",
  11750=>"111000111",
  11751=>"010111111",
  11752=>"000000000",
  11753=>"101111110",
  11754=>"100000000",
  11755=>"100111111",
  11756=>"111111111",
  11757=>"101100110",
  11758=>"111001000",
  11759=>"000000100",
  11760=>"000000000",
  11761=>"000000000",
  11762=>"111111111",
  11763=>"000000000",
  11764=>"000000000",
  11765=>"000000000",
  11766=>"111111111",
  11767=>"110000111",
  11768=>"000000000",
  11769=>"001001011",
  11770=>"001111111",
  11771=>"000111101",
  11772=>"111011111",
  11773=>"110000000",
  11774=>"100110111",
  11775=>"000000000",
  11776=>"111111111",
  11777=>"000110000",
  11778=>"000000000",
  11779=>"000000000",
  11780=>"011111111",
  11781=>"000000000",
  11782=>"000100100",
  11783=>"000000000",
  11784=>"000000000",
  11785=>"100000000",
  11786=>"000000110",
  11787=>"111111111",
  11788=>"000110111",
  11789=>"000000000",
  11790=>"000101100",
  11791=>"111111111",
  11792=>"100011111",
  11793=>"111111001",
  11794=>"000101111",
  11795=>"001000100",
  11796=>"111011011",
  11797=>"111111110",
  11798=>"110110101",
  11799=>"110110100",
  11800=>"111111111",
  11801=>"101001101",
  11802=>"000000000",
  11803=>"000000000",
  11804=>"000000000",
  11805=>"001000000",
  11806=>"011111001",
  11807=>"000000000",
  11808=>"111000000",
  11809=>"110110111",
  11810=>"100100001",
  11811=>"111111111",
  11812=>"000000000",
  11813=>"000000000",
  11814=>"111111001",
  11815=>"111110000",
  11816=>"111111111",
  11817=>"000000000",
  11818=>"111111000",
  11819=>"000110110",
  11820=>"000011000",
  11821=>"000000001",
  11822=>"000000001",
  11823=>"111000010",
  11824=>"110100000",
  11825=>"111111111",
  11826=>"100110111",
  11827=>"000000011",
  11828=>"010010110",
  11829=>"101011111",
  11830=>"000000000",
  11831=>"110010000",
  11832=>"001101111",
  11833=>"010111111",
  11834=>"000000000",
  11835=>"000000110",
  11836=>"000000111",
  11837=>"000101101",
  11838=>"100001001",
  11839=>"000000000",
  11840=>"000000000",
  11841=>"011011111",
  11842=>"011001001",
  11843=>"110110111",
  11844=>"111111111",
  11845=>"111110111",
  11846=>"000110111",
  11847=>"011001000",
  11848=>"011001011",
  11849=>"000000000",
  11850=>"111111011",
  11851=>"000000110",
  11852=>"111001011",
  11853=>"000000000",
  11854=>"111111001",
  11855=>"000110111",
  11856=>"111111111",
  11857=>"010111111",
  11858=>"000000000",
  11859=>"111111111",
  11860=>"000000000",
  11861=>"000111111",
  11862=>"111111111",
  11863=>"000000000",
  11864=>"111111100",
  11865=>"101000101",
  11866=>"100100100",
  11867=>"111111011",
  11868=>"111111111",
  11869=>"110111110",
  11870=>"100000000",
  11871=>"100110110",
  11872=>"010111111",
  11873=>"000100000",
  11874=>"000000000",
  11875=>"111111100",
  11876=>"001011111",
  11877=>"110111111",
  11878=>"101000011",
  11879=>"000000000",
  11880=>"010110010",
  11881=>"111111111",
  11882=>"000000100",
  11883=>"111111110",
  11884=>"111111000",
  11885=>"111111110",
  11886=>"010010111",
  11887=>"111100000",
  11888=>"100000000",
  11889=>"100101111",
  11890=>"000000000",
  11891=>"000111111",
  11892=>"000000000",
  11893=>"001001011",
  11894=>"000000000",
  11895=>"001111110",
  11896=>"000000000",
  11897=>"111111111",
  11898=>"000000000",
  11899=>"111111110",
  11900=>"101111011",
  11901=>"001000000",
  11902=>"011000000",
  11903=>"111000011",
  11904=>"000100111",
  11905=>"110000010",
  11906=>"111000000",
  11907=>"111111111",
  11908=>"000000000",
  11909=>"101110110",
  11910=>"001001011",
  11911=>"110010111",
  11912=>"000100000",
  11913=>"000000001",
  11914=>"111111011",
  11915=>"011010000",
  11916=>"110111111",
  11917=>"110110011",
  11918=>"000110100",
  11919=>"111111011",
  11920=>"111111111",
  11921=>"111101001",
  11922=>"111001000",
  11923=>"000010110",
  11924=>"000100000",
  11925=>"111111111",
  11926=>"000111111",
  11927=>"000000111",
  11928=>"100100000",
  11929=>"111011101",
  11930=>"111010111",
  11931=>"111100101",
  11932=>"111111111",
  11933=>"001001001",
  11934=>"100100000",
  11935=>"000110110",
  11936=>"100100111",
  11937=>"111111111",
  11938=>"011111111",
  11939=>"111010000",
  11940=>"000000111",
  11941=>"110100010",
  11942=>"111110000",
  11943=>"001011110",
  11944=>"111111111",
  11945=>"111111111",
  11946=>"000000000",
  11947=>"011000000",
  11948=>"000000001",
  11949=>"001001001",
  11950=>"111111000",
  11951=>"000100000",
  11952=>"000111111",
  11953=>"110100110",
  11954=>"110111100",
  11955=>"000000000",
  11956=>"101001000",
  11957=>"111111000",
  11958=>"110010010",
  11959=>"111111111",
  11960=>"000000000",
  11961=>"111111100",
  11962=>"111101111",
  11963=>"110110110",
  11964=>"010011011",
  11965=>"000000000",
  11966=>"000000000",
  11967=>"111111111",
  11968=>"000000000",
  11969=>"000000000",
  11970=>"111011001",
  11971=>"000000000",
  11972=>"111111111",
  11973=>"111110110",
  11974=>"000001001",
  11975=>"000000000",
  11976=>"000111111",
  11977=>"001111000",
  11978=>"111111111",
  11979=>"100110100",
  11980=>"000110111",
  11981=>"111110111",
  11982=>"111111111",
  11983=>"010111111",
  11984=>"011011000",
  11985=>"111101101",
  11986=>"100000000",
  11987=>"111111111",
  11988=>"010110111",
  11989=>"111101000",
  11990=>"000000001",
  11991=>"111011000",
  11992=>"011111100",
  11993=>"001111110",
  11994=>"010111111",
  11995=>"000000001",
  11996=>"001001001",
  11997=>"011000000",
  11998=>"000111111",
  11999=>"111111011",
  12000=>"000000011",
  12001=>"001001101",
  12002=>"000000011",
  12003=>"101000000",
  12004=>"000000000",
  12005=>"110111111",
  12006=>"000111111",
  12007=>"000100100",
  12008=>"000000000",
  12009=>"111111110",
  12010=>"100100001",
  12011=>"000010111",
  12012=>"000110111",
  12013=>"111000000",
  12014=>"111111111",
  12015=>"110000111",
  12016=>"000000000",
  12017=>"111110111",
  12018=>"000000000",
  12019=>"111111001",
  12020=>"000000000",
  12021=>"000001001",
  12022=>"000011000",
  12023=>"000111000",
  12024=>"000010011",
  12025=>"111111111",
  12026=>"001111111",
  12027=>"000010000",
  12028=>"000000001",
  12029=>"000011011",
  12030=>"111111111",
  12031=>"000100000",
  12032=>"000000110",
  12033=>"000111111",
  12034=>"000000000",
  12035=>"010000000",
  12036=>"000000101",
  12037=>"000001000",
  12038=>"101001100",
  12039=>"000110111",
  12040=>"000000000",
  12041=>"011111111",
  12042=>"010000110",
  12043=>"011111011",
  12044=>"000001001",
  12045=>"001011110",
  12046=>"011111111",
  12047=>"000011111",
  12048=>"000000010",
  12049=>"001011011",
  12050=>"000110010",
  12051=>"001001000",
  12052=>"000000000",
  12053=>"000000110",
  12054=>"011001011",
  12055=>"000000000",
  12056=>"011000000",
  12057=>"000000100",
  12058=>"111110111",
  12059=>"111011111",
  12060=>"010000110",
  12061=>"101000000",
  12062=>"000000000",
  12063=>"111111111",
  12064=>"110111011",
  12065=>"001111111",
  12066=>"110110000",
  12067=>"111111000",
  12068=>"100101101",
  12069=>"000110111",
  12070=>"011011011",
  12071=>"000000001",
  12072=>"100111001",
  12073=>"110111110",
  12074=>"100100001",
  12075=>"111010001",
  12076=>"000000000",
  12077=>"000000000",
  12078=>"100111000",
  12079=>"000111111",
  12080=>"101001011",
  12081=>"000000111",
  12082=>"011000000",
  12083=>"110010111",
  12084=>"000000000",
  12085=>"001000111",
  12086=>"010010111",
  12087=>"111011111",
  12088=>"000000000",
  12089=>"000000000",
  12090=>"111000000",
  12091=>"001001001",
  12092=>"111111111",
  12093=>"000111111",
  12094=>"000001011",
  12095=>"000000000",
  12096=>"111111111",
  12097=>"111000000",
  12098=>"000100001",
  12099=>"111111111",
  12100=>"111110111",
  12101=>"000111111",
  12102=>"110111111",
  12103=>"001001011",
  12104=>"111111111",
  12105=>"111111000",
  12106=>"111111111",
  12107=>"000111010",
  12108=>"111111111",
  12109=>"000000010",
  12110=>"000100100",
  12111=>"010111111",
  12112=>"100100100",
  12113=>"000000000",
  12114=>"110000010",
  12115=>"111111111",
  12116=>"000000110",
  12117=>"100100000",
  12118=>"000010011",
  12119=>"000000111",
  12120=>"010000000",
  12121=>"100000000",
  12122=>"111101111",
  12123=>"000000000",
  12124=>"111111111",
  12125=>"111111111",
  12126=>"111001001",
  12127=>"111011011",
  12128=>"111111101",
  12129=>"111011000",
  12130=>"100110010",
  12131=>"100101111",
  12132=>"000000000",
  12133=>"111111011",
  12134=>"111111111",
  12135=>"001111011",
  12136=>"101101101",
  12137=>"110110111",
  12138=>"001111111",
  12139=>"000000000",
  12140=>"000001000",
  12141=>"110101111",
  12142=>"100110111",
  12143=>"111111111",
  12144=>"111011000",
  12145=>"111111111",
  12146=>"010000000",
  12147=>"111111110",
  12148=>"000000001",
  12149=>"000000000",
  12150=>"100000000",
  12151=>"110010000",
  12152=>"100110111",
  12153=>"111111111",
  12154=>"111111111",
  12155=>"001000000",
  12156=>"000000000",
  12157=>"111110110",
  12158=>"110110111",
  12159=>"010000101",
  12160=>"100100110",
  12161=>"111111001",
  12162=>"111010000",
  12163=>"001001000",
  12164=>"000000000",
  12165=>"101101111",
  12166=>"000000010",
  12167=>"000000000",
  12168=>"000000111",
  12169=>"011100100",
  12170=>"110110000",
  12171=>"000000001",
  12172=>"111111111",
  12173=>"010011011",
  12174=>"100000000",
  12175=>"000000000",
  12176=>"000000000",
  12177=>"110111101",
  12178=>"101111111",
  12179=>"111011111",
  12180=>"000000000",
  12181=>"000000111",
  12182=>"000110110",
  12183=>"101001111",
  12184=>"000000000",
  12185=>"111010001",
  12186=>"000110000",
  12187=>"000000000",
  12188=>"111100000",
  12189=>"111111111",
  12190=>"111011011",
  12191=>"000000111",
  12192=>"100000000",
  12193=>"111110100",
  12194=>"100111111",
  12195=>"111111111",
  12196=>"110110111",
  12197=>"110110111",
  12198=>"111111110",
  12199=>"011010000",
  12200=>"110100000",
  12201=>"001110111",
  12202=>"000000001",
  12203=>"111001011",
  12204=>"010000000",
  12205=>"000010111",
  12206=>"000000001",
  12207=>"011011000",
  12208=>"111100100",
  12209=>"000000000",
  12210=>"001000000",
  12211=>"000000100",
  12212=>"111100100",
  12213=>"011111100",
  12214=>"000111111",
  12215=>"110110010",
  12216=>"100111111",
  12217=>"000101111",
  12218=>"001001111",
  12219=>"111010000",
  12220=>"000000110",
  12221=>"000110010",
  12222=>"111111111",
  12223=>"001011111",
  12224=>"111111111",
  12225=>"000100100",
  12226=>"111111111",
  12227=>"111011001",
  12228=>"001001101",
  12229=>"001101111",
  12230=>"111111111",
  12231=>"111111011",
  12232=>"000101100",
  12233=>"010011111",
  12234=>"111101111",
  12235=>"111111111",
  12236=>"000010111",
  12237=>"100110111",
  12238=>"110110000",
  12239=>"000111011",
  12240=>"111111111",
  12241=>"010110100",
  12242=>"001001001",
  12243=>"111111001",
  12244=>"110110110",
  12245=>"111111111",
  12246=>"010000000",
  12247=>"011000000",
  12248=>"100101000",
  12249=>"111111111",
  12250=>"001011001",
  12251=>"111000000",
  12252=>"111100111",
  12253=>"111001001",
  12254=>"111111111",
  12255=>"001001001",
  12256=>"111111010",
  12257=>"101111111",
  12258=>"111111111",
  12259=>"011001001",
  12260=>"111111011",
  12261=>"100100000",
  12262=>"001000000",
  12263=>"111000000",
  12264=>"100100111",
  12265=>"000000000",
  12266=>"000000000",
  12267=>"000111111",
  12268=>"110000000",
  12269=>"110110110",
  12270=>"001000110",
  12271=>"111111111",
  12272=>"111000111",
  12273=>"111000000",
  12274=>"000110000",
  12275=>"111111111",
  12276=>"000001001",
  12277=>"011001111",
  12278=>"000000000",
  12279=>"011001100",
  12280=>"000000011",
  12281=>"100100100",
  12282=>"111111111",
  12283=>"011010000",
  12284=>"001001000",
  12285=>"111111111",
  12286=>"000111111",
  12287=>"001001001",
  12288=>"000000010",
  12289=>"110111001",
  12290=>"000110111",
  12291=>"000000000",
  12292=>"101100000",
  12293=>"100110011",
  12294=>"010010111",
  12295=>"111111111",
  12296=>"111100100",
  12297=>"000001111",
  12298=>"000000000",
  12299=>"111111011",
  12300=>"000000000",
  12301=>"111100111",
  12302=>"000100111",
  12303=>"000000110",
  12304=>"111011000",
  12305=>"000111111",
  12306=>"111111010",
  12307=>"110111111",
  12308=>"000000000",
  12309=>"001000000",
  12310=>"000000000",
  12311=>"100000011",
  12312=>"000000100",
  12313=>"000011110",
  12314=>"111111111",
  12315=>"001111111",
  12316=>"001000000",
  12317=>"111111111",
  12318=>"011111110",
  12319=>"011001000",
  12320=>"000000000",
  12321=>"000000000",
  12322=>"011111111",
  12323=>"011001000",
  12324=>"000000000",
  12325=>"000000000",
  12326=>"001011111",
  12327=>"111111111",
  12328=>"001000000",
  12329=>"101000001",
  12330=>"111111010",
  12331=>"111111000",
  12332=>"111111100",
  12333=>"111111011",
  12334=>"000000011",
  12335=>"011000111",
  12336=>"000000000",
  12337=>"000000000",
  12338=>"000010010",
  12339=>"000000000",
  12340=>"101001001",
  12341=>"000111110",
  12342=>"000000000",
  12343=>"100100100",
  12344=>"000000000",
  12345=>"000001000",
  12346=>"000000000",
  12347=>"111111111",
  12348=>"111111001",
  12349=>"000000000",
  12350=>"000100110",
  12351=>"111000000",
  12352=>"101001000",
  12353=>"111111111",
  12354=>"000011111",
  12355=>"000000000",
  12356=>"000000111",
  12357=>"111111111",
  12358=>"000000001",
  12359=>"110111000",
  12360=>"111110110",
  12361=>"110111111",
  12362=>"111111110",
  12363=>"110000000",
  12364=>"000000000",
  12365=>"000000000",
  12366=>"111000000",
  12367=>"000111111",
  12368=>"000011111",
  12369=>"000000000",
  12370=>"010000000",
  12371=>"001011101",
  12372=>"111111111",
  12373=>"001000000",
  12374=>"111101000",
  12375=>"000000100",
  12376=>"000000000",
  12377=>"101000000",
  12378=>"000000111",
  12379=>"001000000",
  12380=>"001000111",
  12381=>"111111000",
  12382=>"000000110",
  12383=>"111111010",
  12384=>"000000001",
  12385=>"111000000",
  12386=>"100000000",
  12387=>"101100111",
  12388=>"000000011",
  12389=>"000000000",
  12390=>"000111111",
  12391=>"011111111",
  12392=>"000111111",
  12393=>"111110111",
  12394=>"001111010",
  12395=>"011011000",
  12396=>"000000111",
  12397=>"111000000",
  12398=>"111111110",
  12399=>"110111111",
  12400=>"001000000",
  12401=>"000000000",
  12402=>"100110110",
  12403=>"000000000",
  12404=>"000000000",
  12405=>"111101111",
  12406=>"001100000",
  12407=>"001000000",
  12408=>"000000100",
  12409=>"111111111",
  12410=>"000000000",
  12411=>"100111000",
  12412=>"111111101",
  12413=>"000000111",
  12414=>"101101111",
  12415=>"000000111",
  12416=>"000000011",
  12417=>"000000111",
  12418=>"111011000",
  12419=>"000000011",
  12420=>"100100011",
  12421=>"000000111",
  12422=>"000000100",
  12423=>"000011000",
  12424=>"000000000",
  12425=>"000000111",
  12426=>"000000000",
  12427=>"000001101",
  12428=>"001100000",
  12429=>"010000011",
  12430=>"111111000",
  12431=>"000000000",
  12432=>"111111111",
  12433=>"000000000",
  12434=>"111000000",
  12435=>"110110000",
  12436=>"000000000",
  12437=>"111111000",
  12438=>"111111111",
  12439=>"110110100",
  12440=>"111001111",
  12441=>"111111111",
  12442=>"111111111",
  12443=>"010111010",
  12444=>"000111001",
  12445=>"111111001",
  12446=>"111111100",
  12447=>"110111000",
  12448=>"000000000",
  12449=>"111110001",
  12450=>"000001010",
  12451=>"000011100",
  12452=>"000001001",
  12453=>"111111111",
  12454=>"111011111",
  12455=>"000100000",
  12456=>"111111111",
  12457=>"000000111",
  12458=>"000000000",
  12459=>"111111100",
  12460=>"001000000",
  12461=>"000000111",
  12462=>"000000111",
  12463=>"010000100",
  12464=>"000000000",
  12465=>"000100000",
  12466=>"110111111",
  12467=>"010000000",
  12468=>"000000000",
  12469=>"011000000",
  12470=>"111000000",
  12471=>"000000001",
  12472=>"111000000",
  12473=>"111111111",
  12474=>"000000101",
  12475=>"011001111",
  12476=>"111011011",
  12477=>"101101111",
  12478=>"000000000",
  12479=>"111110100",
  12480=>"110011000",
  12481=>"010111011",
  12482=>"000110111",
  12483=>"001001001",
  12484=>"011110000",
  12485=>"111111111",
  12486=>"110100111",
  12487=>"000000101",
  12488=>"000111111",
  12489=>"111111111",
  12490=>"101000000",
  12491=>"000000100",
  12492=>"111100100",
  12493=>"100000000",
  12494=>"010011000",
  12495=>"100110111",
  12496=>"000111111",
  12497=>"111111111",
  12498=>"000000111",
  12499=>"110000110",
  12500=>"000000111",
  12501=>"111110100",
  12502=>"111000000",
  12503=>"000000001",
  12504=>"001000000",
  12505=>"000000000",
  12506=>"111000000",
  12507=>"111111001",
  12508=>"111001000",
  12509=>"011111111",
  12510=>"100001000",
  12511=>"111111111",
  12512=>"111111111",
  12513=>"111111000",
  12514=>"000001111",
  12515=>"000000111",
  12516=>"000111111",
  12517=>"111011000",
  12518=>"000110111",
  12519=>"111111011",
  12520=>"111110000",
  12521=>"011111111",
  12522=>"101001000",
  12523=>"111111001",
  12524=>"011011011",
  12525=>"100011000",
  12526=>"111111010",
  12527=>"111101111",
  12528=>"100000001",
  12529=>"000111001",
  12530=>"000000000",
  12531=>"001001111",
  12532=>"111111111",
  12533=>"110111001",
  12534=>"000110111",
  12535=>"111100111",
  12536=>"111000100",
  12537=>"111110010",
  12538=>"000000000",
  12539=>"000000000",
  12540=>"011001001",
  12541=>"111001001",
  12542=>"111011111",
  12543=>"000000000",
  12544=>"000000000",
  12545=>"001010010",
  12546=>"010000000",
  12547=>"010011111",
  12548=>"000000000",
  12549=>"001001101",
  12550=>"111111111",
  12551=>"000111111",
  12552=>"111111110",
  12553=>"111000010",
  12554=>"111111111",
  12555=>"110110000",
  12556=>"111010011",
  12557=>"000001111",
  12558=>"111101001",
  12559=>"000011011",
  12560=>"000111111",
  12561=>"000000000",
  12562=>"100000000",
  12563=>"000101101",
  12564=>"000111111",
  12565=>"010011110",
  12566=>"000100100",
  12567=>"000000000",
  12568=>"111111011",
  12569=>"000110111",
  12570=>"111111000",
  12571=>"000000111",
  12572=>"111000000",
  12573=>"000110111",
  12574=>"010010110",
  12575=>"111111111",
  12576=>"000000111",
  12577=>"111111111",
  12578=>"100110111",
  12579=>"101111111",
  12580=>"111111001",
  12581=>"000111111",
  12582=>"011111001",
  12583=>"000000111",
  12584=>"111011000",
  12585=>"000000000",
  12586=>"111000000",
  12587=>"011111111",
  12588=>"111111111",
  12589=>"011011001",
  12590=>"000000000",
  12591=>"000111011",
  12592=>"011011111",
  12593=>"000000110",
  12594=>"000110111",
  12595=>"111011000",
  12596=>"000000001",
  12597=>"111011111",
  12598=>"100101111",
  12599=>"111111000",
  12600=>"011000110",
  12601=>"111001111",
  12602=>"110110111",
  12603=>"000000111",
  12604=>"111111111",
  12605=>"000000111",
  12606=>"000000000",
  12607=>"111111111",
  12608=>"000000100",
  12609=>"000000000",
  12610=>"001001011",
  12611=>"111111111",
  12612=>"001111111",
  12613=>"111111111",
  12614=>"000000111",
  12615=>"100100000",
  12616=>"000000000",
  12617=>"000000011",
  12618=>"111010101",
  12619=>"000000110",
  12620=>"100110010",
  12621=>"000001000",
  12622=>"111111000",
  12623=>"111001000",
  12624=>"000110110",
  12625=>"010001111",
  12626=>"000011111",
  12627=>"000000000",
  12628=>"000000000",
  12629=>"011010000",
  12630=>"001011000",
  12631=>"111111100",
  12632=>"001001111",
  12633=>"100101101",
  12634=>"001111111",
  12635=>"101101111",
  12636=>"111111110",
  12637=>"000000000",
  12638=>"000000101",
  12639=>"111011000",
  12640=>"000000111",
  12641=>"001000000",
  12642=>"111101111",
  12643=>"111111111",
  12644=>"111100100",
  12645=>"000000000",
  12646=>"110000000",
  12647=>"111101000",
  12648=>"000000111",
  12649=>"000000001",
  12650=>"011011111",
  12651=>"001001111",
  12652=>"000011001",
  12653=>"000000111",
  12654=>"000010111",
  12655=>"000100110",
  12656=>"001001011",
  12657=>"000100111",
  12658=>"000000000",
  12659=>"011001111",
  12660=>"000100100",
  12661=>"111111111",
  12662=>"111001000",
  12663=>"111111000",
  12664=>"111000000",
  12665=>"000000011",
  12666=>"111111111",
  12667=>"111111111",
  12668=>"100111110",
  12669=>"111111111",
  12670=>"000101111",
  12671=>"000000110",
  12672=>"000000111",
  12673=>"111001111",
  12674=>"111111110",
  12675=>"111111111",
  12676=>"011000000",
  12677=>"000000111",
  12678=>"111100000",
  12679=>"000000000",
  12680=>"101001000",
  12681=>"011011011",
  12682=>"010000000",
  12683=>"010000000",
  12684=>"111011000",
  12685=>"010000000",
  12686=>"000000000",
  12687=>"011111111",
  12688=>"111111100",
  12689=>"101101000",
  12690=>"000000001",
  12691=>"111111110",
  12692=>"000000100",
  12693=>"000000011",
  12694=>"101111101",
  12695=>"000000000",
  12696=>"000111111",
  12697=>"000001001",
  12698=>"000000000",
  12699=>"110110110",
  12700=>"111001111",
  12701=>"111101000",
  12702=>"000000101",
  12703=>"000000000",
  12704=>"000000000",
  12705=>"111111000",
  12706=>"011000000",
  12707=>"111001000",
  12708=>"000000000",
  12709=>"000000000",
  12710=>"111111111",
  12711=>"111111111",
  12712=>"000000111",
  12713=>"111111101",
  12714=>"111011000",
  12715=>"001001111",
  12716=>"000000111",
  12717=>"111111011",
  12718=>"110100000",
  12719=>"000000000",
  12720=>"000001111",
  12721=>"001001000",
  12722=>"000110111",
  12723=>"111111010",
  12724=>"000000100",
  12725=>"100000000",
  12726=>"110100100",
  12727=>"110110110",
  12728=>"000110110",
  12729=>"000000000",
  12730=>"000000100",
  12731=>"111111110",
  12732=>"111111111",
  12733=>"001001011",
  12734=>"000000111",
  12735=>"010000001",
  12736=>"111000000",
  12737=>"111111000",
  12738=>"111000101",
  12739=>"011000111",
  12740=>"000000101",
  12741=>"111111100",
  12742=>"101001000",
  12743=>"000000111",
  12744=>"111111101",
  12745=>"110111001",
  12746=>"000000100",
  12747=>"111111000",
  12748=>"000111011",
  12749=>"011000000",
  12750=>"100001111",
  12751=>"111111111",
  12752=>"111000001",
  12753=>"000001011",
  12754=>"111111101",
  12755=>"000011111",
  12756=>"000000000",
  12757=>"101101111",
  12758=>"111111000",
  12759=>"000000011",
  12760=>"000000111",
  12761=>"000000101",
  12762=>"010111111",
  12763=>"001000111",
  12764=>"000110111",
  12765=>"111111110",
  12766=>"001011010",
  12767=>"111110000",
  12768=>"111000000",
  12769=>"000111111",
  12770=>"111010000",
  12771=>"111101100",
  12772=>"000010011",
  12773=>"111111111",
  12774=>"111111000",
  12775=>"111111010",
  12776=>"000110110",
  12777=>"100000000",
  12778=>"000000011",
  12779=>"000000000",
  12780=>"000000000",
  12781=>"000000100",
  12782=>"000111111",
  12783=>"000000111",
  12784=>"000110010",
  12785=>"000001111",
  12786=>"111111000",
  12787=>"100000001",
  12788=>"111000000",
  12789=>"100000000",
  12790=>"111111010",
  12791=>"001011001",
  12792=>"101000001",
  12793=>"000000000",
  12794=>"111110110",
  12795=>"010000010",
  12796=>"111100111",
  12797=>"010100000",
  12798=>"111010011",
  12799=>"000101111",
  12800=>"000000011",
  12801=>"000000000",
  12802=>"101111111",
  12803=>"001000101",
  12804=>"111111011",
  12805=>"000000111",
  12806=>"111001000",
  12807=>"011111111",
  12808=>"111111111",
  12809=>"101000111",
  12810=>"111111111",
  12811=>"111111111",
  12812=>"000110000",
  12813=>"000001000",
  12814=>"010000100",
  12815=>"000000000",
  12816=>"111011111",
  12817=>"010111111",
  12818=>"000100101",
  12819=>"001001111",
  12820=>"111111111",
  12821=>"111111111",
  12822=>"000001001",
  12823=>"110110111",
  12824=>"010110000",
  12825=>"000110100",
  12826=>"000111010",
  12827=>"000011010",
  12828=>"000001000",
  12829=>"111100111",
  12830=>"000000000",
  12831=>"000000001",
  12832=>"111111011",
  12833=>"000011000",
  12834=>"000000001",
  12835=>"010000000",
  12836=>"000000000",
  12837=>"000100000",
  12838=>"111010111",
  12839=>"111100000",
  12840=>"010011110",
  12841=>"100111111",
  12842=>"001000001",
  12843=>"111111100",
  12844=>"010000000",
  12845=>"000000000",
  12846=>"001100101",
  12847=>"111111110",
  12848=>"011011011",
  12849=>"000000101",
  12850=>"000100110",
  12851=>"000000000",
  12852=>"000111111",
  12853=>"111110110",
  12854=>"000111111",
  12855=>"101100100",
  12856=>"111111010",
  12857=>"000011110",
  12858=>"000000000",
  12859=>"000000000",
  12860=>"000101111",
  12861=>"000000000",
  12862=>"000000000",
  12863=>"111111111",
  12864=>"111011000",
  12865=>"100110100",
  12866=>"000000111",
  12867=>"000110000",
  12868=>"111111111",
  12869=>"101111111",
  12870=>"100100000",
  12871=>"111111001",
  12872=>"011011011",
  12873=>"111111111",
  12874=>"011111111",
  12875=>"011011011",
  12876=>"000000100",
  12877=>"110010111",
  12878=>"011000000",
  12879=>"000000000",
  12880=>"111111111",
  12881=>"000100110",
  12882=>"000000000",
  12883=>"100000111",
  12884=>"111111111",
  12885=>"111110110",
  12886=>"111111011",
  12887=>"111111111",
  12888=>"111100110",
  12889=>"111000001",
  12890=>"100000000",
  12891=>"001000000",
  12892=>"010000000",
  12893=>"111111111",
  12894=>"111111000",
  12895=>"111111101",
  12896=>"111111101",
  12897=>"000111000",
  12898=>"111111111",
  12899=>"000000000",
  12900=>"111111100",
  12901=>"000001000",
  12902=>"000111111",
  12903=>"000100101",
  12904=>"000000000",
  12905=>"110100110",
  12906=>"000000000",
  12907=>"100111111",
  12908=>"000000000",
  12909=>"000000010",
  12910=>"000000000",
  12911=>"101101100",
  12912=>"111111111",
  12913=>"100101100",
  12914=>"100100111",
  12915=>"111111000",
  12916=>"000000000",
  12917=>"000111111",
  12918=>"100100000",
  12919=>"010000000",
  12920=>"011011111",
  12921=>"000011111",
  12922=>"000000000",
  12923=>"111100111",
  12924=>"000000000",
  12925=>"100000001",
  12926=>"111111111",
  12927=>"000100111",
  12928=>"111111111",
  12929=>"111111001",
  12930=>"000110111",
  12931=>"001001000",
  12932=>"111011000",
  12933=>"000000000",
  12934=>"000001001",
  12935=>"100000010",
  12936=>"001000100",
  12937=>"111111000",
  12938=>"111000000",
  12939=>"000000011",
  12940=>"111101101",
  12941=>"000000000",
  12942=>"110100100",
  12943=>"000000001",
  12944=>"011001001",
  12945=>"001101111",
  12946=>"000000000",
  12947=>"011011010",
  12948=>"000010000",
  12949=>"111000101",
  12950=>"000000111",
  12951=>"000000000",
  12952=>"111100100",
  12953=>"111111011",
  12954=>"000000000",
  12955=>"000000000",
  12956=>"111111110",
  12957=>"000000000",
  12958=>"000010111",
  12959=>"111111011",
  12960=>"000000000",
  12961=>"000000000",
  12962=>"000100100",
  12963=>"000000000",
  12964=>"000000011",
  12965=>"000000111",
  12966=>"000000000",
  12967=>"110000000",
  12968=>"010010000",
  12969=>"001001000",
  12970=>"111111111",
  12971=>"111111111",
  12972=>"100110110",
  12973=>"000000000",
  12974=>"001000000",
  12975=>"001000000",
  12976=>"000000100",
  12977=>"111111011",
  12978=>"111110000",
  12979=>"000000000",
  12980=>"000000100",
  12981=>"001000000",
  12982=>"101100000",
  12983=>"111111111",
  12984=>"001000000",
  12985=>"001001011",
  12986=>"111010011",
  12987=>"111111001",
  12988=>"111001000",
  12989=>"111011000",
  12990=>"000000000",
  12991=>"101111111",
  12992=>"010000000",
  12993=>"000000000",
  12994=>"000000111",
  12995=>"000110000",
  12996=>"001101111",
  12997=>"011111111",
  12998=>"011000001",
  12999=>"111111111",
  13000=>"111010100",
  13001=>"000111111",
  13002=>"011000000",
  13003=>"111111111",
  13004=>"000000000",
  13005=>"000111111",
  13006=>"111111100",
  13007=>"000000000",
  13008=>"011101111",
  13009=>"000010010",
  13010=>"000100000",
  13011=>"111101101",
  13012=>"011000001",
  13013=>"010010000",
  13014=>"001111111",
  13015=>"100000000",
  13016=>"000000010",
  13017=>"110010100",
  13018=>"111111101",
  13019=>"010010011",
  13020=>"000000000",
  13021=>"000100000",
  13022=>"000000111",
  13023=>"100000110",
  13024=>"000000000",
  13025=>"000000111",
  13026=>"111111111",
  13027=>"000000100",
  13028=>"000101111",
  13029=>"111111110",
  13030=>"011111111",
  13031=>"011000000",
  13032=>"111111000",
  13033=>"001011100",
  13034=>"111111110",
  13035=>"111111010",
  13036=>"000110000",
  13037=>"111110100",
  13038=>"000000000",
  13039=>"111111110",
  13040=>"111000000",
  13041=>"111000000",
  13042=>"000000000",
  13043=>"111100001",
  13044=>"111111111",
  13045=>"010111111",
  13046=>"000100100",
  13047=>"000000100",
  13048=>"000110111",
  13049=>"000000000",
  13050=>"000000000",
  13051=>"111111001",
  13052=>"011101111",
  13053=>"000000110",
  13054=>"000010000",
  13055=>"000000000",
  13056=>"000000000",
  13057=>"011000000",
  13058=>"111101111",
  13059=>"000100111",
  13060=>"000100111",
  13061=>"111100110",
  13062=>"000000000",
  13063=>"111111000",
  13064=>"000000000",
  13065=>"111000000",
  13066=>"111111101",
  13067=>"100110100",
  13068=>"100000000",
  13069=>"111111001",
  13070=>"111111111",
  13071=>"000000000",
  13072=>"100110111",
  13073=>"111111111",
  13074=>"111111111",
  13075=>"011011011",
  13076=>"000000000",
  13077=>"000001001",
  13078=>"101101001",
  13079=>"000111000",
  13080=>"110000110",
  13081=>"111111111",
  13082=>"111111111",
  13083=>"111111111",
  13084=>"101001000",
  13085=>"111100111",
  13086=>"100110111",
  13087=>"000000111",
  13088=>"000000000",
  13089=>"111000000",
  13090=>"000000000",
  13091=>"000000101",
  13092=>"101111111",
  13093=>"110111111",
  13094=>"000011111",
  13095=>"000000101",
  13096=>"000000100",
  13097=>"111111011",
  13098=>"011011000",
  13099=>"111111001",
  13100=>"111111101",
  13101=>"001001111",
  13102=>"000000000",
  13103=>"000000000",
  13104=>"111111111",
  13105=>"111111111",
  13106=>"001000001",
  13107=>"111100111",
  13108=>"111000000",
  13109=>"000000000",
  13110=>"000111111",
  13111=>"011011011",
  13112=>"011111111",
  13113=>"000100100",
  13114=>"000000000",
  13115=>"010100000",
  13116=>"000010011",
  13117=>"000000000",
  13118=>"000001011",
  13119=>"111111001",
  13120=>"000001000",
  13121=>"111111111",
  13122=>"000000111",
  13123=>"011111111",
  13124=>"000000000",
  13125=>"100100110",
  13126=>"111111111",
  13127=>"000000000",
  13128=>"000000000",
  13129=>"111100000",
  13130=>"010000000",
  13131=>"100000000",
  13132=>"100100111",
  13133=>"111111100",
  13134=>"000000001",
  13135=>"011111111",
  13136=>"000000000",
  13137=>"000000000",
  13138=>"111110111",
  13139=>"111010111",
  13140=>"111111111",
  13141=>"000001001",
  13142=>"110010111",
  13143=>"111100100",
  13144=>"111111111",
  13145=>"111000000",
  13146=>"110011000",
  13147=>"000000000",
  13148=>"111111111",
  13149=>"111111111",
  13150=>"000100000",
  13151=>"011011111",
  13152=>"001001011",
  13153=>"111111111",
  13154=>"000000000",
  13155=>"100000111",
  13156=>"110010000",
  13157=>"011001111",
  13158=>"000100111",
  13159=>"110111111",
  13160=>"011011010",
  13161=>"110110010",
  13162=>"000000000",
  13163=>"000110001",
  13164=>"100100000",
  13165=>"010000001",
  13166=>"000000001",
  13167=>"000011000",
  13168=>"111111111",
  13169=>"000000000",
  13170=>"000111001",
  13171=>"011000000",
  13172=>"000000000",
  13173=>"010110000",
  13174=>"000000000",
  13175=>"111111101",
  13176=>"000000000",
  13177=>"000100111",
  13178=>"000000011",
  13179=>"000110010",
  13180=>"100100100",
  13181=>"000000111",
  13182=>"111111111",
  13183=>"000000000",
  13184=>"010001101",
  13185=>"111111111",
  13186=>"111011001",
  13187=>"111101000",
  13188=>"000101111",
  13189=>"000000000",
  13190=>"011000111",
  13191=>"101000101",
  13192=>"001001000",
  13193=>"111111101",
  13194=>"000000000",
  13195=>"001100110",
  13196=>"000101111",
  13197=>"011011011",
  13198=>"111100110",
  13199=>"111111110",
  13200=>"111111111",
  13201=>"111111111",
  13202=>"111001000",
  13203=>"000000100",
  13204=>"111000101",
  13205=>"000000000",
  13206=>"111111001",
  13207=>"110110110",
  13208=>"000000000",
  13209=>"010000000",
  13210=>"000100110",
  13211=>"000000000",
  13212=>"111111010",
  13213=>"001001000",
  13214=>"011110111",
  13215=>"010000000",
  13216=>"111111111",
  13217=>"111110110",
  13218=>"110111000",
  13219=>"110110100",
  13220=>"000000000",
  13221=>"111111111",
  13222=>"111011000",
  13223=>"010111111",
  13224=>"000010000",
  13225=>"100101101",
  13226=>"011111111",
  13227=>"100110111",
  13228=>"111111111",
  13229=>"100000110",
  13230=>"000011111",
  13231=>"010011111",
  13232=>"111111010",
  13233=>"111000000",
  13234=>"000000000",
  13235=>"010100110",
  13236=>"000010000",
  13237=>"111111111",
  13238=>"111111000",
  13239=>"111000000",
  13240=>"000000000",
  13241=>"000000000",
  13242=>"111101111",
  13243=>"100111011",
  13244=>"111001000",
  13245=>"000001001",
  13246=>"100100000",
  13247=>"011011000",
  13248=>"000000000",
  13249=>"101101111",
  13250=>"011010000",
  13251=>"000001111",
  13252=>"111111111",
  13253=>"000110100",
  13254=>"000001000",
  13255=>"001101001",
  13256=>"111111000",
  13257=>"000000000",
  13258=>"111111100",
  13259=>"000000100",
  13260=>"000001000",
  13261=>"111111111",
  13262=>"011010000",
  13263=>"001000010",
  13264=>"000000000",
  13265=>"111111111",
  13266=>"000111110",
  13267=>"000000000",
  13268=>"111111001",
  13269=>"111010000",
  13270=>"000000001",
  13271=>"000010000",
  13272=>"001001000",
  13273=>"000000001",
  13274=>"110111001",
  13275=>"111100000",
  13276=>"111101111",
  13277=>"111100000",
  13278=>"111110000",
  13279=>"010111011",
  13280=>"110100000",
  13281=>"111111111",
  13282=>"011001111",
  13283=>"101101111",
  13284=>"111111111",
  13285=>"001111101",
  13286=>"100000100",
  13287=>"100000101",
  13288=>"111011111",
  13289=>"011111111",
  13290=>"111110000",
  13291=>"001011000",
  13292=>"100111111",
  13293=>"000000000",
  13294=>"100101111",
  13295=>"000000101",
  13296=>"000000000",
  13297=>"111101100",
  13298=>"000011001",
  13299=>"010010110",
  13300=>"111111110",
  13301=>"000000111",
  13302=>"000100000",
  13303=>"010010110",
  13304=>"011111011",
  13305=>"000110000",
  13306=>"001000000",
  13307=>"111000101",
  13308=>"000000000",
  13309=>"111111111",
  13310=>"010000000",
  13311=>"000000001",
  13312=>"101111111",
  13313=>"010000000",
  13314=>"000100100",
  13315=>"000100110",
  13316=>"000001110",
  13317=>"110100000",
  13318=>"000000000",
  13319=>"111111111",
  13320=>"111111111",
  13321=>"000000111",
  13322=>"000000000",
  13323=>"111001011",
  13324=>"000000000",
  13325=>"111111011",
  13326=>"000000011",
  13327=>"111110010",
  13328=>"011111111",
  13329=>"000001000",
  13330=>"111111111",
  13331=>"001000000",
  13332=>"111111111",
  13333=>"001001111",
  13334=>"111111110",
  13335=>"000000110",
  13336=>"000110000",
  13337=>"011111110",
  13338=>"001000101",
  13339=>"011111011",
  13340=>"000110111",
  13341=>"101000000",
  13342=>"001001001",
  13343=>"000000000",
  13344=>"110111000",
  13345=>"000000000",
  13346=>"111100000",
  13347=>"110100000",
  13348=>"000001110",
  13349=>"111110010",
  13350=>"110100000",
  13351=>"000000100",
  13352=>"011111111",
  13353=>"111011001",
  13354=>"001000000",
  13355=>"000000100",
  13356=>"010000000",
  13357=>"111011101",
  13358=>"110111111",
  13359=>"011001001",
  13360=>"100000100",
  13361=>"000000111",
  13362=>"000000100",
  13363=>"000100111",
  13364=>"000000000",
  13365=>"101111111",
  13366=>"100000000",
  13367=>"010111111",
  13368=>"101000011",
  13369=>"110110111",
  13370=>"000000000",
  13371=>"110110111",
  13372=>"111111111",
  13373=>"111111101",
  13374=>"111111111",
  13375=>"111111111",
  13376=>"000000000",
  13377=>"111011111",
  13378=>"110100000",
  13379=>"111111000",
  13380=>"101011111",
  13381=>"001100110",
  13382=>"000000000",
  13383=>"000000000",
  13384=>"011111111",
  13385=>"000000000",
  13386=>"000011111",
  13387=>"001001001",
  13388=>"110110111",
  13389=>"000000000",
  13390=>"000111111",
  13391=>"111101000",
  13392=>"111111111",
  13393=>"110111111",
  13394=>"101101011",
  13395=>"111111111",
  13396=>"110110111",
  13397=>"101000111",
  13398=>"111111111",
  13399=>"000000000",
  13400=>"000101111",
  13401=>"000000000",
  13402=>"111100111",
  13403=>"110000000",
  13404=>"000000111",
  13405=>"111111111",
  13406=>"000001111",
  13407=>"011000000",
  13408=>"000100000",
  13409=>"111110100",
  13410=>"111100000",
  13411=>"111111111",
  13412=>"000111111",
  13413=>"110110100",
  13414=>"000000000",
  13415=>"111111111",
  13416=>"111111011",
  13417=>"001001111",
  13418=>"111011011",
  13419=>"000011111",
  13420=>"011111011",
  13421=>"100100000",
  13422=>"011011111",
  13423=>"001011111",
  13424=>"110110111",
  13425=>"100000000",
  13426=>"111111111",
  13427=>"110111111",
  13428=>"110010010",
  13429=>"000000000",
  13430=>"110111111",
  13431=>"100100111",
  13432=>"110000000",
  13433=>"111101111",
  13434=>"001001111",
  13435=>"000000000",
  13436=>"000000000",
  13437=>"111110111",
  13438=>"111110000",
  13439=>"111111111",
  13440=>"111111111",
  13441=>"111111111",
  13442=>"011000000",
  13443=>"100100010",
  13444=>"000000100",
  13445=>"111111011",
  13446=>"000000110",
  13447=>"011111111",
  13448=>"111111111",
  13449=>"000000111",
  13450=>"100000000",
  13451=>"000000000",
  13452=>"000000000",
  13453=>"110100000",
  13454=>"110110110",
  13455=>"000000000",
  13456=>"111111111",
  13457=>"100100101",
  13458=>"001000000",
  13459=>"000000111",
  13460=>"111101111",
  13461=>"111111111",
  13462=>"000000000",
  13463=>"111011001",
  13464=>"000000000",
  13465=>"111111111",
  13466=>"000000100",
  13467=>"000000000",
  13468=>"111111111",
  13469=>"000000000",
  13470=>"100000100",
  13471=>"000000000",
  13472=>"000000000",
  13473=>"000000000",
  13474=>"000000000",
  13475=>"000100111",
  13476=>"001000000",
  13477=>"111011110",
  13478=>"111100000",
  13479=>"011011111",
  13480=>"110110110",
  13481=>"111111111",
  13482=>"111000000",
  13483=>"000000000",
  13484=>"111111111",
  13485=>"000001000",
  13486=>"001000000",
  13487=>"000111111",
  13488=>"000000111",
  13489=>"100100110",
  13490=>"000000000",
  13491=>"001000101",
  13492=>"010000000",
  13493=>"100110100",
  13494=>"000000000",
  13495=>"000000110",
  13496=>"110000000",
  13497=>"000000000",
  13498=>"000111100",
  13499=>"111111111",
  13500=>"000010011",
  13501=>"111111110",
  13502=>"010110111",
  13503=>"111111111",
  13504=>"000010011",
  13505=>"000100000",
  13506=>"111111111",
  13507=>"011011111",
  13508=>"000000011",
  13509=>"000111110",
  13510=>"110000110",
  13511=>"000101100",
  13512=>"010010000",
  13513=>"000000100",
  13514=>"110111111",
  13515=>"100101101",
  13516=>"000000000",
  13517=>"000111111",
  13518=>"000000110",
  13519=>"101000100",
  13520=>"000000000",
  13521=>"000000001",
  13522=>"110111111",
  13523=>"010111110",
  13524=>"111111111",
  13525=>"001001001",
  13526=>"000000001",
  13527=>"000000000",
  13528=>"000000000",
  13529=>"010011011",
  13530=>"011001001",
  13531=>"111001000",
  13532=>"111111000",
  13533=>"100100111",
  13534=>"000000111",
  13535=>"111111111",
  13536=>"000000000",
  13537=>"111111011",
  13538=>"011000000",
  13539=>"111111111",
  13540=>"100100100",
  13541=>"111111111",
  13542=>"111111111",
  13543=>"001101101",
  13544=>"100111111",
  13545=>"101001110",
  13546=>"110111111",
  13547=>"111111000",
  13548=>"110111111",
  13549=>"000001001",
  13550=>"111111111",
  13551=>"000000000",
  13552=>"001000000",
  13553=>"000111110",
  13554=>"111111111",
  13555=>"101000111",
  13556=>"111110110",
  13557=>"000000000",
  13558=>"100101101",
  13559=>"000000000",
  13560=>"000111111",
  13561=>"000000000",
  13562=>"000000110",
  13563=>"000111111",
  13564=>"011011111",
  13565=>"110111111",
  13566=>"111111111",
  13567=>"000111110",
  13568=>"111111110",
  13569=>"111111111",
  13570=>"000100000",
  13571=>"111111010",
  13572=>"000000000",
  13573=>"111011000",
  13574=>"100111111",
  13575=>"001011011",
  13576=>"000000110",
  13577=>"111000000",
  13578=>"000000000",
  13579=>"100101000",
  13580=>"000000111",
  13581=>"110001111",
  13582=>"101111111",
  13583=>"000000010",
  13584=>"001100100",
  13585=>"001111111",
  13586=>"111100100",
  13587=>"000000000",
  13588=>"011111111",
  13589=>"011001001",
  13590=>"110101111",
  13591=>"000000000",
  13592=>"000000110",
  13593=>"000000100",
  13594=>"000000000",
  13595=>"010110110",
  13596=>"000000100",
  13597=>"110110000",
  13598=>"011000000",
  13599=>"111111000",
  13600=>"110110111",
  13601=>"000000000",
  13602=>"001001001",
  13603=>"011111011",
  13604=>"000000000",
  13605=>"110100101",
  13606=>"000000100",
  13607=>"000001111",
  13608=>"111011000",
  13609=>"100110111",
  13610=>"000000000",
  13611=>"100101100",
  13612=>"111111111",
  13613=>"001001000",
  13614=>"000000000",
  13615=>"111111111",
  13616=>"000000000",
  13617=>"100101111",
  13618=>"111110000",
  13619=>"011011111",
  13620=>"000000000",
  13621=>"111100000",
  13622=>"001101101",
  13623=>"000000000",
  13624=>"100111001",
  13625=>"100111000",
  13626=>"000000000",
  13627=>"000101000",
  13628=>"001001111",
  13629=>"001100110",
  13630=>"000000000",
  13631=>"111111110",
  13632=>"110100110",
  13633=>"000010000",
  13634=>"000000000",
  13635=>"000000100",
  13636=>"000000111",
  13637=>"000000000",
  13638=>"000110000",
  13639=>"000011111",
  13640=>"000000000",
  13641=>"000001000",
  13642=>"010011001",
  13643=>"110100100",
  13644=>"100110110",
  13645=>"011111111",
  13646=>"000000100",
  13647=>"000000000",
  13648=>"111111110",
  13649=>"001000000",
  13650=>"100111101",
  13651=>"000000100",
  13652=>"111111110",
  13653=>"011001001",
  13654=>"110111110",
  13655=>"000000000",
  13656=>"111111111",
  13657=>"000000000",
  13658=>"111110111",
  13659=>"100000110",
  13660=>"111111111",
  13661=>"000000000",
  13662=>"000001011",
  13663=>"000000000",
  13664=>"001001000",
  13665=>"111110111",
  13666=>"000010110",
  13667=>"111111111",
  13668=>"111111110",
  13669=>"001111010",
  13670=>"011111111",
  13671=>"001011111",
  13672=>"001000001",
  13673=>"000000000",
  13674=>"111111111",
  13675=>"110011011",
  13676=>"111111011",
  13677=>"000000000",
  13678=>"111111000",
  13679=>"101101100",
  13680=>"000000000",
  13681=>"000000000",
  13682=>"000000010",
  13683=>"111111111",
  13684=>"001111111",
  13685=>"110100111",
  13686=>"000100100",
  13687=>"001101000",
  13688=>"000000110",
  13689=>"111111011",
  13690=>"111000000",
  13691=>"111111001",
  13692=>"000000100",
  13693=>"000000000",
  13694=>"111111000",
  13695=>"001000000",
  13696=>"001000000",
  13697=>"001111110",
  13698=>"000001011",
  13699=>"000000000",
  13700=>"111111111",
  13701=>"001000000",
  13702=>"100100100",
  13703=>"010000000",
  13704=>"000100100",
  13705=>"100101001",
  13706=>"111000000",
  13707=>"011111111",
  13708=>"000000111",
  13709=>"011111011",
  13710=>"000000000",
  13711=>"000100111",
  13712=>"010000000",
  13713=>"111111110",
  13714=>"000000000",
  13715=>"000011011",
  13716=>"000000111",
  13717=>"000011111",
  13718=>"001000000",
  13719=>"001111110",
  13720=>"000011001",
  13721=>"110100100",
  13722=>"000001011",
  13723=>"001010110",
  13724=>"111011011",
  13725=>"000000000",
  13726=>"000000011",
  13727=>"000100111",
  13728=>"000000000",
  13729=>"011111111",
  13730=>"110111111",
  13731=>"001011111",
  13732=>"110100000",
  13733=>"000000000",
  13734=>"111110100",
  13735=>"000001011",
  13736=>"111111111",
  13737=>"111001000",
  13738=>"000000000",
  13739=>"111111111",
  13740=>"000000010",
  13741=>"001000000",
  13742=>"000001001",
  13743=>"111111111",
  13744=>"111001111",
  13745=>"111111111",
  13746=>"000111000",
  13747=>"000000001",
  13748=>"000000000",
  13749=>"111111111",
  13750=>"111111111",
  13751=>"111111111",
  13752=>"000000010",
  13753=>"011011111",
  13754=>"001000000",
  13755=>"000000000",
  13756=>"111111011",
  13757=>"100000000",
  13758=>"111111101",
  13759=>"000100000",
  13760=>"111111111",
  13761=>"000000000",
  13762=>"000000000",
  13763=>"111111110",
  13764=>"000101011",
  13765=>"000000010",
  13766=>"111001111",
  13767=>"111111111",
  13768=>"000000000",
  13769=>"000000000",
  13770=>"111000101",
  13771=>"111111000",
  13772=>"001011000",
  13773=>"000000000",
  13774=>"011011111",
  13775=>"111100100",
  13776=>"000111111",
  13777=>"000000000",
  13778=>"011111111",
  13779=>"000000111",
  13780=>"100100111",
  13781=>"000000000",
  13782=>"111111111",
  13783=>"000000011",
  13784=>"100100000",
  13785=>"110100101",
  13786=>"000000001",
  13787=>"111010111",
  13788=>"011111111",
  13789=>"001111011",
  13790=>"100000001",
  13791=>"000001011",
  13792=>"111111111",
  13793=>"000011001",
  13794=>"101100000",
  13795=>"100001000",
  13796=>"000000000",
  13797=>"111111010",
  13798=>"000011011",
  13799=>"011011001",
  13800=>"111111111",
  13801=>"000010000",
  13802=>"111111011",
  13803=>"110000000",
  13804=>"000111001",
  13805=>"101100100",
  13806=>"111111100",
  13807=>"000110110",
  13808=>"000000000",
  13809=>"100101001",
  13810=>"111111111",
  13811=>"100100000",
  13812=>"110010010",
  13813=>"010000110",
  13814=>"010110110",
  13815=>"000000000",
  13816=>"111111111",
  13817=>"000000000",
  13818=>"010111111",
  13819=>"011011001",
  13820=>"000011111",
  13821=>"000000000",
  13822=>"000000000",
  13823=>"000000110",
  13824=>"100100001",
  13825=>"000000000",
  13826=>"000001111",
  13827=>"100111111",
  13828=>"110111111",
  13829=>"001000010",
  13830=>"000000111",
  13831=>"000000000",
  13832=>"011011001",
  13833=>"111111000",
  13834=>"111111111",
  13835=>"110111111",
  13836=>"110110100",
  13837=>"100011111",
  13838=>"011111011",
  13839=>"000000000",
  13840=>"001000000",
  13841=>"000000000",
  13842=>"111101111",
  13843=>"000000000",
  13844=>"111111111",
  13845=>"101001011",
  13846=>"111111111",
  13847=>"111111111",
  13848=>"110111110",
  13849=>"000000000",
  13850=>"111000000",
  13851=>"000000011",
  13852=>"111111000",
  13853=>"101000000",
  13854=>"000000000",
  13855=>"110111111",
  13856=>"000000000",
  13857=>"111111111",
  13858=>"111111011",
  13859=>"000000111",
  13860=>"111100000",
  13861=>"000110110",
  13862=>"011000000",
  13863=>"000000101",
  13864=>"000010000",
  13865=>"000000000",
  13866=>"000010111",
  13867=>"111111111",
  13868=>"011001000",
  13869=>"111111111",
  13870=>"000000111",
  13871=>"000110110",
  13872=>"000110111",
  13873=>"000000000",
  13874=>"001011001",
  13875=>"000000110",
  13876=>"111110110",
  13877=>"000000000",
  13878=>"101000000",
  13879=>"000000000",
  13880=>"011000000",
  13881=>"000011011",
  13882=>"111111111",
  13883=>"110011111",
  13884=>"000000000",
  13885=>"111111111",
  13886=>"101000000",
  13887=>"001000001",
  13888=>"111001000",
  13889=>"010011000",
  13890=>"000111111",
  13891=>"001001001",
  13892=>"110110000",
  13893=>"110111111",
  13894=>"111001001",
  13895=>"111111111",
  13896=>"011111100",
  13897=>"001001000",
  13898=>"111101001",
  13899=>"111111011",
  13900=>"000000000",
  13901=>"000000001",
  13902=>"000000011",
  13903=>"101000000",
  13904=>"111111111",
  13905=>"111111111",
  13906=>"000000000",
  13907=>"110110110",
  13908=>"000000000",
  13909=>"110110110",
  13910=>"000000000",
  13911=>"111001000",
  13912=>"011111111",
  13913=>"000000000",
  13914=>"111111100",
  13915=>"001001000",
  13916=>"000000011",
  13917=>"000000000",
  13918=>"110111010",
  13919=>"111111111",
  13920=>"011111111",
  13921=>"110110111",
  13922=>"000000000",
  13923=>"000000000",
  13924=>"111011011",
  13925=>"010000000",
  13926=>"111111000",
  13927=>"000000000",
  13928=>"010111111",
  13929=>"000000000",
  13930=>"000011111",
  13931=>"000111111",
  13932=>"000000000",
  13933=>"010111111",
  13934=>"111000000",
  13935=>"111110110",
  13936=>"010111110",
  13937=>"000000111",
  13938=>"000000001",
  13939=>"111111000",
  13940=>"000000000",
  13941=>"000000111",
  13942=>"111110011",
  13943=>"001000000",
  13944=>"001010000",
  13945=>"000000000",
  13946=>"011111111",
  13947=>"111100100",
  13948=>"111111111",
  13949=>"111101111",
  13950=>"000010111",
  13951=>"011000000",
  13952=>"000111011",
  13953=>"111111111",
  13954=>"111110000",
  13955=>"000011000",
  13956=>"100111111",
  13957=>"111101111",
  13958=>"000010000",
  13959=>"111000000",
  13960=>"111000100",
  13961=>"111111101",
  13962=>"000000000",
  13963=>"000000000",
  13964=>"000000100",
  13965=>"111111111",
  13966=>"000000000",
  13967=>"010011000",
  13968=>"111111111",
  13969=>"111111111",
  13970=>"111111100",
  13971=>"001001000",
  13972=>"000001000",
  13973=>"111111111",
  13974=>"111111111",
  13975=>"111111111",
  13976=>"000000000",
  13977=>"111111111",
  13978=>"000000000",
  13979=>"111111000",
  13980=>"000000000",
  13981=>"000000011",
  13982=>"111111110",
  13983=>"000000000",
  13984=>"111110000",
  13985=>"000010111",
  13986=>"010111111",
  13987=>"000000001",
  13988=>"011011001",
  13989=>"000110110",
  13990=>"111100000",
  13991=>"110111111",
  13992=>"000000000",
  13993=>"000000000",
  13994=>"111000000",
  13995=>"111011000",
  13996=>"111110111",
  13997=>"110110000",
  13998=>"111110000",
  13999=>"000100000",
  14000=>"010111111",
  14001=>"111000000",
  14002=>"001011011",
  14003=>"111111000",
  14004=>"000000101",
  14005=>"101111111",
  14006=>"111111111",
  14007=>"100000011",
  14008=>"001001001",
  14009=>"111111011",
  14010=>"000000001",
  14011=>"001001111",
  14012=>"111111111",
  14013=>"010111100",
  14014=>"100111000",
  14015=>"000000011",
  14016=>"111111111",
  14017=>"000010011",
  14018=>"001000000",
  14019=>"000010111",
  14020=>"001011000",
  14021=>"000000000",
  14022=>"001001000",
  14023=>"000100000",
  14024=>"111111111",
  14025=>"000000000",
  14026=>"110111000",
  14027=>"101101111",
  14028=>"000000001",
  14029=>"000000000",
  14030=>"101101111",
  14031=>"111111111",
  14032=>"111111111",
  14033=>"000000000",
  14034=>"000110111",
  14035=>"111111111",
  14036=>"111110100",
  14037=>"111111111",
  14038=>"100111111",
  14039=>"000000000",
  14040=>"001001001",
  14041=>"111111111",
  14042=>"111111000",
  14043=>"111111001",
  14044=>"111111111",
  14045=>"111100010",
  14046=>"111011001",
  14047=>"011011000",
  14048=>"000000000",
  14049=>"000000010",
  14050=>"000100100",
  14051=>"000000000",
  14052=>"001111111",
  14053=>"000100111",
  14054=>"111111111",
  14055=>"011111111",
  14056=>"111111001",
  14057=>"001011111",
  14058=>"000000000",
  14059=>"100101111",
  14060=>"111111111",
  14061=>"111101111",
  14062=>"000100111",
  14063=>"111111111",
  14064=>"000000000",
  14065=>"111111111",
  14066=>"000000000",
  14067=>"000001111",
  14068=>"000000000",
  14069=>"111111111",
  14070=>"101100100",
  14071=>"000000111",
  14072=>"111111111",
  14073=>"011001000",
  14074=>"000001111",
  14075=>"001111111",
  14076=>"110111100",
  14077=>"001001001",
  14078=>"111101001",
  14079=>"110110100",
  14080=>"100000000",
  14081=>"011001001",
  14082=>"111111001",
  14083=>"010000000",
  14084=>"011011000",
  14085=>"000011011",
  14086=>"111111111",
  14087=>"111111000",
  14088=>"000000000",
  14089=>"000000000",
  14090=>"000000001",
  14091=>"000000100",
  14092=>"001001101",
  14093=>"111011110",
  14094=>"011011100",
  14095=>"000000011",
  14096=>"100111111",
  14097=>"000000000",
  14098=>"111111111",
  14099=>"000011111",
  14100=>"000000000",
  14101=>"000000000",
  14102=>"010011000",
  14103=>"111111000",
  14104=>"000011111",
  14105=>"111111101",
  14106=>"111111111",
  14107=>"111000111",
  14108=>"000000000",
  14109=>"100000100",
  14110=>"111000100",
  14111=>"101100100",
  14112=>"111111101",
  14113=>"111111110",
  14114=>"011000000",
  14115=>"000111111",
  14116=>"000000000",
  14117=>"000000000",
  14118=>"011111111",
  14119=>"000000000",
  14120=>"000000101",
  14121=>"111111111",
  14122=>"011010010",
  14123=>"101101000",
  14124=>"111111111",
  14125=>"001001001",
  14126=>"111111111",
  14127=>"000000000",
  14128=>"000000000",
  14129=>"000000000",
  14130=>"000000000",
  14131=>"000111111",
  14132=>"111110110",
  14133=>"001000100",
  14134=>"000100111",
  14135=>"111000000",
  14136=>"111111000",
  14137=>"000000111",
  14138=>"111111111",
  14139=>"000000000",
  14140=>"100100100",
  14141=>"100011101",
  14142=>"000000000",
  14143=>"000111011",
  14144=>"011011001",
  14145=>"000000000",
  14146=>"000001011",
  14147=>"111111111",
  14148=>"100000000",
  14149=>"110110000",
  14150=>"011000111",
  14151=>"110000000",
  14152=>"000000000",
  14153=>"000000000",
  14154=>"000000000",
  14155=>"111111111",
  14156=>"000000000",
  14157=>"110111111",
  14158=>"001011011",
  14159=>"100100100",
  14160=>"111001011",
  14161=>"000111110",
  14162=>"111111111",
  14163=>"000000000",
  14164=>"111111011",
  14165=>"000111111",
  14166=>"111111111",
  14167=>"000000000",
  14168=>"000000000",
  14169=>"111100000",
  14170=>"111111000",
  14171=>"000000001",
  14172=>"000000000",
  14173=>"111010000",
  14174=>"000001001",
  14175=>"000000000",
  14176=>"000000000",
  14177=>"111000000",
  14178=>"000000000",
  14179=>"000000000",
  14180=>"000000000",
  14181=>"000000000",
  14182=>"000000000",
  14183=>"000000010",
  14184=>"110110110",
  14185=>"000010010",
  14186=>"000111111",
  14187=>"001000000",
  14188=>"110100110",
  14189=>"000111111",
  14190=>"000000111",
  14191=>"000000000",
  14192=>"110111000",
  14193=>"000000011",
  14194=>"000000000",
  14195=>"000000000",
  14196=>"111110000",
  14197=>"000000000",
  14198=>"000000001",
  14199=>"000000000",
  14200=>"000000000",
  14201=>"011001000",
  14202=>"111000111",
  14203=>"111000000",
  14204=>"111111110",
  14205=>"010000000",
  14206=>"101000000",
  14207=>"000000000",
  14208=>"000000000",
  14209=>"011111111",
  14210=>"111111000",
  14211=>"000111011",
  14212=>"001000110",
  14213=>"111101001",
  14214=>"000111111",
  14215=>"001001001",
  14216=>"111111110",
  14217=>"011000000",
  14218=>"000000000",
  14219=>"111101000",
  14220=>"111111111",
  14221=>"111111111",
  14222=>"001001000",
  14223=>"100100111",
  14224=>"000000000",
  14225=>"111111111",
  14226=>"000001111",
  14227=>"111000100",
  14228=>"111111111",
  14229=>"000000000",
  14230=>"110110111",
  14231=>"111111111",
  14232=>"111111111",
  14233=>"111011001",
  14234=>"111111111",
  14235=>"000000000",
  14236=>"101100111",
  14237=>"001111111",
  14238=>"000000000",
  14239=>"000000000",
  14240=>"111111111",
  14241=>"000100000",
  14242=>"101000000",
  14243=>"000000000",
  14244=>"011000000",
  14245=>"111011000",
  14246=>"111011000",
  14247=>"111111110",
  14248=>"000000000",
  14249=>"111110000",
  14250=>"111110000",
  14251=>"101100111",
  14252=>"111110010",
  14253=>"000000000",
  14254=>"111111100",
  14255=>"000000000",
  14256=>"000011001",
  14257=>"000000111",
  14258=>"100100110",
  14259=>"111011000",
  14260=>"011011000",
  14261=>"111111111",
  14262=>"111111001",
  14263=>"001111111",
  14264=>"010011111",
  14265=>"000001111",
  14266=>"111111000",
  14267=>"111111101",
  14268=>"101101111",
  14269=>"100000000",
  14270=>"000000001",
  14271=>"110000000",
  14272=>"000110110",
  14273=>"000000000",
  14274=>"111000000",
  14275=>"000000000",
  14276=>"100110110",
  14277=>"001111111",
  14278=>"110111000",
  14279=>"000000101",
  14280=>"000000110",
  14281=>"000000100",
  14282=>"001001001",
  14283=>"000000000",
  14284=>"001000001",
  14285=>"000000111",
  14286=>"000000111",
  14287=>"000101111",
  14288=>"000000000",
  14289=>"001001011",
  14290=>"110110111",
  14291=>"111111011",
  14292=>"000000000",
  14293=>"111111111",
  14294=>"000100000",
  14295=>"111111001",
  14296=>"000011111",
  14297=>"111111111",
  14298=>"110000000",
  14299=>"000011111",
  14300=>"111111111",
  14301=>"100000000",
  14302=>"000000001",
  14303=>"000000000",
  14304=>"000000000",
  14305=>"111111111",
  14306=>"000000011",
  14307=>"000000000",
  14308=>"111111011",
  14309=>"011000000",
  14310=>"111111010",
  14311=>"000000000",
  14312=>"011011001",
  14313=>"000000000",
  14314=>"100100100",
  14315=>"001000000",
  14316=>"001100000",
  14317=>"111111100",
  14318=>"000001001",
  14319=>"000000000",
  14320=>"000000011",
  14321=>"000000000",
  14322=>"001111111",
  14323=>"000000000",
  14324=>"001011111",
  14325=>"111110100",
  14326=>"000000000",
  14327=>"000000000",
  14328=>"000111111",
  14329=>"111111101",
  14330=>"010010000",
  14331=>"111111000",
  14332=>"011000001",
  14333=>"111001111",
  14334=>"011000000",
  14335=>"001001000",
  14336=>"011011011",
  14337=>"111111111",
  14338=>"000000111",
  14339=>"000000000",
  14340=>"111111111",
  14341=>"110110000",
  14342=>"001000000",
  14343=>"111100111",
  14344=>"111110000",
  14345=>"110100000",
  14346=>"111111111",
  14347=>"100110110",
  14348=>"111101001",
  14349=>"100000000",
  14350=>"000000000",
  14351=>"111111111",
  14352=>"111000000",
  14353=>"000000000",
  14354=>"111111000",
  14355=>"111111111",
  14356=>"111010000",
  14357=>"111001000",
  14358=>"001000111",
  14359=>"000000000",
  14360=>"111110111",
  14361=>"100000000",
  14362=>"111111111",
  14363=>"011011010",
  14364=>"000001001",
  14365=>"111111111",
  14366=>"101001001",
  14367=>"111111110",
  14368=>"000100110",
  14369=>"101111111",
  14370=>"111111100",
  14371=>"000000000",
  14372=>"111111111",
  14373=>"000001001",
  14374=>"110110100",
  14375=>"000000001",
  14376=>"111111111",
  14377=>"111011000",
  14378=>"010100111",
  14379=>"101000000",
  14380=>"000111100",
  14381=>"000001000",
  14382=>"111111111",
  14383=>"111111111",
  14384=>"000000000",
  14385=>"111111000",
  14386=>"011111000",
  14387=>"000110000",
  14388=>"000100110",
  14389=>"000000000",
  14390=>"111111111",
  14391=>"110110000",
  14392=>"000000000",
  14393=>"010000011",
  14394=>"001101100",
  14395=>"111000000",
  14396=>"000000000",
  14397=>"111111111",
  14398=>"000001111",
  14399=>"000000000",
  14400=>"111111111",
  14401=>"100000010",
  14402=>"000000111",
  14403=>"000000000",
  14404=>"111111110",
  14405=>"111111000",
  14406=>"000010110",
  14407=>"011000000",
  14408=>"111011000",
  14409=>"111101111",
  14410=>"000000100",
  14411=>"111110100",
  14412=>"111111111",
  14413=>"000000000",
  14414=>"101111111",
  14415=>"111111000",
  14416=>"110110000",
  14417=>"000100001",
  14418=>"010111101",
  14419=>"001000100",
  14420=>"000110111",
  14421=>"111111111",
  14422=>"000000000",
  14423=>"000110100",
  14424=>"000000000",
  14425=>"000000001",
  14426=>"111011000",
  14427=>"111111000",
  14428=>"000000000",
  14429=>"100111111",
  14430=>"111111111",
  14431=>"000111111",
  14432=>"000000000",
  14433=>"111111111",
  14434=>"100100110",
  14435=>"000000000",
  14436=>"000000000",
  14437=>"111111111",
  14438=>"000001111",
  14439=>"100110000",
  14440=>"111111111",
  14441=>"001111111",
  14442=>"110000000",
  14443=>"111111011",
  14444=>"001000001",
  14445=>"000000000",
  14446=>"111111100",
  14447=>"101000000",
  14448=>"000101000",
  14449=>"000000000",
  14450=>"111100000",
  14451=>"111111110",
  14452=>"110111111",
  14453=>"110110010",
  14454=>"000000000",
  14455=>"110000000",
  14456=>"111111000",
  14457=>"000000000",
  14458=>"000000000",
  14459=>"111111110",
  14460=>"000000100",
  14461=>"000111111",
  14462=>"110000000",
  14463=>"110110000",
  14464=>"000000000",
  14465=>"111011001",
  14466=>"000011011",
  14467=>"000000000",
  14468=>"000000001",
  14469=>"000000111",
  14470=>"000000000",
  14471=>"100000100",
  14472=>"000000000",
  14473=>"110000110",
  14474=>"111011000",
  14475=>"000000011",
  14476=>"111110000",
  14477=>"000000000",
  14478=>"000000110",
  14479=>"000011010",
  14480=>"000100111",
  14481=>"100111111",
  14482=>"010100111",
  14483=>"000011111",
  14484=>"000000111",
  14485=>"111111100",
  14486=>"111111111",
  14487=>"000000100",
  14488=>"000000100",
  14489=>"000000001",
  14490=>"111111110",
  14491=>"001000000",
  14492=>"111011100",
  14493=>"000011000",
  14494=>"000000000",
  14495=>"000000011",
  14496=>"000000000",
  14497=>"111111111",
  14498=>"000001011",
  14499=>"001001000",
  14500=>"000000000",
  14501=>"000000110",
  14502=>"111111101",
  14503=>"110110000",
  14504=>"111100101",
  14505=>"100110100",
  14506=>"100111111",
  14507=>"000000000",
  14508=>"111111111",
  14509=>"001011001",
  14510=>"111111100",
  14511=>"001000100",
  14512=>"101100000",
  14513=>"001001000",
  14514=>"111111111",
  14515=>"111111111",
  14516=>"110110110",
  14517=>"000000100",
  14518=>"111111111",
  14519=>"011011111",
  14520=>"111001001",
  14521=>"000000001",
  14522=>"000000000",
  14523=>"000000000",
  14524=>"010000000",
  14525=>"111111111",
  14526=>"000111111",
  14527=>"111000001",
  14528=>"000000000",
  14529=>"110111000",
  14530=>"111111111",
  14531=>"111111111",
  14532=>"100100111",
  14533=>"000000000",
  14534=>"111111111",
  14535=>"110111101",
  14536=>"000000000",
  14537=>"000000000",
  14538=>"100110000",
  14539=>"000111011",
  14540=>"001001011",
  14541=>"100001001",
  14542=>"111111011",
  14543=>"111111111",
  14544=>"000000000",
  14545=>"000000000",
  14546=>"100100000",
  14547=>"000000000",
  14548=>"111000000",
  14549=>"110110100",
  14550=>"100111111",
  14551=>"100100111",
  14552=>"011000000",
  14553=>"010000000",
  14554=>"110100000",
  14555=>"000000000",
  14556=>"111111111",
  14557=>"110100111",
  14558=>"011111111",
  14559=>"111111101",
  14560=>"111101011",
  14561=>"000000000",
  14562=>"000000000",
  14563=>"011011010",
  14564=>"100111111",
  14565=>"111110010",
  14566=>"101000000",
  14567=>"000000000",
  14568=>"000100111",
  14569=>"000000000",
  14570=>"000000110",
  14571=>"000000000",
  14572=>"111111111",
  14573=>"111111111",
  14574=>"111111111",
  14575=>"000110111",
  14576=>"010001100",
  14577=>"111011101",
  14578=>"000000000",
  14579=>"000000001",
  14580=>"011111110",
  14581=>"000100111",
  14582=>"011110011",
  14583=>"000000001",
  14584=>"000000000",
  14585=>"000000000",
  14586=>"111111011",
  14587=>"000010110",
  14588=>"101101111",
  14589=>"111110110",
  14590=>"011011000",
  14591=>"001001111",
  14592=>"111000010",
  14593=>"110011001",
  14594=>"000000111",
  14595=>"111111111",
  14596=>"111111111",
  14597=>"100110100",
  14598=>"000000000",
  14599=>"101011101",
  14600=>"000000000",
  14601=>"000000111",
  14602=>"111111111",
  14603=>"000000000",
  14604=>"111111111",
  14605=>"110111111",
  14606=>"111111110",
  14607=>"101101100",
  14608=>"110100100",
  14609=>"011000000",
  14610=>"111111111",
  14611=>"000000000",
  14612=>"000000000",
  14613=>"110111010",
  14614=>"000000000",
  14615=>"010000000",
  14616=>"000000000",
  14617=>"000000011",
  14618=>"111010000",
  14619=>"111111100",
  14620=>"100110111",
  14621=>"111111001",
  14622=>"111000000",
  14623=>"111111111",
  14624=>"111100110",
  14625=>"000111111",
  14626=>"101000000",
  14627=>"111111111",
  14628=>"010011111",
  14629=>"010110010",
  14630=>"111111110",
  14631=>"100100000",
  14632=>"110111111",
  14633=>"000000000",
  14634=>"111111100",
  14635=>"000100000",
  14636=>"110111000",
  14637=>"111100000",
  14638=>"000000110",
  14639=>"111111000",
  14640=>"000000000",
  14641=>"110111111",
  14642=>"110100100",
  14643=>"101101111",
  14644=>"000000000",
  14645=>"101100100",
  14646=>"001000000",
  14647=>"000000100",
  14648=>"111111100",
  14649=>"000000000",
  14650=>"000000111",
  14651=>"011001001",
  14652=>"100100000",
  14653=>"000000000",
  14654=>"100000011",
  14655=>"000110111",
  14656=>"111111101",
  14657=>"011111110",
  14658=>"000000000",
  14659=>"000101111",
  14660=>"110100000",
  14661=>"111111000",
  14662=>"100100000",
  14663=>"000000000",
  14664=>"111010000",
  14665=>"110111111",
  14666=>"101000000",
  14667=>"001101111",
  14668=>"010000000",
  14669=>"111111010",
  14670=>"110111111",
  14671=>"001000000",
  14672=>"000000000",
  14673=>"000000000",
  14674=>"000110111",
  14675=>"000000000",
  14676=>"000000000",
  14677=>"011000011",
  14678=>"111111111",
  14679=>"001000000",
  14680=>"100000111",
  14681=>"110111111",
  14682=>"000000000",
  14683=>"011001101",
  14684=>"111111111",
  14685=>"000000000",
  14686=>"000101001",
  14687=>"000000000",
  14688=>"000000001",
  14689=>"000000000",
  14690=>"111111100",
  14691=>"000000110",
  14692=>"111111001",
  14693=>"000000000",
  14694=>"110001000",
  14695=>"000000000",
  14696=>"110110010",
  14697=>"111000000",
  14698=>"111111100",
  14699=>"111011110",
  14700=>"110111110",
  14701=>"110111111",
  14702=>"010100111",
  14703=>"000000000",
  14704=>"110111000",
  14705=>"001001001",
  14706=>"011000000",
  14707=>"011011000",
  14708=>"100000000",
  14709=>"111110000",
  14710=>"111111101",
  14711=>"010000000",
  14712=>"111111111",
  14713=>"111001000",
  14714=>"110111110",
  14715=>"001011011",
  14716=>"000100111",
  14717=>"111111100",
  14718=>"111111110",
  14719=>"111111111",
  14720=>"110111111",
  14721=>"110111000",
  14722=>"111001000",
  14723=>"111111111",
  14724=>"111111000",
  14725=>"000000000",
  14726=>"111111011",
  14727=>"111100100",
  14728=>"000000000",
  14729=>"111111111",
  14730=>"111100010",
  14731=>"111111111",
  14732=>"111111111",
  14733=>"001001001",
  14734=>"000000000",
  14735=>"000000000",
  14736=>"000110111",
  14737=>"111110100",
  14738=>"101101000",
  14739=>"000000000",
  14740=>"000001100",
  14741=>"100100000",
  14742=>"111111111",
  14743=>"001000000",
  14744=>"011001000",
  14745=>"110111111",
  14746=>"000000101",
  14747=>"000000000",
  14748=>"000000000",
  14749=>"000100000",
  14750=>"000000000",
  14751=>"111111110",
  14752=>"111111111",
  14753=>"000000110",
  14754=>"001000000",
  14755=>"110000000",
  14756=>"001000100",
  14757=>"000000000",
  14758=>"000001000",
  14759=>"000000100",
  14760=>"000000000",
  14761=>"000000000",
  14762=>"001000000",
  14763=>"000000000",
  14764=>"110111111",
  14765=>"111111111",
  14766=>"000011111",
  14767=>"111111111",
  14768=>"000000100",
  14769=>"111111100",
  14770=>"000000111",
  14771=>"000000000",
  14772=>"111111111",
  14773=>"110111111",
  14774=>"000000000",
  14775=>"000000000",
  14776=>"111111111",
  14777=>"000000000",
  14778=>"111111100",
  14779=>"001111111",
  14780=>"000001100",
  14781=>"111111111",
  14782=>"111001000",
  14783=>"000000000",
  14784=>"011000000",
  14785=>"001000000",
  14786=>"001011111",
  14787=>"111111111",
  14788=>"111101111",
  14789=>"000000111",
  14790=>"000000001",
  14791=>"000000000",
  14792=>"011000000",
  14793=>"111100000",
  14794=>"000000000",
  14795=>"000000000",
  14796=>"000000010",
  14797=>"001011000",
  14798=>"111000000",
  14799=>"110000000",
  14800=>"000000000",
  14801=>"001001100",
  14802=>"000000000",
  14803=>"110110110",
  14804=>"000000000",
  14805=>"111111111",
  14806=>"000000000",
  14807=>"011011011",
  14808=>"000000000",
  14809=>"100100000",
  14810=>"001111111",
  14811=>"110100100",
  14812=>"111001000",
  14813=>"000100100",
  14814=>"111111111",
  14815=>"100000000",
  14816=>"001001000",
  14817=>"011111111",
  14818=>"010100110",
  14819=>"000000000",
  14820=>"000000010",
  14821=>"111001000",
  14822=>"000000000",
  14823=>"111011000",
  14824=>"000000000",
  14825=>"111111111",
  14826=>"111000000",
  14827=>"111111111",
  14828=>"011011111",
  14829=>"010110100",
  14830=>"000000000",
  14831=>"000000000",
  14832=>"001000111",
  14833=>"000000000",
  14834=>"000000000",
  14835=>"000000000",
  14836=>"111111110",
  14837=>"110110000",
  14838=>"100000111",
  14839=>"000000000",
  14840=>"000000000",
  14841=>"001000000",
  14842=>"000000000",
  14843=>"101111001",
  14844=>"111110100",
  14845=>"000000001",
  14846=>"000000010",
  14847=>"000000111",
  14848=>"000000000",
  14849=>"000000011",
  14850=>"111000000",
  14851=>"111111111",
  14852=>"110111111",
  14853=>"111111111",
  14854=>"000000000",
  14855=>"111100111",
  14856=>"000000000",
  14857=>"000000111",
  14858=>"100000000",
  14859=>"000001111",
  14860=>"111111111",
  14861=>"001001000",
  14862=>"000011011",
  14863=>"100101100",
  14864=>"111111111",
  14865=>"010111111",
  14866=>"000000000",
  14867=>"111111111",
  14868=>"111111111",
  14869=>"111111111",
  14870=>"010111111",
  14871=>"111111110",
  14872=>"111111111",
  14873=>"000000010",
  14874=>"000111111",
  14875=>"000000000",
  14876=>"111111011",
  14877=>"111011000",
  14878=>"000000000",
  14879=>"000000111",
  14880=>"000000011",
  14881=>"111110111",
  14882=>"111111111",
  14883=>"000000000",
  14884=>"000100110",
  14885=>"000000000",
  14886=>"101111111",
  14887=>"000000000",
  14888=>"001000010",
  14889=>"000000001",
  14890=>"111111111",
  14891=>"111111111",
  14892=>"111000000",
  14893=>"100010000",
  14894=>"011011000",
  14895=>"000000000",
  14896=>"111111111",
  14897=>"000000000",
  14898=>"110000000",
  14899=>"000110111",
  14900=>"110110110",
  14901=>"000100110",
  14902=>"111111111",
  14903=>"111101111",
  14904=>"000110000",
  14905=>"011111111",
  14906=>"111111111",
  14907=>"100111011",
  14908=>"001000000",
  14909=>"001000000",
  14910=>"000000000",
  14911=>"000000000",
  14912=>"111111001",
  14913=>"110111111",
  14914=>"111111111",
  14915=>"000101100",
  14916=>"000000000",
  14917=>"001000100",
  14918=>"001001000",
  14919=>"000000000",
  14920=>"111111111",
  14921=>"111111111",
  14922=>"111100111",
  14923=>"011000000",
  14924=>"111011001",
  14925=>"000000000",
  14926=>"010010000",
  14927=>"111001000",
  14928=>"000000100",
  14929=>"111011011",
  14930=>"000010000",
  14931=>"000100000",
  14932=>"111111011",
  14933=>"011011001",
  14934=>"111111111",
  14935=>"111111111",
  14936=>"011011111",
  14937=>"111111111",
  14938=>"101101111",
  14939=>"000100100",
  14940=>"011111010",
  14941=>"000000000",
  14942=>"001001000",
  14943=>"001100000",
  14944=>"000000000",
  14945=>"011111111",
  14946=>"000011011",
  14947=>"111111111",
  14948=>"111111111",
  14949=>"111001001",
  14950=>"111111111",
  14951=>"000000001",
  14952=>"111011000",
  14953=>"001011000",
  14954=>"001111111",
  14955=>"111111111",
  14956=>"000000000",
  14957=>"000000000",
  14958=>"111111111",
  14959=>"000000000",
  14960=>"000000000",
  14961=>"000000000",
  14962=>"111111111",
  14963=>"000110000",
  14964=>"000000000",
  14965=>"111111110",
  14966=>"000110111",
  14967=>"000000000",
  14968=>"000000000",
  14969=>"111111111",
  14970=>"111100000",
  14971=>"000000000",
  14972=>"100100100",
  14973=>"011000100",
  14974=>"000010000",
  14975=>"000111111",
  14976=>"000000000",
  14977=>"011111111",
  14978=>"101100100",
  14979=>"111111111",
  14980=>"000111111",
  14981=>"000111111",
  14982=>"111111110",
  14983=>"111010000",
  14984=>"111111001",
  14985=>"111000000",
  14986=>"111010010",
  14987=>"000000000",
  14988=>"000000011",
  14989=>"000111011",
  14990=>"000000000",
  14991=>"111111111",
  14992=>"000000000",
  14993=>"000000000",
  14994=>"111100100",
  14995=>"111111111",
  14996=>"111111111",
  14997=>"000000100",
  14998=>"000000000",
  14999=>"111111111",
  15000=>"000000000",
  15001=>"000000000",
  15002=>"110101111",
  15003=>"110100100",
  15004=>"111111111",
  15005=>"000000000",
  15006=>"100100110",
  15007=>"111111111",
  15008=>"100100100",
  15009=>"111000000",
  15010=>"000000000",
  15011=>"000111111",
  15012=>"000000000",
  15013=>"011001000",
  15014=>"111101101",
  15015=>"000000000",
  15016=>"001001111",
  15017=>"000000000",
  15018=>"111001000",
  15019=>"000000100",
  15020=>"001011111",
  15021=>"110100101",
  15022=>"011110111",
  15023=>"000100100",
  15024=>"111110111",
  15025=>"000100010",
  15026=>"111111110",
  15027=>"101000000",
  15028=>"111111111",
  15029=>"111111000",
  15030=>"000111111",
  15031=>"011011011",
  15032=>"111111111",
  15033=>"111111000",
  15034=>"011111100",
  15035=>"011100111",
  15036=>"111111111",
  15037=>"000000000",
  15038=>"111111111",
  15039=>"000110000",
  15040=>"000000000",
  15041=>"110000000",
  15042=>"000000000",
  15043=>"111111111",
  15044=>"111111111",
  15045=>"000000000",
  15046=>"011111111",
  15047=>"000110110",
  15048=>"000100100",
  15049=>"001001000",
  15050=>"000000000",
  15051=>"000000000",
  15052=>"111111111",
  15053=>"000111111",
  15054=>"000100100",
  15055=>"011111111",
  15056=>"000000000",
  15057=>"000000000",
  15058=>"001001000",
  15059=>"011011111",
  15060=>"111111011",
  15061=>"000100111",
  15062=>"000000001",
  15063=>"111100111",
  15064=>"011001100",
  15065=>"000000000",
  15066=>"111111111",
  15067=>"011011101",
  15068=>"000000100",
  15069=>"111111011",
  15070=>"000011111",
  15071=>"000000000",
  15072=>"000000000",
  15073=>"000000000",
  15074=>"011000000",
  15075=>"111000111",
  15076=>"111111000",
  15077=>"000000111",
  15078=>"001000001",
  15079=>"111111111",
  15080=>"000000000",
  15081=>"010111111",
  15082=>"000000000",
  15083=>"000000001",
  15084=>"000000000",
  15085=>"000000000",
  15086=>"000000001",
  15087=>"000000000",
  15088=>"111111000",
  15089=>"111111100",
  15090=>"111100000",
  15091=>"000000000",
  15092=>"111111111",
  15093=>"011001001",
  15094=>"100100110",
  15095=>"111111111",
  15096=>"111000000",
  15097=>"000000000",
  15098=>"011110000",
  15099=>"110111111",
  15100=>"000000001",
  15101=>"001001000",
  15102=>"000000100",
  15103=>"111111011",
  15104=>"001101011",
  15105=>"000001000",
  15106=>"000000000",
  15107=>"011111111",
  15108=>"110000000",
  15109=>"000000000",
  15110=>"111111111",
  15111=>"111111111",
  15112=>"000000001",
  15113=>"000000000",
  15114=>"111001100",
  15115=>"011011011",
  15116=>"000000000",
  15117=>"111111110",
  15118=>"000000000",
  15119=>"100000000",
  15120=>"000000000",
  15121=>"000110111",
  15122=>"111111111",
  15123=>"111111111",
  15124=>"000010010",
  15125=>"000000001",
  15126=>"111110110",
  15127=>"011111100",
  15128=>"110100100",
  15129=>"100000000",
  15130=>"101101111",
  15131=>"111100100",
  15132=>"100000000",
  15133=>"111111111",
  15134=>"001000111",
  15135=>"000010111",
  15136=>"000110100",
  15137=>"001001001",
  15138=>"101111100",
  15139=>"111111111",
  15140=>"001001101",
  15141=>"111111111",
  15142=>"000100110",
  15143=>"111111000",
  15144=>"100100000",
  15145=>"000000000",
  15146=>"111111111",
  15147=>"111111000",
  15148=>"000000000",
  15149=>"000000000",
  15150=>"111000111",
  15151=>"000000000",
  15152=>"111111101",
  15153=>"000000000",
  15154=>"000000110",
  15155=>"000011011",
  15156=>"101100100",
  15157=>"000000110",
  15158=>"011111111",
  15159=>"111111111",
  15160=>"010000000",
  15161=>"011111001",
  15162=>"000000000",
  15163=>"001111001",
  15164=>"011001001",
  15165=>"000100100",
  15166=>"111111111",
  15167=>"111111000",
  15168=>"010110000",
  15169=>"101000000",
  15170=>"000000000",
  15171=>"111111111",
  15172=>"001000000",
  15173=>"000000111",
  15174=>"000100000",
  15175=>"000000000",
  15176=>"000000000",
  15177=>"000000000",
  15178=>"111110100",
  15179=>"101110101",
  15180=>"000000000",
  15181=>"111111111",
  15182=>"101000000",
  15183=>"001111110",
  15184=>"000100100",
  15185=>"111110100",
  15186=>"111100100",
  15187=>"000000101",
  15188=>"111111111",
  15189=>"011011011",
  15190=>"000000110",
  15191=>"000100100",
  15192=>"111111000",
  15193=>"100000100",
  15194=>"000000000",
  15195=>"110000001",
  15196=>"101101001",
  15197=>"000000000",
  15198=>"001000001",
  15199=>"110110010",
  15200=>"111111111",
  15201=>"000000000",
  15202=>"000000000",
  15203=>"111101100",
  15204=>"001111111",
  15205=>"000000000",
  15206=>"000000000",
  15207=>"010100111",
  15208=>"111111100",
  15209=>"001011011",
  15210=>"000000000",
  15211=>"100101100",
  15212=>"000111101",
  15213=>"111111111",
  15214=>"001000000",
  15215=>"111111000",
  15216=>"000000000",
  15217=>"000000100",
  15218=>"000000000",
  15219=>"000000000",
  15220=>"000000000",
  15221=>"110000000",
  15222=>"000000111",
  15223=>"000010111",
  15224=>"000000000",
  15225=>"111011000",
  15226=>"000000000",
  15227=>"000011010",
  15228=>"011000000",
  15229=>"000000010",
  15230=>"000000100",
  15231=>"000000000",
  15232=>"000000000",
  15233=>"111100100",
  15234=>"000000001",
  15235=>"000000000",
  15236=>"010011111",
  15237=>"011111011",
  15238=>"011010010",
  15239=>"110111111",
  15240=>"001111110",
  15241=>"000110111",
  15242=>"000000000",
  15243=>"000011000",
  15244=>"111111111",
  15245=>"111111111",
  15246=>"001011111",
  15247=>"001000001",
  15248=>"100101100",
  15249=>"110110110",
  15250=>"011110111",
  15251=>"111111111",
  15252=>"000000000",
  15253=>"000010011",
  15254=>"111111111",
  15255=>"000000000",
  15256=>"000000100",
  15257=>"111001000",
  15258=>"111111110",
  15259=>"011111111",
  15260=>"111111111",
  15261=>"111111111",
  15262=>"000001100",
  15263=>"000000010",
  15264=>"000000000",
  15265=>"011011001",
  15266=>"101111111",
  15267=>"111111111",
  15268=>"001000000",
  15269=>"000000000",
  15270=>"001011000",
  15271=>"110000000",
  15272=>"000000000",
  15273=>"111100100",
  15274=>"000011011",
  15275=>"000000000",
  15276=>"001001011",
  15277=>"011111110",
  15278=>"000011111",
  15279=>"000000000",
  15280=>"010111011",
  15281=>"111111000",
  15282=>"000000000",
  15283=>"111111111",
  15284=>"001011111",
  15285=>"111111111",
  15286=>"000000000",
  15287=>"000000100",
  15288=>"111000101",
  15289=>"011011000",
  15290=>"011011111",
  15291=>"000000000",
  15292=>"111111010",
  15293=>"111111110",
  15294=>"001000110",
  15295=>"111011011",
  15296=>"111111111",
  15297=>"000111111",
  15298=>"111111111",
  15299=>"111111001",
  15300=>"000000111",
  15301=>"000000100",
  15302=>"000000000",
  15303=>"000011000",
  15304=>"000000000",
  15305=>"001000000",
  15306=>"001000000",
  15307=>"111101111",
  15308=>"111110000",
  15309=>"110000000",
  15310=>"111111111",
  15311=>"111001100",
  15312=>"001011011",
  15313=>"101100100",
  15314=>"111001001",
  15315=>"000000000",
  15316=>"000000000",
  15317=>"001001011",
  15318=>"111101000",
  15319=>"111100100",
  15320=>"111111111",
  15321=>"100000000",
  15322=>"001000000",
  15323=>"011111111",
  15324=>"111111111",
  15325=>"000000000",
  15326=>"111111100",
  15327=>"000011111",
  15328=>"000000000",
  15329=>"111111111",
  15330=>"011011000",
  15331=>"000000000",
  15332=>"000101000",
  15333=>"100000011",
  15334=>"000000011",
  15335=>"000000000",
  15336=>"001000000",
  15337=>"011011001",
  15338=>"001010011",
  15339=>"100100000",
  15340=>"101000000",
  15341=>"000100111",
  15342=>"000100111",
  15343=>"000000000",
  15344=>"000000100",
  15345=>"000000000",
  15346=>"111111111",
  15347=>"100000000",
  15348=>"000000000",
  15349=>"010000100",
  15350=>"011101110",
  15351=>"000000100",
  15352=>"000110011",
  15353=>"101101111",
  15354=>"111111111",
  15355=>"111111111",
  15356=>"011001000",
  15357=>"111111111",
  15358=>"111000000",
  15359=>"110111111",
  15360=>"000111111",
  15361=>"000000100",
  15362=>"000000000",
  15363=>"001011111",
  15364=>"000111111",
  15365=>"111110111",
  15366=>"111000000",
  15367=>"111111111",
  15368=>"001001001",
  15369=>"110111011",
  15370=>"100110011",
  15371=>"000110110",
  15372=>"000110110",
  15373=>"111111101",
  15374=>"000000111",
  15375=>"111111111",
  15376=>"000000100",
  15377=>"110011111",
  15378=>"000000010",
  15379=>"111000000",
  15380=>"111011000",
  15381=>"111111111",
  15382=>"000000000",
  15383=>"111111011",
  15384=>"111111111",
  15385=>"111111110",
  15386=>"110000011",
  15387=>"000110000",
  15388=>"000000000",
  15389=>"101111111",
  15390=>"110000000",
  15391=>"111101101",
  15392=>"010000000",
  15393=>"110110000",
  15394=>"000000010",
  15395=>"110000000",
  15396=>"111111111",
  15397=>"000000111",
  15398=>"111111111",
  15399=>"100000000",
  15400=>"111111111",
  15401=>"000000000",
  15402=>"111110111",
  15403=>"111000000",
  15404=>"000000000",
  15405=>"100000100",
  15406=>"110100100",
  15407=>"111011111",
  15408=>"111111111",
  15409=>"000110110",
  15410=>"011011001",
  15411=>"111011111",
  15412=>"110111000",
  15413=>"011011011",
  15414=>"111111111",
  15415=>"111111111",
  15416=>"110010000",
  15417=>"111111111",
  15418=>"000000000",
  15419=>"111111011",
  15420=>"000010111",
  15421=>"100100000",
  15422=>"000000000",
  15423=>"111000000",
  15424=>"000000100",
  15425=>"000111011",
  15426=>"000000000",
  15427=>"111111110",
  15428=>"000000000",
  15429=>"011000100",
  15430=>"111011111",
  15431=>"001001111",
  15432=>"000000000",
  15433=>"101001111",
  15434=>"111111111",
  15435=>"111111111",
  15436=>"111100100",
  15437=>"000001101",
  15438=>"111110000",
  15439=>"111110000",
  15440=>"000000000",
  15441=>"001001001",
  15442=>"010110110",
  15443=>"000001000",
  15444=>"000001001",
  15445=>"000110100",
  15446=>"111100111",
  15447=>"011010011",
  15448=>"111111110",
  15449=>"111101100",
  15450=>"000000000",
  15451=>"101001001",
  15452=>"000000000",
  15453=>"000000001",
  15454=>"000000000",
  15455=>"000000000",
  15456=>"100101111",
  15457=>"000000101",
  15458=>"000000000",
  15459=>"101100110",
  15460=>"001111111",
  15461=>"111000001",
  15462=>"110000000",
  15463=>"000110010",
  15464=>"000000000",
  15465=>"011111011",
  15466=>"111111111",
  15467=>"000000000",
  15468=>"000000000",
  15469=>"110111111",
  15470=>"000000000",
  15471=>"110011111",
  15472=>"000000000",
  15473=>"000001111",
  15474=>"000000001",
  15475=>"011001011",
  15476=>"110000000",
  15477=>"011111111",
  15478=>"000000000",
  15479=>"100100000",
  15480=>"110110110",
  15481=>"111111111",
  15482=>"111111111",
  15483=>"111111111",
  15484=>"000100100",
  15485=>"111111000",
  15486=>"000000000",
  15487=>"111111111",
  15488=>"000000000",
  15489=>"111011111",
  15490=>"011010000",
  15491=>"111111111",
  15492=>"000000000",
  15493=>"000001111",
  15494=>"000100100",
  15495=>"000000000",
  15496=>"011000000",
  15497=>"000100000",
  15498=>"100100000",
  15499=>"000000000",
  15500=>"000000000",
  15501=>"111111111",
  15502=>"101000001",
  15503=>"111111110",
  15504=>"000000000",
  15505=>"111010000",
  15506=>"001111111",
  15507=>"111110110",
  15508=>"000110111",
  15509=>"011110110",
  15510=>"001000000",
  15511=>"111110000",
  15512=>"111111111",
  15513=>"111000000",
  15514=>"111111111",
  15515=>"001001000",
  15516=>"111111111",
  15517=>"001111110",
  15518=>"110000000",
  15519=>"111111111",
  15520=>"000000000",
  15521=>"111111111",
  15522=>"000000000",
  15523=>"011111000",
  15524=>"110111111",
  15525=>"101001000",
  15526=>"000110111",
  15527=>"011111101",
  15528=>"001000000",
  15529=>"110111111",
  15530=>"111011000",
  15531=>"100000000",
  15532=>"000001111",
  15533=>"000001111",
  15534=>"100100000",
  15535=>"000010111",
  15536=>"000000000",
  15537=>"100100101",
  15538=>"111111111",
  15539=>"111111110",
  15540=>"011001000",
  15541=>"000000000",
  15542=>"010000111",
  15543=>"000000000",
  15544=>"111110111",
  15545=>"111011111",
  15546=>"000000000",
  15547=>"111111110",
  15548=>"000000111",
  15549=>"000000000",
  15550=>"111111111",
  15551=>"111010000",
  15552=>"001000001",
  15553=>"111111111",
  15554=>"011010000",
  15555=>"000000000",
  15556=>"111111110",
  15557=>"111111111",
  15558=>"111111100",
  15559=>"000010000",
  15560=>"111111111",
  15561=>"111100100",
  15562=>"110110111",
  15563=>"110000000",
  15564=>"111100000",
  15565=>"011010111",
  15566=>"111111111",
  15567=>"000000100",
  15568=>"111111111",
  15569=>"010110111",
  15570=>"111110111",
  15571=>"111111111",
  15572=>"111111111",
  15573=>"011001000",
  15574=>"000111111",
  15575=>"111111001",
  15576=>"101100100",
  15577=>"000000000",
  15578=>"001000000",
  15579=>"000000001",
  15580=>"111100000",
  15581=>"111111111",
  15582=>"111111111",
  15583=>"000000000",
  15584=>"111111000",
  15585=>"000000000",
  15586=>"000000000",
  15587=>"101111000",
  15588=>"000000110",
  15589=>"111111000",
  15590=>"010000000",
  15591=>"100000000",
  15592=>"101100101",
  15593=>"000000000",
  15594=>"111000110",
  15595=>"000100100",
  15596=>"011000000",
  15597=>"000000000",
  15598=>"111000000",
  15599=>"000100000",
  15600=>"111111111",
  15601=>"111111111",
  15602=>"000000011",
  15603=>"000000011",
  15604=>"000000100",
  15605=>"000000000",
  15606=>"000000000",
  15607=>"000000000",
  15608=>"000000000",
  15609=>"111101000",
  15610=>"000000011",
  15611=>"111111111",
  15612=>"110111001",
  15613=>"001000000",
  15614=>"111000000",
  15615=>"000111010",
  15616=>"011000110",
  15617=>"111110100",
  15618=>"111111111",
  15619=>"000000000",
  15620=>"000000000",
  15621=>"000000000",
  15622=>"000000000",
  15623=>"010010111",
  15624=>"000000000",
  15625=>"100000100",
  15626=>"000000000",
  15627=>"011011000",
  15628=>"111101111",
  15629=>"100111111",
  15630=>"100111111",
  15631=>"000111000",
  15632=>"000000100",
  15633=>"000000010",
  15634=>"111111111",
  15635=>"000100000",
  15636=>"010000000",
  15637=>"000000110",
  15638=>"001000000",
  15639=>"111011010",
  15640=>"111111111",
  15641=>"111111110",
  15642=>"000000111",
  15643=>"111011111",
  15644=>"100001001",
  15645=>"111001000",
  15646=>"010011010",
  15647=>"001000111",
  15648=>"111011111",
  15649=>"111111111",
  15650=>"111111111",
  15651=>"001111111",
  15652=>"011000000",
  15653=>"111111111",
  15654=>"000000100",
  15655=>"010000000",
  15656=>"111111111",
  15657=>"011010000",
  15658=>"001011111",
  15659=>"111111011",
  15660=>"000000000",
  15661=>"101111111",
  15662=>"111111111",
  15663=>"000000000",
  15664=>"000001001",
  15665=>"000000000",
  15666=>"110000000",
  15667=>"000000000",
  15668=>"111111111",
  15669=>"000001001",
  15670=>"000000111",
  15671=>"111100111",
  15672=>"000000000",
  15673=>"000000000",
  15674=>"110000001",
  15675=>"001011011",
  15676=>"111111111",
  15677=>"000000110",
  15678=>"111111111",
  15679=>"010000000",
  15680=>"111111110",
  15681=>"111111111",
  15682=>"111111111",
  15683=>"111111111",
  15684=>"000000011",
  15685=>"001011110",
  15686=>"111000000",
  15687=>"110111111",
  15688=>"000000000",
  15689=>"000000000",
  15690=>"000010010",
  15691=>"101000100",
  15692=>"000000000",
  15693=>"000011111",
  15694=>"000000000",
  15695=>"011011001",
  15696=>"111111111",
  15697=>"001000110",
  15698=>"000000000",
  15699=>"010000000",
  15700=>"000000000",
  15701=>"000010001",
  15702=>"111111111",
  15703=>"100000000",
  15704=>"000011010",
  15705=>"111111111",
  15706=>"111110110",
  15707=>"101111111",
  15708=>"111111010",
  15709=>"011011011",
  15710=>"000000000",
  15711=>"000000000",
  15712=>"111111111",
  15713=>"111100000",
  15714=>"110110000",
  15715=>"110001111",
  15716=>"000000001",
  15717=>"000000000",
  15718=>"111111111",
  15719=>"001001000",
  15720=>"001001001",
  15721=>"001000000",
  15722=>"111111011",
  15723=>"111101111",
  15724=>"000010010",
  15725=>"111011000",
  15726=>"011001011",
  15727=>"111111110",
  15728=>"111100111",
  15729=>"000000000",
  15730=>"000000001",
  15731=>"111110111",
  15732=>"111111101",
  15733=>"000000000",
  15734=>"001101111",
  15735=>"001000011",
  15736=>"011011011",
  15737=>"111111110",
  15738=>"111000001",
  15739=>"111111110",
  15740=>"000000000",
  15741=>"111111000",
  15742=>"010010111",
  15743=>"000001011",
  15744=>"000100110",
  15745=>"100110000",
  15746=>"100100111",
  15747=>"100000000",
  15748=>"111111111",
  15749=>"101101111",
  15750=>"011000111",
  15751=>"111111111",
  15752=>"000000000",
  15753=>"110100000",
  15754=>"100000001",
  15755=>"000000000",
  15756=>"000000111",
  15757=>"111111111",
  15758=>"111011000",
  15759=>"111111111",
  15760=>"000000000",
  15761=>"111111111",
  15762=>"000000010",
  15763=>"111111110",
  15764=>"000000000",
  15765=>"000011000",
  15766=>"000000010",
  15767=>"001001111",
  15768=>"000111111",
  15769=>"000111111",
  15770=>"000000000",
  15771=>"011111111",
  15772=>"111111111",
  15773=>"111000000",
  15774=>"111111111",
  15775=>"111111111",
  15776=>"000000001",
  15777=>"110001001",
  15778=>"000001011",
  15779=>"000000000",
  15780=>"010000111",
  15781=>"111111111",
  15782=>"011000000",
  15783=>"000000000",
  15784=>"000111111",
  15785=>"000000011",
  15786=>"111111111",
  15787=>"001011111",
  15788=>"000000000",
  15789=>"000100100",
  15790=>"000001001",
  15791=>"111111110",
  15792=>"000000000",
  15793=>"111111111",
  15794=>"001000000",
  15795=>"000000001",
  15796=>"000000000",
  15797=>"000000000",
  15798=>"110110111",
  15799=>"000100100",
  15800=>"101101111",
  15801=>"000100111",
  15802=>"000000110",
  15803=>"010000000",
  15804=>"111000000",
  15805=>"000000000",
  15806=>"000000000",
  15807=>"110100000",
  15808=>"111000000",
  15809=>"110110000",
  15810=>"111111111",
  15811=>"011111111",
  15812=>"111001111",
  15813=>"111101111",
  15814=>"100100111",
  15815=>"111111011",
  15816=>"000000011",
  15817=>"110100100",
  15818=>"001111111",
  15819=>"111111111",
  15820=>"111111111",
  15821=>"001111000",
  15822=>"101001011",
  15823=>"111111111",
  15824=>"101000000",
  15825=>"010110011",
  15826=>"100011000",
  15827=>"111011011",
  15828=>"000000000",
  15829=>"000000000",
  15830=>"110100111",
  15831=>"000000000",
  15832=>"111111111",
  15833=>"111110000",
  15834=>"010000110",
  15835=>"110110000",
  15836=>"000110010",
  15837=>"011111111",
  15838=>"111101011",
  15839=>"110110111",
  15840=>"101100100",
  15841=>"100000000",
  15842=>"000000000",
  15843=>"000001000",
  15844=>"010100100",
  15845=>"001011011",
  15846=>"111111111",
  15847=>"111011111",
  15848=>"111011010",
  15849=>"000000111",
  15850=>"000000100",
  15851=>"111111110",
  15852=>"111010010",
  15853=>"100000000",
  15854=>"000000000",
  15855=>"111111111",
  15856=>"100111111",
  15857=>"111010000",
  15858=>"111010110",
  15859=>"111111011",
  15860=>"111011111",
  15861=>"111111111",
  15862=>"000000000",
  15863=>"001000100",
  15864=>"000000000",
  15865=>"011000011",
  15866=>"010111010",
  15867=>"111010000",
  15868=>"000000111",
  15869=>"111111100",
  15870=>"000100110",
  15871=>"111111111",
  15872=>"001111001",
  15873=>"010000001",
  15874=>"110110111",
  15875=>"000110111",
  15876=>"100000110",
  15877=>"010011011",
  15878=>"111111111",
  15879=>"000000000",
  15880=>"000100111",
  15881=>"111111101",
  15882=>"000000000",
  15883=>"000110111",
  15884=>"111111101",
  15885=>"000000010",
  15886=>"001100000",
  15887=>"000000000",
  15888=>"000000000",
  15889=>"000000000",
  15890=>"100000000",
  15891=>"001000000",
  15892=>"111111111",
  15893=>"000110010",
  15894=>"100100110",
  15895=>"001000000",
  15896=>"111111110",
  15897=>"000000000",
  15898=>"010110111",
  15899=>"101100000",
  15900=>"111111111",
  15901=>"111110110",
  15902=>"111010011",
  15903=>"111000000",
  15904=>"000101001",
  15905=>"111111111",
  15906=>"011001000",
  15907=>"111111111",
  15908=>"000000000",
  15909=>"111111101",
  15910=>"011001111",
  15911=>"000000100",
  15912=>"111111111",
  15913=>"000010000",
  15914=>"111111100",
  15915=>"000000000",
  15916=>"000000001",
  15917=>"111111011",
  15918=>"111111111",
  15919=>"110000001",
  15920=>"000000110",
  15921=>"000000000",
  15922=>"001100100",
  15923=>"111111111",
  15924=>"111110110",
  15925=>"011110000",
  15926=>"000000000",
  15927=>"111111111",
  15928=>"100100010",
  15929=>"111110100",
  15930=>"011000000",
  15931=>"010000000",
  15932=>"111111011",
  15933=>"110000000",
  15934=>"101001000",
  15935=>"111111111",
  15936=>"001001011",
  15937=>"110100110",
  15938=>"000110110",
  15939=>"001000000",
  15940=>"100000000",
  15941=>"001001011",
  15942=>"111111111",
  15943=>"111111111",
  15944=>"001111011",
  15945=>"110101111",
  15946=>"000000000",
  15947=>"010000000",
  15948=>"000000011",
  15949=>"000000000",
  15950=>"010000001",
  15951=>"001001000",
  15952=>"000000100",
  15953=>"111111111",
  15954=>"111111111",
  15955=>"111110100",
  15956=>"111111111",
  15957=>"010110110",
  15958=>"111111111",
  15959=>"000101111",
  15960=>"111000000",
  15961=>"011111111",
  15962=>"011110111",
  15963=>"000000000",
  15964=>"111111111",
  15965=>"111111111",
  15966=>"010000000",
  15967=>"111111000",
  15968=>"000000111",
  15969=>"111000000",
  15970=>"111111010",
  15971=>"111111111",
  15972=>"111000000",
  15973=>"111111011",
  15974=>"011000000",
  15975=>"111111111",
  15976=>"110010000",
  15977=>"100111111",
  15978=>"001000000",
  15979=>"000000010",
  15980=>"111110110",
  15981=>"000000000",
  15982=>"111111111",
  15983=>"011011011",
  15984=>"001001011",
  15985=>"000000000",
  15986=>"000000000",
  15987=>"111111000",
  15988=>"000000000",
  15989=>"111011001",
  15990=>"000000000",
  15991=>"111000000",
  15992=>"000000000",
  15993=>"101101111",
  15994=>"100100100",
  15995=>"111111111",
  15996=>"000000000",
  15997=>"000000000",
  15998=>"111111111",
  15999=>"000000000",
  16000=>"111111111",
  16001=>"000000000",
  16002=>"111011111",
  16003=>"111111111",
  16004=>"000000001",
  16005=>"000000011",
  16006=>"111111111",
  16007=>"100001000",
  16008=>"000000000",
  16009=>"110011001",
  16010=>"111111100",
  16011=>"111110110",
  16012=>"111010110",
  16013=>"000000000",
  16014=>"111111111",
  16015=>"110100000",
  16016=>"000000000",
  16017=>"001110100",
  16018=>"000000011",
  16019=>"011111111",
  16020=>"111111111",
  16021=>"000011111",
  16022=>"000001001",
  16023=>"111011011",
  16024=>"111111111",
  16025=>"000000000",
  16026=>"000000000",
  16027=>"111110011",
  16028=>"001001000",
  16029=>"011111111",
  16030=>"001001001",
  16031=>"000000000",
  16032=>"010000000",
  16033=>"111111110",
  16034=>"010010000",
  16035=>"010001000",
  16036=>"000101011",
  16037=>"111111110",
  16038=>"100000000",
  16039=>"001011011",
  16040=>"011011011",
  16041=>"000000000",
  16042=>"000001001",
  16043=>"000000000",
  16044=>"011001000",
  16045=>"111111110",
  16046=>"001000000",
  16047=>"011111000",
  16048=>"010111011",
  16049=>"001001001",
  16050=>"010011011",
  16051=>"100000100",
  16052=>"000000100",
  16053=>"000000000",
  16054=>"001011111",
  16055=>"111110110",
  16056=>"011011011",
  16057=>"111111111",
  16058=>"100101101",
  16059=>"100110111",
  16060=>"111111111",
  16061=>"001001111",
  16062=>"010000000",
  16063=>"000100000",
  16064=>"000111110",
  16065=>"111111010",
  16066=>"000000000",
  16067=>"011010000",
  16068=>"000000000",
  16069=>"111111111",
  16070=>"100001101",
  16071=>"100100110",
  16072=>"000110111",
  16073=>"000111111",
  16074=>"100100110",
  16075=>"100110110",
  16076=>"001001000",
  16077=>"001011000",
  16078=>"111111111",
  16079=>"111111111",
  16080=>"010011111",
  16081=>"000011111",
  16082=>"010000000",
  16083=>"000000000",
  16084=>"111111111",
  16085=>"000001001",
  16086=>"110111111",
  16087=>"110000000",
  16088=>"000101001",
  16089=>"001000000",
  16090=>"000000000",
  16091=>"111110001",
  16092=>"111111111",
  16093=>"111111111",
  16094=>"110000000",
  16095=>"011000000",
  16096=>"000000010",
  16097=>"110110010",
  16098=>"011000000",
  16099=>"111011010",
  16100=>"111111111",
  16101=>"111111011",
  16102=>"100000000",
  16103=>"111100000",
  16104=>"000000000",
  16105=>"100101111",
  16106=>"001000000",
  16107=>"000000000",
  16108=>"111001000",
  16109=>"111111111",
  16110=>"111110101",
  16111=>"000111000",
  16112=>"011000000",
  16113=>"111001000",
  16114=>"000000000",
  16115=>"111111110",
  16116=>"000010110",
  16117=>"110010010",
  16118=>"110000000",
  16119=>"000000011",
  16120=>"111110110",
  16121=>"111001111",
  16122=>"111111111",
  16123=>"110110111",
  16124=>"010011000",
  16125=>"000000000",
  16126=>"000000100",
  16127=>"000000000",
  16128=>"100001101",
  16129=>"010011000",
  16130=>"111111111",
  16131=>"100100100",
  16132=>"000000000",
  16133=>"111111101",
  16134=>"000000110",
  16135=>"011100111",
  16136=>"000000000",
  16137=>"000000000",
  16138=>"010111111",
  16139=>"111100000",
  16140=>"110110110",
  16141=>"111111110",
  16142=>"111111111",
  16143=>"111111111",
  16144=>"111111111",
  16145=>"111001000",
  16146=>"000000000",
  16147=>"010010001",
  16148=>"000000000",
  16149=>"111111111",
  16150=>"101110000",
  16151=>"000100111",
  16152=>"111101000",
  16153=>"001000000",
  16154=>"000100000",
  16155=>"010010000",
  16156=>"010111111",
  16157=>"111010110",
  16158=>"111111011",
  16159=>"111111111",
  16160=>"111111001",
  16161=>"000110111",
  16162=>"111111011",
  16163=>"010000000",
  16164=>"001111111",
  16165=>"111111111",
  16166=>"001011011",
  16167=>"001001001",
  16168=>"011011111",
  16169=>"000000000",
  16170=>"111011001",
  16171=>"000000000",
  16172=>"111110111",
  16173=>"100100000",
  16174=>"111111000",
  16175=>"011101000",
  16176=>"010110010",
  16177=>"111111111",
  16178=>"000011001",
  16179=>"100111111",
  16180=>"110111111",
  16181=>"000011011",
  16182=>"010000000",
  16183=>"111111000",
  16184=>"000110111",
  16185=>"011011111",
  16186=>"100100100",
  16187=>"001010000",
  16188=>"111100111",
  16189=>"000000000",
  16190=>"101101100",
  16191=>"000100000",
  16192=>"111000000",
  16193=>"000000000",
  16194=>"011011010",
  16195=>"100100111",
  16196=>"011011111",
  16197=>"011111110",
  16198=>"000001000",
  16199=>"111111000",
  16200=>"100100000",
  16201=>"111111111",
  16202=>"000000100",
  16203=>"100100100",
  16204=>"111011001",
  16205=>"101111111",
  16206=>"010000000",
  16207=>"000100000",
  16208=>"111110101",
  16209=>"000000000",
  16210=>"111110110",
  16211=>"000000000",
  16212=>"000000000",
  16213=>"111111011",
  16214=>"111111011",
  16215=>"111110110",
  16216=>"011111111",
  16217=>"010011010",
  16218=>"111111111",
  16219=>"000000000",
  16220=>"000000000",
  16221=>"000000000",
  16222=>"000000111",
  16223=>"000000000",
  16224=>"001000010",
  16225=>"111111000",
  16226=>"111100100",
  16227=>"111111111",
  16228=>"000000000",
  16229=>"111111111",
  16230=>"011011111",
  16231=>"010000000",
  16232=>"001000000",
  16233=>"111111110",
  16234=>"111111111",
  16235=>"010010110",
  16236=>"110100100",
  16237=>"100001000",
  16238=>"000000000",
  16239=>"111001111",
  16240=>"001000001",
  16241=>"110111011",
  16242=>"100000001",
  16243=>"111100110",
  16244=>"000000000",
  16245=>"011000000",
  16246=>"011100100",
  16247=>"111110010",
  16248=>"111001000",
  16249=>"111111111",
  16250=>"111111111",
  16251=>"110111111",
  16252=>"000000111",
  16253=>"001000000",
  16254=>"100011001",
  16255=>"000000000",
  16256=>"010010111",
  16257=>"000000000",
  16258=>"000000100",
  16259=>"000000001",
  16260=>"000000001",
  16261=>"010110110",
  16262=>"000101000",
  16263=>"100111111",
  16264=>"100000000",
  16265=>"000000000",
  16266=>"001001011",
  16267=>"100100110",
  16268=>"111100111",
  16269=>"011110000",
  16270=>"111000000",
  16271=>"111111111",
  16272=>"100000000",
  16273=>"111111111",
  16274=>"000000001",
  16275=>"111001111",
  16276=>"011000000",
  16277=>"100100100",
  16278=>"000000000",
  16279=>"000010110",
  16280=>"110111111",
  16281=>"001011111",
  16282=>"011111010",
  16283=>"000000000",
  16284=>"000000000",
  16285=>"000000100",
  16286=>"111111110",
  16287=>"110111111",
  16288=>"000000000",
  16289=>"000000000",
  16290=>"111110111",
  16291=>"100000000",
  16292=>"111111000",
  16293=>"100110011",
  16294=>"111111111",
  16295=>"000000000",
  16296=>"010010111",
  16297=>"010000110",
  16298=>"110000000",
  16299=>"111111000",
  16300=>"010111010",
  16301=>"000000000",
  16302=>"001111111",
  16303=>"111111110",
  16304=>"000000000",
  16305=>"111111111",
  16306=>"001000110",
  16307=>"010000000",
  16308=>"011010000",
  16309=>"011000000",
  16310=>"110000000",
  16311=>"111000100",
  16312=>"110000000",
  16313=>"000000000",
  16314=>"001001100",
  16315=>"000000000",
  16316=>"000011111",
  16317=>"000001001",
  16318=>"110001000",
  16319=>"000000000",
  16320=>"111000000",
  16321=>"000000000",
  16322=>"000000000",
  16323=>"111111111",
  16324=>"111111111",
  16325=>"111000010",
  16326=>"000100000",
  16327=>"110111111",
  16328=>"111001001",
  16329=>"111000110",
  16330=>"000000000",
  16331=>"011000000",
  16332=>"111111111",
  16333=>"111111111",
  16334=>"000000000",
  16335=>"110000011",
  16336=>"111101111",
  16337=>"000000100",
  16338=>"000000000",
  16339=>"000000000",
  16340=>"111110001",
  16341=>"000010000",
  16342=>"001000001",
  16343=>"001000000",
  16344=>"010110000",
  16345=>"011001000",
  16346=>"111001101",
  16347=>"111000000",
  16348=>"000111111",
  16349=>"000000110",
  16350=>"111011000",
  16351=>"110111111",
  16352=>"010001000",
  16353=>"011111101",
  16354=>"110111111",
  16355=>"000000000",
  16356=>"000000000",
  16357=>"000000000",
  16358=>"111111000",
  16359=>"111111111",
  16360=>"111111111",
  16361=>"000010000",
  16362=>"000001001",
  16363=>"001000000",
  16364=>"000001001",
  16365=>"001001011",
  16366=>"100111001",
  16367=>"111001000",
  16368=>"101100000",
  16369=>"010011000",
  16370=>"111111011",
  16371=>"000110110",
  16372=>"111111010",
  16373=>"000000000",
  16374=>"010000000",
  16375=>"000000000",
  16376=>"011110100",
  16377=>"000110110",
  16378=>"000011111",
  16379=>"110111111",
  16380=>"010100000",
  16381=>"011001011",
  16382=>"010111011",
  16383=>"000011011",
  16384=>"001000000",
  16385=>"000000000",
  16386=>"111000001",
  16387=>"100110111",
  16388=>"000000000",
  16389=>"000110000",
  16390=>"001011011",
  16391=>"101000111",
  16392=>"111111000",
  16393=>"111111111",
  16394=>"000000110",
  16395=>"011111000",
  16396=>"000000100",
  16397=>"000000111",
  16398=>"100100111",
  16399=>"000000101",
  16400=>"000001111",
  16401=>"011111111",
  16402=>"110111111",
  16403=>"111000000",
  16404=>"000000000",
  16405=>"111111111",
  16406=>"100101111",
  16407=>"100110111",
  16408=>"111110111",
  16409=>"111101101",
  16410=>"000100111",
  16411=>"001000000",
  16412=>"000100000",
  16413=>"111111001",
  16414=>"111111111",
  16415=>"100011111",
  16416=>"100111111",
  16417=>"111111111",
  16418=>"111111110",
  16419=>"111110110",
  16420=>"000000000",
  16421=>"000000001",
  16422=>"111111101",
  16423=>"100101111",
  16424=>"110111111",
  16425=>"111111000",
  16426=>"000000000",
  16427=>"111010011",
  16428=>"100000001",
  16429=>"111111100",
  16430=>"000001111",
  16431=>"111011001",
  16432=>"110111110",
  16433=>"000001001",
  16434=>"111111011",
  16435=>"111011011",
  16436=>"000001110",
  16437=>"000001000",
  16438=>"111111111",
  16439=>"110110000",
  16440=>"001011000",
  16441=>"110000001",
  16442=>"011111011",
  16443=>"110100110",
  16444=>"100100111",
  16445=>"000000000",
  16446=>"000000100",
  16447=>"011111000",
  16448=>"000000011",
  16449=>"110111111",
  16450=>"011111101",
  16451=>"110110101",
  16452=>"110111011",
  16453=>"011011001",
  16454=>"111000000",
  16455=>"111111111",
  16456=>"111111000",
  16457=>"000001011",
  16458=>"111111010",
  16459=>"111001001",
  16460=>"000000000",
  16461=>"011011001",
  16462=>"110111111",
  16463=>"111101000",
  16464=>"001001001",
  16465=>"110110000",
  16466=>"111111010",
  16467=>"100000100",
  16468=>"000000000",
  16469=>"111111101",
  16470=>"100101111",
  16471=>"100101111",
  16472=>"000000000",
  16473=>"111000000",
  16474=>"000000000",
  16475=>"110110110",
  16476=>"000000000",
  16477=>"111111000",
  16478=>"001001111",
  16479=>"000100000",
  16480=>"111111111",
  16481=>"111111100",
  16482=>"000000000",
  16483=>"000111111",
  16484=>"111111010",
  16485=>"111111111",
  16486=>"111110000",
  16487=>"011001000",
  16488=>"111111000",
  16489=>"000000000",
  16490=>"100000000",
  16491=>"010010000",
  16492=>"000000110",
  16493=>"111111111",
  16494=>"000000100",
  16495=>"000010000",
  16496=>"000000111",
  16497=>"000000101",
  16498=>"110111111",
  16499=>"111111111",
  16500=>"000000011",
  16501=>"111111010",
  16502=>"000000000",
  16503=>"000000000",
  16504=>"111111111",
  16505=>"000000000",
  16506=>"001000000",
  16507=>"000000000",
  16508=>"100100100",
  16509=>"000000011",
  16510=>"000000000",
  16511=>"001011111",
  16512=>"000000000",
  16513=>"111111101",
  16514=>"011111101",
  16515=>"110101111",
  16516=>"111111111",
  16517=>"111000110",
  16518=>"100100000",
  16519=>"000000011",
  16520=>"000000000",
  16521=>"111000000",
  16522=>"010111111",
  16523=>"111011000",
  16524=>"111111111",
  16525=>"101101111",
  16526=>"001000111",
  16527=>"001000000",
  16528=>"100000000",
  16529=>"000000100",
  16530=>"000001000",
  16531=>"001011111",
  16532=>"111011001",
  16533=>"000100100",
  16534=>"111111010",
  16535=>"100100100",
  16536=>"001001101",
  16537=>"000100111",
  16538=>"111011010",
  16539=>"011000000",
  16540=>"010010011",
  16541=>"000000000",
  16542=>"110111110",
  16543=>"011000110",
  16544=>"011000000",
  16545=>"000000000",
  16546=>"011000000",
  16547=>"000010011",
  16548=>"100011000",
  16549=>"011010000",
  16550=>"100100001",
  16551=>"000001111",
  16552=>"111111111",
  16553=>"101111101",
  16554=>"011000000",
  16555=>"011111111",
  16556=>"111111111",
  16557=>"111100100",
  16558=>"100000000",
  16559=>"110111110",
  16560=>"111111111",
  16561=>"000011011",
  16562=>"110111010",
  16563=>"000000000",
  16564=>"100000000",
  16565=>"000000001",
  16566=>"000000101",
  16567=>"001111111",
  16568=>"111111000",
  16569=>"111111111",
  16570=>"000100000",
  16571=>"000000111",
  16572=>"100111111",
  16573=>"100000001",
  16574=>"111000000",
  16575=>"001000000",
  16576=>"000000100",
  16577=>"111000000",
  16578=>"001100101",
  16579=>"000000001",
  16580=>"010111011",
  16581=>"000001111",
  16582=>"110111110",
  16583=>"000100100",
  16584=>"111111011",
  16585=>"001110111",
  16586=>"000000000",
  16587=>"000000000",
  16588=>"101001101",
  16589=>"000000000",
  16590=>"111111111",
  16591=>"000000011",
  16592=>"010011010",
  16593=>"000110110",
  16594=>"000000011",
  16595=>"011001001",
  16596=>"000000000",
  16597=>"111110100",
  16598=>"000000000",
  16599=>"111110100",
  16600=>"111111111",
  16601=>"000000100",
  16602=>"011011111",
  16603=>"111111111",
  16604=>"000000000",
  16605=>"111111111",
  16606=>"111111111",
  16607=>"111111101",
  16608=>"000001111",
  16609=>"110111111",
  16610=>"110100000",
  16611=>"110111000",
  16612=>"000000111",
  16613=>"000010111",
  16614=>"111111110",
  16615=>"111111110",
  16616=>"111111010",
  16617=>"000101001",
  16618=>"111111111",
  16619=>"111111101",
  16620=>"000000000",
  16621=>"000100000",
  16622=>"000000111",
  16623=>"011001111",
  16624=>"001101111",
  16625=>"001111111",
  16626=>"000110111",
  16627=>"100000001",
  16628=>"001001011",
  16629=>"001011011",
  16630=>"000000111",
  16631=>"101000000",
  16632=>"110011000",
  16633=>"000000001",
  16634=>"111101111",
  16635=>"111111111",
  16636=>"000111110",
  16637=>"000111110",
  16638=>"011000000",
  16639=>"111111110",
  16640=>"111111011",
  16641=>"111111111",
  16642=>"001111111",
  16643=>"000000001",
  16644=>"000000100",
  16645=>"011011111",
  16646=>"100000100",
  16647=>"000000101",
  16648=>"000000000",
  16649=>"000000001",
  16650=>"000000000",
  16651=>"001000101",
  16652=>"000000000",
  16653=>"000000000",
  16654=>"000000101",
  16655=>"111111000",
  16656=>"000101101",
  16657=>"000100111",
  16658=>"101111111",
  16659=>"110111111",
  16660=>"010111111",
  16661=>"011111111",
  16662=>"110100100",
  16663=>"010110110",
  16664=>"111111111",
  16665=>"000000011",
  16666=>"110000010",
  16667=>"111111111",
  16668=>"110111100",
  16669=>"110010001",
  16670=>"000000000",
  16671=>"010111111",
  16672=>"000011110",
  16673=>"111110111",
  16674=>"111111000",
  16675=>"111111110",
  16676=>"111011011",
  16677=>"111111111",
  16678=>"010000000",
  16679=>"111111000",
  16680=>"000000000",
  16681=>"111111010",
  16682=>"111111010",
  16683=>"000000000",
  16684=>"011111110",
  16685=>"100111110",
  16686=>"111011111",
  16687=>"000000101",
  16688=>"010000111",
  16689=>"000000000",
  16690=>"111111010",
  16691=>"000000000",
  16692=>"000000000",
  16693=>"000000000",
  16694=>"011000000",
  16695=>"000111111",
  16696=>"111111010",
  16697=>"001000000",
  16698=>"000000000",
  16699=>"011001000",
  16700=>"111111111",
  16701=>"011001111",
  16702=>"000000001",
  16703=>"111111111",
  16704=>"001001001",
  16705=>"110101111",
  16706=>"000000001",
  16707=>"111111111",
  16708=>"000000111",
  16709=>"111111111",
  16710=>"010010001",
  16711=>"111111111",
  16712=>"111101111",
  16713=>"000000011",
  16714=>"001011001",
  16715=>"000000000",
  16716=>"111000000",
  16717=>"000001111",
  16718=>"100100111",
  16719=>"000100100",
  16720=>"100100000",
  16721=>"100001011",
  16722=>"000111111",
  16723=>"111100111",
  16724=>"011000000",
  16725=>"011011001",
  16726=>"100000100",
  16727=>"111110111",
  16728=>"111111111",
  16729=>"000000101",
  16730=>"110111111",
  16731=>"010111111",
  16732=>"110100111",
  16733=>"000000000",
  16734=>"111111111",
  16735=>"111111010",
  16736=>"000000100",
  16737=>"000000000",
  16738=>"111111111",
  16739=>"111101111",
  16740=>"000111111",
  16741=>"100000000",
  16742=>"111000000",
  16743=>"001001011",
  16744=>"001000000",
  16745=>"110000000",
  16746=>"000000111",
  16747=>"011001111",
  16748=>"111111000",
  16749=>"100100000",
  16750=>"001011011",
  16751=>"011011111",
  16752=>"001000000",
  16753=>"111111111",
  16754=>"000000111",
  16755=>"111001000",
  16756=>"000000000",
  16757=>"011001011",
  16758=>"101000001",
  16759=>"000000000",
  16760=>"001001111",
  16761=>"111001001",
  16762=>"111111111",
  16763=>"000000000",
  16764=>"011000000",
  16765=>"111111001",
  16766=>"100100111",
  16767=>"101111111",
  16768=>"100100101",
  16769=>"111111000",
  16770=>"100000011",
  16771=>"011111111",
  16772=>"001001000",
  16773=>"110111111",
  16774=>"111111111",
  16775=>"100110111",
  16776=>"000000000",
  16777=>"111111000",
  16778=>"111111110",
  16779=>"100111110",
  16780=>"100101111",
  16781=>"000100000",
  16782=>"111111110",
  16783=>"110111111",
  16784=>"000000000",
  16785=>"100101111",
  16786=>"110110011",
  16787=>"001100111",
  16788=>"000000110",
  16789=>"010110010",
  16790=>"111111110",
  16791=>"111011000",
  16792=>"000000111",
  16793=>"001001000",
  16794=>"001011111",
  16795=>"100000101",
  16796=>"000000000",
  16797=>"000000000",
  16798=>"111100100",
  16799=>"000000000",
  16800=>"111000000",
  16801=>"111111111",
  16802=>"111100100",
  16803=>"111111000",
  16804=>"111111111",
  16805=>"111100010",
  16806=>"000000000",
  16807=>"111111000",
  16808=>"000010000",
  16809=>"000000111",
  16810=>"110111111",
  16811=>"000000000",
  16812=>"000000111",
  16813=>"101101001",
  16814=>"001000111",
  16815=>"100100000",
  16816=>"000000111",
  16817=>"001111000",
  16818=>"000000000",
  16819=>"000000000",
  16820=>"011000000",
  16821=>"000000000",
  16822=>"001100100",
  16823=>"111111111",
  16824=>"001000001",
  16825=>"000111110",
  16826=>"011000001",
  16827=>"110111111",
  16828=>"001011111",
  16829=>"000000000",
  16830=>"111111111",
  16831=>"111100101",
  16832=>"111111000",
  16833=>"111111010",
  16834=>"000001111",
  16835=>"110000000",
  16836=>"111011111",
  16837=>"000000100",
  16838=>"100000000",
  16839=>"000100000",
  16840=>"111100011",
  16841=>"000000110",
  16842=>"111101111",
  16843=>"000111010",
  16844=>"000000111",
  16845=>"111111111",
  16846=>"000000000",
  16847=>"101101100",
  16848=>"101111111",
  16849=>"000000000",
  16850=>"111111111",
  16851=>"000000111",
  16852=>"111111111",
  16853=>"000000011",
  16854=>"000000010",
  16855=>"010110000",
  16856=>"110100101",
  16857=>"111101010",
  16858=>"100011111",
  16859=>"100111111",
  16860=>"011111111",
  16861=>"111000000",
  16862=>"100110111",
  16863=>"111111111",
  16864=>"111001001",
  16865=>"001001001",
  16866=>"000000101",
  16867=>"000000000",
  16868=>"111111111",
  16869=>"111111101",
  16870=>"000100100",
  16871=>"011111011",
  16872=>"111011111",
  16873=>"000000000",
  16874=>"000100110",
  16875=>"111111000",
  16876=>"110000100",
  16877=>"011011000",
  16878=>"111111111",
  16879=>"000000001",
  16880=>"110011001",
  16881=>"010111100",
  16882=>"111111001",
  16883=>"111001000",
  16884=>"111111110",
  16885=>"000100110",
  16886=>"111111110",
  16887=>"000000000",
  16888=>"100111110",
  16889=>"000000000",
  16890=>"011111011",
  16891=>"111000000",
  16892=>"001111100",
  16893=>"111111111",
  16894=>"000000000",
  16895=>"000100111",
  16896=>"110000100",
  16897=>"001110111",
  16898=>"111111111",
  16899=>"111111101",
  16900=>"011111111",
  16901=>"110100111",
  16902=>"000000000",
  16903=>"000000000",
  16904=>"000111100",
  16905=>"000001001",
  16906=>"111111110",
  16907=>"011011111",
  16908=>"000110010",
  16909=>"111111111",
  16910=>"110010000",
  16911=>"000000000",
  16912=>"111111000",
  16913=>"010110110",
  16914=>"000110111",
  16915=>"000000111",
  16916=>"110010000",
  16917=>"100000111",
  16918=>"000000000",
  16919=>"001001011",
  16920=>"110100111",
  16921=>"011110100",
  16922=>"111001000",
  16923=>"000110011",
  16924=>"000000001",
  16925=>"111110000",
  16926=>"111001000",
  16927=>"001011000",
  16928=>"000010010",
  16929=>"111111111",
  16930=>"111111110",
  16931=>"000001101",
  16932=>"111100110",
  16933=>"100110110",
  16934=>"000000000",
  16935=>"100000000",
  16936=>"111001000",
  16937=>"000101000",
  16938=>"000000110",
  16939=>"000000000",
  16940=>"110111111",
  16941=>"111011111",
  16942=>"110111111",
  16943=>"000100111",
  16944=>"111111011",
  16945=>"000000000",
  16946=>"010000100",
  16947=>"111011111",
  16948=>"100100000",
  16949=>"000100111",
  16950=>"000000011",
  16951=>"011110110",
  16952=>"111111111",
  16953=>"101100000",
  16954=>"111101101",
  16955=>"000001011",
  16956=>"111001000",
  16957=>"111111110",
  16958=>"000000001",
  16959=>"000000001",
  16960=>"100011000",
  16961=>"111111000",
  16962=>"001000100",
  16963=>"100000000",
  16964=>"000000110",
  16965=>"000000010",
  16966=>"111111111",
  16967=>"111111111",
  16968=>"100110110",
  16969=>"000000000",
  16970=>"000000000",
  16971=>"011011111",
  16972=>"111000000",
  16973=>"000100000",
  16974=>"000001101",
  16975=>"111001001",
  16976=>"000110110",
  16977=>"000000000",
  16978=>"110111111",
  16979=>"100001100",
  16980=>"000111111",
  16981=>"111111000",
  16982=>"111111111",
  16983=>"000000000",
  16984=>"001101001",
  16985=>"000000100",
  16986=>"100111111",
  16987=>"000001001",
  16988=>"111111111",
  16989=>"011001001",
  16990=>"111111101",
  16991=>"001000000",
  16992=>"000000110",
  16993=>"001011000",
  16994=>"111111001",
  16995=>"000000000",
  16996=>"100111111",
  16997=>"000010000",
  16998=>"100100111",
  16999=>"111011001",
  17000=>"111111111",
  17001=>"111100000",
  17002=>"110110110",
  17003=>"111011111",
  17004=>"000000000",
  17005=>"000000000",
  17006=>"000000110",
  17007=>"111111000",
  17008=>"000000000",
  17009=>"110110101",
  17010=>"100100101",
  17011=>"111110000",
  17012=>"101111111",
  17013=>"001000000",
  17014=>"001000000",
  17015=>"100111111",
  17016=>"000000000",
  17017=>"100100011",
  17018=>"111111101",
  17019=>"111100100",
  17020=>"111111101",
  17021=>"010111110",
  17022=>"000000001",
  17023=>"000000000",
  17024=>"000010110",
  17025=>"111100100",
  17026=>"000000000",
  17027=>"100000000",
  17028=>"001101111",
  17029=>"110111111",
  17030=>"110000000",
  17031=>"001111111",
  17032=>"001111111",
  17033=>"001111011",
  17034=>"111111111",
  17035=>"000110110",
  17036=>"100000111",
  17037=>"100101111",
  17038=>"111111110",
  17039=>"110011000",
  17040=>"000000000",
  17041=>"010010000",
  17042=>"001000001",
  17043=>"100000000",
  17044=>"001000000",
  17045=>"111111101",
  17046=>"111110111",
  17047=>"111101111",
  17048=>"111110111",
  17049=>"000000000",
  17050=>"000000001",
  17051=>"111111111",
  17052=>"000110100",
  17053=>"111100000",
  17054=>"011111110",
  17055=>"000000011",
  17056=>"011011100",
  17057=>"110101111",
  17058=>"111000000",
  17059=>"111111111",
  17060=>"000000000",
  17061=>"101111111",
  17062=>"000000000",
  17063=>"000011011",
  17064=>"000100111",
  17065=>"000000000",
  17066=>"000000000",
  17067=>"111000111",
  17068=>"111111011",
  17069=>"100000000",
  17070=>"110111111",
  17071=>"110010000",
  17072=>"000100110",
  17073=>"100001101",
  17074=>"001111111",
  17075=>"111111000",
  17076=>"000001011",
  17077=>"000000101",
  17078=>"000000100",
  17079=>"000110110",
  17080=>"111111011",
  17081=>"000000000",
  17082=>"000000000",
  17083=>"000110000",
  17084=>"001001001",
  17085=>"110110010",
  17086=>"000000101",
  17087=>"011000000",
  17088=>"001011111",
  17089=>"000011011",
  17090=>"000000000",
  17091=>"000000000",
  17092=>"000000000",
  17093=>"000000000",
  17094=>"010010111",
  17095=>"100100110",
  17096=>"000000000",
  17097=>"111111000",
  17098=>"001111000",
  17099=>"000000000",
  17100=>"111111001",
  17101=>"101001001",
  17102=>"000011100",
  17103=>"100110110",
  17104=>"111111111",
  17105=>"111100110",
  17106=>"011111111",
  17107=>"110110100",
  17108=>"101100111",
  17109=>"110110000",
  17110=>"100100111",
  17111=>"000011000",
  17112=>"111111111",
  17113=>"100111111",
  17114=>"001011001",
  17115=>"111111111",
  17116=>"110010010",
  17117=>"001001001",
  17118=>"011111111",
  17119=>"111111110",
  17120=>"111111111",
  17121=>"000000000",
  17122=>"100000000",
  17123=>"111110111",
  17124=>"000011111",
  17125=>"000000110",
  17126=>"001001101",
  17127=>"000000001",
  17128=>"000000100",
  17129=>"111111111",
  17130=>"110110000",
  17131=>"001000000",
  17132=>"000001111",
  17133=>"111101111",
  17134=>"111000001",
  17135=>"000000000",
  17136=>"111110111",
  17137=>"000000111",
  17138=>"111000111",
  17139=>"110110111",
  17140=>"000111100",
  17141=>"000000000",
  17142=>"110100100",
  17143=>"101000000",
  17144=>"000110111",
  17145=>"111111111",
  17146=>"110100000",
  17147=>"111111111",
  17148=>"110110110",
  17149=>"111100100",
  17150=>"100101001",
  17151=>"000000000",
  17152=>"000000000",
  17153=>"010000000",
  17154=>"000000000",
  17155=>"110110111",
  17156=>"000000100",
  17157=>"111111111",
  17158=>"000000111",
  17159=>"011000100",
  17160=>"111111101",
  17161=>"000111111",
  17162=>"111111111",
  17163=>"111110001",
  17164=>"000000000",
  17165=>"000000000",
  17166=>"100111111",
  17167=>"000000111",
  17168=>"001100101",
  17169=>"110000000",
  17170=>"001000000",
  17171=>"001000001",
  17172=>"000110101",
  17173=>"000000100",
  17174=>"000000000",
  17175=>"001011111",
  17176=>"111111011",
  17177=>"000110111",
  17178=>"000110000",
  17179=>"011111111",
  17180=>"011011001",
  17181=>"000000101",
  17182=>"110111110",
  17183=>"111110111",
  17184=>"100000001",
  17185=>"000100100",
  17186=>"000000001",
  17187=>"101011000",
  17188=>"000011011",
  17189=>"111000110",
  17190=>"111111111",
  17191=>"110000110",
  17192=>"000101001",
  17193=>"111110010",
  17194=>"101100100",
  17195=>"000001011",
  17196=>"011000000",
  17197=>"000110111",
  17198=>"000101111",
  17199=>"010111111",
  17200=>"111111111",
  17201=>"000000110",
  17202=>"001010111",
  17203=>"001001000",
  17204=>"111111000",
  17205=>"000000110",
  17206=>"000000001",
  17207=>"011000000",
  17208=>"100000000",
  17209=>"101000000",
  17210=>"000000000",
  17211=>"000000000",
  17212=>"111101100",
  17213=>"111111001",
  17214=>"111101001",
  17215=>"111000000",
  17216=>"111011111",
  17217=>"011111110",
  17218=>"011111111",
  17219=>"000000000",
  17220=>"111101001",
  17221=>"000000000",
  17222=>"000110011",
  17223=>"011111111",
  17224=>"000000000",
  17225=>"111000000",
  17226=>"001110110",
  17227=>"000000000",
  17228=>"111111111",
  17229=>"101000000",
  17230=>"111111111",
  17231=>"011111101",
  17232=>"110110111",
  17233=>"111111111",
  17234=>"000000000",
  17235=>"100100110",
  17236=>"111111111",
  17237=>"111111111",
  17238=>"000000111",
  17239=>"111000100",
  17240=>"011000111",
  17241=>"111111111",
  17242=>"100000000",
  17243=>"111110111",
  17244=>"011110000",
  17245=>"111111111",
  17246=>"000000000",
  17247=>"000100110",
  17248=>"000111111",
  17249=>"000000000",
  17250=>"011010011",
  17251=>"111111111",
  17252=>"000000000",
  17253=>"000000000",
  17254=>"101000000",
  17255=>"000010000",
  17256=>"000010001",
  17257=>"011000000",
  17258=>"111111111",
  17259=>"001011000",
  17260=>"100111111",
  17261=>"000110000",
  17262=>"000000000",
  17263=>"001000000",
  17264=>"000100011",
  17265=>"111111000",
  17266=>"000000100",
  17267=>"001111111",
  17268=>"100110100",
  17269=>"000001000",
  17270=>"000100011",
  17271=>"111001001",
  17272=>"110110110",
  17273=>"100000000",
  17274=>"111110000",
  17275=>"001000000",
  17276=>"001001111",
  17277=>"111111111",
  17278=>"111111110",
  17279=>"001001001",
  17280=>"000000000",
  17281=>"111111111",
  17282=>"000000100",
  17283=>"000000110",
  17284=>"101111111",
  17285=>"111110110",
  17286=>"111000110",
  17287=>"000000001",
  17288=>"000111111",
  17289=>"000001100",
  17290=>"110010010",
  17291=>"000000100",
  17292=>"111111111",
  17293=>"111111101",
  17294=>"000000000",
  17295=>"000000011",
  17296=>"000000000",
  17297=>"000000110",
  17298=>"000000000",
  17299=>"011011011",
  17300=>"111101111",
  17301=>"000000000",
  17302=>"111111011",
  17303=>"110101111",
  17304=>"111000111",
  17305=>"001000001",
  17306=>"111111111",
  17307=>"111001011",
  17308=>"001011000",
  17309=>"001111101",
  17310=>"111111110",
  17311=>"000001000",
  17312=>"000000000",
  17313=>"000011010",
  17314=>"000000000",
  17315=>"101001111",
  17316=>"111111010",
  17317=>"111101001",
  17318=>"000000000",
  17319=>"000000111",
  17320=>"000000111",
  17321=>"110111001",
  17322=>"000111111",
  17323=>"000000000",
  17324=>"000000000",
  17325=>"001001000",
  17326=>"000000000",
  17327=>"000000000",
  17328=>"111000000",
  17329=>"000111111",
  17330=>"100110110",
  17331=>"000000011",
  17332=>"111111111",
  17333=>"010110111",
  17334=>"000010000",
  17335=>"100000011",
  17336=>"110000111",
  17337=>"111001000",
  17338=>"000100101",
  17339=>"000100010",
  17340=>"111001011",
  17341=>"010010111",
  17342=>"000000111",
  17343=>"000111000",
  17344=>"111110000",
  17345=>"111111111",
  17346=>"000000000",
  17347=>"100000000",
  17348=>"001111001",
  17349=>"111111001",
  17350=>"000000000",
  17351=>"000110110",
  17352=>"000000111",
  17353=>"111100100",
  17354=>"000000111",
  17355=>"000000111",
  17356=>"111001011",
  17357=>"111111000",
  17358=>"000001011",
  17359=>"000000111",
  17360=>"000000111",
  17361=>"000000000",
  17362=>"000000000",
  17363=>"111111111",
  17364=>"001011001",
  17365=>"000000000",
  17366=>"111111000",
  17367=>"001011001",
  17368=>"000000000",
  17369=>"010000100",
  17370=>"111111011",
  17371=>"000110110",
  17372=>"000001111",
  17373=>"000000000",
  17374=>"111101111",
  17375=>"000000000",
  17376=>"110111001",
  17377=>"000000000",
  17378=>"000111111",
  17379=>"000000000",
  17380=>"111111010",
  17381=>"001011011",
  17382=>"000000011",
  17383=>"111111111",
  17384=>"100100000",
  17385=>"111000111",
  17386=>"000000001",
  17387=>"010000000",
  17388=>"010110100",
  17389=>"111111111",
  17390=>"111001111",
  17391=>"000000000",
  17392=>"111000000",
  17393=>"000000010",
  17394=>"000101101",
  17395=>"000100000",
  17396=>"100100000",
  17397=>"000101111",
  17398=>"000111111",
  17399=>"011001001",
  17400=>"111001000",
  17401=>"000010110",
  17402=>"000110110",
  17403=>"111111111",
  17404=>"001000000",
  17405=>"111111001",
  17406=>"000000000",
  17407=>"001001001",
  17408=>"000000001",
  17409=>"000100000",
  17410=>"111111111",
  17411=>"000111111",
  17412=>"111110000",
  17413=>"101000000",
  17414=>"111111111",
  17415=>"111111111",
  17416=>"000000000",
  17417=>"001000000",
  17418=>"101001001",
  17419=>"101000101",
  17420=>"110000000",
  17421=>"111111000",
  17422=>"000100000",
  17423=>"011111000",
  17424=>"110110110",
  17425=>"001111111",
  17426=>"110111010",
  17427=>"001100001",
  17428=>"000000111",
  17429=>"101000000",
  17430=>"100001101",
  17431=>"111111111",
  17432=>"111111111",
  17433=>"000001111",
  17434=>"000000000",
  17435=>"000000101",
  17436=>"111011111",
  17437=>"111111111",
  17438=>"110110111",
  17439=>"000000000",
  17440=>"000110110",
  17441=>"100000000",
  17442=>"110111010",
  17443=>"000000000",
  17444=>"111001011",
  17445=>"001111111",
  17446=>"000000000",
  17447=>"000000000",
  17448=>"001001001",
  17449=>"000000101",
  17450=>"001000101",
  17451=>"111111011",
  17452=>"110000000",
  17453=>"110111111",
  17454=>"101000001",
  17455=>"000000101",
  17456=>"001010111",
  17457=>"111111000",
  17458=>"111111001",
  17459=>"000000101",
  17460=>"110010000",
  17461=>"100100000",
  17462=>"110111010",
  17463=>"000000001",
  17464=>"111110000",
  17465=>"000100101",
  17466=>"111111110",
  17467=>"111111111",
  17468=>"000000101",
  17469=>"111111111",
  17470=>"001000000",
  17471=>"010011001",
  17472=>"011111111",
  17473=>"000000111",
  17474=>"110111101",
  17475=>"110000001",
  17476=>"110110000",
  17477=>"001011000",
  17478=>"000001111",
  17479=>"111111111",
  17480=>"111111111",
  17481=>"000000000",
  17482=>"100000111",
  17483=>"100100111",
  17484=>"111111001",
  17485=>"111111111",
  17486=>"000000010",
  17487=>"000001111",
  17488=>"000000000",
  17489=>"010011000",
  17490=>"111011011",
  17491=>"000001000",
  17492=>"000001000",
  17493=>"100110100",
  17494=>"110110100",
  17495=>"011111111",
  17496=>"110111010",
  17497=>"111101111",
  17498=>"111111111",
  17499=>"110000000",
  17500=>"111111111",
  17501=>"000000000",
  17502=>"110110111",
  17503=>"011011001",
  17504=>"111111010",
  17505=>"000100111",
  17506=>"000000110",
  17507=>"000000000",
  17508=>"111111000",
  17509=>"011000110",
  17510=>"011001111",
  17511=>"010010000",
  17512=>"010111000",
  17513=>"000000110",
  17514=>"000000000",
  17515=>"000000010",
  17516=>"110100100",
  17517=>"111111111",
  17518=>"001111100",
  17519=>"000000000",
  17520=>"110110000",
  17521=>"000000000",
  17522=>"000011011",
  17523=>"000000100",
  17524=>"000100111",
  17525=>"111110010",
  17526=>"000000111",
  17527=>"111111111",
  17528=>"001000000",
  17529=>"000001001",
  17530=>"111000000",
  17531=>"001001011",
  17532=>"100100100",
  17533=>"000000001",
  17534=>"100000000",
  17535=>"000000000",
  17536=>"100101110",
  17537=>"111110111",
  17538=>"010010110",
  17539=>"000000000",
  17540=>"000000111",
  17541=>"111100110",
  17542=>"110000000",
  17543=>"111001001",
  17544=>"001110000",
  17545=>"000000111",
  17546=>"111101000",
  17547=>"001100111",
  17548=>"000100111",
  17549=>"011111001",
  17550=>"111111111",
  17551=>"011000000",
  17552=>"000001001",
  17553=>"000000001",
  17554=>"010100010",
  17555=>"001001101",
  17556=>"110110111",
  17557=>"100000000",
  17558=>"101000101",
  17559=>"101000100",
  17560=>"001001101",
  17561=>"010111111",
  17562=>"010000110",
  17563=>"000000001",
  17564=>"110110110",
  17565=>"111000101",
  17566=>"111111111",
  17567=>"111111111",
  17568=>"000000000",
  17569=>"100000000",
  17570=>"011111000",
  17571=>"111111101",
  17572=>"100000100",
  17573=>"111111000",
  17574=>"000000001",
  17575=>"000000000",
  17576=>"000000110",
  17577=>"000001111",
  17578=>"100000111",
  17579=>"000000000",
  17580=>"011111111",
  17581=>"100100101",
  17582=>"110000111",
  17583=>"001101111",
  17584=>"111111010",
  17585=>"000000001",
  17586=>"111111010",
  17587=>"111101001",
  17588=>"110000000",
  17589=>"111100100",
  17590=>"000000011",
  17591=>"110111111",
  17592=>"011111011",
  17593=>"111001111",
  17594=>"111001000",
  17595=>"000110110",
  17596=>"000000000",
  17597=>"000000111",
  17598=>"000000000",
  17599=>"000000000",
  17600=>"101001111",
  17601=>"111000000",
  17602=>"111111111",
  17603=>"111111000",
  17604=>"001001101",
  17605=>"000000110",
  17606=>"000010111",
  17607=>"111001111",
  17608=>"010111111",
  17609=>"000000100",
  17610=>"001111001",
  17611=>"111100110",
  17612=>"010010000",
  17613=>"000011011",
  17614=>"000000011",
  17615=>"111111111",
  17616=>"000000000",
  17617=>"000000000",
  17618=>"110111011",
  17619=>"000000100",
  17620=>"111001001",
  17621=>"000000000",
  17622=>"000000000",
  17623=>"000000101",
  17624=>"000000000",
  17625=>"111111110",
  17626=>"111111111",
  17627=>"000110000",
  17628=>"000111111",
  17629=>"000010111",
  17630=>"000110110",
  17631=>"000000000",
  17632=>"001001111",
  17633=>"000000110",
  17634=>"010110000",
  17635=>"111110010",
  17636=>"100110100",
  17637=>"001001001",
  17638=>"111111101",
  17639=>"111111111",
  17640=>"101111111",
  17641=>"111110000",
  17642=>"110111000",
  17643=>"000000110",
  17644=>"000000111",
  17645=>"000000000",
  17646=>"111000101",
  17647=>"111111111",
  17648=>"111001001",
  17649=>"011111100",
  17650=>"111111111",
  17651=>"000000000",
  17652=>"011111111",
  17653=>"111010000",
  17654=>"100001000",
  17655=>"110111000",
  17656=>"011111111",
  17657=>"101111111",
  17658=>"110010000",
  17659=>"001101111",
  17660=>"001001011",
  17661=>"101001011",
  17662=>"000000100",
  17663=>"110000111",
  17664=>"000000000",
  17665=>"100000000",
  17666=>"110000000",
  17667=>"000000101",
  17668=>"111111110",
  17669=>"000000000",
  17670=>"000000000",
  17671=>"000000101",
  17672=>"111111111",
  17673=>"000111111",
  17674=>"000000111",
  17675=>"111111000",
  17676=>"000000000",
  17677=>"011111101",
  17678=>"000000000",
  17679=>"011101110",
  17680=>"000001000",
  17681=>"001111111",
  17682=>"111000010",
  17683=>"010110111",
  17684=>"001001001",
  17685=>"111111111",
  17686=>"001011011",
  17687=>"111011011",
  17688=>"000111001",
  17689=>"111100000",
  17690=>"000000111",
  17691=>"110110000",
  17692=>"000000000",
  17693=>"000000000",
  17694=>"000000000",
  17695=>"011111111",
  17696=>"111111001",
  17697=>"100000000",
  17698=>"111111110",
  17699=>"000000100",
  17700=>"001011011",
  17701=>"001000000",
  17702=>"111001000",
  17703=>"000010110",
  17704=>"111111100",
  17705=>"111111000",
  17706=>"110111010",
  17707=>"000000111",
  17708=>"010000111",
  17709=>"100001111",
  17710=>"001000000",
  17711=>"000000000",
  17712=>"000000000",
  17713=>"011010000",
  17714=>"000000001",
  17715=>"000010010",
  17716=>"000000000",
  17717=>"111100000",
  17718=>"111000001",
  17719=>"100110000",
  17720=>"000010000",
  17721=>"100000111",
  17722=>"001000101",
  17723=>"010000000",
  17724=>"000000110",
  17725=>"110001001",
  17726=>"111111111",
  17727=>"000000111",
  17728=>"011011001",
  17729=>"011001011",
  17730=>"001001101",
  17731=>"011011001",
  17732=>"110110000",
  17733=>"000000000",
  17734=>"111110110",
  17735=>"000000000",
  17736=>"101001111",
  17737=>"111000000",
  17738=>"000101111",
  17739=>"100001001",
  17740=>"000000000",
  17741=>"000000000",
  17742=>"010010111",
  17743=>"000001000",
  17744=>"011101111",
  17745=>"000000101",
  17746=>"000000000",
  17747=>"000000110",
  17748=>"111000000",
  17749=>"000010001",
  17750=>"110110100",
  17751=>"111111111",
  17752=>"111111111",
  17753=>"000000111",
  17754=>"010000000",
  17755=>"010110110",
  17756=>"000000111",
  17757=>"011010111",
  17758=>"110000000",
  17759=>"000100100",
  17760=>"101001101",
  17761=>"000000000",
  17762=>"111111011",
  17763=>"100000000",
  17764=>"000011011",
  17765=>"010000000",
  17766=>"100100110",
  17767=>"001000111",
  17768=>"000000101",
  17769=>"111010110",
  17770=>"000000111",
  17771=>"110100111",
  17772=>"110110100",
  17773=>"101100000",
  17774=>"111111111",
  17775=>"001001111",
  17776=>"000100000",
  17777=>"111111000",
  17778=>"000000000",
  17779=>"011111000",
  17780=>"110100100",
  17781=>"111111010",
  17782=>"000000001",
  17783=>"100101111",
  17784=>"111000111",
  17785=>"111111101",
  17786=>"111111111",
  17787=>"011010100",
  17788=>"110100101",
  17789=>"000000000",
  17790=>"101101101",
  17791=>"001000001",
  17792=>"011111001",
  17793=>"000000011",
  17794=>"100010111",
  17795=>"000000000",
  17796=>"000010111",
  17797=>"000111110",
  17798=>"000011011",
  17799=>"101000111",
  17800=>"100000000",
  17801=>"000000000",
  17802=>"000000000",
  17803=>"000110000",
  17804=>"001111111",
  17805=>"000010000",
  17806=>"000000111",
  17807=>"000110110",
  17808=>"001000001",
  17809=>"110110000",
  17810=>"000111101",
  17811=>"001001100",
  17812=>"111111111",
  17813=>"000010010",
  17814=>"010110110",
  17815=>"100100000",
  17816=>"000000111",
  17817=>"011010000",
  17818=>"111001111",
  17819=>"100000000",
  17820=>"000110110",
  17821=>"111001001",
  17822=>"001000000",
  17823=>"111110000",
  17824=>"000000100",
  17825=>"011011011",
  17826=>"111000000",
  17827=>"000000100",
  17828=>"111111000",
  17829=>"111101101",
  17830=>"000001000",
  17831=>"000010001",
  17832=>"001101101",
  17833=>"100111111",
  17834=>"000000010",
  17835=>"000000000",
  17836=>"100000110",
  17837=>"011110100",
  17838=>"000000001",
  17839=>"110110100",
  17840=>"000001111",
  17841=>"000111010",
  17842=>"101000000",
  17843=>"000000000",
  17844=>"000111111",
  17845=>"111111111",
  17846=>"111110100",
  17847=>"000000100",
  17848=>"000000000",
  17849=>"111111011",
  17850=>"010000000",
  17851=>"111111110",
  17852=>"000000000",
  17853=>"001011111",
  17854=>"000100000",
  17855=>"000000000",
  17856=>"111111000",
  17857=>"111111111",
  17858=>"000000010",
  17859=>"000001000",
  17860=>"000010111",
  17861=>"101001101",
  17862=>"000000000",
  17863=>"101111011",
  17864=>"000000111",
  17865=>"100000111",
  17866=>"101001100",
  17867=>"111111111",
  17868=>"010001000",
  17869=>"001011111",
  17870=>"000000000",
  17871=>"100000000",
  17872=>"000011001",
  17873=>"101111111",
  17874=>"000110000",
  17875=>"001001001",
  17876=>"010010001",
  17877=>"000000000",
  17878=>"000110110",
  17879=>"111111011",
  17880=>"000000100",
  17881=>"000000000",
  17882=>"001001000",
  17883=>"100000110",
  17884=>"101000000",
  17885=>"000000110",
  17886=>"011111000",
  17887=>"100000001",
  17888=>"001101111",
  17889=>"001000000",
  17890=>"000111111",
  17891=>"101101101",
  17892=>"100001000",
  17893=>"000001000",
  17894=>"111011000",
  17895=>"110100111",
  17896=>"101100101",
  17897=>"111010000",
  17898=>"000000000",
  17899=>"000001001",
  17900=>"000000000",
  17901=>"000111000",
  17902=>"101100111",
  17903=>"010111111",
  17904=>"001000000",
  17905=>"110110000",
  17906=>"111111111",
  17907=>"000000000",
  17908=>"000010110",
  17909=>"101000101",
  17910=>"001001001",
  17911=>"001101101",
  17912=>"110110000",
  17913=>"001000100",
  17914=>"110000000",
  17915=>"100000001",
  17916=>"111011000",
  17917=>"000110110",
  17918=>"001111111",
  17919=>"000000101",
  17920=>"011000000",
  17921=>"111011001",
  17922=>"111001001",
  17923=>"101001111",
  17924=>"111111111",
  17925=>"111111010",
  17926=>"000000000",
  17927=>"111001111",
  17928=>"100100101",
  17929=>"110110000",
  17930=>"000010110",
  17931=>"011011011",
  17932=>"100110110",
  17933=>"111111000",
  17934=>"100111011",
  17935=>"111111111",
  17936=>"000000101",
  17937=>"111110000",
  17938=>"111111100",
  17939=>"000000111",
  17940=>"001000001",
  17941=>"111011001",
  17942=>"111111111",
  17943=>"001000000",
  17944=>"111111111",
  17945=>"100111111",
  17946=>"010011111",
  17947=>"111111111",
  17948=>"110111111",
  17949=>"011011111",
  17950=>"110100100",
  17951=>"111111101",
  17952=>"111111100",
  17953=>"001100111",
  17954=>"111111111",
  17955=>"000111111",
  17956=>"111110000",
  17957=>"111111111",
  17958=>"000000000",
  17959=>"111111111",
  17960=>"100100011",
  17961=>"001000000",
  17962=>"011011011",
  17963=>"001111101",
  17964=>"111111000",
  17965=>"000000000",
  17966=>"001001011",
  17967=>"000001011",
  17968=>"000000000",
  17969=>"000000000",
  17970=>"101111111",
  17971=>"000111100",
  17972=>"011011111",
  17973=>"010000000",
  17974=>"111111111",
  17975=>"111111000",
  17976=>"000000111",
  17977=>"111111010",
  17978=>"111111111",
  17979=>"111100101",
  17980=>"000000100",
  17981=>"000000000",
  17982=>"101000000",
  17983=>"001001111",
  17984=>"111111010",
  17985=>"010000000",
  17986=>"000000001",
  17987=>"000101111",
  17988=>"010011001",
  17989=>"111111110",
  17990=>"000010000",
  17991=>"000000001",
  17992=>"001000000",
  17993=>"101001011",
  17994=>"000000101",
  17995=>"110000001",
  17996=>"001001001",
  17997=>"100000010",
  17998=>"101110100",
  17999=>"111111111",
  18000=>"110100000",
  18001=>"111111001",
  18002=>"111111111",
  18003=>"000000110",
  18004=>"111000000",
  18005=>"000101111",
  18006=>"110111110",
  18007=>"111111110",
  18008=>"001001000",
  18009=>"100000101",
  18010=>"101111111",
  18011=>"110000000",
  18012=>"111110100",
  18013=>"001000101",
  18014=>"011001111",
  18015=>"011001100",
  18016=>"000011010",
  18017=>"001000100",
  18018=>"111111111",
  18019=>"111001001",
  18020=>"111111111",
  18021=>"110111011",
  18022=>"001001001",
  18023=>"101111101",
  18024=>"010111111",
  18025=>"011000000",
  18026=>"000000111",
  18027=>"000110011",
  18028=>"000000000",
  18029=>"000000000",
  18030=>"101101101",
  18031=>"000110110",
  18032=>"111111111",
  18033=>"001111111",
  18034=>"111111111",
  18035=>"100011001",
  18036=>"010010000",
  18037=>"110111111",
  18038=>"100000101",
  18039=>"000111111",
  18040=>"000000110",
  18041=>"001000000",
  18042=>"011111111",
  18043=>"100100000",
  18044=>"100100100",
  18045=>"000000000",
  18046=>"000000000",
  18047=>"010010010",
  18048=>"111100000",
  18049=>"111111111",
  18050=>"011001000",
  18051=>"011010000",
  18052=>"000000011",
  18053=>"111000111",
  18054=>"011011111",
  18055=>"000001001",
  18056=>"110111011",
  18057=>"000111111",
  18058=>"000000000",
  18059=>"000101000",
  18060=>"111011110",
  18061=>"011101000",
  18062=>"111111111",
  18063=>"111111110",
  18064=>"101101111",
  18065=>"000000000",
  18066=>"000000000",
  18067=>"111111110",
  18068=>"000000111",
  18069=>"111000000",
  18070=>"111001101",
  18071=>"000000000",
  18072=>"100101101",
  18073=>"111111111",
  18074=>"000000000",
  18075=>"111101111",
  18076=>"001001000",
  18077=>"110110110",
  18078=>"111111111",
  18079=>"001010110",
  18080=>"000000000",
  18081=>"100111101",
  18082=>"111111111",
  18083=>"111000000",
  18084=>"110001000",
  18085=>"111111111",
  18086=>"101111110",
  18087=>"111110100",
  18088=>"000000000",
  18089=>"111100110",
  18090=>"110000000",
  18091=>"111001001",
  18092=>"101100100",
  18093=>"001000001",
  18094=>"000000000",
  18095=>"000000111",
  18096=>"000000000",
  18097=>"101100000",
  18098=>"011111111",
  18099=>"111111111",
  18100=>"000000000",
  18101=>"110111000",
  18102=>"111110110",
  18103=>"001101101",
  18104=>"111111001",
  18105=>"000000000",
  18106=>"011111000",
  18107=>"000000000",
  18108=>"000000000",
  18109=>"111111010",
  18110=>"000000000",
  18111=>"100100111",
  18112=>"111111111",
  18113=>"000000000",
  18114=>"111111111",
  18115=>"111111111",
  18116=>"001001001",
  18117=>"000000000",
  18118=>"111001001",
  18119=>"111110100",
  18120=>"110111111",
  18121=>"011111111",
  18122=>"100100111",
  18123=>"000000000",
  18124=>"111111111",
  18125=>"011011010",
  18126=>"000001001",
  18127=>"000000110",
  18128=>"001000000",
  18129=>"000000111",
  18130=>"111111000",
  18131=>"011000000",
  18132=>"100000000",
  18133=>"000001001",
  18134=>"000000000",
  18135=>"111110110",
  18136=>"111111111",
  18137=>"000000001",
  18138=>"110110000",
  18139=>"000000111",
  18140=>"001000000",
  18141=>"000010111",
  18142=>"110111101",
  18143=>"001000001",
  18144=>"000000000",
  18145=>"010000000",
  18146=>"111000000",
  18147=>"100100000",
  18148=>"000100111",
  18149=>"001001011",
  18150=>"000010000",
  18151=>"011011111",
  18152=>"011011001",
  18153=>"100110111",
  18154=>"110100100",
  18155=>"000111111",
  18156=>"110000101",
  18157=>"111111111",
  18158=>"111000000",
  18159=>"000000101",
  18160=>"000000000",
  18161=>"000000000",
  18162=>"000000000",
  18163=>"000000101",
  18164=>"111111011",
  18165=>"100110111",
  18166=>"111111001",
  18167=>"011111011",
  18168=>"010000000",
  18169=>"111111111",
  18170=>"000111000",
  18171=>"000010000",
  18172=>"011011001",
  18173=>"000000001",
  18174=>"011100000",
  18175=>"111111111",
  18176=>"001111111",
  18177=>"000000000",
  18178=>"000000000",
  18179=>"111001001",
  18180=>"111111111",
  18181=>"100100110",
  18182=>"111110100",
  18183=>"010110111",
  18184=>"010000000",
  18185=>"011000001",
  18186=>"111111001",
  18187=>"000000000",
  18188=>"111111010",
  18189=>"000000000",
  18190=>"000000010",
  18191=>"000000000",
  18192=>"111111011",
  18193=>"010111111",
  18194=>"100100111",
  18195=>"001111100",
  18196=>"110101000",
  18197=>"000000000",
  18198=>"111011100",
  18199=>"000000000",
  18200=>"111111000",
  18201=>"100000000",
  18202=>"000000000",
  18203=>"110100000",
  18204=>"100001001",
  18205=>"111011011",
  18206=>"000000000",
  18207=>"000000111",
  18208=>"111011001",
  18209=>"001000011",
  18210=>"000001000",
  18211=>"100111010",
  18212=>"110011011",
  18213=>"010111111",
  18214=>"111111111",
  18215=>"100110111",
  18216=>"001000111",
  18217=>"111101000",
  18218=>"000000001",
  18219=>"000000000",
  18220=>"000110000",
  18221=>"000001001",
  18222=>"111100111",
  18223=>"111111111",
  18224=>"110110110",
  18225=>"010010110",
  18226=>"001001000",
  18227=>"111111111",
  18228=>"010110010",
  18229=>"001001011",
  18230=>"110110011",
  18231=>"000000100",
  18232=>"010011011",
  18233=>"000000000",
  18234=>"101000101",
  18235=>"000000000",
  18236=>"000010011",
  18237=>"011111010",
  18238=>"011001111",
  18239=>"000000111",
  18240=>"100000000",
  18241=>"111111110",
  18242=>"110111000",
  18243=>"000001000",
  18244=>"111111111",
  18245=>"000000000",
  18246=>"011000000",
  18247=>"000000000",
  18248=>"001000000",
  18249=>"011111111",
  18250=>"110111111",
  18251=>"011011111",
  18252=>"110000000",
  18253=>"010000000",
  18254=>"000000000",
  18255=>"111111100",
  18256=>"111000000",
  18257=>"110111111",
  18258=>"111111111",
  18259=>"011000001",
  18260=>"010010000",
  18261=>"011011011",
  18262=>"000000000",
  18263=>"111111101",
  18264=>"100100000",
  18265=>"000111111",
  18266=>"000000110",
  18267=>"000000000",
  18268=>"111111111",
  18269=>"111011000",
  18270=>"000000100",
  18271=>"011111110",
  18272=>"011011001",
  18273=>"101000110",
  18274=>"111100100",
  18275=>"001000000",
  18276=>"001001000",
  18277=>"000000000",
  18278=>"000000011",
  18279=>"001000000",
  18280=>"100100110",
  18281=>"000001011",
  18282=>"111111111",
  18283=>"010111111",
  18284=>"000100000",
  18285=>"010111111",
  18286=>"111111000",
  18287=>"111000000",
  18288=>"111111111",
  18289=>"000000000",
  18290=>"000000111",
  18291=>"111111011",
  18292=>"000000000",
  18293=>"000000000",
  18294=>"110100000",
  18295=>"111111001",
  18296=>"000000000",
  18297=>"101000000",
  18298=>"111111001",
  18299=>"111111111",
  18300=>"000100000",
  18301=>"000000111",
  18302=>"110000000",
  18303=>"111000000",
  18304=>"111110100",
  18305=>"000010111",
  18306=>"111111111",
  18307=>"000000000",
  18308=>"111111111",
  18309=>"110100000",
  18310=>"111110111",
  18311=>"000010111",
  18312=>"111000101",
  18313=>"111111001",
  18314=>"111111011",
  18315=>"000011011",
  18316=>"111001001",
  18317=>"100110110",
  18318=>"010111000",
  18319=>"000000000",
  18320=>"111101111",
  18321=>"011001011",
  18322=>"111111110",
  18323=>"000000000",
  18324=>"111011000",
  18325=>"000010000",
  18326=>"111111000",
  18327=>"000000011",
  18328=>"010111111",
  18329=>"001111111",
  18330=>"000000001",
  18331=>"011111011",
  18332=>"000000000",
  18333=>"111000100",
  18334=>"010110111",
  18335=>"000011010",
  18336=>"000100000",
  18337=>"111000100",
  18338=>"111110100",
  18339=>"110111111",
  18340=>"101101001",
  18341=>"011011011",
  18342=>"111111111",
  18343=>"110010000",
  18344=>"111111000",
  18345=>"111000000",
  18346=>"111111111",
  18347=>"000010110",
  18348=>"111111000",
  18349=>"000001001",
  18350=>"001110111",
  18351=>"000000100",
  18352=>"101000111",
  18353=>"000010000",
  18354=>"000000100",
  18355=>"111111111",
  18356=>"011110110",
  18357=>"000000111",
  18358=>"000000111",
  18359=>"000000000",
  18360=>"000000000",
  18361=>"111111100",
  18362=>"110111000",
  18363=>"111000000",
  18364=>"000000000",
  18365=>"000001011",
  18366=>"000000000",
  18367=>"001000000",
  18368=>"100100001",
  18369=>"111111001",
  18370=>"010111111",
  18371=>"111111000",
  18372=>"000100000",
  18373=>"101101001",
  18374=>"111110010",
  18375=>"011011011",
  18376=>"000000000",
  18377=>"000100100",
  18378=>"101111111",
  18379=>"000000111",
  18380=>"010000000",
  18381=>"001001001",
  18382=>"111111001",
  18383=>"001000111",
  18384=>"001000100",
  18385=>"011111011",
  18386=>"000000111",
  18387=>"111111011",
  18388=>"000000001",
  18389=>"000000000",
  18390=>"111100000",
  18391=>"011011011",
  18392=>"100100111",
  18393=>"000000111",
  18394=>"000000000",
  18395=>"111000000",
  18396=>"111000000",
  18397=>"011011111",
  18398=>"100100111",
  18399=>"001001101",
  18400=>"000010000",
  18401=>"000000000",
  18402=>"000000000",
  18403=>"000100100",
  18404=>"001001000",
  18405=>"111011000",
  18406=>"111111001",
  18407=>"110111111",
  18408=>"000000000",
  18409=>"110110000",
  18410=>"000001010",
  18411=>"011000011",
  18412=>"000000100",
  18413=>"000100110",
  18414=>"101101101",
  18415=>"010111111",
  18416=>"000000110",
  18417=>"000000100",
  18418=>"000000000",
  18419=>"111111111",
  18420=>"111111110",
  18421=>"001000000",
  18422=>"111111010",
  18423=>"000000000",
  18424=>"000111111",
  18425=>"111101000",
  18426=>"000000000",
  18427=>"000000100",
  18428=>"000000000",
  18429=>"000000000",
  18430=>"000000101",
  18431=>"000000000",
  18432=>"110000000",
  18433=>"111000000",
  18434=>"111111111",
  18435=>"110110110",
  18436=>"011010111",
  18437=>"000000111",
  18438=>"111111101",
  18439=>"111110111",
  18440=>"000000000",
  18441=>"111111111",
  18442=>"110110110",
  18443=>"011111111",
  18444=>"111100111",
  18445=>"001001011",
  18446=>"000000111",
  18447=>"001001001",
  18448=>"000100111",
  18449=>"010110000",
  18450=>"111110111",
  18451=>"000000001",
  18452=>"001000011",
  18453=>"111011111",
  18454=>"111101011",
  18455=>"111110110",
  18456=>"000000111",
  18457=>"001000000",
  18458=>"101111111",
  18459=>"111100000",
  18460=>"111001111",
  18461=>"100110111",
  18462=>"000110111",
  18463=>"001101100",
  18464=>"000100111",
  18465=>"110110111",
  18466=>"111100001",
  18467=>"000000111",
  18468=>"000000001",
  18469=>"101001111",
  18470=>"110110011",
  18471=>"111111000",
  18472=>"001000111",
  18473=>"000001000",
  18474=>"001001111",
  18475=>"001001111",
  18476=>"000000000",
  18477=>"111111100",
  18478=>"000101111",
  18479=>"100100100",
  18480=>"110100000",
  18481=>"001100100",
  18482=>"000100000",
  18483=>"000000000",
  18484=>"000000101",
  18485=>"000000000",
  18486=>"111101111",
  18487=>"111001001",
  18488=>"111010001",
  18489=>"000100111",
  18490=>"001101111",
  18491=>"111101100",
  18492=>"000000111",
  18493=>"100110110",
  18494=>"000000000",
  18495=>"000000000",
  18496=>"001001001",
  18497=>"000000000",
  18498=>"001001111",
  18499=>"101111101",
  18500=>"000000000",
  18501=>"001001111",
  18502=>"000000000",
  18503=>"111101111",
  18504=>"110110110",
  18505=>"101101111",
  18506=>"011011010",
  18507=>"111111000",
  18508=>"110110000",
  18509=>"111111111",
  18510=>"000000101",
  18511=>"111001101",
  18512=>"111001000",
  18513=>"001001111",
  18514=>"010000000",
  18515=>"000110110",
  18516=>"001101111",
  18517=>"111111111",
  18518=>"000000000",
  18519=>"111111111",
  18520=>"000000111",
  18521=>"111101111",
  18522=>"111100000",
  18523=>"000000110",
  18524=>"111111111",
  18525=>"001000111",
  18526=>"001000100",
  18527=>"100110111",
  18528=>"100110110",
  18529=>"110100100",
  18530=>"000000111",
  18531=>"000111110",
  18532=>"110110010",
  18533=>"111111111",
  18534=>"000000111",
  18535=>"111001101",
  18536=>"100111111",
  18537=>"011111111",
  18538=>"001001111",
  18539=>"001000101",
  18540=>"000000001",
  18541=>"111111001",
  18542=>"111010010",
  18543=>"110110000",
  18544=>"000000000",
  18545=>"110110111",
  18546=>"000100110",
  18547=>"000000000",
  18548=>"001001111",
  18549=>"111111111",
  18550=>"000000111",
  18551=>"111011011",
  18552=>"111111111",
  18553=>"111111000",
  18554=>"001001111",
  18555=>"111111111",
  18556=>"100100100",
  18557=>"000000000",
  18558=>"000000000",
  18559=>"110111000",
  18560=>"001000110",
  18561=>"101100000",
  18562=>"001000000",
  18563=>"100100111",
  18564=>"000001001",
  18565=>"111111011",
  18566=>"000110000",
  18567=>"000000000",
  18568=>"001000001",
  18569=>"001001011",
  18570=>"000000110",
  18571=>"010010110",
  18572=>"000000001",
  18573=>"001000001",
  18574=>"111001111",
  18575=>"000000001",
  18576=>"001001111",
  18577=>"100111111",
  18578=>"000000000",
  18579=>"000001001",
  18580=>"000000001",
  18581=>"101000001",
  18582=>"111111000",
  18583=>"100100101",
  18584=>"000000001",
  18585=>"111111011",
  18586=>"110111111",
  18587=>"000000000",
  18588=>"001001111",
  18589=>"011111110",
  18590=>"110110000",
  18591=>"011111011",
  18592=>"111110111",
  18593=>"001111111",
  18594=>"000000111",
  18595=>"000010000",
  18596=>"011001001",
  18597=>"111011011",
  18598=>"110111111",
  18599=>"011111011",
  18600=>"000000000",
  18601=>"000111001",
  18602=>"101110100",
  18603=>"000000110",
  18604=>"111111111",
  18605=>"100110110",
  18606=>"001001111",
  18607=>"111011000",
  18608=>"110110000",
  18609=>"000010000",
  18610=>"111111011",
  18611=>"111111000",
  18612=>"111101111",
  18613=>"001001001",
  18614=>"001001001",
  18615=>"111111101",
  18616=>"001000000",
  18617=>"111011000",
  18618=>"011001001",
  18619=>"001001011",
  18620=>"001101111",
  18621=>"011000000",
  18622=>"000001000",
  18623=>"000000001",
  18624=>"111111111",
  18625=>"111110111",
  18626=>"010000001",
  18627=>"111111100",
  18628=>"000011110",
  18629=>"001000000",
  18630=>"001001111",
  18631=>"110110000",
  18632=>"001000110",
  18633=>"000000111",
  18634=>"000001111",
  18635=>"001000101",
  18636=>"000001111",
  18637=>"111111101",
  18638=>"101101100",
  18639=>"011000000",
  18640=>"000000101",
  18641=>"111111111",
  18642=>"101111000",
  18643=>"110010000",
  18644=>"101000011",
  18645=>"000000011",
  18646=>"000000000",
  18647=>"001001111",
  18648=>"000000000",
  18649=>"000000111",
  18650=>"111101000",
  18651=>"111010010",
  18652=>"111000010",
  18653=>"101101111",
  18654=>"101111100",
  18655=>"000101111",
  18656=>"000000000",
  18657=>"000010110",
  18658=>"111111111",
  18659=>"001000100",
  18660=>"100000001",
  18661=>"000000010",
  18662=>"001000110",
  18663=>"000000001",
  18664=>"110110000",
  18665=>"000001111",
  18666=>"100110100",
  18667=>"111110100",
  18668=>"011101001",
  18669=>"111001000",
  18670=>"000001111",
  18671=>"111111000",
  18672=>"111111111",
  18673=>"101111111",
  18674=>"111111111",
  18675=>"001001110",
  18676=>"111111111",
  18677=>"011010110",
  18678=>"111111001",
  18679=>"111111111",
  18680=>"000001111",
  18681=>"001000100",
  18682=>"000010000",
  18683=>"100010000",
  18684=>"110111111",
  18685=>"000000011",
  18686=>"111100101",
  18687=>"001001011",
  18688=>"001110000",
  18689=>"001001011",
  18690=>"000110000",
  18691=>"111111011",
  18692=>"000000000",
  18693=>"000001011",
  18694=>"111011010",
  18695=>"110110110",
  18696=>"110110000",
  18697=>"000000000",
  18698=>"100100101",
  18699=>"100101111",
  18700=>"000000111",
  18701=>"000001101",
  18702=>"000001101",
  18703=>"000000000",
  18704=>"001010111",
  18705=>"101101111",
  18706=>"000000111",
  18707=>"000001001",
  18708=>"000001111",
  18709=>"000111111",
  18710=>"100000000",
  18711=>"000001111",
  18712=>"111111111",
  18713=>"111111000",
  18714=>"000001001",
  18715=>"111111111",
  18716=>"000000001",
  18717=>"000000000",
  18718=>"011001011",
  18719=>"110000000",
  18720=>"111011000",
  18721=>"110101111",
  18722=>"000000111",
  18723=>"110110000",
  18724=>"111010000",
  18725=>"111010000",
  18726=>"000000101",
  18727=>"110010000",
  18728=>"000000000",
  18729=>"010011001",
  18730=>"000100111",
  18731=>"100000000",
  18732=>"000000000",
  18733=>"001111010",
  18734=>"111000000",
  18735=>"000001001",
  18736=>"000110011",
  18737=>"000000000",
  18738=>"111111010",
  18739=>"000000100",
  18740=>"111111000",
  18741=>"000000000",
  18742=>"000000011",
  18743=>"000000000",
  18744=>"000000100",
  18745=>"000110101",
  18746=>"101101111",
  18747=>"111111001",
  18748=>"111110110",
  18749=>"001000111",
  18750=>"011000001",
  18751=>"111111111",
  18752=>"001001001",
  18753=>"001111111",
  18754=>"000110110",
  18755=>"000000100",
  18756=>"111111001",
  18757=>"110111100",
  18758=>"111101101",
  18759=>"000001001",
  18760=>"011000001",
  18761=>"111111000",
  18762=>"000000110",
  18763=>"110100001",
  18764=>"111101000",
  18765=>"000111111",
  18766=>"011000000",
  18767=>"000110000",
  18768=>"001001111",
  18769=>"000000000",
  18770=>"000000100",
  18771=>"000000110",
  18772=>"000111110",
  18773=>"011011011",
  18774=>"001001111",
  18775=>"101001111",
  18776=>"001011010",
  18777=>"010000000",
  18778=>"000000000",
  18779=>"001001111",
  18780=>"111111111",
  18781=>"000111111",
  18782=>"000000111",
  18783=>"000000110",
  18784=>"000001111",
  18785=>"000001111",
  18786=>"001111110",
  18787=>"000001111",
  18788=>"011111100",
  18789=>"100110110",
  18790=>"000011000",
  18791=>"110110111",
  18792=>"100110110",
  18793=>"011000000",
  18794=>"000000111",
  18795=>"100110110",
  18796=>"110110100",
  18797=>"111000111",
  18798=>"011011111",
  18799=>"000000000",
  18800=>"101001011",
  18801=>"000000000",
  18802=>"111111111",
  18803=>"111000011",
  18804=>"111111111",
  18805=>"111111111",
  18806=>"000010000",
  18807=>"111111100",
  18808=>"111001111",
  18809=>"000000000",
  18810=>"000000111",
  18811=>"110110111",
  18812=>"000000111",
  18813=>"000000001",
  18814=>"111111111",
  18815=>"000000001",
  18816=>"000110111",
  18817=>"110100000",
  18818=>"100111101",
  18819=>"000001111",
  18820=>"111111111",
  18821=>"010111100",
  18822=>"001000000",
  18823=>"000000000",
  18824=>"001001001",
  18825=>"111111101",
  18826=>"110110000",
  18827=>"111000000",
  18828=>"001001001",
  18829=>"001000111",
  18830=>"110110111",
  18831=>"111111110",
  18832=>"010111000",
  18833=>"111111111",
  18834=>"000111111",
  18835=>"111111111",
  18836=>"101110000",
  18837=>"000000000",
  18838=>"000000111",
  18839=>"000100101",
  18840=>"001011111",
  18841=>"000000000",
  18842=>"110110010",
  18843=>"001001000",
  18844=>"001011111",
  18845=>"000000000",
  18846=>"000001000",
  18847=>"111111111",
  18848=>"000000000",
  18849=>"111011000",
  18850=>"100111111",
  18851=>"000010000",
  18852=>"001001101",
  18853=>"000000000",
  18854=>"111110000",
  18855=>"100110110",
  18856=>"000000000",
  18857=>"111111111",
  18858=>"111111111",
  18859=>"100000111",
  18860=>"000010010",
  18861=>"110110010",
  18862=>"111111111",
  18863=>"001001011",
  18864=>"111111110",
  18865=>"000000000",
  18866=>"111111111",
  18867=>"110100100",
  18868=>"000000000",
  18869=>"000010111",
  18870=>"001001101",
  18871=>"111011011",
  18872=>"000000000",
  18873=>"110110110",
  18874=>"100000000",
  18875=>"111110000",
  18876=>"111110011",
  18877=>"110000000",
  18878=>"000000111",
  18879=>"111110011",
  18880=>"000000000",
  18881=>"110100100",
  18882=>"010111000",
  18883=>"110000000",
  18884=>"111111111",
  18885=>"111011010",
  18886=>"101100000",
  18887=>"100000111",
  18888=>"000000100",
  18889=>"000000001",
  18890=>"101101111",
  18891=>"011111111",
  18892=>"110000000",
  18893=>"111111111",
  18894=>"000000000",
  18895=>"000001111",
  18896=>"000010000",
  18897=>"101101111",
  18898=>"111110110",
  18899=>"000100111",
  18900=>"111111110",
  18901=>"111111111",
  18902=>"000110111",
  18903=>"000000100",
  18904=>"000000000",
  18905=>"110100111",
  18906=>"100000000",
  18907=>"001000000",
  18908=>"000000111",
  18909=>"001001001",
  18910=>"111111000",
  18911=>"111100110",
  18912=>"001000000",
  18913=>"111110111",
  18914=>"000101000",
  18915=>"001001111",
  18916=>"001111111",
  18917=>"011001111",
  18918=>"000000011",
  18919=>"111000000",
  18920=>"000000001",
  18921=>"000000111",
  18922=>"000000000",
  18923=>"000011111",
  18924=>"010000000",
  18925=>"001001001",
  18926=>"000110111",
  18927=>"101001111",
  18928=>"000000000",
  18929=>"111111101",
  18930=>"100111101",
  18931=>"000000011",
  18932=>"111001110",
  18933=>"111100100",
  18934=>"000000100",
  18935=>"110110000",
  18936=>"111111111",
  18937=>"001011001",
  18938=>"000100000",
  18939=>"000000100",
  18940=>"000000001",
  18941=>"001000000",
  18942=>"111111111",
  18943=>"111111111",
  18944=>"000000110",
  18945=>"000100100",
  18946=>"000000000",
  18947=>"000010101",
  18948=>"001111111",
  18949=>"101100000",
  18950=>"101001001",
  18951=>"000000000",
  18952=>"000000000",
  18953=>"000000000",
  18954=>"001001000",
  18955=>"000001000",
  18956=>"111101000",
  18957=>"100000010",
  18958=>"101000100",
  18959=>"111111111",
  18960=>"111001011",
  18961=>"101000000",
  18962=>"111111111",
  18963=>"000000001",
  18964=>"101111111",
  18965=>"001000100",
  18966=>"110010010",
  18967=>"001011001",
  18968=>"000100100",
  18969=>"110001001",
  18970=>"000000000",
  18971=>"111111101",
  18972=>"101001101",
  18973=>"000000000",
  18974=>"000110110",
  18975=>"011011111",
  18976=>"101111111",
  18977=>"001000000",
  18978=>"001101101",
  18979=>"011111110",
  18980=>"111000000",
  18981=>"100111111",
  18982=>"000111000",
  18983=>"000000000",
  18984=>"101100000",
  18985=>"010111011",
  18986=>"000000000",
  18987=>"111111011",
  18988=>"101000000",
  18989=>"011000000",
  18990=>"111111111",
  18991=>"000000000",
  18992=>"000111111",
  18993=>"111111111",
  18994=>"100000000",
  18995=>"110111111",
  18996=>"000001001",
  18997=>"111011011",
  18998=>"001001001",
  18999=>"110100000",
  19000=>"001101111",
  19001=>"100100111",
  19002=>"111111111",
  19003=>"010110110",
  19004=>"111101100",
  19005=>"111111111",
  19006=>"110100000",
  19007=>"000000000",
  19008=>"111000111",
  19009=>"011011001",
  19010=>"111111111",
  19011=>"000000000",
  19012=>"000000100",
  19013=>"111111110",
  19014=>"111100000",
  19015=>"000001101",
  19016=>"011101100",
  19017=>"111111000",
  19018=>"001001001",
  19019=>"001001001",
  19020=>"000010000",
  19021=>"111000100",
  19022=>"000111101",
  19023=>"000000000",
  19024=>"111111000",
  19025=>"110000000",
  19026=>"000000000",
  19027=>"000001001",
  19028=>"111101111",
  19029=>"000000011",
  19030=>"111110010",
  19031=>"111000011",
  19032=>"000000111",
  19033=>"100000000",
  19034=>"101101000",
  19035=>"001000000",
  19036=>"101111100",
  19037=>"000000000",
  19038=>"111011000",
  19039=>"111111111",
  19040=>"011101111",
  19041=>"110101111",
  19042=>"101001001",
  19043=>"000000000",
  19044=>"111110000",
  19045=>"111110000",
  19046=>"000000000",
  19047=>"000000000",
  19048=>"000000111",
  19049=>"111111111",
  19050=>"000001011",
  19051=>"000100100",
  19052=>"011001000",
  19053=>"111111111",
  19054=>"111010110",
  19055=>"110110011",
  19056=>"111011011",
  19057=>"111111111",
  19058=>"000000000",
  19059=>"000011000",
  19060=>"000001011",
  19061=>"001001111",
  19062=>"000010000",
  19063=>"101101111",
  19064=>"101000000",
  19065=>"111111111",
  19066=>"000000100",
  19067=>"011110111",
  19068=>"110110110",
  19069=>"000000000",
  19070=>"111111111",
  19071=>"000000000",
  19072=>"000000000",
  19073=>"011111111",
  19074=>"111011000",
  19075=>"110111111",
  19076=>"111100101",
  19077=>"111111111",
  19078=>"001000001",
  19079=>"100111111",
  19080=>"000000000",
  19081=>"110100000",
  19082=>"100111110",
  19083=>"111111111",
  19084=>"000000000",
  19085=>"000000000",
  19086=>"011110110",
  19087=>"000000000",
  19088=>"000000000",
  19089=>"000001001",
  19090=>"111000000",
  19091=>"000011111",
  19092=>"000000100",
  19093=>"101100100",
  19094=>"000000111",
  19095=>"000000000",
  19096=>"001001001",
  19097=>"110011111",
  19098=>"000000000",
  19099=>"000000000",
  19100=>"100101001",
  19101=>"111000000",
  19102=>"100100111",
  19103=>"000000000",
  19104=>"111111111",
  19105=>"100100000",
  19106=>"100100100",
  19107=>"001111111",
  19108=>"001001001",
  19109=>"111101100",
  19110=>"111111010",
  19111=>"111111000",
  19112=>"000000000",
  19113=>"111111111",
  19114=>"000000000",
  19115=>"110101000",
  19116=>"000000000",
  19117=>"100110111",
  19118=>"000000000",
  19119=>"101111111",
  19120=>"110110111",
  19121=>"001000001",
  19122=>"100110100",
  19123=>"000000000",
  19124=>"111111111",
  19125=>"111111011",
  19126=>"000000000",
  19127=>"010111111",
  19128=>"001001011",
  19129=>"000000000",
  19130=>"000000000",
  19131=>"111001000",
  19132=>"000000111",
  19133=>"000000000",
  19134=>"111111111",
  19135=>"111111110",
  19136=>"000000000",
  19137=>"111111011",
  19138=>"001011011",
  19139=>"000000000",
  19140=>"000000111",
  19141=>"000000000",
  19142=>"000000000",
  19143=>"001000010",
  19144=>"111111111",
  19145=>"111111100",
  19146=>"101000100",
  19147=>"111000000",
  19148=>"000000000",
  19149=>"011101101",
  19150=>"111100111",
  19151=>"111111111",
  19152=>"110110100",
  19153=>"000000000",
  19154=>"111100100",
  19155=>"001000111",
  19156=>"000000000",
  19157=>"111111111",
  19158=>"111010000",
  19159=>"001000000",
  19160=>"000000000",
  19161=>"001100100",
  19162=>"000000000",
  19163=>"000000000",
  19164=>"111111111",
  19165=>"111110100",
  19166=>"111111000",
  19167=>"000001001",
  19168=>"111111111",
  19169=>"000000000",
  19170=>"010110110",
  19171=>"111111100",
  19172=>"110100100",
  19173=>"000001000",
  19174=>"100100111",
  19175=>"000101111",
  19176=>"001000000",
  19177=>"111101101",
  19178=>"001000001",
  19179=>"111000000",
  19180=>"000001010",
  19181=>"111110110",
  19182=>"000000111",
  19183=>"000000000",
  19184=>"001111111",
  19185=>"111111111",
  19186=>"111100000",
  19187=>"100000011",
  19188=>"011011111",
  19189=>"110100100",
  19190=>"011101111",
  19191=>"000010011",
  19192=>"000000100",
  19193=>"000000000",
  19194=>"111111111",
  19195=>"011111000",
  19196=>"000100111",
  19197=>"001001000",
  19198=>"111111111",
  19199=>"001000100",
  19200=>"000000000",
  19201=>"001001001",
  19202=>"111111111",
  19203=>"111111111",
  19204=>"000000000",
  19205=>"001001111",
  19206=>"000000000",
  19207=>"111111111",
  19208=>"101111111",
  19209=>"000000000",
  19210=>"100111000",
  19211=>"000000000",
  19212=>"000100111",
  19213=>"000000000",
  19214=>"111111110",
  19215=>"001001101",
  19216=>"001111111",
  19217=>"000000000",
  19218=>"000000011",
  19219=>"001101001",
  19220=>"111111111",
  19221=>"111100100",
  19222=>"111111111",
  19223=>"111100111",
  19224=>"111111111",
  19225=>"111111111",
  19226=>"100000000",
  19227=>"100110111",
  19228=>"111001101",
  19229=>"000111111",
  19230=>"000000000",
  19231=>"111111100",
  19232=>"000000001",
  19233=>"000000110",
  19234=>"111000000",
  19235=>"001101111",
  19236=>"111010010",
  19237=>"100100000",
  19238=>"000000000",
  19239=>"000001000",
  19240=>"000000011",
  19241=>"111000000",
  19242=>"101101111",
  19243=>"100100100",
  19244=>"111101111",
  19245=>"000000000",
  19246=>"111011000",
  19247=>"000000000",
  19248=>"101100000",
  19249=>"000001001",
  19250=>"111101100",
  19251=>"000100000",
  19252=>"111111111",
  19253=>"011001111",
  19254=>"000000110",
  19255=>"111111111",
  19256=>"000000000",
  19257=>"000000000",
  19258=>"100100100",
  19259=>"001000100",
  19260=>"000000000",
  19261=>"000000011",
  19262=>"000000000",
  19263=>"100000000",
  19264=>"000001111",
  19265=>"000000000",
  19266=>"111111101",
  19267=>"000000110",
  19268=>"001000000",
  19269=>"100100000",
  19270=>"111111111",
  19271=>"100000000",
  19272=>"111110110",
  19273=>"111100000",
  19274=>"000000111",
  19275=>"110000000",
  19276=>"000000000",
  19277=>"000011111",
  19278=>"111001000",
  19279=>"000000000",
  19280=>"000100100",
  19281=>"101000110",
  19282=>"001001001",
  19283=>"100100111",
  19284=>"001000000",
  19285=>"011001001",
  19286=>"111001001",
  19287=>"111110111",
  19288=>"111111111",
  19289=>"111111111",
  19290=>"111111111",
  19291=>"011000110",
  19292=>"000000111",
  19293=>"000000000",
  19294=>"000111111",
  19295=>"000000000",
  19296=>"000000000",
  19297=>"000000011",
  19298=>"000001001",
  19299=>"111001101",
  19300=>"000000010",
  19301=>"100100111",
  19302=>"000000000",
  19303=>"001000000",
  19304=>"100001001",
  19305=>"111000000",
  19306=>"111111111",
  19307=>"111110000",
  19308=>"111111111",
  19309=>"101111101",
  19310=>"000001001",
  19311=>"001001001",
  19312=>"000111111",
  19313=>"000000000",
  19314=>"111111111",
  19315=>"110110010",
  19316=>"111100100",
  19317=>"101100100",
  19318=>"111000000",
  19319=>"110111111",
  19320=>"111101111",
  19321=>"000000110",
  19322=>"111111111",
  19323=>"000001000",
  19324=>"111111111",
  19325=>"000000000",
  19326=>"000100100",
  19327=>"000000000",
  19328=>"000001101",
  19329=>"000000000",
  19330=>"111111111",
  19331=>"111111111",
  19332=>"111111100",
  19333=>"111111000",
  19334=>"000001111",
  19335=>"000000110",
  19336=>"000100111",
  19337=>"011001110",
  19338=>"001011110",
  19339=>"000000000",
  19340=>"111111111",
  19341=>"110110110",
  19342=>"000100100",
  19343=>"000111010",
  19344=>"001000000",
  19345=>"111010000",
  19346=>"000111111",
  19347=>"000000000",
  19348=>"010111111",
  19349=>"011011000",
  19350=>"111111110",
  19351=>"000001011",
  19352=>"000110111",
  19353=>"101111111",
  19354=>"000000001",
  19355=>"100100011",
  19356=>"000000000",
  19357=>"001110010",
  19358=>"111011010",
  19359=>"111111111",
  19360=>"111111111",
  19361=>"000000010",
  19362=>"101001001",
  19363=>"000011111",
  19364=>"001001001",
  19365=>"111111111",
  19366=>"111111101",
  19367=>"000000000",
  19368=>"011111110",
  19369=>"000000100",
  19370=>"111111111",
  19371=>"101111111",
  19372=>"000000000",
  19373=>"001001111",
  19374=>"100000000",
  19375=>"110111111",
  19376=>"111011111",
  19377=>"000110111",
  19378=>"100011000",
  19379=>"111111111",
  19380=>"111111101",
  19381=>"110110000",
  19382=>"000100100",
  19383=>"000111111",
  19384=>"000000000",
  19385=>"110110100",
  19386=>"000000000",
  19387=>"100100000",
  19388=>"000111111",
  19389=>"000110011",
  19390=>"111111111",
  19391=>"111100111",
  19392=>"000000000",
  19393=>"000000000",
  19394=>"111111110",
  19395=>"000100000",
  19396=>"100101111",
  19397=>"110110111",
  19398=>"000000000",
  19399=>"010111111",
  19400=>"000000111",
  19401=>"000000011",
  19402=>"000000010",
  19403=>"000000000",
  19404=>"110100111",
  19405=>"100000000",
  19406=>"100100000",
  19407=>"000111111",
  19408=>"000110110",
  19409=>"011111001",
  19410=>"000100110",
  19411=>"010000000",
  19412=>"111111001",
  19413=>"001110000",
  19414=>"010000110",
  19415=>"000000000",
  19416=>"111111111",
  19417=>"000000000",
  19418=>"000000000",
  19419=>"100000000",
  19420=>"001000000",
  19421=>"111111000",
  19422=>"000001000",
  19423=>"011001001",
  19424=>"000000000",
  19425=>"111000000",
  19426=>"000110111",
  19427=>"111111111",
  19428=>"000000000",
  19429=>"010000000",
  19430=>"111111111",
  19431=>"111111101",
  19432=>"000000000",
  19433=>"000000000",
  19434=>"000111111",
  19435=>"000000000",
  19436=>"111111111",
  19437=>"000110111",
  19438=>"000001011",
  19439=>"101000000",
  19440=>"111000110",
  19441=>"111111111",
  19442=>"000000110",
  19443=>"000000000",
  19444=>"000011000",
  19445=>"000010011",
  19446=>"000000000",
  19447=>"000000000",
  19448=>"000000000",
  19449=>"110111111",
  19450=>"111001111",
  19451=>"100000100",
  19452=>"000001000",
  19453=>"000000000",
  19454=>"111111111",
  19455=>"000000000",
  19456=>"111111010",
  19457=>"000000000",
  19458=>"000111111",
  19459=>"000000000",
  19460=>"111111111",
  19461=>"011011111",
  19462=>"111010111",
  19463=>"000000011",
  19464=>"011000111",
  19465=>"001000000",
  19466=>"000011011",
  19467=>"011000000",
  19468=>"101000000",
  19469=>"000000000",
  19470=>"000101111",
  19471=>"111111011",
  19472=>"000000000",
  19473=>"111111111",
  19474=>"111011000",
  19475=>"000110110",
  19476=>"000000110",
  19477=>"101000001",
  19478=>"000000000",
  19479=>"111111110",
  19480=>"100000000",
  19481=>"111011111",
  19482=>"001011000",
  19483=>"111101111",
  19484=>"111111111",
  19485=>"110110000",
  19486=>"111100100",
  19487=>"000100000",
  19488=>"110110000",
  19489=>"100000000",
  19490=>"000000010",
  19491=>"011111111",
  19492=>"011111001",
  19493=>"111001001",
  19494=>"000000001",
  19495=>"010010000",
  19496=>"111111111",
  19497=>"000111111",
  19498=>"000110111",
  19499=>"011111000",
  19500=>"111111111",
  19501=>"000000010",
  19502=>"010000000",
  19503=>"100000000",
  19504=>"000000011",
  19505=>"000100110",
  19506=>"110110110",
  19507=>"001000110",
  19508=>"011111111",
  19509=>"110111111",
  19510=>"000000000",
  19511=>"111111111",
  19512=>"100100111",
  19513=>"110110110",
  19514=>"111111100",
  19515=>"110110000",
  19516=>"111101111",
  19517=>"110000000",
  19518=>"000001000",
  19519=>"100111111",
  19520=>"100110111",
  19521=>"101111110",
  19522=>"000110010",
  19523=>"010111111",
  19524=>"110111000",
  19525=>"011110110",
  19526=>"011111011",
  19527=>"101111111",
  19528=>"110010000",
  19529=>"111101101",
  19530=>"000000111",
  19531=>"101101101",
  19532=>"110111111",
  19533=>"111101111",
  19534=>"001000101",
  19535=>"000100000",
  19536=>"111111000",
  19537=>"111111111",
  19538=>"000000000",
  19539=>"000001101",
  19540=>"001100000",
  19541=>"000100111",
  19542=>"111111111",
  19543=>"000100111",
  19544=>"000000001",
  19545=>"111111000",
  19546=>"000000001",
  19547=>"111111111",
  19548=>"111001111",
  19549=>"110000000",
  19550=>"000000001",
  19551=>"000000000",
  19552=>"111000000",
  19553=>"110111111",
  19554=>"000000000",
  19555=>"000000111",
  19556=>"010010111",
  19557=>"000000000",
  19558=>"000000111",
  19559=>"111111111",
  19560=>"000000000",
  19561=>"011000000",
  19562=>"010111111",
  19563=>"000000000",
  19564=>"000000000",
  19565=>"000000000",
  19566=>"110000110",
  19567=>"101000000",
  19568=>"111111111",
  19569=>"011110100",
  19570=>"101101111",
  19571=>"000111111",
  19572=>"100111100",
  19573=>"000010000",
  19574=>"001111111",
  19575=>"000110000",
  19576=>"000100100",
  19577=>"010111110",
  19578=>"001001010",
  19579=>"000000100",
  19580=>"101111000",
  19581=>"010110111",
  19582=>"011000000",
  19583=>"000000000",
  19584=>"000000000",
  19585=>"111111111",
  19586=>"011111111",
  19587=>"000000000",
  19588=>"001111111",
  19589=>"111100111",
  19590=>"110111110",
  19591=>"111000000",
  19592=>"100101001",
  19593=>"111111111",
  19594=>"000000000",
  19595=>"110110000",
  19596=>"111111001",
  19597=>"001000000",
  19598=>"111010111",
  19599=>"110110111",
  19600=>"110100100",
  19601=>"111111111",
  19602=>"001000101",
  19603=>"000111111",
  19604=>"111111011",
  19605=>"111000000",
  19606=>"000000100",
  19607=>"000101111",
  19608=>"000000000",
  19609=>"111011001",
  19610=>"110011111",
  19611=>"111110111",
  19612=>"100111001",
  19613=>"000001000",
  19614=>"011101100",
  19615=>"010000000",
  19616=>"001111111",
  19617=>"111111011",
  19618=>"000000110",
  19619=>"110011111",
  19620=>"100000110",
  19621=>"100101100",
  19622=>"000011000",
  19623=>"111101111",
  19624=>"000111001",
  19625=>"110000111",
  19626=>"110111000",
  19627=>"111000000",
  19628=>"111111111",
  19629=>"011101001",
  19630=>"101001000",
  19631=>"111010000",
  19632=>"000000000",
  19633=>"111000000",
  19634=>"010111111",
  19635=>"111000000",
  19636=>"111000000",
  19637=>"111111000",
  19638=>"110100111",
  19639=>"011011000",
  19640=>"111101111",
  19641=>"111111111",
  19642=>"110000001",
  19643=>"000001011",
  19644=>"000000000",
  19645=>"001111001",
  19646=>"000000011",
  19647=>"011111111",
  19648=>"111000000",
  19649=>"111011110",
  19650=>"010000000",
  19651=>"000000000",
  19652=>"000000000",
  19653=>"000110111",
  19654=>"100111111",
  19655=>"000000000",
  19656=>"000000000",
  19657=>"000000111",
  19658=>"110110111",
  19659=>"111000000",
  19660=>"111111100",
  19661=>"010110110",
  19662=>"001001111",
  19663=>"000000000",
  19664=>"011000000",
  19665=>"111111111",
  19666=>"111111011",
  19667=>"010010000",
  19668=>"111111111",
  19669=>"100000000",
  19670=>"011010000",
  19671=>"111111111",
  19672=>"111111000",
  19673=>"000000000",
  19674=>"000000000",
  19675=>"001000000",
  19676=>"001000000",
  19677=>"111000000",
  19678=>"000110111",
  19679=>"111101111",
  19680=>"000000000",
  19681=>"000011011",
  19682=>"011111111",
  19683=>"100110111",
  19684=>"111110100",
  19685=>"111111111",
  19686=>"010000000",
  19687=>"111111111",
  19688=>"001000000",
  19689=>"000110111",
  19690=>"001011010",
  19691=>"111101111",
  19692=>"110100111",
  19693=>"000110110",
  19694=>"000000000",
  19695=>"000000000",
  19696=>"111111111",
  19697=>"111110100",
  19698=>"111001000",
  19699=>"000000000",
  19700=>"111000000",
  19701=>"001000001",
  19702=>"111111000",
  19703=>"000000000",
  19704=>"000000000",
  19705=>"100111001",
  19706=>"000000111",
  19707=>"111111111",
  19708=>"100100000",
  19709=>"111011001",
  19710=>"111111110",
  19711=>"111000000",
  19712=>"100000000",
  19713=>"101001111",
  19714=>"111111111",
  19715=>"111111100",
  19716=>"001000000",
  19717=>"111111111",
  19718=>"000000100",
  19719=>"001001111",
  19720=>"110110111",
  19721=>"000011010",
  19722=>"110010011",
  19723=>"110110111",
  19724=>"001001111",
  19725=>"111111110",
  19726=>"000001001",
  19727=>"111000000",
  19728=>"111000000",
  19729=>"111000000",
  19730=>"111000000",
  19731=>"101001111",
  19732=>"000000001",
  19733=>"011000000",
  19734=>"111111000",
  19735=>"000000000",
  19736=>"010010111",
  19737=>"100000100",
  19738=>"100000000",
  19739=>"100000100",
  19740=>"011100000",
  19741=>"111111111",
  19742=>"111111111",
  19743=>"111001001",
  19744=>"111111101",
  19745=>"111001110",
  19746=>"001100000",
  19747=>"100000110",
  19748=>"000000000",
  19749=>"000000000",
  19750=>"000000011",
  19751=>"000000000",
  19752=>"000000000",
  19753=>"011010011",
  19754=>"000001011",
  19755=>"000000111",
  19756=>"110111111",
  19757=>"001001000",
  19758=>"000000011",
  19759=>"110011011",
  19760=>"010111111",
  19761=>"000000000",
  19762=>"100111111",
  19763=>"000111111",
  19764=>"000000000",
  19765=>"001000000",
  19766=>"000001001",
  19767=>"000111111",
  19768=>"111000000",
  19769=>"111000000",
  19770=>"111111100",
  19771=>"000000000",
  19772=>"110110110",
  19773=>"011000011",
  19774=>"110100000",
  19775=>"000000000",
  19776=>"111111001",
  19777=>"110010000",
  19778=>"000111001",
  19779=>"111110010",
  19780=>"000111111",
  19781=>"000000000",
  19782=>"000000000",
  19783=>"111111001",
  19784=>"010000010",
  19785=>"000000000",
  19786=>"101110111",
  19787=>"011111111",
  19788=>"000000001",
  19789=>"000000111",
  19790=>"000000000",
  19791=>"110111111",
  19792=>"011000100",
  19793=>"001000000",
  19794=>"111011111",
  19795=>"111111111",
  19796=>"000000000",
  19797=>"011001000",
  19798=>"111000010",
  19799=>"111011011",
  19800=>"000000001",
  19801=>"000010010",
  19802=>"111111011",
  19803=>"111111000",
  19804=>"000010110",
  19805=>"111111111",
  19806=>"000000000",
  19807=>"011011011",
  19808=>"000000110",
  19809=>"111000111",
  19810=>"111111011",
  19811=>"111111111",
  19812=>"110110000",
  19813=>"000000011",
  19814=>"111110000",
  19815=>"001001000",
  19816=>"110110110",
  19817=>"000000000",
  19818=>"000000000",
  19819=>"111111111",
  19820=>"111010000",
  19821=>"110000011",
  19822=>"011001001",
  19823=>"000000111",
  19824=>"011111111",
  19825=>"111000000",
  19826=>"111111111",
  19827=>"011001011",
  19828=>"111111111",
  19829=>"000001010",
  19830=>"000111111",
  19831=>"111111000",
  19832=>"000000000",
  19833=>"111111111",
  19834=>"111111111",
  19835=>"101000000",
  19836=>"000010111",
  19837=>"011000000",
  19838=>"001000000",
  19839=>"000000000",
  19840=>"111001111",
  19841=>"101111111",
  19842=>"000010011",
  19843=>"010000000",
  19844=>"110110000",
  19845=>"000000000",
  19846=>"000101110",
  19847=>"001000000",
  19848=>"000000100",
  19849=>"111111111",
  19850=>"111111110",
  19851=>"011000000",
  19852=>"111001111",
  19853=>"100111111",
  19854=>"000000000",
  19855=>"000000000",
  19856=>"111111111",
  19857=>"011010000",
  19858=>"011011010",
  19859=>"111111011",
  19860=>"000000111",
  19861=>"111110110",
  19862=>"001101111",
  19863=>"111111111",
  19864=>"101000000",
  19865=>"111111010",
  19866=>"000001111",
  19867=>"110111111",
  19868=>"001001111",
  19869=>"010000000",
  19870=>"111000110",
  19871=>"111000100",
  19872=>"111010000",
  19873=>"110100100",
  19874=>"100000111",
  19875=>"000000110",
  19876=>"000000000",
  19877=>"110110111",
  19878=>"000000111",
  19879=>"000000100",
  19880=>"000000000",
  19881=>"001001001",
  19882=>"101000111",
  19883=>"000001011",
  19884=>"001111000",
  19885=>"001011010",
  19886=>"110110000",
  19887=>"000000000",
  19888=>"110110000",
  19889=>"111111111",
  19890=>"111001011",
  19891=>"010000011",
  19892=>"111111011",
  19893=>"000001111",
  19894=>"000001001",
  19895=>"111111110",
  19896=>"000010100",
  19897=>"010000111",
  19898=>"000000000",
  19899=>"111111000",
  19900=>"000000000",
  19901=>"111011011",
  19902=>"001001111",
  19903=>"100111110",
  19904=>"000000100",
  19905=>"000000000",
  19906=>"111111111",
  19907=>"000111111",
  19908=>"100111111",
  19909=>"111011111",
  19910=>"111111000",
  19911=>"111000001",
  19912=>"111111110",
  19913=>"110111100",
  19914=>"001111111",
  19915=>"011001111",
  19916=>"000000000",
  19917=>"000001011",
  19918=>"000000000",
  19919=>"111111111",
  19920=>"111111111",
  19921=>"111111111",
  19922=>"011011000",
  19923=>"100000111",
  19924=>"000000000",
  19925=>"111001111",
  19926=>"110111111",
  19927=>"100100100",
  19928=>"000000110",
  19929=>"111111111",
  19930=>"110111111",
  19931=>"100000000",
  19932=>"011111110",
  19933=>"101000100",
  19934=>"000000000",
  19935=>"100100100",
  19936=>"111000001",
  19937=>"111111111",
  19938=>"000000000",
  19939=>"111111111",
  19940=>"000000011",
  19941=>"111101101",
  19942=>"100001011",
  19943=>"000000001",
  19944=>"101111111",
  19945=>"000000000",
  19946=>"100000000",
  19947=>"011011000",
  19948=>"000000001",
  19949=>"011011001",
  19950=>"101101111",
  19951=>"001001001",
  19952=>"111111111",
  19953=>"011111110",
  19954=>"011001000",
  19955=>"011000101",
  19956=>"000111000",
  19957=>"110111110",
  19958=>"000111111",
  19959=>"100111111",
  19960=>"111111011",
  19961=>"111100100",
  19962=>"001000000",
  19963=>"011011111",
  19964=>"110110111",
  19965=>"001100111",
  19966=>"000000000",
  19967=>"100110100",
  19968=>"111111111",
  19969=>"111101011",
  19970=>"000000101",
  19971=>"000100110",
  19972=>"000000001",
  19973=>"100100111",
  19974=>"111111110",
  19975=>"000000000",
  19976=>"000000100",
  19977=>"100100110",
  19978=>"010111111",
  19979=>"100000001",
  19980=>"000000000",
  19981=>"111000000",
  19982=>"000000000",
  19983=>"111111111",
  19984=>"000000001",
  19985=>"110110110",
  19986=>"000000000",
  19987=>"111111111",
  19988=>"100100100",
  19989=>"100100100",
  19990=>"000000010",
  19991=>"100000001",
  19992=>"110111111",
  19993=>"001000000",
  19994=>"111111000",
  19995=>"111111000",
  19996=>"001011111",
  19997=>"111000001",
  19998=>"111011001",
  19999=>"111111110",
  20000=>"000001111",
  20001=>"100000000",
  20002=>"111100000",
  20003=>"111110000",
  20004=>"111111111",
  20005=>"000000011",
  20006=>"111111111",
  20007=>"000101000",
  20008=>"111111111",
  20009=>"110111111",
  20010=>"000000000",
  20011=>"000000010",
  20012=>"111001001",
  20013=>"000100000",
  20014=>"000000000",
  20015=>"101000000",
  20016=>"111111111",
  20017=>"111111111",
  20018=>"101100000",
  20019=>"111111011",
  20020=>"101101101",
  20021=>"100000000",
  20022=>"001111001",
  20023=>"000000100",
  20024=>"000001001",
  20025=>"000000000",
  20026=>"111101100",
  20027=>"010010000",
  20028=>"000000000",
  20029=>"000000000",
  20030=>"000000101",
  20031=>"111111000",
  20032=>"011011011",
  20033=>"000000010",
  20034=>"001111111",
  20035=>"110000000",
  20036=>"111111111",
  20037=>"000000000",
  20038=>"100100111",
  20039=>"111111111",
  20040=>"101001101",
  20041=>"111111111",
  20042=>"000000000",
  20043=>"001000111",
  20044=>"000110110",
  20045=>"000001001",
  20046=>"000110111",
  20047=>"111011001",
  20048=>"111111100",
  20049=>"111111111",
  20050=>"110110111",
  20051=>"000000000",
  20052=>"000000000",
  20053=>"111111011",
  20054=>"111101111",
  20055=>"000000000",
  20056=>"000000000",
  20057=>"000000111",
  20058=>"001110000",
  20059=>"111111111",
  20060=>"000000111",
  20061=>"011000000",
  20062=>"000000000",
  20063=>"111111111",
  20064=>"111111100",
  20065=>"000000111",
  20066=>"111111111",
  20067=>"110000000",
  20068=>"110000010",
  20069=>"111011010",
  20070=>"111100111",
  20071=>"111000001",
  20072=>"001001000",
  20073=>"000011111",
  20074=>"111111000",
  20075=>"000000100",
  20076=>"000000000",
  20077=>"101000000",
  20078=>"000111111",
  20079=>"110110111",
  20080=>"001111111",
  20081=>"111101111",
  20082=>"111111111",
  20083=>"111100101",
  20084=>"000000000",
  20085=>"101000000",
  20086=>"000000111",
  20087=>"000000000",
  20088=>"001000000",
  20089=>"111111111",
  20090=>"101111101",
  20091=>"000000010",
  20092=>"100100000",
  20093=>"011101111",
  20094=>"100000000",
  20095=>"111111111",
  20096=>"000000000",
  20097=>"000010010",
  20098=>"111111111",
  20099=>"000100100",
  20100=>"111111111",
  20101=>"111101000",
  20102=>"101000110",
  20103=>"000000001",
  20104=>"111000000",
  20105=>"011000000",
  20106=>"000100101",
  20107=>"000000000",
  20108=>"111111101",
  20109=>"111111111",
  20110=>"111110000",
  20111=>"111100110",
  20112=>"100000000",
  20113=>"000000000",
  20114=>"000001111",
  20115=>"111101101",
  20116=>"111000000",
  20117=>"000000000",
  20118=>"000000000",
  20119=>"001001101",
  20120=>"001000000",
  20121=>"000000011",
  20122=>"111000000",
  20123=>"011111001",
  20124=>"100000000",
  20125=>"011000111",
  20126=>"111101111",
  20127=>"000000000",
  20128=>"111101111",
  20129=>"011011101",
  20130=>"001000000",
  20131=>"000000000",
  20132=>"000111111",
  20133=>"111111110",
  20134=>"111111111",
  20135=>"111111000",
  20136=>"000000111",
  20137=>"110110010",
  20138=>"111000100",
  20139=>"100000111",
  20140=>"111111000",
  20141=>"001000000",
  20142=>"000000111",
  20143=>"000100000",
  20144=>"110110110",
  20145=>"100000001",
  20146=>"111111011",
  20147=>"001000000",
  20148=>"111111111",
  20149=>"000000001",
  20150=>"111111111",
  20151=>"100111111",
  20152=>"111101111",
  20153=>"110010000",
  20154=>"000000000",
  20155=>"110101100",
  20156=>"100011001",
  20157=>"110100100",
  20158=>"111111111",
  20159=>"111111111",
  20160=>"000000000",
  20161=>"001001001",
  20162=>"111111100",
  20163=>"000000000",
  20164=>"111111111",
  20165=>"001001001",
  20166=>"000100110",
  20167=>"100000001",
  20168=>"000011011",
  20169=>"000001011",
  20170=>"000000001",
  20171=>"111100100",
  20172=>"100000101",
  20173=>"010011011",
  20174=>"101100001",
  20175=>"000000111",
  20176=>"000000000",
  20177=>"000000001",
  20178=>"111001000",
  20179=>"111001000",
  20180=>"001011001",
  20181=>"110111111",
  20182=>"000000010",
  20183=>"000000101",
  20184=>"000000000",
  20185=>"100100111",
  20186=>"111100111",
  20187=>"111111010",
  20188=>"111011101",
  20189=>"000000000",
  20190=>"111111111",
  20191=>"000000000",
  20192=>"000111111",
  20193=>"000000000",
  20194=>"111111000",
  20195=>"000111111",
  20196=>"000000010",
  20197=>"111111111",
  20198=>"101000100",
  20199=>"000000110",
  20200=>"000110110",
  20201=>"111111111",
  20202=>"100100110",
  20203=>"001000000",
  20204=>"111111111",
  20205=>"000000000",
  20206=>"000000100",
  20207=>"000000110",
  20208=>"000000000",
  20209=>"000000000",
  20210=>"001000000",
  20211=>"001000101",
  20212=>"110110010",
  20213=>"100110111",
  20214=>"110110110",
  20215=>"111111111",
  20216=>"111000000",
  20217=>"001000000",
  20218=>"110110110",
  20219=>"000000000",
  20220=>"101101111",
  20221=>"000000101",
  20222=>"000111111",
  20223=>"100000000",
  20224=>"000000000",
  20225=>"000000001",
  20226=>"100000000",
  20227=>"111111110",
  20228=>"111000000",
  20229=>"000000000",
  20230=>"111111110",
  20231=>"111011101",
  20232=>"111111111",
  20233=>"111000000",
  20234=>"101101101",
  20235=>"000000011",
  20236=>"000000000",
  20237=>"000000000",
  20238=>"000000000",
  20239=>"100000000",
  20240=>"000011111",
  20241=>"001001111",
  20242=>"000000000",
  20243=>"000000001",
  20244=>"000000000",
  20245=>"111111111",
  20246=>"001001000",
  20247=>"111111000",
  20248=>"101111111",
  20249=>"000100000",
  20250=>"000111111",
  20251=>"110000000",
  20252=>"110100100",
  20253=>"111101111",
  20254=>"000000000",
  20255=>"111110111",
  20256=>"001000001",
  20257=>"000000000",
  20258=>"111010000",
  20259=>"000000001",
  20260=>"111111000",
  20261=>"111110100",
  20262=>"100000000",
  20263=>"000000001",
  20264=>"000000011",
  20265=>"100111001",
  20266=>"100101001",
  20267=>"000100000",
  20268=>"111111111",
  20269=>"000000000",
  20270=>"000000000",
  20271=>"000000000",
  20272=>"111111110",
  20273=>"000000000",
  20274=>"111111111",
  20275=>"000100000",
  20276=>"000010000",
  20277=>"000100101",
  20278=>"000000001",
  20279=>"111111111",
  20280=>"000000000",
  20281=>"111111111",
  20282=>"000000111",
  20283=>"000000001",
  20284=>"001001101",
  20285=>"101111110",
  20286=>"000000000",
  20287=>"000000000",
  20288=>"000000000",
  20289=>"001111111",
  20290=>"000000111",
  20291=>"010111111",
  20292=>"111111111",
  20293=>"011011001",
  20294=>"001001001",
  20295=>"010110110",
  20296=>"000000000",
  20297=>"111111100",
  20298=>"111111001",
  20299=>"101101101",
  20300=>"000000000",
  20301=>"000000000",
  20302=>"100001111",
  20303=>"100000000",
  20304=>"101000000",
  20305=>"000000000",
  20306=>"000010111",
  20307=>"000000000",
  20308=>"111001111",
  20309=>"001001001",
  20310=>"000000010",
  20311=>"001101111",
  20312=>"111111111",
  20313=>"111111111",
  20314=>"011111111",
  20315=>"000110111",
  20316=>"000001111",
  20317=>"111111111",
  20318=>"110111111",
  20319=>"111111111",
  20320=>"000000000",
  20321=>"001001001",
  20322=>"100110000",
  20323=>"100111111",
  20324=>"000100000",
  20325=>"101001001",
  20326=>"000000000",
  20327=>"000000010",
  20328=>"100100100",
  20329=>"001000111",
  20330=>"000000111",
  20331=>"111101111",
  20332=>"000000110",
  20333=>"001001111",
  20334=>"111101111",
  20335=>"010111000",
  20336=>"000000000",
  20337=>"000010000",
  20338=>"000111111",
  20339=>"100000011",
  20340=>"110100000",
  20341=>"111000000",
  20342=>"011001111",
  20343=>"111111000",
  20344=>"000000011",
  20345=>"000000000",
  20346=>"110010000",
  20347=>"000000100",
  20348=>"000000110",
  20349=>"111111111",
  20350=>"001001000",
  20351=>"000000011",
  20352=>"111011011",
  20353=>"011011011",
  20354=>"000000000",
  20355=>"000100111",
  20356=>"111111111",
  20357=>"000110110",
  20358=>"000110110",
  20359=>"000000100",
  20360=>"000000000",
  20361=>"111000000",
  20362=>"110111111",
  20363=>"000010000",
  20364=>"110111111",
  20365=>"000000000",
  20366=>"111011001",
  20367=>"110000011",
  20368=>"000000010",
  20369=>"111111111",
  20370=>"000000000",
  20371=>"101001000",
  20372=>"111000000",
  20373=>"010010000",
  20374=>"111111111",
  20375=>"110110100",
  20376=>"111111100",
  20377=>"111111111",
  20378=>"010000000",
  20379=>"111111111",
  20380=>"100100110",
  20381=>"111110111",
  20382=>"010001001",
  20383=>"000000000",
  20384=>"000000000",
  20385=>"000000001",
  20386=>"000000111",
  20387=>"000000000",
  20388=>"000001111",
  20389=>"111111111",
  20390=>"000000110",
  20391=>"000000111",
  20392=>"110000000",
  20393=>"100000001",
  20394=>"000000100",
  20395=>"000000001",
  20396=>"010100100",
  20397=>"101000000",
  20398=>"000100111",
  20399=>"100111111",
  20400=>"000000000",
  20401=>"000001111",
  20402=>"000000000",
  20403=>"111000000",
  20404=>"111111111",
  20405=>"111111111",
  20406=>"001101111",
  20407=>"111111111",
  20408=>"000000000",
  20409=>"000010111",
  20410=>"111101111",
  20411=>"001111111",
  20412=>"111111110",
  20413=>"011001001",
  20414=>"000000000",
  20415=>"000000000",
  20416=>"011111110",
  20417=>"111111111",
  20418=>"000000000",
  20419=>"000000111",
  20420=>"000100101",
  20421=>"000000110",
  20422=>"000100000",
  20423=>"000110100",
  20424=>"000000000",
  20425=>"111111111",
  20426=>"000101100",
  20427=>"101000000",
  20428=>"110111000",
  20429=>"001000000",
  20430=>"000000000",
  20431=>"000000100",
  20432=>"000000000",
  20433=>"000000000",
  20434=>"111111111",
  20435=>"111110000",
  20436=>"001000000",
  20437=>"000010111",
  20438=>"111111111",
  20439=>"001011010",
  20440=>"111111111",
  20441=>"000000001",
  20442=>"000000000",
  20443=>"111111111",
  20444=>"011011011",
  20445=>"111000000",
  20446=>"111111111",
  20447=>"000000000",
  20448=>"001001010",
  20449=>"111111111",
  20450=>"000000000",
  20451=>"111111111",
  20452=>"101111111",
  20453=>"011010010",
  20454=>"111111110",
  20455=>"000000000",
  20456=>"111111111",
  20457=>"000000000",
  20458=>"111111111",
  20459=>"110111111",
  20460=>"111000010",
  20461=>"100111000",
  20462=>"000000110",
  20463=>"000001011",
  20464=>"000000101",
  20465=>"111011011",
  20466=>"111001111",
  20467=>"001000111",
  20468=>"101101111",
  20469=>"110000000",
  20470=>"111111111",
  20471=>"001011111",
  20472=>"111111111",
  20473=>"100000100",
  20474=>"111111111",
  20475=>"101000100",
  20476=>"101100000",
  20477=>"111111100",
  20478=>"000000000",
  20479=>"111001111",
  20480=>"000000000",
  20481=>"110000000",
  20482=>"111111111",
  20483=>"111111111",
  20484=>"111111111",
  20485=>"000000011",
  20486=>"000110111",
  20487=>"111111111",
  20488=>"000000111",
  20489=>"111111000",
  20490=>"111001001",
  20491=>"001000000",
  20492=>"111111000",
  20493=>"000000000",
  20494=>"111111011",
  20495=>"011111111",
  20496=>"000000010",
  20497=>"111000000",
  20498=>"111101001",
  20499=>"000000000",
  20500=>"001000000",
  20501=>"111111111",
  20502=>"000000000",
  20503=>"001001001",
  20504=>"111111110",
  20505=>"100111111",
  20506=>"100001111",
  20507=>"010000000",
  20508=>"110000000",
  20509=>"111111001",
  20510=>"111001001",
  20511=>"000000000",
  20512=>"111111111",
  20513=>"110111110",
  20514=>"000000111",
  20515=>"010111000",
  20516=>"111000000",
  20517=>"111110100",
  20518=>"000000000",
  20519=>"000000111",
  20520=>"000000000",
  20521=>"111110000",
  20522=>"101111111",
  20523=>"111111001",
  20524=>"000000001",
  20525=>"000001111",
  20526=>"000000011",
  20527=>"011011001",
  20528=>"011111110",
  20529=>"000000000",
  20530=>"111111111",
  20531=>"000100011",
  20532=>"111111111",
  20533=>"111000110",
  20534=>"111000000",
  20535=>"011011100",
  20536=>"111111111",
  20537=>"000000000",
  20538=>"111111111",
  20539=>"111101111",
  20540=>"111000000",
  20541=>"111111000",
  20542=>"110010000",
  20543=>"011000001",
  20544=>"111011011",
  20545=>"000000000",
  20546=>"000111111",
  20547=>"111111111",
  20548=>"111110000",
  20549=>"000011011",
  20550=>"111111000",
  20551=>"111001000",
  20552=>"011011000",
  20553=>"111111111",
  20554=>"110100111",
  20555=>"111111010",
  20556=>"100110111",
  20557=>"000000000",
  20558=>"000010111",
  20559=>"000010110",
  20560=>"000000000",
  20561=>"111111001",
  20562=>"000000000",
  20563=>"011110110",
  20564=>"000001001",
  20565=>"000000110",
  20566=>"001000001",
  20567=>"001011001",
  20568=>"111111111",
  20569=>"111111111",
  20570=>"000000000",
  20571=>"110110110",
  20572=>"000000111",
  20573=>"111111111",
  20574=>"111111111",
  20575=>"111111100",
  20576=>"111111111",
  20577=>"000000000",
  20578=>"011011001",
  20579=>"000110100",
  20580=>"111111111",
  20581=>"001001111",
  20582=>"001000000",
  20583=>"111111001",
  20584=>"111111111",
  20585=>"101000111",
  20586=>"000000111",
  20587=>"000001011",
  20588=>"010110000",
  20589=>"111111000",
  20590=>"000000000",
  20591=>"001000000",
  20592=>"100000111",
  20593=>"000011111",
  20594=>"010000000",
  20595=>"111111111",
  20596=>"110000000",
  20597=>"111111111",
  20598=>"111111111",
  20599=>"111111111",
  20600=>"111011001",
  20601=>"000000000",
  20602=>"101101111",
  20603=>"100000000",
  20604=>"110110000",
  20605=>"111111111",
  20606=>"000000000",
  20607=>"011001001",
  20608=>"111111111",
  20609=>"000000000",
  20610=>"011000000",
  20611=>"000000001",
  20612=>"000000000",
  20613=>"001000111",
  20614=>"001001000",
  20615=>"100000000",
  20616=>"101000000",
  20617=>"000111111",
  20618=>"000000000",
  20619=>"101000000",
  20620=>"000000000",
  20621=>"000000000",
  20622=>"100001011",
  20623=>"111111000",
  20624=>"000000000",
  20625=>"000000000",
  20626=>"000000000",
  20627=>"100101100",
  20628=>"111001000",
  20629=>"111010001",
  20630=>"000111111",
  20631=>"100111100",
  20632=>"000000000",
  20633=>"111000000",
  20634=>"000000000",
  20635=>"000000000",
  20636=>"000000000",
  20637=>"111111111",
  20638=>"010011111",
  20639=>"011101111",
  20640=>"001001000",
  20641=>"111011011",
  20642=>"000111111",
  20643=>"000110110",
  20644=>"000000000",
  20645=>"111111111",
  20646=>"101101111",
  20647=>"111101100",
  20648=>"000010000",
  20649=>"100101000",
  20650=>"111111111",
  20651=>"001001011",
  20652=>"001001000",
  20653=>"000100111",
  20654=>"000000001",
  20655=>"000000001",
  20656=>"111111000",
  20657=>"011011111",
  20658=>"111111000",
  20659=>"001101101",
  20660=>"001101111",
  20661=>"010111111",
  20662=>"000000101",
  20663=>"000110111",
  20664=>"111110100",
  20665=>"111111111",
  20666=>"001001011",
  20667=>"011000000",
  20668=>"111001000",
  20669=>"010110111",
  20670=>"000000111",
  20671=>"000000000",
  20672=>"111111000",
  20673=>"111001111",
  20674=>"010111011",
  20675=>"111000000",
  20676=>"111011000",
  20677=>"111001000",
  20678=>"000000000",
  20679=>"000000000",
  20680=>"101000001",
  20681=>"110000000",
  20682=>"000000000",
  20683=>"000000000",
  20684=>"001001110",
  20685=>"111111111",
  20686=>"111111111",
  20687=>"000000000",
  20688=>"000000000",
  20689=>"000000000",
  20690=>"000000111",
  20691=>"000000000",
  20692=>"000000001",
  20693=>"110000100",
  20694=>"111000000",
  20695=>"000000000",
  20696=>"111111111",
  20697=>"000011111",
  20698=>"111111100",
  20699=>"001000000",
  20700=>"110000000",
  20701=>"100000001",
  20702=>"000000000",
  20703=>"111111111",
  20704=>"110000000",
  20705=>"000000010",
  20706=>"111111010",
  20707=>"000000000",
  20708=>"111011111",
  20709=>"100111111",
  20710=>"110110000",
  20711=>"000000111",
  20712=>"101000000",
  20713=>"111111101",
  20714=>"101110000",
  20715=>"011001000",
  20716=>"000000000",
  20717=>"111100000",
  20718=>"111000000",
  20719=>"111011111",
  20720=>"000000100",
  20721=>"111111111",
  20722=>"111111011",
  20723=>"000000010",
  20724=>"000000110",
  20725=>"111111110",
  20726=>"100100110",
  20727=>"111111111",
  20728=>"111111100",
  20729=>"000000000",
  20730=>"011010010",
  20731=>"111111111",
  20732=>"111110110",
  20733=>"001000000",
  20734=>"000000000",
  20735=>"111111100",
  20736=>"111000000",
  20737=>"111111000",
  20738=>"000000011",
  20739=>"000100111",
  20740=>"111111111",
  20741=>"111111111",
  20742=>"001000000",
  20743=>"101000000",
  20744=>"110110001",
  20745=>"000000000",
  20746=>"101100000",
  20747=>"111111000",
  20748=>"000000000",
  20749=>"001111011",
  20750=>"110111001",
  20751=>"001001000",
  20752=>"111000000",
  20753=>"000011111",
  20754=>"000000111",
  20755=>"111111111",
  20756=>"000000000",
  20757=>"111111111",
  20758=>"011000000",
  20759=>"000000000",
  20760=>"011011111",
  20761=>"111111111",
  20762=>"111100000",
  20763=>"111111111",
  20764=>"001000000",
  20765=>"000000000",
  20766=>"000000011",
  20767=>"110111001",
  20768=>"111111000",
  20769=>"000000000",
  20770=>"000011000",
  20771=>"000000000",
  20772=>"111111111",
  20773=>"011011111",
  20774=>"001000001",
  20775=>"000000000",
  20776=>"111111111",
  20777=>"001001111",
  20778=>"000111111",
  20779=>"000000000",
  20780=>"010010000",
  20781=>"111111011",
  20782=>"000000101",
  20783=>"000100000",
  20784=>"010000000",
  20785=>"011111111",
  20786=>"111111000",
  20787=>"000000000",
  20788=>"111000000",
  20789=>"111101000",
  20790=>"000000000",
  20791=>"111001001",
  20792=>"111111111",
  20793=>"111001111",
  20794=>"000111111",
  20795=>"111111111",
  20796=>"011011001",
  20797=>"011000000",
  20798=>"001111111",
  20799=>"000000001",
  20800=>"000000000",
  20801=>"000000000",
  20802=>"011111111",
  20803=>"000100110",
  20804=>"000000000",
  20805=>"111111100",
  20806=>"111101100",
  20807=>"111110100",
  20808=>"111101100",
  20809=>"000000011",
  20810=>"110011001",
  20811=>"011111110",
  20812=>"000000111",
  20813=>"100111111",
  20814=>"000000001",
  20815=>"101101111",
  20816=>"111111110",
  20817=>"000000011",
  20818=>"111111111",
  20819=>"110110111",
  20820=>"100000000",
  20821=>"011011000",
  20822=>"000111111",
  20823=>"001000000",
  20824=>"000100111",
  20825=>"000010110",
  20826=>"111000000",
  20827=>"000011111",
  20828=>"000000000",
  20829=>"000010110",
  20830=>"000000111",
  20831=>"000000100",
  20832=>"000000101",
  20833=>"000000111",
  20834=>"111111110",
  20835=>"100000000",
  20836=>"111111111",
  20837=>"000011011",
  20838=>"000000000",
  20839=>"000000000",
  20840=>"100100000",
  20841=>"111000000",
  20842=>"111000000",
  20843=>"110110000",
  20844=>"111101000",
  20845=>"111101000",
  20846=>"000000110",
  20847=>"000111111",
  20848=>"000000110",
  20849=>"000011111",
  20850=>"000000111",
  20851=>"000111011",
  20852=>"111111010",
  20853=>"111000111",
  20854=>"000000000",
  20855=>"000000000",
  20856=>"000000111",
  20857=>"000000000",
  20858=>"000000000",
  20859=>"000001001",
  20860=>"001000000",
  20861=>"011111111",
  20862=>"011111001",
  20863=>"000000111",
  20864=>"111111111",
  20865=>"111111000",
  20866=>"110110110",
  20867=>"100110011",
  20868=>"111011111",
  20869=>"010010000",
  20870=>"011000000",
  20871=>"111000000",
  20872=>"100000100",
  20873=>"000000000",
  20874=>"100111111",
  20875=>"100100010",
  20876=>"100100100",
  20877=>"000110110",
  20878=>"111110000",
  20879=>"000110010",
  20880=>"001000000",
  20881=>"010100111",
  20882=>"111111111",
  20883=>"000000000",
  20884=>"000000111",
  20885=>"111000000",
  20886=>"000000010",
  20887=>"111111111",
  20888=>"111011000",
  20889=>"111111111",
  20890=>"000001111",
  20891=>"011111111",
  20892=>"001111110",
  20893=>"011111111",
  20894=>"100001000",
  20895=>"111111111",
  20896=>"111111111",
  20897=>"110001000",
  20898=>"010010000",
  20899=>"011111001",
  20900=>"001001001",
  20901=>"111111111",
  20902=>"111000111",
  20903=>"111100000",
  20904=>"011000000",
  20905=>"000000001",
  20906=>"000000000",
  20907=>"000000000",
  20908=>"000000000",
  20909=>"000000000",
  20910=>"000000000",
  20911=>"000000111",
  20912=>"101111111",
  20913=>"111001000",
  20914=>"000000000",
  20915=>"111101001",
  20916=>"000110100",
  20917=>"000000111",
  20918=>"000000111",
  20919=>"000000000",
  20920=>"010000000",
  20921=>"001000000",
  20922=>"000000011",
  20923=>"011001111",
  20924=>"111111011",
  20925=>"111100000",
  20926=>"000001001",
  20927=>"000000000",
  20928=>"000000111",
  20929=>"100100000",
  20930=>"111111111",
  20931=>"011000100",
  20932=>"111000000",
  20933=>"011001000",
  20934=>"000111111",
  20935=>"001001000",
  20936=>"000000000",
  20937=>"100101111",
  20938=>"000000110",
  20939=>"111000000",
  20940=>"010000000",
  20941=>"111110000",
  20942=>"101000000",
  20943=>"000111111",
  20944=>"111000000",
  20945=>"000000000",
  20946=>"111111111",
  20947=>"100101111",
  20948=>"000000111",
  20949=>"111000000",
  20950=>"000000000",
  20951=>"111001001",
  20952=>"111000100",
  20953=>"111000000",
  20954=>"111111111",
  20955=>"001001001",
  20956=>"000000000",
  20957=>"000000001",
  20958=>"111000000",
  20959=>"000111111",
  20960=>"101001000",
  20961=>"111111111",
  20962=>"000111111",
  20963=>"000110000",
  20964=>"111111111",
  20965=>"000001111",
  20966=>"000000000",
  20967=>"000000000",
  20968=>"111111111",
  20969=>"111000000",
  20970=>"000000000",
  20971=>"000000111",
  20972=>"000000000",
  20973=>"101101101",
  20974=>"000100001",
  20975=>"111001000",
  20976=>"100100000",
  20977=>"000111111",
  20978=>"000000001",
  20979=>"111111000",
  20980=>"001001010",
  20981=>"000111111",
  20982=>"000000100",
  20983=>"001001001",
  20984=>"111111000",
  20985=>"001001000",
  20986=>"111000000",
  20987=>"001001001",
  20988=>"111001100",
  20989=>"001000000",
  20990=>"111011011",
  20991=>"000000100",
  20992=>"111001001",
  20993=>"000000000",
  20994=>"111111110",
  20995=>"010011011",
  20996=>"000000000",
  20997=>"100101000",
  20998=>"111000011",
  20999=>"001111111",
  21000=>"110111000",
  21001=>"110111111",
  21002=>"101101101",
  21003=>"010000001",
  21004=>"100000111",
  21005=>"000000101",
  21006=>"000001001",
  21007=>"101000111",
  21008=>"001001001",
  21009=>"111111111",
  21010=>"111111111",
  21011=>"000111111",
  21012=>"110111111",
  21013=>"010000101",
  21014=>"111001111",
  21015=>"011110100",
  21016=>"000000001",
  21017=>"100100010",
  21018=>"000000101",
  21019=>"110111111",
  21020=>"001111111",
  21021=>"111111111",
  21022=>"100000001",
  21023=>"000000001",
  21024=>"000000001",
  21025=>"110111111",
  21026=>"100100000",
  21027=>"111100000",
  21028=>"000000101",
  21029=>"110110010",
  21030=>"110000111",
  21031=>"000000111",
  21032=>"001000101",
  21033=>"010011000",
  21034=>"000000000",
  21035=>"101101111",
  21036=>"000001000",
  21037=>"011001000",
  21038=>"001111111",
  21039=>"000000101",
  21040=>"001001111",
  21041=>"001001111",
  21042=>"110111010",
  21043=>"010110010",
  21044=>"111101111",
  21045=>"100000100",
  21046=>"111000000",
  21047=>"000000111",
  21048=>"000000000",
  21049=>"001001011",
  21050=>"111111000",
  21051=>"111111110",
  21052=>"101101101",
  21053=>"111000000",
  21054=>"111111111",
  21055=>"000000000",
  21056=>"111111111",
  21057=>"001110111",
  21058=>"111010000",
  21059=>"000000000",
  21060=>"100000000",
  21061=>"001000110",
  21062=>"000000000",
  21063=>"101111111",
  21064=>"110110110",
  21065=>"000100111",
  21066=>"000000000",
  21067=>"000001001",
  21068=>"000011001",
  21069=>"010000000",
  21070=>"100110000",
  21071=>"110111111",
  21072=>"111111010",
  21073=>"001000100",
  21074=>"111000110",
  21075=>"001001101",
  21076=>"111000000",
  21077=>"000000000",
  21078=>"101001010",
  21079=>"100001111",
  21080=>"000011111",
  21081=>"001001001",
  21082=>"110000000",
  21083=>"110111010",
  21084=>"010010010",
  21085=>"000000111",
  21086=>"000000101",
  21087=>"000100100",
  21088=>"011001000",
  21089=>"000000000",
  21090=>"100100110",
  21091=>"000101000",
  21092=>"000000000",
  21093=>"000000010",
  21094=>"000000110",
  21095=>"000000000",
  21096=>"000000000",
  21097=>"000001111",
  21098=>"010010111",
  21099=>"010100110",
  21100=>"101000100",
  21101=>"110010000",
  21102=>"111110111",
  21103=>"000110110",
  21104=>"000000000",
  21105=>"001001000",
  21106=>"101111101",
  21107=>"000000000",
  21108=>"001000111",
  21109=>"110111111",
  21110=>"000001000",
  21111=>"111111111",
  21112=>"000111111",
  21113=>"001111111",
  21114=>"010010000",
  21115=>"010000010",
  21116=>"100110111",
  21117=>"000001111",
  21118=>"111111000",
  21119=>"000000000",
  21120=>"111000000",
  21121=>"100000111",
  21122=>"000001000",
  21123=>"001001111",
  21124=>"101001001",
  21125=>"110000001",
  21126=>"110100000",
  21127=>"100001001",
  21128=>"000111111",
  21129=>"000000000",
  21130=>"000001000",
  21131=>"000000111",
  21132=>"111110001",
  21133=>"000000101",
  21134=>"111111111",
  21135=>"110000000",
  21136=>"100000000",
  21137=>"001001000",
  21138=>"100111111",
  21139=>"000000000",
  21140=>"001000011",
  21141=>"000010000",
  21142=>"000000111",
  21143=>"100000111",
  21144=>"001001111",
  21145=>"000001111",
  21146=>"000000101",
  21147=>"001011000",
  21148=>"111010111",
  21149=>"000110000",
  21150=>"000000110",
  21151=>"010001011",
  21152=>"111100110",
  21153=>"111001000",
  21154=>"111111110",
  21155=>"110000000",
  21156=>"111110010",
  21157=>"111000011",
  21158=>"000010000",
  21159=>"011000000",
  21160=>"000000000",
  21161=>"000001000",
  21162=>"010010000",
  21163=>"000000000",
  21164=>"101111111",
  21165=>"100111100",
  21166=>"100000010",
  21167=>"000100100",
  21168=>"111000111",
  21169=>"000000100",
  21170=>"111111110",
  21171=>"011001011",
  21172=>"000110011",
  21173=>"001001001",
  21174=>"000000111",
  21175=>"000000000",
  21176=>"111111111",
  21177=>"111111101",
  21178=>"000100100",
  21179=>"000001000",
  21180=>"110111010",
  21181=>"110110111",
  21182=>"000111111",
  21183=>"101001111",
  21184=>"111001000",
  21185=>"111111110",
  21186=>"001000000",
  21187=>"100000000",
  21188=>"001000000",
  21189=>"000101111",
  21190=>"011010110",
  21191=>"111111010",
  21192=>"000011011",
  21193=>"000001100",
  21194=>"000000100",
  21195=>"111001001",
  21196=>"110000000",
  21197=>"111011000",
  21198=>"111110110",
  21199=>"000011111",
  21200=>"111100000",
  21201=>"111111111",
  21202=>"000111000",
  21203=>"010011011",
  21204=>"111111111",
  21205=>"110000001",
  21206=>"000000000",
  21207=>"001000000",
  21208=>"111111000",
  21209=>"010000110",
  21210=>"111111111",
  21211=>"110100111",
  21212=>"110100101",
  21213=>"000000000",
  21214=>"111000000",
  21215=>"101001001",
  21216=>"111000000",
  21217=>"000000000",
  21218=>"000000110",
  21219=>"111110000",
  21220=>"000000000",
  21221=>"010111011",
  21222=>"010000010",
  21223=>"000001001",
  21224=>"011011000",
  21225=>"000111000",
  21226=>"111111011",
  21227=>"111111010",
  21228=>"111001000",
  21229=>"111010000",
  21230=>"001101101",
  21231=>"100111000",
  21232=>"111101111",
  21233=>"011000001",
  21234=>"000000000",
  21235=>"000001111",
  21236=>"111001001",
  21237=>"011011001",
  21238=>"111010001",
  21239=>"100000000",
  21240=>"011111111",
  21241=>"111111111",
  21242=>"001001000",
  21243=>"101111101",
  21244=>"001110110",
  21245=>"110000000",
  21246=>"010010000",
  21247=>"111000000",
  21248=>"111001001",
  21249=>"000001001",
  21250=>"000100110",
  21251=>"111000000",
  21252=>"000000001",
  21253=>"000000000",
  21254=>"010010111",
  21255=>"111000000",
  21256=>"100000111",
  21257=>"111111001",
  21258=>"000111110",
  21259=>"111000000",
  21260=>"001000111",
  21261=>"111111111",
  21262=>"111111011",
  21263=>"111100000",
  21264=>"000010000",
  21265=>"110001000",
  21266=>"000000000",
  21267=>"110100111",
  21268=>"000111111",
  21269=>"000000000",
  21270=>"110111000",
  21271=>"111000000",
  21272=>"111110010",
  21273=>"000000111",
  21274=>"110111111",
  21275=>"000000001",
  21276=>"000110111",
  21277=>"000001111",
  21278=>"011111111",
  21279=>"110100000",
  21280=>"000100100",
  21281=>"101000000",
  21282=>"110110110",
  21283=>"111111111",
  21284=>"010111111",
  21285=>"000001100",
  21286=>"100110100",
  21287=>"011111111",
  21288=>"000110101",
  21289=>"011011011",
  21290=>"000000000",
  21291=>"000000101",
  21292=>"111100110",
  21293=>"000000111",
  21294=>"100011000",
  21295=>"000011011",
  21296=>"000000111",
  21297=>"111111110",
  21298=>"001111111",
  21299=>"000000110",
  21300=>"111111000",
  21301=>"110111111",
  21302=>"000000000",
  21303=>"100000000",
  21304=>"000110111",
  21305=>"000111101",
  21306=>"010010000",
  21307=>"111111011",
  21308=>"100000000",
  21309=>"101000000",
  21310=>"000001111",
  21311=>"111111110",
  21312=>"001001001",
  21313=>"001000000",
  21314=>"001000110",
  21315=>"011011000",
  21316=>"101000101",
  21317=>"111111000",
  21318=>"111111111",
  21319=>"110111111",
  21320=>"000000000",
  21321=>"000000000",
  21322=>"000000000",
  21323=>"000100000",
  21324=>"000000001",
  21325=>"000000111",
  21326=>"111111111",
  21327=>"011110110",
  21328=>"111000000",
  21329=>"000000111",
  21330=>"111111111",
  21331=>"001000111",
  21332=>"000000001",
  21333=>"000000000",
  21334=>"000000000",
  21335=>"001000111",
  21336=>"111111110",
  21337=>"010010000",
  21338=>"111101100",
  21339=>"001001101",
  21340=>"010111010",
  21341=>"000011111",
  21342=>"001011000",
  21343=>"000000111",
  21344=>"110110000",
  21345=>"111000001",
  21346=>"111100100",
  21347=>"000101101",
  21348=>"110100110",
  21349=>"100000001",
  21350=>"111111111",
  21351=>"111111000",
  21352=>"001001111",
  21353=>"100111000",
  21354=>"001001000",
  21355=>"111111111",
  21356=>"010000000",
  21357=>"111000010",
  21358=>"001011001",
  21359=>"001000100",
  21360=>"000001000",
  21361=>"111001111",
  21362=>"000010111",
  21363=>"111001001",
  21364=>"111111001",
  21365=>"111001010",
  21366=>"000000010",
  21367=>"111110000",
  21368=>"000000000",
  21369=>"000100110",
  21370=>"001000101",
  21371=>"110111110",
  21372=>"111111111",
  21373=>"111000111",
  21374=>"110110110",
  21375=>"111110000",
  21376=>"100100111",
  21377=>"000001000",
  21378=>"100000001",
  21379=>"000010010",
  21380=>"000110000",
  21381=>"001000000",
  21382=>"010111111",
  21383=>"011011000",
  21384=>"000011000",
  21385=>"111111000",
  21386=>"000000000",
  21387=>"011011001",
  21388=>"000000000",
  21389=>"111111011",
  21390=>"100000010",
  21391=>"011011001",
  21392=>"111111000",
  21393=>"101101101",
  21394=>"001011111",
  21395=>"010000000",
  21396=>"010110111",
  21397=>"000000010",
  21398=>"110110110",
  21399=>"111101100",
  21400=>"010111111",
  21401=>"010000000",
  21402=>"000001111",
  21403=>"000111111",
  21404=>"000000100",
  21405=>"111001111",
  21406=>"110000111",
  21407=>"000100111",
  21408=>"001000001",
  21409=>"001001000",
  21410=>"111000111",
  21411=>"000000000",
  21412=>"000000000",
  21413=>"111111111",
  21414=>"000000000",
  21415=>"101111000",
  21416=>"000101111",
  21417=>"000101110",
  21418=>"100101101",
  21419=>"111001101",
  21420=>"000010000",
  21421=>"000001111",
  21422=>"111111010",
  21423=>"110010010",
  21424=>"111110000",
  21425=>"001000111",
  21426=>"110111011",
  21427=>"100000010",
  21428=>"100000000",
  21429=>"000000000",
  21430=>"111111111",
  21431=>"000001000",
  21432=>"010110110",
  21433=>"110111111",
  21434=>"011000011",
  21435=>"010010111",
  21436=>"000000000",
  21437=>"000000111",
  21438=>"000000000",
  21439=>"100001101",
  21440=>"010110010",
  21441=>"001111000",
  21442=>"011111001",
  21443=>"111000000",
  21444=>"100000110",
  21445=>"110101111",
  21446=>"000000111",
  21447=>"000110100",
  21448=>"010000000",
  21449=>"110000111",
  21450=>"000000100",
  21451=>"000000001",
  21452=>"000000111",
  21453=>"110000010",
  21454=>"100000000",
  21455=>"000000101",
  21456=>"000111000",
  21457=>"000000000",
  21458=>"110000010",
  21459=>"000100110",
  21460=>"101101011",
  21461=>"110000111",
  21462=>"011111111",
  21463=>"111000000",
  21464=>"100000100",
  21465=>"111001111",
  21466=>"100000000",
  21467=>"110110110",
  21468=>"010110111",
  21469=>"000100100",
  21470=>"111111000",
  21471=>"110010010",
  21472=>"101000000",
  21473=>"111111111",
  21474=>"000000001",
  21475=>"101000000",
  21476=>"010111100",
  21477=>"000000111",
  21478=>"000000000",
  21479=>"001001000",
  21480=>"111001100",
  21481=>"110100101",
  21482=>"010111111",
  21483=>"011011011",
  21484=>"000000000",
  21485=>"111111011",
  21486=>"101111111",
  21487=>"001001101",
  21488=>"010000000",
  21489=>"111111110",
  21490=>"100000000",
  21491=>"000011001",
  21492=>"001011111",
  21493=>"111111000",
  21494=>"100000000",
  21495=>"110110100",
  21496=>"011010000",
  21497=>"011110000",
  21498=>"100110111",
  21499=>"001001111",
  21500=>"010011111",
  21501=>"110000110",
  21502=>"110111110",
  21503=>"001111111",
  21504=>"000000000",
  21505=>"000000000",
  21506=>"000000101",
  21507=>"111111100",
  21508=>"000000000",
  21509=>"111011000",
  21510=>"111111110",
  21511=>"000000000",
  21512=>"011111111",
  21513=>"111001000",
  21514=>"000000000",
  21515=>"110111111",
  21516=>"010110110",
  21517=>"101101100",
  21518=>"111111000",
  21519=>"000000111",
  21520=>"000000000",
  21521=>"111111110",
  21522=>"000111111",
  21523=>"001001111",
  21524=>"000001001",
  21525=>"000000000",
  21526=>"000000001",
  21527=>"011011011",
  21528=>"111111000",
  21529=>"011011001",
  21530=>"111101111",
  21531=>"101001001",
  21532=>"000000000",
  21533=>"001000111",
  21534=>"000011111",
  21535=>"000111111",
  21536=>"001000100",
  21537=>"000000001",
  21538=>"000010000",
  21539=>"000000000",
  21540=>"000000000",
  21541=>"000000000",
  21542=>"111111111",
  21543=>"011000000",
  21544=>"011111101",
  21545=>"000001111",
  21546=>"000000000",
  21547=>"111111110",
  21548=>"000000111",
  21549=>"000100000",
  21550=>"011000000",
  21551=>"001000001",
  21552=>"001000011",
  21553=>"110110110",
  21554=>"000001000",
  21555=>"000110100",
  21556=>"011001011",
  21557=>"000000100",
  21558=>"100000000",
  21559=>"000000000",
  21560=>"111110100",
  21561=>"000110111",
  21562=>"000110010",
  21563=>"001010111",
  21564=>"000000111",
  21565=>"001001011",
  21566=>"011111101",
  21567=>"000000111",
  21568=>"000000000",
  21569=>"000000001",
  21570=>"000000000",
  21571=>"111111011",
  21572=>"110010000",
  21573=>"110000000",
  21574=>"111111111",
  21575=>"111101101",
  21576=>"000001011",
  21577=>"000011011",
  21578=>"000000000",
  21579=>"111111011",
  21580=>"010000001",
  21581=>"000000100",
  21582=>"000000010",
  21583=>"111111110",
  21584=>"000000000",
  21585=>"111011001",
  21586=>"111111000",
  21587=>"000000000",
  21588=>"110110110",
  21589=>"000000011",
  21590=>"000000011",
  21591=>"000000000",
  21592=>"111111111",
  21593=>"000000111",
  21594=>"000000000",
  21595=>"111111110",
  21596=>"101101111",
  21597=>"001000001",
  21598=>"010010111",
  21599=>"111111111",
  21600=>"000000000",
  21601=>"000000000",
  21602=>"110000111",
  21603=>"000000000",
  21604=>"111111111",
  21605=>"111111111",
  21606=>"111011010",
  21607=>"110000110",
  21608=>"011111000",
  21609=>"001001011",
  21610=>"001001100",
  21611=>"000001111",
  21612=>"011011000",
  21613=>"000000101",
  21614=>"000011000",
  21615=>"010011010",
  21616=>"111111010",
  21617=>"101000000",
  21618=>"011001101",
  21619=>"000000110",
  21620=>"111110000",
  21621=>"111111111",
  21622=>"000000111",
  21623=>"010011111",
  21624=>"001000000",
  21625=>"000000000",
  21626=>"000011111",
  21627=>"000000000",
  21628=>"100110000",
  21629=>"000000000",
  21630=>"000000011",
  21631=>"111111111",
  21632=>"000100111",
  21633=>"000000011",
  21634=>"010000000",
  21635=>"100101100",
  21636=>"101000000",
  21637=>"000000000",
  21638=>"111100000",
  21639=>"000000001",
  21640=>"111111100",
  21641=>"000000000",
  21642=>"100111111",
  21643=>"001111110",
  21644=>"111011011",
  21645=>"111111000",
  21646=>"000111111",
  21647=>"111111000",
  21648=>"000000000",
  21649=>"111110110",
  21650=>"111000000",
  21651=>"000000000",
  21652=>"000000100",
  21653=>"111111111",
  21654=>"001111111",
  21655=>"111001000",
  21656=>"001011111",
  21657=>"000000000",
  21658=>"011010110",
  21659=>"000000000",
  21660=>"010000000",
  21661=>"000000000",
  21662=>"111111111",
  21663=>"011111111",
  21664=>"000000111",
  21665=>"000000001",
  21666=>"111110000",
  21667=>"000010110",
  21668=>"000011111",
  21669=>"000001001",
  21670=>"111000111",
  21671=>"111101101",
  21672=>"111011001",
  21673=>"000000000",
  21674=>"011000110",
  21675=>"111111111",
  21676=>"110110110",
  21677=>"111111111",
  21678=>"000010111",
  21679=>"001111111",
  21680=>"111110110",
  21681=>"100100100",
  21682=>"111111111",
  21683=>"110000000",
  21684=>"000000111",
  21685=>"110110111",
  21686=>"000000000",
  21687=>"000000100",
  21688=>"000000111",
  21689=>"000001001",
  21690=>"100000011",
  21691=>"011011111",
  21692=>"001111001",
  21693=>"111111000",
  21694=>"100000000",
  21695=>"000000001",
  21696=>"000000000",
  21697=>"000001001",
  21698=>"000011111",
  21699=>"111111111",
  21700=>"001001111",
  21701=>"001101111",
  21702=>"001001001",
  21703=>"101000101",
  21704=>"011110110",
  21705=>"011001101",
  21706=>"111111011",
  21707=>"000011000",
  21708=>"001111111",
  21709=>"000011011",
  21710=>"000000000",
  21711=>"111111010",
  21712=>"000100000",
  21713=>"011110010",
  21714=>"110110110",
  21715=>"111011000",
  21716=>"111110000",
  21717=>"111111000",
  21718=>"011011011",
  21719=>"000000010",
  21720=>"000111111",
  21721=>"100000000",
  21722=>"000000000",
  21723=>"000111111",
  21724=>"111111111",
  21725=>"111111101",
  21726=>"111111111",
  21727=>"000000100",
  21728=>"111100111",
  21729=>"111111111",
  21730=>"111111111",
  21731=>"100101111",
  21732=>"000000001",
  21733=>"011011011",
  21734=>"110110101",
  21735=>"011111111",
  21736=>"000001100",
  21737=>"101101100",
  21738=>"111110110",
  21739=>"000001001",
  21740=>"111010000",
  21741=>"111111111",
  21742=>"110101000",
  21743=>"000000000",
  21744=>"100111111",
  21745=>"110000100",
  21746=>"111111111",
  21747=>"111000000",
  21748=>"111111110",
  21749=>"111111111",
  21750=>"000000001",
  21751=>"111111001",
  21752=>"010000000",
  21753=>"000000001",
  21754=>"110000110",
  21755=>"011111111",
  21756=>"110110110",
  21757=>"000000000",
  21758=>"100111101",
  21759=>"110010000",
  21760=>"000000000",
  21761=>"001001101",
  21762=>"000000101",
  21763=>"100111100",
  21764=>"000111111",
  21765=>"110110010",
  21766=>"000000011",
  21767=>"000010000",
  21768=>"000000000",
  21769=>"000000000",
  21770=>"111001000",
  21771=>"111001111",
  21772=>"001001001",
  21773=>"111111001",
  21774=>"000000011",
  21775=>"001011111",
  21776=>"000000000",
  21777=>"000000110",
  21778=>"001000001",
  21779=>"000000000",
  21780=>"000000100",
  21781=>"000000000",
  21782=>"000000000",
  21783=>"000000001",
  21784=>"111111011",
  21785=>"111111111",
  21786=>"000001001",
  21787=>"110010110",
  21788=>"110110110",
  21789=>"111000000",
  21790=>"000010000",
  21791=>"000000001",
  21792=>"000010110",
  21793=>"011011000",
  21794=>"000000000",
  21795=>"101001001",
  21796=>"110110110",
  21797=>"000000110",
  21798=>"111111011",
  21799=>"111111111",
  21800=>"111111111",
  21801=>"111111010",
  21802=>"000000010",
  21803=>"011000000",
  21804=>"010001101",
  21805=>"111111111",
  21806=>"100010010",
  21807=>"000100111",
  21808=>"000000010",
  21809=>"011011001",
  21810=>"110000000",
  21811=>"110111111",
  21812=>"001010000",
  21813=>"011111111",
  21814=>"000000000",
  21815=>"111111111",
  21816=>"001000111",
  21817=>"111001001",
  21818=>"110111000",
  21819=>"001111111",
  21820=>"110000000",
  21821=>"111111110",
  21822=>"100100000",
  21823=>"100000000",
  21824=>"000100000",
  21825=>"111111111",
  21826=>"001011111",
  21827=>"000000000",
  21828=>"000000001",
  21829=>"001000000",
  21830=>"111111111",
  21831=>"000001011",
  21832=>"111111111",
  21833=>"110110010",
  21834=>"100111001",
  21835=>"010000000",
  21836=>"111110100",
  21837=>"000000111",
  21838=>"000000100",
  21839=>"111111111",
  21840=>"111111111",
  21841=>"111000011",
  21842=>"111111111",
  21843=>"111111101",
  21844=>"000000110",
  21845=>"001011001",
  21846=>"110011000",
  21847=>"000001011",
  21848=>"111111111",
  21849=>"111011000",
  21850=>"011110000",
  21851=>"111111111",
  21852=>"000000001",
  21853=>"000111111",
  21854=>"000000000",
  21855=>"011001111",
  21856=>"000000000",
  21857=>"101110110",
  21858=>"110110000",
  21859=>"001000101",
  21860=>"111111111",
  21861=>"000000000",
  21862=>"000100001",
  21863=>"111111111",
  21864=>"011001001",
  21865=>"111001111",
  21866=>"000111000",
  21867=>"011111111",
  21868=>"000000000",
  21869=>"111001011",
  21870=>"100110000",
  21871=>"110100000",
  21872=>"000100111",
  21873=>"000110100",
  21874=>"111111111",
  21875=>"011011011",
  21876=>"000000100",
  21877=>"000000111",
  21878=>"111011000",
  21879=>"111001000",
  21880=>"100000000",
  21881=>"111111111",
  21882=>"000000111",
  21883=>"110000000",
  21884=>"000010110",
  21885=>"111111010",
  21886=>"111111000",
  21887=>"111111111",
  21888=>"000000000",
  21889=>"000000010",
  21890=>"110000000",
  21891=>"111111111",
  21892=>"111111111",
  21893=>"011111000",
  21894=>"111111110",
  21895=>"001011011",
  21896=>"100000000",
  21897=>"111111111",
  21898=>"111111011",
  21899=>"001001001",
  21900=>"101101111",
  21901=>"111111111",
  21902=>"000000110",
  21903=>"000000001",
  21904=>"100000100",
  21905=>"000000011",
  21906=>"111111111",
  21907=>"111000000",
  21908=>"000000000",
  21909=>"000010110",
  21910=>"111011000",
  21911=>"111011000",
  21912=>"000110111",
  21913=>"110000010",
  21914=>"101100111",
  21915=>"111111100",
  21916=>"111111111",
  21917=>"011000000",
  21918=>"100001111",
  21919=>"011011011",
  21920=>"010000100",
  21921=>"010010100",
  21922=>"000001111",
  21923=>"111111111",
  21924=>"111111100",
  21925=>"010110111",
  21926=>"111111111",
  21927=>"010010011",
  21928=>"000000000",
  21929=>"110000000",
  21930=>"110000000",
  21931=>"111110000",
  21932=>"100101111",
  21933=>"001000000",
  21934=>"000111111",
  21935=>"011000100",
  21936=>"000111111",
  21937=>"000000000",
  21938=>"000000111",
  21939=>"111111111",
  21940=>"001000000",
  21941=>"001001001",
  21942=>"011111100",
  21943=>"110010000",
  21944=>"000000000",
  21945=>"000000000",
  21946=>"000000000",
  21947=>"001101100",
  21948=>"111010000",
  21949=>"001001111",
  21950=>"000000000",
  21951=>"100111111",
  21952=>"000100000",
  21953=>"111101111",
  21954=>"111111111",
  21955=>"100010111",
  21956=>"111111110",
  21957=>"000000110",
  21958=>"001001111",
  21959=>"000000000",
  21960=>"111001111",
  21961=>"100100111",
  21962=>"001000000",
  21963=>"111101110",
  21964=>"000000000",
  21965=>"000000000",
  21966=>"111111010",
  21967=>"000100111",
  21968=>"000000000",
  21969=>"100000110",
  21970=>"111111111",
  21971=>"000000111",
  21972=>"111111101",
  21973=>"111011100",
  21974=>"000000000",
  21975=>"000111111",
  21976=>"111111011",
  21977=>"000000111",
  21978=>"000000000",
  21979=>"111111111",
  21980=>"001001011",
  21981=>"011010011",
  21982=>"000000100",
  21983=>"100100111",
  21984=>"000001111",
  21985=>"111111010",
  21986=>"000011000",
  21987=>"111111011",
  21988=>"110000000",
  21989=>"111011001",
  21990=>"111111111",
  21991=>"111111111",
  21992=>"001001011",
  21993=>"111111101",
  21994=>"100000111",
  21995=>"110011100",
  21996=>"001000000",
  21997=>"111011000",
  21998=>"000001001",
  21999=>"111111010",
  22000=>"000000111",
  22001=>"111001011",
  22002=>"111110111",
  22003=>"001000000",
  22004=>"111010110",
  22005=>"111000111",
  22006=>"000000100",
  22007=>"000001001",
  22008=>"111010000",
  22009=>"011011000",
  22010=>"111111111",
  22011=>"011111011",
  22012=>"000000000",
  22013=>"011000000",
  22014=>"100010010",
  22015=>"110111111",
  22016=>"111111100",
  22017=>"111000011",
  22018=>"010000111",
  22019=>"111111000",
  22020=>"001000000",
  22021=>"000000000",
  22022=>"010110111",
  22023=>"111111111",
  22024=>"111111111",
  22025=>"110000000",
  22026=>"111111000",
  22027=>"011000000",
  22028=>"000001011",
  22029=>"000110111",
  22030=>"111110110",
  22031=>"011010111",
  22032=>"111111111",
  22033=>"000000010",
  22034=>"000110110",
  22035=>"011111111",
  22036=>"111100111",
  22037=>"000000001",
  22038=>"000000100",
  22039=>"001001001",
  22040=>"111110000",
  22041=>"001000011",
  22042=>"000000000",
  22043=>"000000000",
  22044=>"111111111",
  22045=>"000000000",
  22046=>"001000011",
  22047=>"100001110",
  22048=>"000000000",
  22049=>"111111110",
  22050=>"111011111",
  22051=>"111000000",
  22052=>"111110110",
  22053=>"010110111",
  22054=>"011101111",
  22055=>"111001001",
  22056=>"111111111",
  22057=>"000000000",
  22058=>"000000111",
  22059=>"010000010",
  22060=>"001000000",
  22061=>"001011111",
  22062=>"011011110",
  22063=>"111111111",
  22064=>"111011000",
  22065=>"101100111",
  22066=>"011101000",
  22067=>"111111111",
  22068=>"000110110",
  22069=>"011010000",
  22070=>"111111111",
  22071=>"111011110",
  22072=>"000101111",
  22073=>"111111111",
  22074=>"000000000",
  22075=>"000000000",
  22076=>"111111000",
  22077=>"000000000",
  22078=>"010111011",
  22079=>"001000000",
  22080=>"111110110",
  22081=>"000100111",
  22082=>"100111111",
  22083=>"111000111",
  22084=>"010011001",
  22085=>"000010010",
  22086=>"111111000",
  22087=>"111111111",
  22088=>"000111111",
  22089=>"001101111",
  22090=>"000000000",
  22091=>"111110111",
  22092=>"111111110",
  22093=>"100000000",
  22094=>"011000000",
  22095=>"000000000",
  22096=>"000000000",
  22097=>"111111011",
  22098=>"110010110",
  22099=>"101111110",
  22100=>"000000000",
  22101=>"111111111",
  22102=>"111101111",
  22103=>"000000000",
  22104=>"001001001",
  22105=>"000000000",
  22106=>"000000100",
  22107=>"111111000",
  22108=>"110111111",
  22109=>"001101100",
  22110=>"000000000",
  22111=>"010110110",
  22112=>"000110110",
  22113=>"011000000",
  22114=>"000100100",
  22115=>"000000111",
  22116=>"111101111",
  22117=>"111110001",
  22118=>"000000000",
  22119=>"000000100",
  22120=>"000000111",
  22121=>"111000000",
  22122=>"111110100",
  22123=>"000100110",
  22124=>"101111111",
  22125=>"111111111",
  22126=>"000000000",
  22127=>"100110010",
  22128=>"000000000",
  22129=>"101101111",
  22130=>"000000000",
  22131=>"000001000",
  22132=>"111111111",
  22133=>"000000011",
  22134=>"111111000",
  22135=>"011011001",
  22136=>"000000011",
  22137=>"111111111",
  22138=>"110100110",
  22139=>"011000000",
  22140=>"110110100",
  22141=>"000111111",
  22142=>"110100000",
  22143=>"000000000",
  22144=>"000000000",
  22145=>"111010010",
  22146=>"100110000",
  22147=>"111110111",
  22148=>"111111111",
  22149=>"111111100",
  22150=>"111111111",
  22151=>"111111001",
  22152=>"111010011",
  22153=>"110110110",
  22154=>"001001011",
  22155=>"100001111",
  22156=>"111111111",
  22157=>"000000000",
  22158=>"111100000",
  22159=>"111111111",
  22160=>"111011111",
  22161=>"000000000",
  22162=>"000000110",
  22163=>"000010000",
  22164=>"001000110",
  22165=>"111111111",
  22166=>"000001011",
  22167=>"000000000",
  22168=>"111111011",
  22169=>"111111111",
  22170=>"111111111",
  22171=>"000000000",
  22172=>"000000000",
  22173=>"000011111",
  22174=>"011001111",
  22175=>"000000110",
  22176=>"000011110",
  22177=>"000000000",
  22178=>"111111101",
  22179=>"111010010",
  22180=>"101101100",
  22181=>"100100110",
  22182=>"111011000",
  22183=>"111111001",
  22184=>"111000000",
  22185=>"111000101",
  22186=>"000111111",
  22187=>"001001001",
  22188=>"111100010",
  22189=>"011011011",
  22190=>"111111011",
  22191=>"111011111",
  22192=>"111011011",
  22193=>"100000000",
  22194=>"110100111",
  22195=>"000000000",
  22196=>"111111110",
  22197=>"000000000",
  22198=>"000000111",
  22199=>"111111111",
  22200=>"000001001",
  22201=>"011111111",
  22202=>"100000000",
  22203=>"000000111",
  22204=>"001011000",
  22205=>"111111010",
  22206=>"111111111",
  22207=>"111111111",
  22208=>"111111110",
  22209=>"000000100",
  22210=>"000001111",
  22211=>"110000011",
  22212=>"111001000",
  22213=>"001011011",
  22214=>"111000000",
  22215=>"000001000",
  22216=>"011011111",
  22217=>"011111111",
  22218=>"000000000",
  22219=>"000110110",
  22220=>"000011111",
  22221=>"110111000",
  22222=>"000000110",
  22223=>"111111111",
  22224=>"110000101",
  22225=>"000000101",
  22226=>"110000011",
  22227=>"000000000",
  22228=>"111111010",
  22229=>"111110111",
  22230=>"011000000",
  22231=>"111111111",
  22232=>"001000100",
  22233=>"000000000",
  22234=>"111010000",
  22235=>"000000111",
  22236=>"011001111",
  22237=>"111111110",
  22238=>"110111110",
  22239=>"001001000",
  22240=>"111110100",
  22241=>"111111000",
  22242=>"111111010",
  22243=>"111111000",
  22244=>"110111111",
  22245=>"100000000",
  22246=>"000100111",
  22247=>"110000000",
  22248=>"001000000",
  22249=>"111111111",
  22250=>"001000001",
  22251=>"000000000",
  22252=>"111111111",
  22253=>"000000000",
  22254=>"111111111",
  22255=>"000000000",
  22256=>"000000111",
  22257=>"000000111",
  22258=>"000111111",
  22259=>"000000001",
  22260=>"000000000",
  22261=>"011011000",
  22262=>"001000110",
  22263=>"101000000",
  22264=>"101111111",
  22265=>"001000000",
  22266=>"111111111",
  22267=>"111100000",
  22268=>"110110110",
  22269=>"011001000",
  22270=>"111111110",
  22271=>"111111111",
  22272=>"000000000",
  22273=>"010111110",
  22274=>"111110000",
  22275=>"110000110",
  22276=>"000000000",
  22277=>"111000000",
  22278=>"000000000",
  22279=>"000000100",
  22280=>"000000100",
  22281=>"111111111",
  22282=>"111000000",
  22283=>"000000010",
  22284=>"011101111",
  22285=>"000000000",
  22286=>"000000000",
  22287=>"000110111",
  22288=>"000000001",
  22289=>"111110110",
  22290=>"000000000",
  22291=>"110000000",
  22292=>"000111111",
  22293=>"000000000",
  22294=>"011011000",
  22295=>"111111111",
  22296=>"111110000",
  22297=>"111000110",
  22298=>"000011111",
  22299=>"011000000",
  22300=>"111111111",
  22301=>"011011011",
  22302=>"000110111",
  22303=>"100000000",
  22304=>"111110100",
  22305=>"000111111",
  22306=>"001100110",
  22307=>"111101000",
  22308=>"000110010",
  22309=>"111111000",
  22310=>"111111011",
  22311=>"000100100",
  22312=>"111111111",
  22313=>"000000000",
  22314=>"000111101",
  22315=>"000100110",
  22316=>"000110000",
  22317=>"111000000",
  22318=>"000000111",
  22319=>"001001101",
  22320=>"001000000",
  22321=>"111111111",
  22322=>"011001111",
  22323=>"111111110",
  22324=>"000001101",
  22325=>"111110000",
  22326=>"111001111",
  22327=>"001111111",
  22328=>"001111011",
  22329=>"111111011",
  22330=>"000000111",
  22331=>"000110000",
  22332=>"111110110",
  22333=>"111001101",
  22334=>"000101111",
  22335=>"000001000",
  22336=>"001000111",
  22337=>"111000111",
  22338=>"001001111",
  22339=>"100100000",
  22340=>"110111111",
  22341=>"011000000",
  22342=>"000000000",
  22343=>"111111111",
  22344=>"000100111",
  22345=>"000000000",
  22346=>"000000001",
  22347=>"000101111",
  22348=>"010010010",
  22349=>"111111110",
  22350=>"001000000",
  22351=>"000000001",
  22352=>"011011000",
  22353=>"100100111",
  22354=>"000000111",
  22355=>"000000111",
  22356=>"011000000",
  22357=>"111011011",
  22358=>"111000000",
  22359=>"000000000",
  22360=>"111111000",
  22361=>"111111111",
  22362=>"000000001",
  22363=>"000000000",
  22364=>"001000001",
  22365=>"010000000",
  22366=>"000000000",
  22367=>"111111100",
  22368=>"110100111",
  22369=>"000000001",
  22370=>"011011100",
  22371=>"000000000",
  22372=>"110111111",
  22373=>"000000000",
  22374=>"000000000",
  22375=>"000000000",
  22376=>"001000000",
  22377=>"000000000",
  22378=>"111111111",
  22379=>"011011111",
  22380=>"111111000",
  22381=>"100111111",
  22382=>"110111111",
  22383=>"110000110",
  22384=>"000000011",
  22385=>"110111110",
  22386=>"000000000",
  22387=>"111000100",
  22388=>"110111000",
  22389=>"000100100",
  22390=>"111001011",
  22391=>"000100111",
  22392=>"000000000",
  22393=>"111000001",
  22394=>"011010011",
  22395=>"111011111",
  22396=>"111111111",
  22397=>"111111011",
  22398=>"111011011",
  22399=>"000000111",
  22400=>"000110000",
  22401=>"111011011",
  22402=>"100111111",
  22403=>"111011111",
  22404=>"111111011",
  22405=>"000000101",
  22406=>"111100100",
  22407=>"111011001",
  22408=>"111011000",
  22409=>"111111111",
  22410=>"111111111",
  22411=>"111110000",
  22412=>"000001011",
  22413=>"010100001",
  22414=>"011011001",
  22415=>"011011001",
  22416=>"000000100",
  22417=>"010000000",
  22418=>"011010101",
  22419=>"111111111",
  22420=>"000000111",
  22421=>"000100000",
  22422=>"111000001",
  22423=>"111000000",
  22424=>"000001001",
  22425=>"111111000",
  22426=>"110000000",
  22427=>"000000010",
  22428=>"111111110",
  22429=>"111111111",
  22430=>"011111111",
  22431=>"000111110",
  22432=>"110111111",
  22433=>"000001111",
  22434=>"111111111",
  22435=>"010000110",
  22436=>"111111010",
  22437=>"111110000",
  22438=>"000000001",
  22439=>"111111111",
  22440=>"100110111",
  22441=>"001000100",
  22442=>"001000011",
  22443=>"001001111",
  22444=>"111111110",
  22445=>"000000000",
  22446=>"001111110",
  22447=>"000001011",
  22448=>"000000000",
  22449=>"000111111",
  22450=>"001011111",
  22451=>"111110110",
  22452=>"001000011",
  22453=>"011000100",
  22454=>"001011111",
  22455=>"000000000",
  22456=>"110001111",
  22457=>"110110111",
  22458=>"110010111",
  22459=>"011111111",
  22460=>"111111111",
  22461=>"110000100",
  22462=>"111110000",
  22463=>"000010111",
  22464=>"000000000",
  22465=>"000110111",
  22466=>"111111111",
  22467=>"111111111",
  22468=>"001001001",
  22469=>"111111111",
  22470=>"011000100",
  22471=>"000000000",
  22472=>"110100000",
  22473=>"000000000",
  22474=>"111001100",
  22475=>"000000010",
  22476=>"100000110",
  22477=>"111111001",
  22478=>"110011011",
  22479=>"111111111",
  22480=>"000000011",
  22481=>"111100111",
  22482=>"000000001",
  22483=>"111111111",
  22484=>"111111111",
  22485=>"000100000",
  22486=>"000000000",
  22487=>"101111111",
  22488=>"111011111",
  22489=>"000001111",
  22490=>"000000111",
  22491=>"011111110",
  22492=>"011111111",
  22493=>"011011001",
  22494=>"111000000",
  22495=>"100110111",
  22496=>"000000000",
  22497=>"000000000",
  22498=>"110010000",
  22499=>"110110111",
  22500=>"001111111",
  22501=>"001111111",
  22502=>"001000000",
  22503=>"110111010",
  22504=>"011000000",
  22505=>"111011111",
  22506=>"101001001",
  22507=>"011000000",
  22508=>"000000001",
  22509=>"011100101",
  22510=>"001000000",
  22511=>"111000000",
  22512=>"110100111",
  22513=>"000000110",
  22514=>"111011000",
  22515=>"000110111",
  22516=>"111000000",
  22517=>"010100100",
  22518=>"111011011",
  22519=>"110110010",
  22520=>"000000000",
  22521=>"011001101",
  22522=>"000000001",
  22523=>"000111111",
  22524=>"011000111",
  22525=>"010011111",
  22526=>"011111111",
  22527=>"000000011",
  22528=>"000010111",
  22529=>"000000111",
  22530=>"100111111",
  22531=>"111000000",
  22532=>"000001011",
  22533=>"000001011",
  22534=>"111111111",
  22535=>"000000000",
  22536=>"000000111",
  22537=>"000011000",
  22538=>"000000000",
  22539=>"111111000",
  22540=>"110111111",
  22541=>"000001000",
  22542=>"000000000",
  22543=>"111111111",
  22544=>"101111000",
  22545=>"110111111",
  22546=>"111111000",
  22547=>"111111110",
  22548=>"111111111",
  22549=>"111111111",
  22550=>"000000111",
  22551=>"000000111",
  22552=>"111000111",
  22553=>"000000000",
  22554=>"110111111",
  22555=>"000110111",
  22556=>"111000000",
  22557=>"000111111",
  22558=>"011001001",
  22559=>"000000111",
  22560=>"110000110",
  22561=>"110111001",
  22562=>"111111011",
  22563=>"111011001",
  22564=>"001111110",
  22565=>"111111111",
  22566=>"111111110",
  22567=>"000110111",
  22568=>"000000000",
  22569=>"111110010",
  22570=>"111111000",
  22571=>"101000000",
  22572=>"111101111",
  22573=>"111111111",
  22574=>"000111000",
  22575=>"000000000",
  22576=>"000000000",
  22577=>"111010000",
  22578=>"100100000",
  22579=>"110111111",
  22580=>"110010000",
  22581=>"100011000",
  22582=>"101000000",
  22583=>"111111000",
  22584=>"000100110",
  22585=>"000101010",
  22586=>"111111111",
  22587=>"111110100",
  22588=>"001001000",
  22589=>"000111001",
  22590=>"000000000",
  22591=>"110000111",
  22592=>"111111111",
  22593=>"010110110",
  22594=>"111000000",
  22595=>"000000000",
  22596=>"111111111",
  22597=>"111001001",
  22598=>"111100000",
  22599=>"000000000",
  22600=>"100111111",
  22601=>"000000110",
  22602=>"000000100",
  22603=>"000111111",
  22604=>"000001000",
  22605=>"000111111",
  22606=>"011111111",
  22607=>"000111111",
  22608=>"111111111",
  22609=>"010111010",
  22610=>"000000000",
  22611=>"000100110",
  22612=>"000111111",
  22613=>"000000001",
  22614=>"000000100",
  22615=>"000111111",
  22616=>"001111111",
  22617=>"111000101",
  22618=>"001111111",
  22619=>"000000110",
  22620=>"000000001",
  22621=>"000000000",
  22622=>"111111100",
  22623=>"011010100",
  22624=>"000000000",
  22625=>"111110000",
  22626=>"000000010",
  22627=>"110000000",
  22628=>"000110000",
  22629=>"000111111",
  22630=>"000000100",
  22631=>"111001000",
  22632=>"111111000",
  22633=>"111111100",
  22634=>"111101001",
  22635=>"111111001",
  22636=>"000000000",
  22637=>"000000000",
  22638=>"011111000",
  22639=>"000000011",
  22640=>"000110111",
  22641=>"110111111",
  22642=>"011111000",
  22643=>"100101000",
  22644=>"011000000",
  22645=>"101001011",
  22646=>"111111000",
  22647=>"000000001",
  22648=>"100110111",
  22649=>"101101111",
  22650=>"011111111",
  22651=>"000100110",
  22652=>"000111110",
  22653=>"000000000",
  22654=>"000000010",
  22655=>"010000000",
  22656=>"000011111",
  22657=>"000000000",
  22658=>"000011111",
  22659=>"000010001",
  22660=>"110000000",
  22661=>"000001111",
  22662=>"111101111",
  22663=>"000000100",
  22664=>"111011001",
  22665=>"111110000",
  22666=>"000000000",
  22667=>"111111111",
  22668=>"000000000",
  22669=>"111111111",
  22670=>"111111000",
  22671=>"111111111",
  22672=>"000000000",
  22673=>"010000111",
  22674=>"111111111",
  22675=>"101111111",
  22676=>"000000111",
  22677=>"001100000",
  22678=>"111111111",
  22679=>"000000111",
  22680=>"100000111",
  22681=>"111111111",
  22682=>"000000000",
  22683=>"000000111",
  22684=>"111000000",
  22685=>"110011101",
  22686=>"000000001",
  22687=>"111000111",
  22688=>"001001111",
  22689=>"111000000",
  22690=>"001000000",
  22691=>"101000111",
  22692=>"100111111",
  22693=>"000111011",
  22694=>"111111111",
  22695=>"000011000",
  22696=>"000111111",
  22697=>"111111111",
  22698=>"000001111",
  22699=>"001000111",
  22700=>"000000000",
  22701=>"110111111",
  22702=>"000100000",
  22703=>"000000110",
  22704=>"000000000",
  22705=>"000000000",
  22706=>"111111111",
  22707=>"111111111",
  22708=>"100111110",
  22709=>"111000000",
  22710=>"000000000",
  22711=>"000000000",
  22712=>"000111111",
  22713=>"111110111",
  22714=>"111111111",
  22715=>"000001001",
  22716=>"111111111",
  22717=>"000001111",
  22718=>"111111000",
  22719=>"000001000",
  22720=>"111111111",
  22721=>"111001111",
  22722=>"000101000",
  22723=>"000111000",
  22724=>"000111111",
  22725=>"111111111",
  22726=>"111101001",
  22727=>"000000000",
  22728=>"111000110",
  22729=>"000001001",
  22730=>"110000001",
  22731=>"111000000",
  22732=>"111111111",
  22733=>"000000111",
  22734=>"010111111",
  22735=>"100100000",
  22736=>"000000000",
  22737=>"001011111",
  22738=>"000000000",
  22739=>"000000111",
  22740=>"100000110",
  22741=>"111111011",
  22742=>"111111111",
  22743=>"000000111",
  22744=>"000000000",
  22745=>"000001000",
  22746=>"000000111",
  22747=>"000000000",
  22748=>"000000100",
  22749=>"000100110",
  22750=>"000000000",
  22751=>"100100000",
  22752=>"000000000",
  22753=>"111111110",
  22754=>"000011111",
  22755=>"110111111",
  22756=>"001000000",
  22757=>"100000000",
  22758=>"000001011",
  22759=>"111111111",
  22760=>"111111111",
  22761=>"000000000",
  22762=>"000110100",
  22763=>"000000000",
  22764=>"010000000",
  22765=>"000000111",
  22766=>"111111011",
  22767=>"111111111",
  22768=>"111111111",
  22769=>"111100100",
  22770=>"001101111",
  22771=>"000000101",
  22772=>"111000000",
  22773=>"110110111",
  22774=>"001110000",
  22775=>"111001000",
  22776=>"111111010",
  22777=>"000000000",
  22778=>"000000000",
  22779=>"000000000",
  22780=>"100100111",
  22781=>"000000100",
  22782=>"111101000",
  22783=>"101101000",
  22784=>"111111000",
  22785=>"101101111",
  22786=>"000000000",
  22787=>"101100111",
  22788=>"001000000",
  22789=>"011001000",
  22790=>"000000111",
  22791=>"011111111",
  22792=>"000000111",
  22793=>"010110000",
  22794=>"111111000",
  22795=>"011111111",
  22796=>"111111111",
  22797=>"000000000",
  22798=>"000101111",
  22799=>"001000010",
  22800=>"101100111",
  22801=>"111000000",
  22802=>"000000000",
  22803=>"101000000",
  22804=>"101000000",
  22805=>"000000111",
  22806=>"110110111",
  22807=>"111111000",
  22808=>"111111000",
  22809=>"000000111",
  22810=>"110111000",
  22811=>"111001001",
  22812=>"011011011",
  22813=>"111111111",
  22814=>"111111011",
  22815=>"000000111",
  22816=>"000011000",
  22817=>"111111011",
  22818=>"111111000",
  22819=>"000000101",
  22820=>"000000111",
  22821=>"111001000",
  22822=>"110001111",
  22823=>"010111011",
  22824=>"100101000",
  22825=>"000111110",
  22826=>"111111110",
  22827=>"000000011",
  22828=>"111111111",
  22829=>"000000000",
  22830=>"111000111",
  22831=>"100000101",
  22832=>"111111000",
  22833=>"000000000",
  22834=>"000001000",
  22835=>"000000000",
  22836=>"110001011",
  22837=>"001000000",
  22838=>"000100100",
  22839=>"110000111",
  22840=>"000100111",
  22841=>"111101100",
  22842=>"100111111",
  22843=>"111001000",
  22844=>"111111100",
  22845=>"000100100",
  22846=>"111111111",
  22847=>"111000000",
  22848=>"001000000",
  22849=>"000000000",
  22850=>"010111100",
  22851=>"001111000",
  22852=>"000000100",
  22853=>"000000001",
  22854=>"000000000",
  22855=>"111100110",
  22856=>"000000000",
  22857=>"000000011",
  22858=>"000000111",
  22859=>"000100110",
  22860=>"111000000",
  22861=>"111111000",
  22862=>"000001101",
  22863=>"110110110",
  22864=>"100100101",
  22865=>"111111011",
  22866=>"010100111",
  22867=>"000000000",
  22868=>"111111111",
  22869=>"011011011",
  22870=>"100111111",
  22871=>"111111010",
  22872=>"000000000",
  22873=>"111111111",
  22874=>"000000111",
  22875=>"111111111",
  22876=>"110000111",
  22877=>"000000000",
  22878=>"111010000",
  22879=>"111001000",
  22880=>"001000000",
  22881=>"000000000",
  22882=>"110000000",
  22883=>"100000111",
  22884=>"000000000",
  22885=>"000000000",
  22886=>"111000001",
  22887=>"000000000",
  22888=>"001001000",
  22889=>"000111111",
  22890=>"111111000",
  22891=>"000000000",
  22892=>"110111110",
  22893=>"111110110",
  22894=>"111001111",
  22895=>"100111111",
  22896=>"100000111",
  22897=>"000011001",
  22898=>"110100111",
  22899=>"100100110",
  22900=>"000111011",
  22901=>"000000000",
  22902=>"000101100",
  22903=>"000010111",
  22904=>"000111111",
  22905=>"000000011",
  22906=>"100000000",
  22907=>"000100111",
  22908=>"001001001",
  22909=>"001000000",
  22910=>"000000000",
  22911=>"111101111",
  22912=>"100011111",
  22913=>"111111111",
  22914=>"111100000",
  22915=>"110111111",
  22916=>"111000011",
  22917=>"110111111",
  22918=>"100000100",
  22919=>"111111000",
  22920=>"111111000",
  22921=>"000000000",
  22922=>"000000001",
  22923=>"111111111",
  22924=>"101000000",
  22925=>"000000000",
  22926=>"111111111",
  22927=>"111111000",
  22928=>"000000111",
  22929=>"000000000",
  22930=>"111111111",
  22931=>"000000000",
  22932=>"001000000",
  22933=>"000111000",
  22934=>"011111011",
  22935=>"000001001",
  22936=>"111000000",
  22937=>"111000101",
  22938=>"111111111",
  22939=>"100100000",
  22940=>"100000000",
  22941=>"111110111",
  22942=>"111000000",
  22943=>"000000000",
  22944=>"111111111",
  22945=>"000110100",
  22946=>"000110111",
  22947=>"001001001",
  22948=>"100000111",
  22949=>"111111111",
  22950=>"000000010",
  22951=>"000011000",
  22952=>"111110111",
  22953=>"000001001",
  22954=>"110011001",
  22955=>"111000000",
  22956=>"000000000",
  22957=>"000000000",
  22958=>"111101010",
  22959=>"000000000",
  22960=>"000000111",
  22961=>"111111110",
  22962=>"000000100",
  22963=>"111000000",
  22964=>"000000000",
  22965=>"000000111",
  22966=>"000000111",
  22967=>"100000110",
  22968=>"100111111",
  22969=>"011111111",
  22970=>"001111111",
  22971=>"000111000",
  22972=>"111011111",
  22973=>"110011111",
  22974=>"111000110",
  22975=>"110111111",
  22976=>"010110111",
  22977=>"000000000",
  22978=>"000010000",
  22979=>"010110111",
  22980=>"000111100",
  22981=>"100000111",
  22982=>"000000000",
  22983=>"000100000",
  22984=>"111100110",
  22985=>"111111000",
  22986=>"000000101",
  22987=>"000000110",
  22988=>"111100000",
  22989=>"000000000",
  22990=>"111111000",
  22991=>"111000000",
  22992=>"011011000",
  22993=>"101100100",
  22994=>"111111001",
  22995=>"000000000",
  22996=>"000000000",
  22997=>"111111001",
  22998=>"100111000",
  22999=>"110110100",
  23000=>"101000000",
  23001=>"011011011",
  23002=>"111111000",
  23003=>"000000000",
  23004=>"110000000",
  23005=>"000000100",
  23006=>"000000011",
  23007=>"101111000",
  23008=>"111000000",
  23009=>"001000000",
  23010=>"111000000",
  23011=>"111111001",
  23012=>"000000011",
  23013=>"000001111",
  23014=>"001111000",
  23015=>"010110000",
  23016=>"000000111",
  23017=>"000000011",
  23018=>"000000100",
  23019=>"111111100",
  23020=>"000000111",
  23021=>"011001111",
  23022=>"000111001",
  23023=>"111111100",
  23024=>"000001100",
  23025=>"111001100",
  23026=>"000010111",
  23027=>"110111111",
  23028=>"111111111",
  23029=>"101000100",
  23030=>"000000000",
  23031=>"000000000",
  23032=>"100100111",
  23033=>"111101111",
  23034=>"110111000",
  23035=>"000000000",
  23036=>"111111111",
  23037=>"111111111",
  23038=>"111111111",
  23039=>"001111111",
  23040=>"100001011",
  23041=>"001000000",
  23042=>"100101001",
  23043=>"100100101",
  23044=>"011001111",
  23045=>"000111000",
  23046=>"101000011",
  23047=>"111100000",
  23048=>"011011000",
  23049=>"110000000",
  23050=>"000000111",
  23051=>"111111111",
  23052=>"000000110",
  23053=>"100001001",
  23054=>"100111111",
  23055=>"111101001",
  23056=>"111111010",
  23057=>"000111111",
  23058=>"101101101",
  23059=>"110111111",
  23060=>"101111111",
  23061=>"111111000",
  23062=>"000000001",
  23063=>"000011111",
  23064=>"000010110",
  23065=>"100000001",
  23066=>"111111111",
  23067=>"100110100",
  23068=>"110100001",
  23069=>"000000001",
  23070=>"001001001",
  23071=>"111111111",
  23072=>"001001000",
  23073=>"001111111",
  23074=>"111111111",
  23075=>"111001011",
  23076=>"111111111",
  23077=>"111111111",
  23078=>"000100100",
  23079=>"100100111",
  23080=>"111000111",
  23081=>"001000000",
  23082=>"000101111",
  23083=>"111100000",
  23084=>"110111111",
  23085=>"100110101",
  23086=>"111001111",
  23087=>"110000000",
  23088=>"000000000",
  23089=>"101001001",
  23090=>"000000000",
  23091=>"100100100",
  23092=>"000011000",
  23093=>"111111001",
  23094=>"000000101",
  23095=>"000000000",
  23096=>"001001001",
  23097=>"111111111",
  23098=>"000000000",
  23099=>"110111110",
  23100=>"111111111",
  23101=>"000000000",
  23102=>"011011000",
  23103=>"100000101",
  23104=>"011111100",
  23105=>"111010000",
  23106=>"100000100",
  23107=>"111010010",
  23108=>"001001011",
  23109=>"111111000",
  23110=>"000000000",
  23111=>"000000111",
  23112=>"111111011",
  23113=>"000000111",
  23114=>"111111111",
  23115=>"111111100",
  23116=>"000000111",
  23117=>"111000111",
  23118=>"000000000",
  23119=>"111111111",
  23120=>"111001000",
  23121=>"111111110",
  23122=>"111111111",
  23123=>"000000000",
  23124=>"101000001",
  23125=>"000111011",
  23126=>"000000001",
  23127=>"111001000",
  23128=>"011011000",
  23129=>"001000000",
  23130=>"111101111",
  23131=>"000000000",
  23132=>"111001101",
  23133=>"010110110",
  23134=>"111000000",
  23135=>"111011011",
  23136=>"001000000",
  23137=>"111111001",
  23138=>"111111000",
  23139=>"011111111",
  23140=>"011010111",
  23141=>"000000111",
  23142=>"111000000",
  23143=>"100100110",
  23144=>"110111111",
  23145=>"000000000",
  23146=>"111111000",
  23147=>"000000000",
  23148=>"000000000",
  23149=>"100000000",
  23150=>"110111111",
  23151=>"111111111",
  23152=>"000000111",
  23153=>"001110100",
  23154=>"111111111",
  23155=>"111111111",
  23156=>"000000000",
  23157=>"000110111",
  23158=>"011111000",
  23159=>"000000000",
  23160=>"101111000",
  23161=>"111111111",
  23162=>"001000000",
  23163=>"100000111",
  23164=>"000111110",
  23165=>"000000000",
  23166=>"111000000",
  23167=>"010000110",
  23168=>"111110000",
  23169=>"111101000",
  23170=>"111111111",
  23171=>"000100100",
  23172=>"000000000",
  23173=>"111000001",
  23174=>"000000000",
  23175=>"111111000",
  23176=>"110000000",
  23177=>"011111101",
  23178=>"111010000",
  23179=>"111111011",
  23180=>"111001000",
  23181=>"111111000",
  23182=>"101111111",
  23183=>"000111001",
  23184=>"011011000",
  23185=>"111001000",
  23186=>"111110010",
  23187=>"011101101",
  23188=>"000000000",
  23189=>"000000110",
  23190=>"100111111",
  23191=>"111111100",
  23192=>"100000000",
  23193=>"111000111",
  23194=>"111000000",
  23195=>"111111000",
  23196=>"000011000",
  23197=>"000110111",
  23198=>"111111111",
  23199=>"111111111",
  23200=>"111110111",
  23201=>"000000000",
  23202=>"100110111",
  23203=>"000000000",
  23204=>"111000001",
  23205=>"000000011",
  23206=>"111010010",
  23207=>"011100000",
  23208=>"000000010",
  23209=>"001101000",
  23210=>"100000001",
  23211=>"000000000",
  23212=>"111111111",
  23213=>"000000000",
  23214=>"001000000",
  23215=>"001101111",
  23216=>"000000011",
  23217=>"110110110",
  23218=>"111011111",
  23219=>"001001000",
  23220=>"000000000",
  23221=>"000000110",
  23222=>"111111111",
  23223=>"111111000",
  23224=>"111111111",
  23225=>"111111111",
  23226=>"111000000",
  23227=>"000000000",
  23228=>"110111111",
  23229=>"000000110",
  23230=>"110000111",
  23231=>"000111111",
  23232=>"000000111",
  23233=>"001001100",
  23234=>"000111111",
  23235=>"000010000",
  23236=>"111111111",
  23237=>"000000111",
  23238=>"000111011",
  23239=>"000000111",
  23240=>"000000110",
  23241=>"111111111",
  23242=>"111111111",
  23243=>"110110110",
  23244=>"110111111",
  23245=>"000001001",
  23246=>"000000000",
  23247=>"000000000",
  23248=>"101111010",
  23249=>"011011111",
  23250=>"100111111",
  23251=>"111111111",
  23252=>"101000001",
  23253=>"111111111",
  23254=>"010010000",
  23255=>"000000000",
  23256=>"000000111",
  23257=>"000011000",
  23258=>"000000000",
  23259=>"000000000",
  23260=>"000000000",
  23261=>"110111111",
  23262=>"000000000",
  23263=>"000000000",
  23264=>"111000000",
  23265=>"000000011",
  23266=>"000000011",
  23267=>"111111001",
  23268=>"111011001",
  23269=>"000000000",
  23270=>"111000000",
  23271=>"000011001",
  23272=>"111101101",
  23273=>"111001000",
  23274=>"000110111",
  23275=>"000000000",
  23276=>"000111111",
  23277=>"001000000",
  23278=>"000001111",
  23279=>"111111000",
  23280=>"000001000",
  23281=>"100111110",
  23282=>"110110110",
  23283=>"000000110",
  23284=>"000000000",
  23285=>"111111000",
  23286=>"000011011",
  23287=>"110000010",
  23288=>"110111111",
  23289=>"000000000",
  23290=>"000011111",
  23291=>"010111000",
  23292=>"000100100",
  23293=>"011000000",
  23294=>"000000001",
  23295=>"000000000",
  23296=>"111111111",
  23297=>"001001000",
  23298=>"111111111",
  23299=>"111111111",
  23300=>"000000001",
  23301=>"001000000",
  23302=>"000000000",
  23303=>"011000000",
  23304=>"000000110",
  23305=>"111101111",
  23306=>"111000000",
  23307=>"100000011",
  23308=>"000000000",
  23309=>"000000000",
  23310=>"000000000",
  23311=>"111001001",
  23312=>"000000000",
  23313=>"100001111",
  23314=>"111000000",
  23315=>"010010010",
  23316=>"111111011",
  23317=>"000011000",
  23318=>"001001101",
  23319=>"000000010",
  23320=>"111111100",
  23321=>"111111001",
  23322=>"101101000",
  23323=>"000000011",
  23324=>"011010010",
  23325=>"111111000",
  23326=>"000000000",
  23327=>"111000011",
  23328=>"000110010",
  23329=>"011111111",
  23330=>"111111111",
  23331=>"000000111",
  23332=>"001001000",
  23333=>"111111111",
  23334=>"100100000",
  23335=>"000000100",
  23336=>"111111111",
  23337=>"000000000",
  23338=>"000000000",
  23339=>"111111111",
  23340=>"111110111",
  23341=>"110110111",
  23342=>"000000000",
  23343=>"001000000",
  23344=>"001110111",
  23345=>"000000000",
  23346=>"110111101",
  23347=>"000001000",
  23348=>"000101101",
  23349=>"111100000",
  23350=>"111000000",
  23351=>"111001000",
  23352=>"010111111",
  23353=>"000100000",
  23354=>"000000010",
  23355=>"000000111",
  23356=>"000000000",
  23357=>"000000100",
  23358=>"111111111",
  23359=>"100100101",
  23360=>"001000000",
  23361=>"111010111",
  23362=>"110110110",
  23363=>"111110111",
  23364=>"000000100",
  23365=>"110010111",
  23366=>"000000001",
  23367=>"000110111",
  23368=>"000000000",
  23369=>"110100000",
  23370=>"111101000",
  23371=>"011111111",
  23372=>"001000111",
  23373=>"000010110",
  23374=>"111111111",
  23375=>"111111110",
  23376=>"000000001",
  23377=>"111000111",
  23378=>"111000000",
  23379=>"111011001",
  23380=>"011000000",
  23381=>"001001011",
  23382=>"101001101",
  23383=>"111111000",
  23384=>"000000000",
  23385=>"111011000",
  23386=>"111111111",
  23387=>"111101100",
  23388=>"111000000",
  23389=>"000111111",
  23390=>"111000000",
  23391=>"000000000",
  23392=>"000100000",
  23393=>"111111111",
  23394=>"000000000",
  23395=>"111010000",
  23396=>"110110000",
  23397=>"000001111",
  23398=>"110111111",
  23399=>"000000000",
  23400=>"110111110",
  23401=>"110111111",
  23402=>"000000101",
  23403=>"111111111",
  23404=>"000000000",
  23405=>"000000000",
  23406=>"000000100",
  23407=>"111110111",
  23408=>"000011111",
  23409=>"000001011",
  23410=>"100111111",
  23411=>"111111100",
  23412=>"000000000",
  23413=>"000111111",
  23414=>"000000001",
  23415=>"000000010",
  23416=>"000000111",
  23417=>"110111001",
  23418=>"110111111",
  23419=>"100100110",
  23420=>"111111111",
  23421=>"111100000",
  23422=>"000000111",
  23423=>"111101100",
  23424=>"100110110",
  23425=>"000000000",
  23426=>"011011001",
  23427=>"111100100",
  23428=>"000100100",
  23429=>"110010110",
  23430=>"111111001",
  23431=>"001000000",
  23432=>"001000001",
  23433=>"000111000",
  23434=>"100100100",
  23435=>"000000011",
  23436=>"000101111",
  23437=>"001111111",
  23438=>"011011111",
  23439=>"111111111",
  23440=>"000000000",
  23441=>"000000000",
  23442=>"000000000",
  23443=>"100000000",
  23444=>"001101011",
  23445=>"000010110",
  23446=>"111111111",
  23447=>"000000000",
  23448=>"000000111",
  23449=>"000011111",
  23450=>"100111000",
  23451=>"000000000",
  23452=>"100000111",
  23453=>"111111000",
  23454=>"101001001",
  23455=>"000000000",
  23456=>"001001111",
  23457=>"101000000",
  23458=>"001001000",
  23459=>"111001001",
  23460=>"100101011",
  23461=>"000000100",
  23462=>"100000000",
  23463=>"000000000",
  23464=>"111111100",
  23465=>"000000000",
  23466=>"010011111",
  23467=>"001001111",
  23468=>"000000000",
  23469=>"101011001",
  23470=>"111111111",
  23471=>"111111111",
  23472=>"000000111",
  23473=>"010110000",
  23474=>"111111111",
  23475=>"000110111",
  23476=>"111000000",
  23477=>"000111011",
  23478=>"111111111",
  23479=>"101100000",
  23480=>"111111110",
  23481=>"110010000",
  23482=>"000001111",
  23483=>"100000000",
  23484=>"110000000",
  23485=>"100000111",
  23486=>"001001100",
  23487=>"000000100",
  23488=>"000110000",
  23489=>"111111111",
  23490=>"111111111",
  23491=>"000000000",
  23492=>"111101100",
  23493=>"111011011",
  23494=>"000000000",
  23495=>"011010000",
  23496=>"110000000",
  23497=>"110111111",
  23498=>"000000000",
  23499=>"000011011",
  23500=>"111110111",
  23501=>"001000000",
  23502=>"100001000",
  23503=>"110000001",
  23504=>"111011000",
  23505=>"000000000",
  23506=>"110000000",
  23507=>"111111111",
  23508=>"111110011",
  23509=>"111101101",
  23510=>"000000111",
  23511=>"000000000",
  23512=>"101001111",
  23513=>"111111111",
  23514=>"001000000",
  23515=>"111111111",
  23516=>"111111111",
  23517=>"011000000",
  23518=>"111111011",
  23519=>"000000000",
  23520=>"000000000",
  23521=>"000000000",
  23522=>"111111100",
  23523=>"101100100",
  23524=>"111111001",
  23525=>"111111111",
  23526=>"000000001",
  23527=>"111101000",
  23528=>"100000000",
  23529=>"010111010",
  23530=>"111001001",
  23531=>"000000000",
  23532=>"111111111",
  23533=>"111000000",
  23534=>"000000110",
  23535=>"100111111",
  23536=>"111101000",
  23537=>"000001000",
  23538=>"100111111",
  23539=>"000111111",
  23540=>"000000000",
  23541=>"111111100",
  23542=>"000000000",
  23543=>"001100100",
  23544=>"011010000",
  23545=>"100000000",
  23546=>"000011111",
  23547=>"110110111",
  23548=>"111111001",
  23549=>"011001000",
  23550=>"000000000",
  23551=>"111111111",
  23552=>"110110000",
  23553=>"011000001",
  23554=>"101111110",
  23555=>"000000011",
  23556=>"001011001",
  23557=>"010011011",
  23558=>"000000000",
  23559=>"000000000",
  23560=>"100111111",
  23561=>"111110100",
  23562=>"110000000",
  23563=>"000000001",
  23564=>"111111100",
  23565=>"111111111",
  23566=>"100100100",
  23567=>"111111111",
  23568=>"000000000",
  23569=>"110110110",
  23570=>"000000100",
  23571=>"000000000",
  23572=>"111000111",
  23573=>"011111110",
  23574=>"111111111",
  23575=>"011011111",
  23576=>"110000111",
  23577=>"100110111",
  23578=>"011011111",
  23579=>"111011001",
  23580=>"000001111",
  23581=>"110001001",
  23582=>"100110100",
  23583=>"110110110",
  23584=>"000111111",
  23585=>"000000000",
  23586=>"101100001",
  23587=>"111111111",
  23588=>"000000000",
  23589=>"011010000",
  23590=>"011111000",
  23591=>"110110110",
  23592=>"110000000",
  23593=>"000000000",
  23594=>"000010111",
  23595=>"000000100",
  23596=>"111111111",
  23597=>"000000000",
  23598=>"000000000",
  23599=>"000011011",
  23600=>"000000000",
  23601=>"001000000",
  23602=>"111111111",
  23603=>"000000000",
  23604=>"111111111",
  23605=>"111111011",
  23606=>"111001111",
  23607=>"001000100",
  23608=>"100110100",
  23609=>"000111001",
  23610=>"000000000",
  23611=>"110000000",
  23612=>"100110111",
  23613=>"111000111",
  23614=>"110111111",
  23615=>"001000001",
  23616=>"010011111",
  23617=>"001111111",
  23618=>"110000000",
  23619=>"000000000",
  23620=>"010000010",
  23621=>"000100100",
  23622=>"111000000",
  23623=>"011001000",
  23624=>"000110110",
  23625=>"111100111",
  23626=>"000000000",
  23627=>"100100100",
  23628=>"100111111",
  23629=>"000000111",
  23630=>"000010110",
  23631=>"111111111",
  23632=>"111101000",
  23633=>"110111111",
  23634=>"010000101",
  23635=>"000000100",
  23636=>"000010011",
  23637=>"011111111",
  23638=>"000000011",
  23639=>"000001001",
  23640=>"010000000",
  23641=>"111111111",
  23642=>"111000110",
  23643=>"111111111",
  23644=>"111111111",
  23645=>"111111111",
  23646=>"000000100",
  23647=>"111111111",
  23648=>"100110110",
  23649=>"111101111",
  23650=>"000101111",
  23651=>"000000001",
  23652=>"000000111",
  23653=>"000110111",
  23654=>"000110110",
  23655=>"111111101",
  23656=>"011111111",
  23657=>"001000100",
  23658=>"000000000",
  23659=>"111111111",
  23660=>"000100000",
  23661=>"000000000",
  23662=>"011011001",
  23663=>"111111011",
  23664=>"000000000",
  23665=>"000000000",
  23666=>"001001001",
  23667=>"110010111",
  23668=>"111111111",
  23669=>"001110100",
  23670=>"001001111",
  23671=>"011111000",
  23672=>"000000000",
  23673=>"011000000",
  23674=>"000000000",
  23675=>"000000000",
  23676=>"110110100",
  23677=>"000000000",
  23678=>"000000000",
  23679=>"000000000",
  23680=>"111111111",
  23681=>"010110000",
  23682=>"111111111",
  23683=>"000000000",
  23684=>"000001000",
  23685=>"001000000",
  23686=>"111100100",
  23687=>"000000001",
  23688=>"100000000",
  23689=>"111111111",
  23690=>"110000000",
  23691=>"111111101",
  23692=>"110111111",
  23693=>"111111111",
  23694=>"110111111",
  23695=>"111111011",
  23696=>"111111111",
  23697=>"111011000",
  23698=>"000000101",
  23699=>"110111000",
  23700=>"000000000",
  23701=>"111111111",
  23702=>"111111000",
  23703=>"111110000",
  23704=>"111001000",
  23705=>"100110111",
  23706=>"110110111",
  23707=>"000000000",
  23708=>"000000000",
  23709=>"000011111",
  23710=>"000001111",
  23711=>"000000000",
  23712=>"000000000",
  23713=>"111000000",
  23714=>"110000000",
  23715=>"111001001",
  23716=>"000001011",
  23717=>"000000111",
  23718=>"011001011",
  23719=>"111111101",
  23720=>"111111111",
  23721=>"000001100",
  23722=>"011111000",
  23723=>"111001111",
  23724=>"000011011",
  23725=>"001101100",
  23726=>"000001101",
  23727=>"011011111",
  23728=>"011011111",
  23729=>"000000100",
  23730=>"111111011",
  23731=>"000000001",
  23732=>"010100110",
  23733=>"000000000",
  23734=>"000000001",
  23735=>"000000000",
  23736=>"110000000",
  23737=>"000000000",
  23738=>"000000001",
  23739=>"111111110",
  23740=>"000000000",
  23741=>"100100000",
  23742=>"111111110",
  23743=>"111111111",
  23744=>"111111111",
  23745=>"111111111",
  23746=>"010000100",
  23747=>"000000000",
  23748=>"001111111",
  23749=>"000001001",
  23750=>"000000100",
  23751=>"000110110",
  23752=>"000011011",
  23753=>"111001111",
  23754=>"111011111",
  23755=>"000000000",
  23756=>"101101011",
  23757=>"011110011",
  23758=>"111100000",
  23759=>"000000000",
  23760=>"000000000",
  23761=>"000000001",
  23762=>"100100000",
  23763=>"000000100",
  23764=>"110000000",
  23765=>"110001101",
  23766=>"000000000",
  23767=>"111110000",
  23768=>"111111111",
  23769=>"000000111",
  23770=>"000010000",
  23771=>"000000100",
  23772=>"001000000",
  23773=>"111010111",
  23774=>"111111111",
  23775=>"000111111",
  23776=>"001011011",
  23777=>"001100111",
  23778=>"000011111",
  23779=>"001000000",
  23780=>"011001000",
  23781=>"111011011",
  23782=>"000111111",
  23783=>"110111001",
  23784=>"000000110",
  23785=>"000001000",
  23786=>"000000000",
  23787=>"000000000",
  23788=>"111111111",
  23789=>"111110111",
  23790=>"000111111",
  23791=>"001000000",
  23792=>"111111100",
  23793=>"111111111",
  23794=>"001000000",
  23795=>"000000101",
  23796=>"011110000",
  23797=>"111111111",
  23798=>"111011011",
  23799=>"111111011",
  23800=>"000000111",
  23801=>"111111011",
  23802=>"000000000",
  23803=>"100000000",
  23804=>"111011111",
  23805=>"100000001",
  23806=>"000000000",
  23807=>"000000110",
  23808=>"111111001",
  23809=>"111111111",
  23810=>"000000000",
  23811=>"111111111",
  23812=>"000000000",
  23813=>"000000101",
  23814=>"000000000",
  23815=>"111111111",
  23816=>"000000000",
  23817=>"111011011",
  23818=>"111111111",
  23819=>"100000111",
  23820=>"000000000",
  23821=>"000000000",
  23822=>"000100110",
  23823=>"110110110",
  23824=>"100000000",
  23825=>"111001100",
  23826=>"111110111",
  23827=>"100000001",
  23828=>"111111000",
  23829=>"111111111",
  23830=>"111111111",
  23831=>"111111110",
  23832=>"110010000",
  23833=>"111111011",
  23834=>"101001000",
  23835=>"000000000",
  23836=>"111111111",
  23837=>"000000000",
  23838=>"111111111",
  23839=>"111111111",
  23840=>"011001000",
  23841=>"111011000",
  23842=>"000100111",
  23843=>"111111111",
  23844=>"101111111",
  23845=>"000001001",
  23846=>"111111111",
  23847=>"000010000",
  23848=>"000000000",
  23849=>"011111111",
  23850=>"011011111",
  23851=>"111111111",
  23852=>"111111111",
  23853=>"110110110",
  23854=>"000000000",
  23855=>"000000000",
  23856=>"110111100",
  23857=>"111110111",
  23858=>"111110001",
  23859=>"000000000",
  23860=>"110000100",
  23861=>"000000000",
  23862=>"100001000",
  23863=>"111111111",
  23864=>"000000000",
  23865=>"000000000",
  23866=>"000000100",
  23867=>"111111111",
  23868=>"110110111",
  23869=>"011000000",
  23870=>"100111111",
  23871=>"100100000",
  23872=>"000010111",
  23873=>"000000000",
  23874=>"011001101",
  23875=>"111111010",
  23876=>"001001000",
  23877=>"111111111",
  23878=>"000000000",
  23879=>"001000000",
  23880=>"111111111",
  23881=>"100110000",
  23882=>"000000001",
  23883=>"011111111",
  23884=>"111000000",
  23885=>"100111111",
  23886=>"111111101",
  23887=>"110111111",
  23888=>"011011001",
  23889=>"000000000",
  23890=>"000000000",
  23891=>"111111111",
  23892=>"100100111",
  23893=>"011111000",
  23894=>"111111001",
  23895=>"111111111",
  23896=>"000000000",
  23897=>"111111111",
  23898=>"000000000",
  23899=>"011000000",
  23900=>"111111111",
  23901=>"111111111",
  23902=>"000000000",
  23903=>"100111011",
  23904=>"000000001",
  23905=>"100000000",
  23906=>"000001000",
  23907=>"111001011",
  23908=>"110111111",
  23909=>"000000000",
  23910=>"001000000",
  23911=>"111111111",
  23912=>"001111111",
  23913=>"111000011",
  23914=>"110110110",
  23915=>"111011001",
  23916=>"111111110",
  23917=>"010111111",
  23918=>"111111111",
  23919=>"100000000",
  23920=>"000000000",
  23921=>"000000000",
  23922=>"010011000",
  23923=>"100100000",
  23924=>"011000000",
  23925=>"000000001",
  23926=>"000000110",
  23927=>"111101111",
  23928=>"111100111",
  23929=>"110111111",
  23930=>"111111111",
  23931=>"000000000",
  23932=>"001000000",
  23933=>"111111111",
  23934=>"000000000",
  23935=>"000000000",
  23936=>"000100111",
  23937=>"111111000",
  23938=>"000000000",
  23939=>"111000000",
  23940=>"111111111",
  23941=>"111111111",
  23942=>"111101100",
  23943=>"111011011",
  23944=>"000000110",
  23945=>"000010111",
  23946=>"111000000",
  23947=>"000000000",
  23948=>"111111111",
  23949=>"101101111",
  23950=>"110111111",
  23951=>"110111111",
  23952=>"111110000",
  23953=>"000110111",
  23954=>"000000000",
  23955=>"111111111",
  23956=>"000000000",
  23957=>"000100000",
  23958=>"001111111",
  23959=>"111111110",
  23960=>"000000000",
  23961=>"111001000",
  23962=>"100100111",
  23963=>"111111111",
  23964=>"000000000",
  23965=>"000111111",
  23966=>"000000000",
  23967=>"000000110",
  23968=>"100100000",
  23969=>"001001100",
  23970=>"001001001",
  23971=>"000100110",
  23972=>"111111111",
  23973=>"000000000",
  23974=>"000010110",
  23975=>"111111111",
  23976=>"000000001",
  23977=>"011001001",
  23978=>"111110110",
  23979=>"000000100",
  23980=>"000000000",
  23981=>"111001001",
  23982=>"111111111",
  23983=>"111111111",
  23984=>"111111111",
  23985=>"000100111",
  23986=>"111111101",
  23987=>"111000111",
  23988=>"001000001",
  23989=>"000000000",
  23990=>"110110111",
  23991=>"000000000",
  23992=>"111111110",
  23993=>"111000000",
  23994=>"111010010",
  23995=>"000000000",
  23996=>"111111111",
  23997=>"111111111",
  23998=>"000000000",
  23999=>"111111111",
  24000=>"111111111",
  24001=>"100001111",
  24002=>"000000000",
  24003=>"000100111",
  24004=>"111111111",
  24005=>"000101111",
  24006=>"110110000",
  24007=>"000000000",
  24008=>"111001101",
  24009=>"111111111",
  24010=>"000000100",
  24011=>"111111111",
  24012=>"111110000",
  24013=>"010111011",
  24014=>"111011001",
  24015=>"111111111",
  24016=>"110110000",
  24017=>"111110111",
  24018=>"111111011",
  24019=>"001111000",
  24020=>"001001001",
  24021=>"111111111",
  24022=>"111111111",
  24023=>"000000001",
  24024=>"111111111",
  24025=>"000011001",
  24026=>"110000001",
  24027=>"111111101",
  24028=>"000000000",
  24029=>"110111111",
  24030=>"100111011",
  24031=>"111111111",
  24032=>"111111111",
  24033=>"011000000",
  24034=>"110101111",
  24035=>"110111111",
  24036=>"000011011",
  24037=>"100000000",
  24038=>"000000000",
  24039=>"111111100",
  24040=>"110011001",
  24041=>"000000000",
  24042=>"011001001",
  24043=>"000001000",
  24044=>"001000000",
  24045=>"000000100",
  24046=>"000000000",
  24047=>"000111011",
  24048=>"000000000",
  24049=>"000000101",
  24050=>"011000000",
  24051=>"000011011",
  24052=>"000001000",
  24053=>"111111111",
  24054=>"000000000",
  24055=>"100110110",
  24056=>"111011111",
  24057=>"110111010",
  24058=>"000000111",
  24059=>"000000000",
  24060=>"111111111",
  24061=>"010001011",
  24062=>"111111000",
  24063=>"111000000",
  24064=>"000000000",
  24065=>"011011111",
  24066=>"101000111",
  24067=>"001011000",
  24068=>"011011001",
  24069=>"010010011",
  24070=>"000000000",
  24071=>"111111111",
  24072=>"000000000",
  24073=>"111111111",
  24074=>"111111111",
  24075=>"111111000",
  24076=>"111111111",
  24077=>"011111111",
  24078=>"000000000",
  24079=>"111111111",
  24080=>"111111111",
  24081=>"111111111",
  24082=>"000000000",
  24083=>"111101101",
  24084=>"100110111",
  24085=>"000000000",
  24086=>"111111111",
  24087=>"101001001",
  24088=>"011011111",
  24089=>"000111101",
  24090=>"111111111",
  24091=>"100000000",
  24092=>"111111111",
  24093=>"111011001",
  24094=>"000001001",
  24095=>"001001111",
  24096=>"110000000",
  24097=>"111000110",
  24098=>"111111001",
  24099=>"111111010",
  24100=>"000011111",
  24101=>"111111110",
  24102=>"000011011",
  24103=>"000000000",
  24104=>"000000000",
  24105=>"000000000",
  24106=>"111101101",
  24107=>"000000000",
  24108=>"101111111",
  24109=>"100000000",
  24110=>"010001011",
  24111=>"111011011",
  24112=>"000000000",
  24113=>"111111111",
  24114=>"111111111",
  24115=>"000000000",
  24116=>"111111000",
  24117=>"111111100",
  24118=>"000000000",
  24119=>"111111011",
  24120=>"101111111",
  24121=>"111111000",
  24122=>"000000000",
  24123=>"000111110",
  24124=>"100000000",
  24125=>"000000000",
  24126=>"111111111",
  24127=>"111111111",
  24128=>"000000000",
  24129=>"111111011",
  24130=>"000000000",
  24131=>"001001000",
  24132=>"000001000",
  24133=>"100110110",
  24134=>"111000001",
  24135=>"001101111",
  24136=>"001111011",
  24137=>"000000000",
  24138=>"111111111",
  24139=>"001000000",
  24140=>"000000111",
  24141=>"111011000",
  24142=>"000000000",
  24143=>"011000100",
  24144=>"011111111",
  24145=>"111111000",
  24146=>"001011011",
  24147=>"000000000",
  24148=>"011011001",
  24149=>"000000110",
  24150=>"111111110",
  24151=>"011000010",
  24152=>"001001001",
  24153=>"000000000",
  24154=>"101011110",
  24155=>"001000000",
  24156=>"111111111",
  24157=>"010110111",
  24158=>"111101100",
  24159=>"000000001",
  24160=>"000000000",
  24161=>"000000000",
  24162=>"000000000",
  24163=>"110110011",
  24164=>"111110100",
  24165=>"000000001",
  24166=>"111111001",
  24167=>"111000000",
  24168=>"000000000",
  24169=>"111111111",
  24170=>"001000000",
  24171=>"111111111",
  24172=>"011001000",
  24173=>"111000000",
  24174=>"000000101",
  24175=>"000000000",
  24176=>"110000111",
  24177=>"000100100",
  24178=>"000000001",
  24179=>"000000111",
  24180=>"111111111",
  24181=>"000001000",
  24182=>"000000000",
  24183=>"111111000",
  24184=>"111111111",
  24185=>"111111111",
  24186=>"001000001",
  24187=>"001011111",
  24188=>"000000001",
  24189=>"000001111",
  24190=>"000000000",
  24191=>"001001101",
  24192=>"000000000",
  24193=>"111111110",
  24194=>"000000000",
  24195=>"101101110",
  24196=>"111110111",
  24197=>"100000100",
  24198=>"000110000",
  24199=>"010000000",
  24200=>"000000000",
  24201=>"010000000",
  24202=>"111010111",
  24203=>"000011111",
  24204=>"000000000",
  24205=>"110110000",
  24206=>"000000000",
  24207=>"000100110",
  24208=>"000000111",
  24209=>"011001111",
  24210=>"011111111",
  24211=>"111011001",
  24212=>"000000100",
  24213=>"001000110",
  24214=>"010111111",
  24215=>"111101100",
  24216=>"001111111",
  24217=>"000111000",
  24218=>"111000000",
  24219=>"010000000",
  24220=>"111111111",
  24221=>"111011001",
  24222=>"011011000",
  24223=>"111110000",
  24224=>"000000000",
  24225=>"000000000",
  24226=>"010111110",
  24227=>"111111111",
  24228=>"001001001",
  24229=>"011111110",
  24230=>"111111111",
  24231=>"011001100",
  24232=>"000010000",
  24233=>"001001000",
  24234=>"000000000",
  24235=>"000000000",
  24236=>"011111100",
  24237=>"111111110",
  24238=>"011010111",
  24239=>"000000000",
  24240=>"111111111",
  24241=>"001011001",
  24242=>"111111110",
  24243=>"111110100",
  24244=>"111111111",
  24245=>"110100100",
  24246=>"111111111",
  24247=>"000000110",
  24248=>"111000000",
  24249=>"111111111",
  24250=>"111011010",
  24251=>"011110110",
  24252=>"000000000",
  24253=>"000000111",
  24254=>"000000000",
  24255=>"001000000",
  24256=>"001011011",
  24257=>"111111111",
  24258=>"111111111",
  24259=>"111111111",
  24260=>"000000000",
  24261=>"000100000",
  24262=>"111111000",
  24263=>"111111111",
  24264=>"000001000",
  24265=>"111111111",
  24266=>"000000000",
  24267=>"111111111",
  24268=>"001000100",
  24269=>"000000000",
  24270=>"111111111",
  24271=>"001000000",
  24272=>"000110100",
  24273=>"011000000",
  24274=>"111111111",
  24275=>"001000000",
  24276=>"000000000",
  24277=>"001001000",
  24278=>"110111111",
  24279=>"000000000",
  24280=>"111111000",
  24281=>"000011110",
  24282=>"110000000",
  24283=>"000000111",
  24284=>"001111111",
  24285=>"000001111",
  24286=>"111110111",
  24287=>"000000000",
  24288=>"100000110",
  24289=>"000000000",
  24290=>"111111111",
  24291=>"000000110",
  24292=>"000000010",
  24293=>"110110100",
  24294=>"000000000",
  24295=>"001000101",
  24296=>"111111111",
  24297=>"001001001",
  24298=>"110111111",
  24299=>"001110000",
  24300=>"111111101",
  24301=>"111000000",
  24302=>"111011001",
  24303=>"111000000",
  24304=>"001111001",
  24305=>"000111111",
  24306=>"111111111",
  24307=>"000010000",
  24308=>"000000000",
  24309=>"111111110",
  24310=>"011001001",
  24311=>"111111000",
  24312=>"000101111",
  24313=>"110100111",
  24314=>"000000000",
  24315=>"000000000",
  24316=>"001001001",
  24317=>"111011100",
  24318=>"011111111",
  24319=>"001000000",
  24320=>"001010000",
  24321=>"111111111",
  24322=>"000000000",
  24323=>"000100100",
  24324=>"000000110",
  24325=>"000110110",
  24326=>"100101000",
  24327=>"000000111",
  24328=>"110111111",
  24329=>"111111111",
  24330=>"000011000",
  24331=>"001011000",
  24332=>"110110110",
  24333=>"111111010",
  24334=>"000000000",
  24335=>"111101101",
  24336=>"000110111",
  24337=>"110010100",
  24338=>"000000000",
  24339=>"000010010",
  24340=>"011011110",
  24341=>"111100111",
  24342=>"001000000",
  24343=>"000001111",
  24344=>"011011111",
  24345=>"111111111",
  24346=>"001011000",
  24347=>"111111110",
  24348=>"010011110",
  24349=>"000000000",
  24350=>"110111110",
  24351=>"000010111",
  24352=>"000100100",
  24353=>"000010111",
  24354=>"000000000",
  24355=>"000001000",
  24356=>"000111111",
  24357=>"000000101",
  24358=>"000000100",
  24359=>"000000101",
  24360=>"000000000",
  24361=>"110110000",
  24362=>"111111111",
  24363=>"100000000",
  24364=>"100000000",
  24365=>"111111100",
  24366=>"011111111",
  24367=>"001000001",
  24368=>"011011000",
  24369=>"111111000",
  24370=>"000000000",
  24371=>"000000111",
  24372=>"001001011",
  24373=>"011001000",
  24374=>"000000100",
  24375=>"111011111",
  24376=>"000000000",
  24377=>"100001111",
  24378=>"001000000",
  24379=>"000111111",
  24380=>"000000000",
  24381=>"000010110",
  24382=>"111011111",
  24383=>"000000000",
  24384=>"001000000",
  24385=>"111111101",
  24386=>"111111101",
  24387=>"000000000",
  24388=>"000011000",
  24389=>"000100001",
  24390=>"111111111",
  24391=>"000111111",
  24392=>"111111001",
  24393=>"011000000",
  24394=>"011111111",
  24395=>"000001001",
  24396=>"000000000",
  24397=>"111111100",
  24398=>"000111111",
  24399=>"000011011",
  24400=>"000100000",
  24401=>"001000000",
  24402=>"001001011",
  24403=>"000000000",
  24404=>"110111111",
  24405=>"111111011",
  24406=>"000000000",
  24407=>"000000000",
  24408=>"111111111",
  24409=>"111111111",
  24410=>"010000000",
  24411=>"000000000",
  24412=>"000000100",
  24413=>"000000000",
  24414=>"111011111",
  24415=>"000000000",
  24416=>"000001010",
  24417=>"000001111",
  24418=>"101100100",
  24419=>"111111111",
  24420=>"000001001",
  24421=>"001000000",
  24422=>"111111111",
  24423=>"111111000",
  24424=>"000000000",
  24425=>"000000000",
  24426=>"111001001",
  24427=>"000000000",
  24428=>"011111111",
  24429=>"111000000",
  24430=>"111111100",
  24431=>"000000000",
  24432=>"111111101",
  24433=>"011011011",
  24434=>"111111111",
  24435=>"110111111",
  24436=>"000000000",
  24437=>"000001000",
  24438=>"111111111",
  24439=>"111000110",
  24440=>"000000110",
  24441=>"110110111",
  24442=>"001111111",
  24443=>"100000000",
  24444=>"000000110",
  24445=>"000000000",
  24446=>"000101111",
  24447=>"000000000",
  24448=>"000000000",
  24449=>"000011111",
  24450=>"011111111",
  24451=>"111111111",
  24452=>"111111111",
  24453=>"000000000",
  24454=>"000000000",
  24455=>"000000111",
  24456=>"000000000",
  24457=>"001001000",
  24458=>"000000000",
  24459=>"111101111",
  24460=>"011111000",
  24461=>"100101111",
  24462=>"000000000",
  24463=>"000000000",
  24464=>"100111110",
  24465=>"000111111",
  24466=>"110111101",
  24467=>"000000011",
  24468=>"000000000",
  24469=>"000000000",
  24470=>"000011111",
  24471=>"000000000",
  24472=>"000110110",
  24473=>"000000001",
  24474=>"001111000",
  24475=>"111111111",
  24476=>"000000000",
  24477=>"010111000",
  24478=>"010000000",
  24479=>"000000000",
  24480=>"010010000",
  24481=>"010000110",
  24482=>"000000000",
  24483=>"000000000",
  24484=>"111111110",
  24485=>"110111111",
  24486=>"000000111",
  24487=>"111111111",
  24488=>"000000000",
  24489=>"000000000",
  24490=>"101001000",
  24491=>"001000000",
  24492=>"000000000",
  24493=>"111111111",
  24494=>"000000001",
  24495=>"000000111",
  24496=>"111111101",
  24497=>"111111111",
  24498=>"110011111",
  24499=>"000011110",
  24500=>"100000111",
  24501=>"100000000",
  24502=>"011011111",
  24503=>"010011111",
  24504=>"000000000",
  24505=>"111111111",
  24506=>"111010000",
  24507=>"011111111",
  24508=>"000000000",
  24509=>"100000100",
  24510=>"100000000",
  24511=>"001001000",
  24512=>"111111110",
  24513=>"100110110",
  24514=>"010010110",
  24515=>"110111111",
  24516=>"011001000",
  24517=>"011011001",
  24518=>"000000000",
  24519=>"100110111",
  24520=>"000011000",
  24521=>"111111110",
  24522=>"000111010",
  24523=>"000000000",
  24524=>"000000000",
  24525=>"001001000",
  24526=>"111111111",
  24527=>"000000010",
  24528=>"100000000",
  24529=>"100110110",
  24530=>"000000000",
  24531=>"111111111",
  24532=>"000110110",
  24533=>"010011000",
  24534=>"000000000",
  24535=>"110111111",
  24536=>"000000100",
  24537=>"011011000",
  24538=>"111111111",
  24539=>"111111111",
  24540=>"010010111",
  24541=>"001000000",
  24542=>"111111111",
  24543=>"000000000",
  24544=>"111110100",
  24545=>"111111100",
  24546=>"111111011",
  24547=>"000000000",
  24548=>"011111111",
  24549=>"111101000",
  24550=>"000000000",
  24551=>"000110110",
  24552=>"000011111",
  24553=>"111001011",
  24554=>"011110111",
  24555=>"010000100",
  24556=>"010000011",
  24557=>"101000000",
  24558=>"111111111",
  24559=>"111000000",
  24560=>"000000000",
  24561=>"000000000",
  24562=>"000000000",
  24563=>"000000000",
  24564=>"111111111",
  24565=>"000000000",
  24566=>"001000000",
  24567=>"111111111",
  24568=>"000100000",
  24569=>"000000001",
  24570=>"001001111",
  24571=>"000000000",
  24572=>"000000000",
  24573=>"010000111",
  24574=>"011111111",
  24575=>"100110111",
  24576=>"011110010",
  24577=>"000000010",
  24578=>"011111111",
  24579=>"000100101",
  24580=>"011110000",
  24581=>"111000101",
  24582=>"000000001",
  24583=>"110111111",
  24584=>"111111110",
  24585=>"001001001",
  24586=>"000110110",
  24587=>"100100000",
  24588=>"100111001",
  24589=>"111111111",
  24590=>"101100111",
  24591=>"000011111",
  24592=>"111001000",
  24593=>"000111110",
  24594=>"100100000",
  24595=>"000100000",
  24596=>"000000001",
  24597=>"101000100",
  24598=>"111111001",
  24599=>"000000100",
  24600=>"111101000",
  24601=>"100111000",
  24602=>"111110100",
  24603=>"111001001",
  24604=>"000000111",
  24605=>"100111001",
  24606=>"110110000",
  24607=>"111000110",
  24608=>"110110010",
  24609=>"111011010",
  24610=>"000000010",
  24611=>"111001000",
  24612=>"000000000",
  24613=>"111111111",
  24614=>"111011111",
  24615=>"000000000",
  24616=>"001001111",
  24617=>"000000000",
  24618=>"000000010",
  24619=>"111001001",
  24620=>"000111110",
  24621=>"000000000",
  24622=>"000000000",
  24623=>"111000000",
  24624=>"011111110",
  24625=>"000000101",
  24626=>"111001000",
  24627=>"111111111",
  24628=>"111111000",
  24629=>"100000000",
  24630=>"000000000",
  24631=>"001001011",
  24632=>"111111110",
  24633=>"111100001",
  24634=>"000000000",
  24635=>"000010011",
  24636=>"001001000",
  24637=>"111111111",
  24638=>"000110011",
  24639=>"000000111",
  24640=>"000001111",
  24641=>"001000111",
  24642=>"000000000",
  24643=>"000000000",
  24644=>"111011000",
  24645=>"001011011",
  24646=>"000000111",
  24647=>"111001000",
  24648=>"111111100",
  24649=>"101101000",
  24650=>"111111011",
  24651=>"010010111",
  24652=>"111110110",
  24653=>"101111111",
  24654=>"001000000",
  24655=>"111001011",
  24656=>"110000011",
  24657=>"111111111",
  24658=>"100000000",
  24659=>"000000110",
  24660=>"000111111",
  24661=>"000000101",
  24662=>"000000100",
  24663=>"000000010",
  24664=>"111000010",
  24665=>"111101101",
  24666=>"111011110",
  24667=>"001001001",
  24668=>"000000010",
  24669=>"111111111",
  24670=>"010000000",
  24671=>"111011011",
  24672=>"010010010",
  24673=>"111000001",
  24674=>"010110000",
  24675=>"011111111",
  24676=>"001001100",
  24677=>"111111110",
  24678=>"111111011",
  24679=>"111111111",
  24680=>"001000111",
  24681=>"000000010",
  24682=>"100001111",
  24683=>"111111111",
  24684=>"001001000",
  24685=>"000000000",
  24686=>"000000001",
  24687=>"101111111",
  24688=>"001000000",
  24689=>"000100111",
  24690=>"000000000",
  24691=>"100000110",
  24692=>"010000111",
  24693=>"000000001",
  24694=>"000110111",
  24695=>"000000000",
  24696=>"000000001",
  24697=>"100000001",
  24698=>"000000100",
  24699=>"100101111",
  24700=>"001101001",
  24701=>"000000000",
  24702=>"000000000",
  24703=>"000100000",
  24704=>"000000000",
  24705=>"111110111",
  24706=>"111011000",
  24707=>"000000001",
  24708=>"111111011",
  24709=>"101101111",
  24710=>"000000000",
  24711=>"000000111",
  24712=>"111111001",
  24713=>"111101000",
  24714=>"000000000",
  24715=>"100000011",
  24716=>"000000000",
  24717=>"101111111",
  24718=>"111111110",
  24719=>"000000000",
  24720=>"111111111",
  24721=>"111011111",
  24722=>"001000000",
  24723=>"000100110",
  24724=>"000000101",
  24725=>"000001010",
  24726=>"100110111",
  24727=>"000000001",
  24728=>"001011111",
  24729=>"000110111",
  24730=>"111111010",
  24731=>"011010110",
  24732=>"111000000",
  24733=>"100110001",
  24734=>"000001000",
  24735=>"111111111",
  24736=>"110100100",
  24737=>"000000001",
  24738=>"000001111",
  24739=>"111110010",
  24740=>"111011111",
  24741=>"000000000",
  24742=>"000000101",
  24743=>"110100100",
  24744=>"111100001",
  24745=>"001101111",
  24746=>"111100100",
  24747=>"111000000",
  24748=>"011000001",
  24749=>"001001011",
  24750=>"001001000",
  24751=>"111111010",
  24752=>"000110000",
  24753=>"001100000",
  24754=>"111111111",
  24755=>"111001000",
  24756=>"111111111",
  24757=>"110100000",
  24758=>"000000000",
  24759=>"011011111",
  24760=>"111110111",
  24761=>"001111111",
  24762=>"000000001",
  24763=>"111011011",
  24764=>"111001111",
  24765=>"001001001",
  24766=>"100110010",
  24767=>"000010000",
  24768=>"100100000",
  24769=>"111111010",
  24770=>"101000001",
  24771=>"111111111",
  24772=>"111111111",
  24773=>"010111010",
  24774=>"000001111",
  24775=>"010000000",
  24776=>"000000000",
  24777=>"110111111",
  24778=>"001011111",
  24779=>"000000000",
  24780=>"101101101",
  24781=>"001011111",
  24782=>"001001011",
  24783=>"000001001",
  24784=>"000000000",
  24785=>"000000000",
  24786=>"000011011",
  24787=>"000000000",
  24788=>"100001111",
  24789=>"111111111",
  24790=>"111111110",
  24791=>"000000000",
  24792=>"000000001",
  24793=>"011001011",
  24794=>"101101111",
  24795=>"111100000",
  24796=>"111111111",
  24797=>"110111000",
  24798=>"111110110",
  24799=>"111111111",
  24800=>"000000100",
  24801=>"000000110",
  24802=>"000000000",
  24803=>"100000000",
  24804=>"000000010",
  24805=>"000000000",
  24806=>"000000000",
  24807=>"111010000",
  24808=>"000000000",
  24809=>"010000110",
  24810=>"000000000",
  24811=>"111111011",
  24812=>"111111110",
  24813=>"111111111",
  24814=>"110111010",
  24815=>"000000111",
  24816=>"000000000",
  24817=>"111111111",
  24818=>"111111111",
  24819=>"011000110",
  24820=>"000000000",
  24821=>"111111110",
  24822=>"000110010",
  24823=>"111111111",
  24824=>"000100110",
  24825=>"000000000",
  24826=>"000000100",
  24827=>"100110100",
  24828=>"001001001",
  24829=>"001011111",
  24830=>"000000100",
  24831=>"111001001",
  24832=>"111001001",
  24833=>"000001000",
  24834=>"000000011",
  24835=>"111111111",
  24836=>"000000001",
  24837=>"011000000",
  24838=>"000111111",
  24839=>"000010100",
  24840=>"000000001",
  24841=>"011011000",
  24842=>"111111111",
  24843=>"110110110",
  24844=>"101101101",
  24845=>"111010000",
  24846=>"111111111",
  24847=>"101101000",
  24848=>"100100110",
  24849=>"111111000",
  24850=>"000101101",
  24851=>"000000000",
  24852=>"111110000",
  24853=>"000000000",
  24854=>"110111001",
  24855=>"111110010",
  24856=>"111111111",
  24857=>"100010000",
  24858=>"010110000",
  24859=>"010011001",
  24860=>"111111111",
  24861=>"011000000",
  24862=>"111111111",
  24863=>"111111011",
  24864=>"000111111",
  24865=>"111110000",
  24866=>"000111011",
  24867=>"011001111",
  24868=>"111111111",
  24869=>"011011111",
  24870=>"111100000",
  24871=>"110010111",
  24872=>"111111000",
  24873=>"111111010",
  24874=>"100000000",
  24875=>"111111111",
  24876=>"010010111",
  24877=>"001001001",
  24878=>"000000000",
  24879=>"000000000",
  24880=>"000000000",
  24881=>"000000000",
  24882=>"111001011",
  24883=>"110110111",
  24884=>"000000000",
  24885=>"111110111",
  24886=>"000000000",
  24887=>"000000000",
  24888=>"000000000",
  24889=>"101101101",
  24890=>"011000000",
  24891=>"000000011",
  24892=>"000000000",
  24893=>"000011111",
  24894=>"111111111",
  24895=>"111111011",
  24896=>"000001111",
  24897=>"111111000",
  24898=>"000000001",
  24899=>"000001011",
  24900=>"011001100",
  24901=>"111111111",
  24902=>"001001001",
  24903=>"000010000",
  24904=>"000000000",
  24905=>"000000010",
  24906=>"111011000",
  24907=>"100110110",
  24908=>"100000000",
  24909=>"110111110",
  24910=>"111110010",
  24911=>"000000001",
  24912=>"011111111",
  24913=>"111110110",
  24914=>"000000000",
  24915=>"000000000",
  24916=>"100000000",
  24917=>"011011001",
  24918=>"100000000",
  24919=>"000000100",
  24920=>"001011111",
  24921=>"000000000",
  24922=>"111000000",
  24923=>"110110100",
  24924=>"000101000",
  24925=>"000000001",
  24926=>"000000001",
  24927=>"011001000",
  24928=>"000000100",
  24929=>"011001001",
  24930=>"111111011",
  24931=>"001001100",
  24932=>"111111000",
  24933=>"111111111",
  24934=>"000000111",
  24935=>"111111111",
  24936=>"001001011",
  24937=>"010000001",
  24938=>"110110000",
  24939=>"000000000",
  24940=>"111110110",
  24941=>"000000001",
  24942=>"101000000",
  24943=>"111010000",
  24944=>"111111111",
  24945=>"000000000",
  24946=>"111001101",
  24947=>"000000001",
  24948=>"000000000",
  24949=>"011011001",
  24950=>"101100100",
  24951=>"110000000",
  24952=>"000001001",
  24953=>"000000111",
  24954=>"111111001",
  24955=>"111010000",
  24956=>"110000010",
  24957=>"000000000",
  24958=>"111111010",
  24959=>"001000000",
  24960=>"000000000",
  24961=>"010111111",
  24962=>"110110110",
  24963=>"001010011",
  24964=>"111111111",
  24965=>"001001001",
  24966=>"000001111",
  24967=>"111111111",
  24968=>"000001001",
  24969=>"111111101",
  24970=>"011111111",
  24971=>"011000000",
  24972=>"101101111",
  24973=>"000000001",
  24974=>"010000100",
  24975=>"000110010",
  24976=>"011010000",
  24977=>"100000000",
  24978=>"000000000",
  24979=>"000000000",
  24980=>"001000010",
  24981=>"000000000",
  24982=>"100000000",
  24983=>"111011111",
  24984=>"110001011",
  24985=>"000000011",
  24986=>"001101111",
  24987=>"111111101",
  24988=>"000000101",
  24989=>"111111111",
  24990=>"000000000",
  24991=>"000000011",
  24992=>"111111100",
  24993=>"111111000",
  24994=>"011000101",
  24995=>"000111111",
  24996=>"000000100",
  24997=>"000000000",
  24998=>"111111111",
  24999=>"111110111",
  25000=>"000010000",
  25001=>"111110110",
  25002=>"000000000",
  25003=>"000000000",
  25004=>"000000000",
  25005=>"100101001",
  25006=>"111110111",
  25007=>"000000000",
  25008=>"111001101",
  25009=>"100100000",
  25010=>"111110010",
  25011=>"111100000",
  25012=>"110110100",
  25013=>"000000000",
  25014=>"111111111",
  25015=>"111110100",
  25016=>"001001011",
  25017=>"110110111",
  25018=>"001011010",
  25019=>"001001001",
  25020=>"000111111",
  25021=>"111111111",
  25022=>"000000001",
  25023=>"100110100",
  25024=>"000000111",
  25025=>"000000011",
  25026=>"011000000",
  25027=>"000000000",
  25028=>"111111111",
  25029=>"111111111",
  25030=>"000000000",
  25031=>"000110111",
  25032=>"111101111",
  25033=>"000000000",
  25034=>"000000111",
  25035=>"011111001",
  25036=>"000000000",
  25037=>"111111111",
  25038=>"001001000",
  25039=>"100110111",
  25040=>"000000000",
  25041=>"111111111",
  25042=>"000000000",
  25043=>"000000111",
  25044=>"111110000",
  25045=>"000000000",
  25046=>"010000000",
  25047=>"011011111",
  25048=>"111101001",
  25049=>"001000001",
  25050=>"110010000",
  25051=>"000111111",
  25052=>"000000000",
  25053=>"010110000",
  25054=>"000001000",
  25055=>"100100100",
  25056=>"000100110",
  25057=>"000000000",
  25058=>"000000000",
  25059=>"101000000",
  25060=>"111111000",
  25061=>"111111110",
  25062=>"000000111",
  25063=>"000101111",
  25064=>"000000101",
  25065=>"000000110",
  25066=>"000001000",
  25067=>"000101111",
  25068=>"000000001",
  25069=>"000101110",
  25070=>"111111001",
  25071=>"000110000",
  25072=>"000000000",
  25073=>"000000000",
  25074=>"000111111",
  25075=>"111111011",
  25076=>"110111011",
  25077=>"000000000",
  25078=>"111111111",
  25079=>"110110000",
  25080=>"011111100",
  25081=>"011001001",
  25082=>"000110111",
  25083=>"101000001",
  25084=>"000101000",
  25085=>"010000001",
  25086=>"010100101",
  25087=>"000000000",
  25088=>"111101100",
  25089=>"101111111",
  25090=>"110111111",
  25091=>"000000000",
  25092=>"011011001",
  25093=>"000000000",
  25094=>"011001011",
  25095=>"111111111",
  25096=>"111111111",
  25097=>"000000010",
  25098=>"111111111",
  25099=>"011000011",
  25100=>"111111110",
  25101=>"000000111",
  25102=>"001001111",
  25103=>"000001001",
  25104=>"110001001",
  25105=>"000000011",
  25106=>"111100000",
  25107=>"111111000",
  25108=>"110110010",
  25109=>"110111110",
  25110=>"111111111",
  25111=>"110111111",
  25112=>"000000100",
  25113=>"000000000",
  25114=>"010110110",
  25115=>"000100000",
  25116=>"110111111",
  25117=>"110000000",
  25118=>"001001000",
  25119=>"111111011",
  25120=>"000001000",
  25121=>"111111111",
  25122=>"000000100",
  25123=>"100001111",
  25124=>"111110010",
  25125=>"111000000",
  25126=>"000000000",
  25127=>"001001111",
  25128=>"000000000",
  25129=>"010010000",
  25130=>"111111111",
  25131=>"000000000",
  25132=>"001000111",
  25133=>"000001001",
  25134=>"001111110",
  25135=>"111111000",
  25136=>"100100000",
  25137=>"000000111",
  25138=>"111101001",
  25139=>"000111110",
  25140=>"000000010",
  25141=>"011111111",
  25142=>"111111000",
  25143=>"011000100",
  25144=>"111111110",
  25145=>"101000111",
  25146=>"000000000",
  25147=>"000000000",
  25148=>"000000000",
  25149=>"000001110",
  25150=>"111111111",
  25151=>"000000101",
  25152=>"100100111",
  25153=>"000010010",
  25154=>"101001111",
  25155=>"000000000",
  25156=>"000001111",
  25157=>"011111111",
  25158=>"111100000",
  25159=>"111111111",
  25160=>"111111111",
  25161=>"000000100",
  25162=>"000001001",
  25163=>"111011111",
  25164=>"000000000",
  25165=>"000010000",
  25166=>"010001000",
  25167=>"111100111",
  25168=>"111011111",
  25169=>"000110111",
  25170=>"111111000",
  25171=>"100111111",
  25172=>"000010000",
  25173=>"101111111",
  25174=>"101100000",
  25175=>"100100111",
  25176=>"100000000",
  25177=>"000000000",
  25178=>"110010000",
  25179=>"111111111",
  25180=>"000000001",
  25181=>"110000101",
  25182=>"010001111",
  25183=>"111111110",
  25184=>"000000000",
  25185=>"000000111",
  25186=>"000110000",
  25187=>"111001111",
  25188=>"111111111",
  25189=>"111111111",
  25190=>"000000000",
  25191=>"000110111",
  25192=>"000000011",
  25193=>"111111111",
  25194=>"111100110",
  25195=>"111011011",
  25196=>"110110110",
  25197=>"111111111",
  25198=>"111111110",
  25199=>"100000000",
  25200=>"000010000",
  25201=>"000000000",
  25202=>"000100111",
  25203=>"100100000",
  25204=>"111111000",
  25205=>"000000111",
  25206=>"111111110",
  25207=>"011010111",
  25208=>"000100111",
  25209=>"110100100",
  25210=>"000111111",
  25211=>"000000000",
  25212=>"000100110",
  25213=>"011111011",
  25214=>"000000111",
  25215=>"000000000",
  25216=>"000000000",
  25217=>"111111110",
  25218=>"110000011",
  25219=>"111111101",
  25220=>"000111111",
  25221=>"000000001",
  25222=>"000001001",
  25223=>"111000000",
  25224=>"111001000",
  25225=>"000001001",
  25226=>"001000001",
  25227=>"000000000",
  25228=>"000001111",
  25229=>"101101001",
  25230=>"001001111",
  25231=>"000001000",
  25232=>"110000011",
  25233=>"110110110",
  25234=>"111011011",
  25235=>"001111111",
  25236=>"000100000",
  25237=>"010000000",
  25238=>"111111111",
  25239=>"111111111",
  25240=>"001011111",
  25241=>"111111111",
  25242=>"111111111",
  25243=>"000000000",
  25244=>"000000000",
  25245=>"011011011",
  25246=>"111000000",
  25247=>"111101000",
  25248=>"100100000",
  25249=>"000000000",
  25250=>"000000000",
  25251=>"011011011",
  25252=>"011011111",
  25253=>"010010011",
  25254=>"000000000",
  25255=>"000001111",
  25256=>"000000000",
  25257=>"111110111",
  25258=>"000000000",
  25259=>"110110110",
  25260=>"000000111",
  25261=>"000100001",
  25262=>"000100011",
  25263=>"011111111",
  25264=>"111111000",
  25265=>"000000000",
  25266=>"111000111",
  25267=>"000000000",
  25268=>"010000000",
  25269=>"111011000",
  25270=>"000000001",
  25271=>"000000000",
  25272=>"111111111",
  25273=>"000000111",
  25274=>"100111111",
  25275=>"011011111",
  25276=>"111111111",
  25277=>"010000100",
  25278=>"000000000",
  25279=>"110101001",
  25280=>"001000000",
  25281=>"111111100",
  25282=>"011000000",
  25283=>"111011000",
  25284=>"000000101",
  25285=>"110111111",
  25286=>"000000110",
  25287=>"101111001",
  25288=>"010000000",
  25289=>"111001000",
  25290=>"101100001",
  25291=>"000001111",
  25292=>"001000001",
  25293=>"000000100",
  25294=>"111000000",
  25295=>"000000000",
  25296=>"011100000",
  25297=>"000001001",
  25298=>"111011011",
  25299=>"110111111",
  25300=>"001101101",
  25301=>"110100111",
  25302=>"111111111",
  25303=>"111111111",
  25304=>"111111111",
  25305=>"011000000",
  25306=>"000000000",
  25307=>"111111111",
  25308=>"111111111",
  25309=>"111111110",
  25310=>"000111111",
  25311=>"111110100",
  25312=>"000000000",
  25313=>"000000000",
  25314=>"111111111",
  25315=>"001001011",
  25316=>"111111100",
  25317=>"111111001",
  25318=>"100000000",
  25319=>"001000100",
  25320=>"111111111",
  25321=>"001000111",
  25322=>"000011011",
  25323=>"000000101",
  25324=>"111111111",
  25325=>"000001111",
  25326=>"000000111",
  25327=>"111111111",
  25328=>"000000000",
  25329=>"011001111",
  25330=>"011001000",
  25331=>"111110000",
  25332=>"111101000",
  25333=>"111111111",
  25334=>"000001001",
  25335=>"110110111",
  25336=>"000000000",
  25337=>"110110111",
  25338=>"111110111",
  25339=>"000001001",
  25340=>"111111111",
  25341=>"001000111",
  25342=>"110000000",
  25343=>"000010010",
  25344=>"111011111",
  25345=>"110110110",
  25346=>"101000000",
  25347=>"000000000",
  25348=>"000000100",
  25349=>"000110110",
  25350=>"000000000",
  25351=>"111111111",
  25352=>"110110111",
  25353=>"000000000",
  25354=>"111111111",
  25355=>"111100100",
  25356=>"001001111",
  25357=>"000000110",
  25358=>"110111111",
  25359=>"111111010",
  25360=>"011111101",
  25361=>"010110000",
  25362=>"111111111",
  25363=>"011011011",
  25364=>"111101000",
  25365=>"000001111",
  25366=>"111111101",
  25367=>"000000000",
  25368=>"001001111",
  25369=>"001111011",
  25370=>"111000011",
  25371=>"011110110",
  25372=>"001001001",
  25373=>"000000000",
  25374=>"111111111",
  25375=>"110100110",
  25376=>"001000111",
  25377=>"110110110",
  25378=>"110100000",
  25379=>"000000010",
  25380=>"000001111",
  25381=>"011111011",
  25382=>"011111111",
  25383=>"000000000",
  25384=>"111111111",
  25385=>"110111111",
  25386=>"000000100",
  25387=>"000000000",
  25388=>"000100110",
  25389=>"111111111",
  25390=>"000000111",
  25391=>"011000011",
  25392=>"000000000",
  25393=>"110110111",
  25394=>"100000000",
  25395=>"100110110",
  25396=>"111001011",
  25397=>"110110100",
  25398=>"110110000",
  25399=>"110111111",
  25400=>"000000111",
  25401=>"000000100",
  25402=>"000000000",
  25403=>"111110110",
  25404=>"111111111",
  25405=>"000000000",
  25406=>"100100000",
  25407=>"001111001",
  25408=>"000000000",
  25409=>"000000000",
  25410=>"111111111",
  25411=>"101111000",
  25412=>"101110111",
  25413=>"100100110",
  25414=>"000000000",
  25415=>"111111111",
  25416=>"100000000",
  25417=>"000000000",
  25418=>"000001011",
  25419=>"000100100",
  25420=>"111111000",
  25421=>"111111111",
  25422=>"111000100",
  25423=>"111111111",
  25424=>"111011111",
  25425=>"111111111",
  25426=>"111111111",
  25427=>"000000000",
  25428=>"000000000",
  25429=>"011011011",
  25430=>"111111111",
  25431=>"000000000",
  25432=>"111101001",
  25433=>"111111111",
  25434=>"001000011",
  25435=>"011011111",
  25436=>"011011111",
  25437=>"000111111",
  25438=>"111111001",
  25439=>"000000111",
  25440=>"111111011",
  25441=>"100110000",
  25442=>"001110100",
  25443=>"000000000",
  25444=>"000110111",
  25445=>"000000000",
  25446=>"000000111",
  25447=>"111111111",
  25448=>"000001001",
  25449=>"101100111",
  25450=>"111111010",
  25451=>"111111111",
  25452=>"100000100",
  25453=>"100111111",
  25454=>"110010000",
  25455=>"100000000",
  25456=>"000000000",
  25457=>"111111111",
  25458=>"000000000",
  25459=>"111111111",
  25460=>"110111011",
  25461=>"101111000",
  25462=>"111111111",
  25463=>"000000100",
  25464=>"111101100",
  25465=>"000000011",
  25466=>"110110111",
  25467=>"000000000",
  25468=>"000000001",
  25469=>"000000100",
  25470=>"000000000",
  25471=>"111111111",
  25472=>"110110110",
  25473=>"100111101",
  25474=>"010111111",
  25475=>"000000000",
  25476=>"110000110",
  25477=>"001001001",
  25478=>"000000100",
  25479=>"100101101",
  25480=>"111111111",
  25481=>"100101001",
  25482=>"111111000",
  25483=>"111000000",
  25484=>"100000000",
  25485=>"001001111",
  25486=>"111111111",
  25487=>"111011001",
  25488=>"000000000",
  25489=>"000000100",
  25490=>"110111110",
  25491=>"110111111",
  25492=>"111110110",
  25493=>"000010000",
  25494=>"000000100",
  25495=>"001001001",
  25496=>"100111110",
  25497=>"000000000",
  25498=>"000000000",
  25499=>"111111110",
  25500=>"111000000",
  25501=>"000000000",
  25502=>"000000111",
  25503=>"111111111",
  25504=>"000010110",
  25505=>"110110110",
  25506=>"111001010",
  25507=>"000000011",
  25508=>"001111111",
  25509=>"100000001",
  25510=>"000000000",
  25511=>"111111111",
  25512=>"011001000",
  25513=>"111111111",
  25514=>"000000000",
  25515=>"111000000",
  25516=>"000111111",
  25517=>"100011011",
  25518=>"000000100",
  25519=>"100100111",
  25520=>"111000111",
  25521=>"111111111",
  25522=>"001001011",
  25523=>"100000111",
  25524=>"100000110",
  25525=>"011111110",
  25526=>"111111111",
  25527=>"001000000",
  25528=>"000111111",
  25529=>"111111111",
  25530=>"000000000",
  25531=>"111111011",
  25532=>"111111111",
  25533=>"001100111",
  25534=>"011000000",
  25535=>"001011110",
  25536=>"001000000",
  25537=>"110010000",
  25538=>"111111111",
  25539=>"100000000",
  25540=>"111111111",
  25541=>"100000000",
  25542=>"100100000",
  25543=>"000000000",
  25544=>"111111111",
  25545=>"100111111",
  25546=>"000100000",
  25547=>"111111111",
  25548=>"000000000",
  25549=>"111110000",
  25550=>"101111011",
  25551=>"111111110",
  25552=>"011011001",
  25553=>"001001001",
  25554=>"000001111",
  25555=>"100101111",
  25556=>"001001001",
  25557=>"111011000",
  25558=>"111110000",
  25559=>"111101011",
  25560=>"001000111",
  25561=>"111001000",
  25562=>"111111111",
  25563=>"111111000",
  25564=>"000100111",
  25565=>"010001001",
  25566=>"111111011",
  25567=>"111111111",
  25568=>"000000111",
  25569=>"101111000",
  25570=>"111111111",
  25571=>"000000000",
  25572=>"111111111",
  25573=>"000000000",
  25574=>"000000011",
  25575=>"110010011",
  25576=>"000000010",
  25577=>"000000000",
  25578=>"000100110",
  25579=>"001001000",
  25580=>"011000010",
  25581=>"000010000",
  25582=>"111110110",
  25583=>"011111111",
  25584=>"111111111",
  25585=>"000000000",
  25586=>"111001000",
  25587=>"110111111",
  25588=>"000000111",
  25589=>"000000000",
  25590=>"100000000",
  25591=>"100001000",
  25592=>"011000000",
  25593=>"100100000",
  25594=>"111111111",
  25595=>"110111110",
  25596=>"110000000",
  25597=>"111111111",
  25598=>"000000000",
  25599=>"001001101",
  25600=>"000000000",
  25601=>"000000000",
  25602=>"111111111",
  25603=>"000000111",
  25604=>"011111111",
  25605=>"111111001",
  25606=>"111111010",
  25607=>"101000000",
  25608=>"100100000",
  25609=>"001000001",
  25610=>"111111101",
  25611=>"111110000",
  25612=>"000110010",
  25613=>"000000000",
  25614=>"000100000",
  25615=>"011011111",
  25616=>"000000000",
  25617=>"010111101",
  25618=>"111111111",
  25619=>"001000000",
  25620=>"111111101",
  25621=>"111000111",
  25622=>"111111111",
  25623=>"001001100",
  25624=>"000000000",
  25625=>"011011011",
  25626=>"100000000",
  25627=>"111111011",
  25628=>"000000000",
  25629=>"111111100",
  25630=>"000001111",
  25631=>"000000000",
  25632=>"011111111",
  25633=>"100111011",
  25634=>"110110110",
  25635=>"001000111",
  25636=>"000001111",
  25637=>"000000000",
  25638=>"000001101",
  25639=>"111111111",
  25640=>"001001000",
  25641=>"110110010",
  25642=>"101111111",
  25643=>"000000000",
  25644=>"111111011",
  25645=>"101100000",
  25646=>"000000000",
  25647=>"100100110",
  25648=>"111111000",
  25649=>"000100000",
  25650=>"100100001",
  25651=>"001011001",
  25652=>"100100000",
  25653=>"110110010",
  25654=>"111101111",
  25655=>"110111111",
  25656=>"011000000",
  25657=>"000000011",
  25658=>"001000101",
  25659=>"111111111",
  25660=>"101001101",
  25661=>"011000100",
  25662=>"111110000",
  25663=>"000000000",
  25664=>"111110000",
  25665=>"000000000",
  25666=>"000000101",
  25667=>"100110111",
  25668=>"000000100",
  25669=>"011111111",
  25670=>"001101001",
  25671=>"111111111",
  25672=>"100101100",
  25673=>"001000101",
  25674=>"001001000",
  25675=>"000000001",
  25676=>"000101000",
  25677=>"000000000",
  25678=>"101111111",
  25679=>"101000000",
  25680=>"000000001",
  25681=>"101111111",
  25682=>"001001000",
  25683=>"000000000",
  25684=>"000001000",
  25685=>"000000000",
  25686=>"000000000",
  25687=>"111111111",
  25688=>"101000000",
  25689=>"101101111",
  25690=>"111111111",
  25691=>"110100100",
  25692=>"000011100",
  25693=>"000000000",
  25694=>"100100110",
  25695=>"001001000",
  25696=>"110000000",
  25697=>"110110110",
  25698=>"010011010",
  25699=>"000110110",
  25700=>"110000000",
  25701=>"111111111",
  25702=>"000000001",
  25703=>"110000000",
  25704=>"000111111",
  25705=>"111111111",
  25706=>"111011011",
  25707=>"000111111",
  25708=>"110000000",
  25709=>"000000000",
  25710=>"111111001",
  25711=>"000000111",
  25712=>"000000000",
  25713=>"111011000",
  25714=>"111100000",
  25715=>"000000111",
  25716=>"000000000",
  25717=>"010111111",
  25718=>"111111110",
  25719=>"000000001",
  25720=>"000000100",
  25721=>"000000100",
  25722=>"000000000",
  25723=>"101101100",
  25724=>"100110110",
  25725=>"000001111",
  25726=>"000000000",
  25727=>"110110101",
  25728=>"111111111",
  25729=>"110000000",
  25730=>"111111111",
  25731=>"101101000",
  25732=>"010000001",
  25733=>"111111111",
  25734=>"111110100",
  25735=>"000000110",
  25736=>"000000111",
  25737=>"101000111",
  25738=>"010010000",
  25739=>"000000000",
  25740=>"000011111",
  25741=>"111110000",
  25742=>"000011111",
  25743=>"110110101",
  25744=>"000000101",
  25745=>"000000000",
  25746=>"100100000",
  25747=>"011011110",
  25748=>"010000000",
  25749=>"111110110",
  25750=>"000000000",
  25751=>"001000100",
  25752=>"000000001",
  25753=>"111111010",
  25754=>"000001111",
  25755=>"111111111",
  25756=>"000000001",
  25757=>"000000000",
  25758=>"111101111",
  25759=>"000000111",
  25760=>"111011101",
  25761=>"111100000",
  25762=>"111111000",
  25763=>"000011011",
  25764=>"000000000",
  25765=>"111111111",
  25766=>"001001100",
  25767=>"011000000",
  25768=>"000111111",
  25769=>"000000000",
  25770=>"001000000",
  25771=>"111111111",
  25772=>"101111111",
  25773=>"100101100",
  25774=>"111111000",
  25775=>"111110110",
  25776=>"111111111",
  25777=>"111111111",
  25778=>"010111111",
  25779=>"011101001",
  25780=>"100100100",
  25781=>"100000000",
  25782=>"000011001",
  25783=>"000000001",
  25784=>"111111111",
  25785=>"000011011",
  25786=>"000000000",
  25787=>"100001001",
  25788=>"111101101",
  25789=>"111111111",
  25790=>"110100100",
  25791=>"000010010",
  25792=>"010111011",
  25793=>"001000001",
  25794=>"101111111",
  25795=>"010110000",
  25796=>"111111001",
  25797=>"000000111",
  25798=>"000000001",
  25799=>"110001000",
  25800=>"111111111",
  25801=>"000000000",
  25802=>"111111000",
  25803=>"101000000",
  25804=>"111111001",
  25805=>"111110111",
  25806=>"111111111",
  25807=>"111110100",
  25808=>"101011010",
  25809=>"101001011",
  25810=>"111111001",
  25811=>"111110110",
  25812=>"100000001",
  25813=>"110111111",
  25814=>"101000000",
  25815=>"111111111",
  25816=>"000000000",
  25817=>"111001111",
  25818=>"111100101",
  25819=>"111111001",
  25820=>"000111111",
  25821=>"111111111",
  25822=>"000000001",
  25823=>"110010000",
  25824=>"001001111",
  25825=>"001001000",
  25826=>"110000111",
  25827=>"111111111",
  25828=>"000101001",
  25829=>"001001000",
  25830=>"100100100",
  25831=>"111111111",
  25832=>"000000100",
  25833=>"000110000",
  25834=>"001001001",
  25835=>"111111000",
  25836=>"000000000",
  25837=>"000111111",
  25838=>"100110111",
  25839=>"010111111",
  25840=>"001000000",
  25841=>"111111111",
  25842=>"000001011",
  25843=>"000000000",
  25844=>"011010110",
  25845=>"101000000",
  25846=>"000000000",
  25847=>"111111111",
  25848=>"000000001",
  25849=>"000000000",
  25850=>"010011011",
  25851=>"011111111",
  25852=>"110110010",
  25853=>"000000000",
  25854=>"000000000",
  25855=>"100001001",
  25856=>"111111111",
  25857=>"111111000",
  25858=>"111111111",
  25859=>"010000000",
  25860=>"101100000",
  25861=>"111011000",
  25862=>"111001001",
  25863=>"111000000",
  25864=>"000001111",
  25865=>"000000000",
  25866=>"000000111",
  25867=>"000000000",
  25868=>"001000011",
  25869=>"100000000",
  25870=>"111111111",
  25871=>"111110000",
  25872=>"000111111",
  25873=>"010101111",
  25874=>"111101111",
  25875=>"100111111",
  25876=>"000011111",
  25877=>"000000000",
  25878=>"100000000",
  25879=>"000000000",
  25880=>"000000000",
  25881=>"010111111",
  25882=>"000000000",
  25883=>"110110111",
  25884=>"000111101",
  25885=>"110111111",
  25886=>"000000000",
  25887=>"010010111",
  25888=>"011011011",
  25889=>"100110110",
  25890=>"011011001",
  25891=>"001001111",
  25892=>"001111111",
  25893=>"010111111",
  25894=>"000000100",
  25895=>"100111111",
  25896=>"000000100",
  25897=>"011111111",
  25898=>"110111000",
  25899=>"000000000",
  25900=>"011010000",
  25901=>"001001011",
  25902=>"000000000",
  25903=>"110111111",
  25904=>"000000000",
  25905=>"000000000",
  25906=>"111111111",
  25907=>"010010000",
  25908=>"111111000",
  25909=>"000011000",
  25910=>"001111111",
  25911=>"000101111",
  25912=>"000000010",
  25913=>"111111111",
  25914=>"000000000",
  25915=>"111100000",
  25916=>"001011011",
  25917=>"111111111",
  25918=>"000011110",
  25919=>"000101111",
  25920=>"000000000",
  25921=>"000001101",
  25922=>"000000000",
  25923=>"111000000",
  25924=>"110111010",
  25925=>"001011111",
  25926=>"000000100",
  25927=>"110110010",
  25928=>"000000101",
  25929=>"110110000",
  25930=>"111111101",
  25931=>"000000000",
  25932=>"111111111",
  25933=>"111000100",
  25934=>"000000001",
  25935=>"000000001",
  25936=>"001001111",
  25937=>"000001001",
  25938=>"000000111",
  25939=>"110010110",
  25940=>"000111000",
  25941=>"001011011",
  25942=>"110110000",
  25943=>"111111111",
  25944=>"111111000",
  25945=>"001001000",
  25946=>"111111000",
  25947=>"011111111",
  25948=>"000000000",
  25949=>"000000100",
  25950=>"011111111",
  25951=>"111011000",
  25952=>"000000000",
  25953=>"100111111",
  25954=>"111000000",
  25955=>"111101111",
  25956=>"110110010",
  25957=>"000000000",
  25958=>"111000000",
  25959=>"001111111",
  25960=>"100100100",
  25961=>"111111010",
  25962=>"000000000",
  25963=>"111000001",
  25964=>"010011000",
  25965=>"110111111",
  25966=>"000000000",
  25967=>"000000000",
  25968=>"110011011",
  25969=>"011011000",
  25970=>"110000000",
  25971=>"011011011",
  25972=>"011011000",
  25973=>"111001000",
  25974=>"000001000",
  25975=>"111001000",
  25976=>"000000000",
  25977=>"111111010",
  25978=>"111000000",
  25979=>"000111111",
  25980=>"110010010",
  25981=>"000000001",
  25982=>"111110111",
  25983=>"010011011",
  25984=>"110111111",
  25985=>"000000001",
  25986=>"000101111",
  25987=>"111000000",
  25988=>"111111000",
  25989=>"011111111",
  25990=>"111111000",
  25991=>"000110111",
  25992=>"001000000",
  25993=>"000000000",
  25994=>"011000000",
  25995=>"111011000",
  25996=>"111011111",
  25997=>"011010000",
  25998=>"111111011",
  25999=>"111111111",
  26000=>"000000000",
  26001=>"111111110",
  26002=>"111111001",
  26003=>"100100110",
  26004=>"000000110",
  26005=>"000000000",
  26006=>"000000000",
  26007=>"000000000",
  26008=>"111000000",
  26009=>"110110111",
  26010=>"111111011",
  26011=>"101000001",
  26012=>"110111111",
  26013=>"000000000",
  26014=>"101000000",
  26015=>"111110000",
  26016=>"111000110",
  26017=>"001100100",
  26018=>"110100101",
  26019=>"111111001",
  26020=>"100000001",
  26021=>"000000011",
  26022=>"101111001",
  26023=>"110110100",
  26024=>"000000001",
  26025=>"000000100",
  26026=>"111111111",
  26027=>"000000000",
  26028=>"000000001",
  26029=>"111000000",
  26030=>"111111001",
  26031=>"000000001",
  26032=>"110111111",
  26033=>"110110000",
  26034=>"111100000",
  26035=>"111100000",
  26036=>"110111011",
  26037=>"111000110",
  26038=>"011001100",
  26039=>"111111111",
  26040=>"000000010",
  26041=>"010011001",
  26042=>"111111111",
  26043=>"001001111",
  26044=>"010100000",
  26045=>"111111111",
  26046=>"111111111",
  26047=>"100010000",
  26048=>"001001011",
  26049=>"100100110",
  26050=>"000000000",
  26051=>"110111111",
  26052=>"111111011",
  26053=>"110010000",
  26054=>"110111000",
  26055=>"000000111",
  26056=>"000000000",
  26057=>"000000011",
  26058=>"101001000",
  26059=>"111000000",
  26060=>"000000000",
  26061=>"110100111",
  26062=>"111110100",
  26063=>"111111101",
  26064=>"000000000",
  26065=>"011111111",
  26066=>"100110111",
  26067=>"000000000",
  26068=>"111111001",
  26069=>"011111111",
  26070=>"000000111",
  26071=>"000010000",
  26072=>"001111000",
  26073=>"111111000",
  26074=>"000000111",
  26075=>"100000000",
  26076=>"001011001",
  26077=>"111001000",
  26078=>"000000100",
  26079=>"111111000",
  26080=>"000000001",
  26081=>"110000000",
  26082=>"000000111",
  26083=>"000001001",
  26084=>"000000000",
  26085=>"000000000",
  26086=>"100000000",
  26087=>"000000000",
  26088=>"100011001",
  26089=>"111111111",
  26090=>"010010011",
  26091=>"101101101",
  26092=>"101001101",
  26093=>"000000000",
  26094=>"000100100",
  26095=>"000000000",
  26096=>"110111000",
  26097=>"111111111",
  26098=>"001001101",
  26099=>"000000000",
  26100=>"011010000",
  26101=>"110000010",
  26102=>"000000000",
  26103=>"100000000",
  26104=>"000111111",
  26105=>"011001001",
  26106=>"111001000",
  26107=>"111001001",
  26108=>"000000000",
  26109=>"111111111",
  26110=>"111111000",
  26111=>"000000010",
  26112=>"111111111",
  26113=>"000000000",
  26114=>"001001101",
  26115=>"111111111",
  26116=>"111111111",
  26117=>"000011011",
  26118=>"111111111",
  26119=>"000000000",
  26120=>"000000011",
  26121=>"000111111",
  26122=>"111111111",
  26123=>"101001000",
  26124=>"111110110",
  26125=>"101000111",
  26126=>"100111111",
  26127=>"110000000",
  26128=>"001111000",
  26129=>"011110110",
  26130=>"001101111",
  26131=>"000000000",
  26132=>"000000000",
  26133=>"110000000",
  26134=>"111111110",
  26135=>"111001000",
  26136=>"110001111",
  26137=>"111111111",
  26138=>"001111111",
  26139=>"110101101",
  26140=>"111111111",
  26141=>"111111011",
  26142=>"110111111",
  26143=>"111110000",
  26144=>"001001000",
  26145=>"111111111",
  26146=>"111110110",
  26147=>"111001001",
  26148=>"000000000",
  26149=>"000000000",
  26150=>"111001001",
  26151=>"000011001",
  26152=>"001111111",
  26153=>"000000000",
  26154=>"001000011",
  26155=>"111000000",
  26156=>"000111111",
  26157=>"000010000",
  26158=>"111100100",
  26159=>"000000100",
  26160=>"111111111",
  26161=>"111111111",
  26162=>"000000100",
  26163=>"110111111",
  26164=>"111111100",
  26165=>"111111111",
  26166=>"111101101",
  26167=>"000000001",
  26168=>"000000111",
  26169=>"000001001",
  26170=>"111110111",
  26171=>"111111001",
  26172=>"000100111",
  26173=>"101100111",
  26174=>"001000000",
  26175=>"111111111",
  26176=>"111111111",
  26177=>"110100111",
  26178=>"000000111",
  26179=>"000011111",
  26180=>"111011111",
  26181=>"000010110",
  26182=>"000000101",
  26183=>"000000000",
  26184=>"111111100",
  26185=>"000000111",
  26186=>"000000000",
  26187=>"111111000",
  26188=>"001000011",
  26189=>"100100111",
  26190=>"111111111",
  26191=>"111101111",
  26192=>"011111111",
  26193=>"001000100",
  26194=>"000111111",
  26195=>"000000100",
  26196=>"000001001",
  26197=>"101111110",
  26198=>"000000001",
  26199=>"000101111",
  26200=>"111110000",
  26201=>"000000001",
  26202=>"110111000",
  26203=>"010111111",
  26204=>"110111111",
  26205=>"000000001",
  26206=>"000000000",
  26207=>"111011000",
  26208=>"011000010",
  26209=>"111111111",
  26210=>"000101111",
  26211=>"110111111",
  26212=>"000110110",
  26213=>"111111111",
  26214=>"000000000",
  26215=>"000000000",
  26216=>"111011011",
  26217=>"000000000",
  26218=>"100100001",
  26219=>"100100000",
  26220=>"000000000",
  26221=>"000000000",
  26222=>"000000000",
  26223=>"101111111",
  26224=>"000111100",
  26225=>"110110011",
  26226=>"011011111",
  26227=>"011111111",
  26228=>"000100000",
  26229=>"000100111",
  26230=>"000000110",
  26231=>"000000000",
  26232=>"000000001",
  26233=>"001000000",
  26234=>"100000000",
  26235=>"111111111",
  26236=>"000000100",
  26237=>"000000000",
  26238=>"100101111",
  26239=>"111011010",
  26240=>"100000001",
  26241=>"000010000",
  26242=>"110010010",
  26243=>"000111111",
  26244=>"100100001",
  26245=>"011111111",
  26246=>"000001101",
  26247=>"011000111",
  26248=>"111100101",
  26249=>"001000100",
  26250=>"000111111",
  26251=>"111111111",
  26252=>"000000000",
  26253=>"111111001",
  26254=>"111001000",
  26255=>"111111110",
  26256=>"000000000",
  26257=>"110110111",
  26258=>"001011100",
  26259=>"000110111",
  26260=>"000000000",
  26261=>"000000000",
  26262=>"000000000",
  26263=>"111111100",
  26264=>"000000000",
  26265=>"000000111",
  26266=>"111111111",
  26267=>"001000001",
  26268=>"000000000",
  26269=>"111001100",
  26270=>"000000000",
  26271=>"111111111",
  26272=>"110111000",
  26273=>"111000111",
  26274=>"010011111",
  26275=>"001001001",
  26276=>"111001000",
  26277=>"100100100",
  26278=>"000000111",
  26279=>"011011111",
  26280=>"000011000",
  26281=>"000000000",
  26282=>"000000000",
  26283=>"000000000",
  26284=>"000000000",
  26285=>"100100100",
  26286=>"111111111",
  26287=>"111110000",
  26288=>"000110110",
  26289=>"111111101",
  26290=>"111111111",
  26291=>"110000111",
  26292=>"000101111",
  26293=>"000000100",
  26294=>"000000000",
  26295=>"111110010",
  26296=>"000000000",
  26297=>"111111000",
  26298=>"000000000",
  26299=>"111111000",
  26300=>"001001001",
  26301=>"000000110",
  26302=>"100111100",
  26303=>"010000000",
  26304=>"111111111",
  26305=>"000001111",
  26306=>"111111111",
  26307=>"000000000",
  26308=>"000000000",
  26309=>"001000000",
  26310=>"111101111",
  26311=>"001001001",
  26312=>"000000000",
  26313=>"001001001",
  26314=>"111111111",
  26315=>"011000000",
  26316=>"000000111",
  26317=>"111000000",
  26318=>"000000111",
  26319=>"000000000",
  26320=>"111111111",
  26321=>"111111111",
  26322=>"000000100",
  26323=>"000000000",
  26324=>"111000000",
  26325=>"001110100",
  26326=>"000000000",
  26327=>"001111111",
  26328=>"111110000",
  26329=>"000000111",
  26330=>"111111111",
  26331=>"011111001",
  26332=>"000000100",
  26333=>"101001000",
  26334=>"000000100",
  26335=>"000000001",
  26336=>"111111111",
  26337=>"000001001",
  26338=>"011111111",
  26339=>"000000000",
  26340=>"111001001",
  26341=>"011011101",
  26342=>"110111011",
  26343=>"000000001",
  26344=>"111111111",
  26345=>"000000100",
  26346=>"110001111",
  26347=>"000000000",
  26348=>"000001001",
  26349=>"110000000",
  26350=>"000000000",
  26351=>"000000000",
  26352=>"011000000",
  26353=>"111111111",
  26354=>"110110010",
  26355=>"001000101",
  26356=>"111111111",
  26357=>"111110000",
  26358=>"011011011",
  26359=>"111111111",
  26360=>"111111111",
  26361=>"000000000",
  26362=>"000001000",
  26363=>"111111010",
  26364=>"100100101",
  26365=>"011011111",
  26366=>"000000000",
  26367=>"100100111",
  26368=>"001000000",
  26369=>"000000000",
  26370=>"110010011",
  26371=>"000000100",
  26372=>"000000000",
  26373=>"000100111",
  26374=>"001000000",
  26375=>"000001111",
  26376=>"100111111",
  26377=>"111001000",
  26378=>"100001001",
  26379=>"000000000",
  26380=>"101000000",
  26381=>"001100000",
  26382=>"011111111",
  26383=>"000111111",
  26384=>"011001011",
  26385=>"111111110",
  26386=>"111100001",
  26387=>"000000000",
  26388=>"101000101",
  26389=>"110111111",
  26390=>"100110110",
  26391=>"000000000",
  26392=>"111000000",
  26393=>"000000000",
  26394=>"000001000",
  26395=>"000000001",
  26396=>"000000100",
  26397=>"011010000",
  26398=>"000000000",
  26399=>"011010000",
  26400=>"000111111",
  26401=>"111111111",
  26402=>"000000000",
  26403=>"000000000",
  26404=>"000011111",
  26405=>"111000000",
  26406=>"000000101",
  26407=>"110000110",
  26408=>"111111111",
  26409=>"000000000",
  26410=>"011110110",
  26411=>"001011000",
  26412=>"000000001",
  26413=>"111011001",
  26414=>"000100111",
  26415=>"111100111",
  26416=>"111011011",
  26417=>"111111001",
  26418=>"000000111",
  26419=>"000000011",
  26420=>"010111011",
  26421=>"000000000",
  26422=>"000000000",
  26423=>"000000100",
  26424=>"000000000",
  26425=>"000000111",
  26426=>"000000000",
  26427=>"000011010",
  26428=>"001101100",
  26429=>"000000000",
  26430=>"111011000",
  26431=>"111100101",
  26432=>"000000100",
  26433=>"000101001",
  26434=>"000100111",
  26435=>"000000000",
  26436=>"111111111",
  26437=>"000000111",
  26438=>"001011001",
  26439=>"000001111",
  26440=>"000000000",
  26441=>"011001111",
  26442=>"110010111",
  26443=>"100000000",
  26444=>"001000101",
  26445=>"000110010",
  26446=>"000000001",
  26447=>"011010011",
  26448=>"001001111",
  26449=>"110111111",
  26450=>"000000000",
  26451=>"000000000",
  26452=>"000000000",
  26453=>"011011000",
  26454=>"000111111",
  26455=>"011001011",
  26456=>"000000000",
  26457=>"000000101",
  26458=>"000000000",
  26459=>"111111000",
  26460=>"111111100",
  26461=>"111111111",
  26462=>"010000000",
  26463=>"111111111",
  26464=>"111111111",
  26465=>"111001100",
  26466=>"000100100",
  26467=>"101111111",
  26468=>"001101111",
  26469=>"001000000",
  26470=>"111111111",
  26471=>"011111111",
  26472=>"001000000",
  26473=>"110110000",
  26474=>"000011011",
  26475=>"000100100",
  26476=>"110011001",
  26477=>"011000000",
  26478=>"110010010",
  26479=>"011000010",
  26480=>"000000111",
  26481=>"100110110",
  26482=>"001000000",
  26483=>"110110111",
  26484=>"000110000",
  26485=>"001100111",
  26486=>"011111001",
  26487=>"000000011",
  26488=>"000011111",
  26489=>"000000110",
  26490=>"111111000",
  26491=>"000000000",
  26492=>"111110001",
  26493=>"111111111",
  26494=>"000010001",
  26495=>"111000000",
  26496=>"011001001",
  26497=>"111111111",
  26498=>"111111101",
  26499=>"000000010",
  26500=>"111111111",
  26501=>"111111001",
  26502=>"110111100",
  26503=>"011011000",
  26504=>"100101111",
  26505=>"100011111",
  26506=>"111011001",
  26507=>"111111011",
  26508=>"111111111",
  26509=>"101111111",
  26510=>"101101101",
  26511=>"111111111",
  26512=>"000000000",
  26513=>"100111111",
  26514=>"011000100",
  26515=>"000000111",
  26516=>"110000000",
  26517=>"010010000",
  26518=>"000000000",
  26519=>"100110111",
  26520=>"101000000",
  26521=>"011011111",
  26522=>"111111111",
  26523=>"111111100",
  26524=>"001101101",
  26525=>"011111111",
  26526=>"000101001",
  26527=>"111111111",
  26528=>"110111111",
  26529=>"011110100",
  26530=>"111100001",
  26531=>"000000000",
  26532=>"111111111",
  26533=>"011111111",
  26534=>"111001101",
  26535=>"000000111",
  26536=>"110010111",
  26537=>"000001011",
  26538=>"000000010",
  26539=>"000000101",
  26540=>"000000001",
  26541=>"011011000",
  26542=>"000111000",
  26543=>"000000100",
  26544=>"110100100",
  26545=>"111011011",
  26546=>"000000111",
  26547=>"000111000",
  26548=>"001000100",
  26549=>"000000000",
  26550=>"000000101",
  26551=>"011000100",
  26552=>"000100000",
  26553=>"111111000",
  26554=>"000000000",
  26555=>"101001001",
  26556=>"111000111",
  26557=>"111011111",
  26558=>"010000100",
  26559=>"111110110",
  26560=>"000000101",
  26561=>"001101111",
  26562=>"001000111",
  26563=>"000000000",
  26564=>"000111111",
  26565=>"011011111",
  26566=>"000000101",
  26567=>"011111111",
  26568=>"101000000",
  26569=>"111111111",
  26570=>"000001101",
  26571=>"111101011",
  26572=>"110100000",
  26573=>"011111111",
  26574=>"011111111",
  26575=>"111110010",
  26576=>"000100110",
  26577=>"111111111",
  26578=>"100000000",
  26579=>"000000000",
  26580=>"111111110",
  26581=>"111111111",
  26582=>"111111001",
  26583=>"111110100",
  26584=>"110111111",
  26585=>"111100001",
  26586=>"000111111",
  26587=>"001001000",
  26588=>"001111111",
  26589=>"000000000",
  26590=>"000000111",
  26591=>"111111001",
  26592=>"001111111",
  26593=>"000000000",
  26594=>"010000000",
  26595=>"000100101",
  26596=>"111111111",
  26597=>"100000000",
  26598=>"111100101",
  26599=>"000000000",
  26600=>"000001001",
  26601=>"000000000",
  26602=>"000010010",
  26603=>"111101111",
  26604=>"100100111",
  26605=>"001100100",
  26606=>"000101101",
  26607=>"111001000",
  26608=>"000100100",
  26609=>"000000100",
  26610=>"111111111",
  26611=>"000000000",
  26612=>"000000111",
  26613=>"111111111",
  26614=>"000000000",
  26615=>"011111100",
  26616=>"000000000",
  26617=>"111101111",
  26618=>"000000111",
  26619=>"101000000",
  26620=>"001011111",
  26621=>"110111111",
  26622=>"000001101",
  26623=>"000000100",
  26624=>"000010111",
  26625=>"011000000",
  26626=>"101111111",
  26627=>"111111000",
  26628=>"001001101",
  26629=>"000001111",
  26630=>"000000100",
  26631=>"000000100",
  26632=>"000000000",
  26633=>"000111111",
  26634=>"100101100",
  26635=>"010010110",
  26636=>"001000110",
  26637=>"001011000",
  26638=>"010000111",
  26639=>"000000000",
  26640=>"111000000",
  26641=>"111111011",
  26642=>"110111111",
  26643=>"101111111",
  26644=>"000000111",
  26645=>"111000000",
  26646=>"111110000",
  26647=>"111111111",
  26648=>"111111011",
  26649=>"111111000",
  26650=>"111111111",
  26651=>"111111000",
  26652=>"000111111",
  26653=>"000111111",
  26654=>"000000010",
  26655=>"000000000",
  26656=>"000000110",
  26657=>"110111111",
  26658=>"111110111",
  26659=>"111011000",
  26660=>"010010000",
  26661=>"011011000",
  26662=>"101001000",
  26663=>"000000000",
  26664=>"000000110",
  26665=>"000110000",
  26666=>"111111111",
  26667=>"100111111",
  26668=>"000000000",
  26669=>"111100011",
  26670=>"101100001",
  26671=>"111110010",
  26672=>"000010111",
  26673=>"000000111",
  26674=>"110011001",
  26675=>"100011111",
  26676=>"100111111",
  26677=>"011001001",
  26678=>"110000011",
  26679=>"111110111",
  26680=>"000000000",
  26681=>"000001111",
  26682=>"000000001",
  26683=>"111000000",
  26684=>"000000000",
  26685=>"100000111",
  26686=>"111111111",
  26687=>"000000000",
  26688=>"000000100",
  26689=>"100001111",
  26690=>"101111111",
  26691=>"000100111",
  26692=>"110110111",
  26693=>"000000000",
  26694=>"000000000",
  26695=>"111100111",
  26696=>"110111111",
  26697=>"000000101",
  26698=>"000011000",
  26699=>"110000100",
  26700=>"000111111",
  26701=>"011000111",
  26702=>"000000111",
  26703=>"101000111",
  26704=>"101001001",
  26705=>"111001001",
  26706=>"000100000",
  26707=>"000110111",
  26708=>"000000000",
  26709=>"000000000",
  26710=>"000111111",
  26711=>"000000000",
  26712=>"000000111",
  26713=>"000000110",
  26714=>"001101111",
  26715=>"011001001",
  26716=>"000000000",
  26717=>"000110111",
  26718=>"111111111",
  26719=>"110111110",
  26720=>"111111000",
  26721=>"000000111",
  26722=>"111001001",
  26723=>"000111011",
  26724=>"000000100",
  26725=>"111000000",
  26726=>"111100111",
  26727=>"010111100",
  26728=>"111100000",
  26729=>"111100100",
  26730=>"000001011",
  26731=>"110110110",
  26732=>"111011011",
  26733=>"100000000",
  26734=>"111111111",
  26735=>"000110111",
  26736=>"000000000",
  26737=>"011100111",
  26738=>"000111111",
  26739=>"111011111",
  26740=>"011001000",
  26741=>"001011111",
  26742=>"111111000",
  26743=>"000000111",
  26744=>"000000111",
  26745=>"000000000",
  26746=>"101100100",
  26747=>"000000001",
  26748=>"010011111",
  26749=>"110111111",
  26750=>"111110111",
  26751=>"000100000",
  26752=>"000001000",
  26753=>"000000000",
  26754=>"111111110",
  26755=>"000000110",
  26756=>"000000000",
  26757=>"000100111",
  26758=>"001000000",
  26759=>"111111111",
  26760=>"000000000",
  26761=>"000000000",
  26762=>"111111111",
  26763=>"111111110",
  26764=>"000100100",
  26765=>"111110111",
  26766=>"011000101",
  26767=>"001000010",
  26768=>"000000111",
  26769=>"000001001",
  26770=>"000000000",
  26771=>"101001000",
  26772=>"000000000",
  26773=>"111111101",
  26774=>"000000000",
  26775=>"111000000",
  26776=>"000101111",
  26777=>"000000111",
  26778=>"001001001",
  26779=>"010110010",
  26780=>"111000000",
  26781=>"000000000",
  26782=>"011010111",
  26783=>"000000000",
  26784=>"000010100",
  26785=>"101000000",
  26786=>"111111000",
  26787=>"111111111",
  26788=>"111011001",
  26789=>"111110000",
  26790=>"111111111",
  26791=>"001111100",
  26792=>"000000101",
  26793=>"000010110",
  26794=>"000000111",
  26795=>"010000100",
  26796=>"000111111",
  26797=>"000110111",
  26798=>"110111111",
  26799=>"111100000",
  26800=>"000000101",
  26801=>"100100101",
  26802=>"111111100",
  26803=>"000000111",
  26804=>"000000000",
  26805=>"000100111",
  26806=>"000000111",
  26807=>"111111111",
  26808=>"111001001",
  26809=>"000101111",
  26810=>"111100001",
  26811=>"101100101",
  26812=>"111001000",
  26813=>"011011111",
  26814=>"101100000",
  26815=>"010011000",
  26816=>"000000000",
  26817=>"000000111",
  26818=>"000000000",
  26819=>"010111111",
  26820=>"000000000",
  26821=>"000000000",
  26822=>"000100110",
  26823=>"011111101",
  26824=>"000111100",
  26825=>"000000101",
  26826=>"100001111",
  26827=>"111111110",
  26828=>"000000000",
  26829=>"011111111",
  26830=>"111100111",
  26831=>"000100110",
  26832=>"100000011",
  26833=>"111101100",
  26834=>"000000000",
  26835=>"000000111",
  26836=>"011011011",
  26837=>"101001011",
  26838=>"111111000",
  26839=>"010000001",
  26840=>"111111000",
  26841=>"000000010",
  26842=>"000000011",
  26843=>"000011000",
  26844=>"111000001",
  26845=>"000100111",
  26846=>"111111110",
  26847=>"000000000",
  26848=>"000000000",
  26849=>"000000100",
  26850=>"000100100",
  26851=>"111111111",
  26852=>"111111000",
  26853=>"110110110",
  26854=>"111100000",
  26855=>"111111000",
  26856=>"010000000",
  26857=>"011001101",
  26858=>"111111101",
  26859=>"110100100",
  26860=>"111101001",
  26861=>"000000000",
  26862=>"010000000",
  26863=>"000000000",
  26864=>"000110111",
  26865=>"000110000",
  26866=>"110100000",
  26867=>"001011000",
  26868=>"111111111",
  26869=>"001001001",
  26870=>"011011000",
  26871=>"111111111",
  26872=>"000000101",
  26873=>"000000101",
  26874=>"000100111",
  26875=>"000110111",
  26876=>"111101011",
  26877=>"001001001",
  26878=>"000011111",
  26879=>"111111111",
  26880=>"111010010",
  26881=>"011111111",
  26882=>"100100111",
  26883=>"010000000",
  26884=>"111001000",
  26885=>"000000011",
  26886=>"111111111",
  26887=>"000000111",
  26888=>"111111111",
  26889=>"000000000",
  26890=>"000000011",
  26891=>"111111000",
  26892=>"001001111",
  26893=>"001111111",
  26894=>"111111111",
  26895=>"001000000",
  26896=>"000000100",
  26897=>"111111110",
  26898=>"111001011",
  26899=>"000000000",
  26900=>"000001011",
  26901=>"000000001",
  26902=>"111011001",
  26903=>"000000000",
  26904=>"100110100",
  26905=>"111011000",
  26906=>"001101111",
  26907=>"000100100",
  26908=>"111111110",
  26909=>"000000011",
  26910=>"111110111",
  26911=>"111000001",
  26912=>"000000011",
  26913=>"100111001",
  26914=>"000000111",
  26915=>"001100101",
  26916=>"011111011",
  26917=>"111000000",
  26918=>"111111001",
  26919=>"000000110",
  26920=>"000001000",
  26921=>"000000000",
  26922=>"111000111",
  26923=>"000000000",
  26924=>"101000000",
  26925=>"000001110",
  26926=>"000000000",
  26927=>"000000101",
  26928=>"110011100",
  26929=>"000111111",
  26930=>"111101111",
  26931=>"000000000",
  26932=>"001111111",
  26933=>"000000000",
  26934=>"111111000",
  26935=>"000000000",
  26936=>"110111000",
  26937=>"111000000",
  26938=>"000011111",
  26939=>"000000000",
  26940=>"111111110",
  26941=>"111101000",
  26942=>"010010011",
  26943=>"000000110",
  26944=>"000000000",
  26945=>"111000000",
  26946=>"000000010",
  26947=>"000000000",
  26948=>"110000100",
  26949=>"000000111",
  26950=>"010000000",
  26951=>"111111111",
  26952=>"111110111",
  26953=>"111110000",
  26954=>"000000101",
  26955=>"001101111",
  26956=>"011000000",
  26957=>"000000000",
  26958=>"100111111",
  26959=>"000001011",
  26960=>"100100110",
  26961=>"000000000",
  26962=>"011001111",
  26963=>"111001001",
  26964=>"111111111",
  26965=>"000000101",
  26966=>"001000000",
  26967=>"111111000",
  26968=>"101101111",
  26969=>"001001101",
  26970=>"000011111",
  26971=>"101111000",
  26972=>"010010111",
  26973=>"000000000",
  26974=>"000000000",
  26975=>"101111111",
  26976=>"000000000",
  26977=>"000010110",
  26978=>"000001111",
  26979=>"000000100",
  26980=>"110110111",
  26981=>"000001000",
  26982=>"010111010",
  26983=>"000000000",
  26984=>"011111111",
  26985=>"000000000",
  26986=>"000000000",
  26987=>"111101000",
  26988=>"000010000",
  26989=>"111100101",
  26990=>"010110111",
  26991=>"000000000",
  26992=>"001001000",
  26993=>"000000000",
  26994=>"101111011",
  26995=>"000000001",
  26996=>"111111111",
  26997=>"000000001",
  26998=>"011111111",
  26999=>"010111111",
  27000=>"000111111",
  27001=>"000010000",
  27002=>"011011000",
  27003=>"001001111",
  27004=>"111111000",
  27005=>"111000000",
  27006=>"000001000",
  27007=>"000000000",
  27008=>"011010000",
  27009=>"000000001",
  27010=>"011111100",
  27011=>"001000000",
  27012=>"111001110",
  27013=>"101000000",
  27014=>"000000000",
  27015=>"000000000",
  27016=>"000001111",
  27017=>"111100100",
  27018=>"000000000",
  27019=>"111111000",
  27020=>"111011111",
  27021=>"111111111",
  27022=>"000000111",
  27023=>"111111001",
  27024=>"011011000",
  27025=>"110000110",
  27026=>"000100110",
  27027=>"111111001",
  27028=>"000000000",
  27029=>"000000000",
  27030=>"001001001",
  27031=>"000001011",
  27032=>"111100000",
  27033=>"011001101",
  27034=>"111111111",
  27035=>"111000000",
  27036=>"111011111",
  27037=>"000110111",
  27038=>"000000100",
  27039=>"000000111",
  27040=>"000000111",
  27041=>"000100111",
  27042=>"101010000",
  27043=>"111111111",
  27044=>"111111011",
  27045=>"100000000",
  27046=>"000101111",
  27047=>"010110000",
  27048=>"000000000",
  27049=>"111111110",
  27050=>"111111111",
  27051=>"000001111",
  27052=>"111000101",
  27053=>"000101000",
  27054=>"000000000",
  27055=>"101111111",
  27056=>"000000000",
  27057=>"010000000",
  27058=>"000111111",
  27059=>"111111010",
  27060=>"101001000",
  27061=>"100100100",
  27062=>"001000110",
  27063=>"111111111",
  27064=>"110000000",
  27065=>"111111111",
  27066=>"111100100",
  27067=>"000000111",
  27068=>"101101111",
  27069=>"111001000",
  27070=>"000100000",
  27071=>"001001011",
  27072=>"110111110",
  27073=>"101101111",
  27074=>"000000000",
  27075=>"111111111",
  27076=>"101101111",
  27077=>"000000000",
  27078=>"010111000",
  27079=>"111111111",
  27080=>"111111111",
  27081=>"000000100",
  27082=>"000000001",
  27083=>"000000110",
  27084=>"111000111",
  27085=>"111111000",
  27086=>"111111011",
  27087=>"011111000",
  27088=>"000000111",
  27089=>"100100111",
  27090=>"111111000",
  27091=>"011001110",
  27092=>"011011111",
  27093=>"101100100",
  27094=>"000101111",
  27095=>"111111011",
  27096=>"000000000",
  27097=>"000111111",
  27098=>"000000000",
  27099=>"000101111",
  27100=>"111111011",
  27101=>"001011000",
  27102=>"111111111",
  27103=>"001001001",
  27104=>"000100111",
  27105=>"000011001",
  27106=>"100000111",
  27107=>"000110110",
  27108=>"111011011",
  27109=>"011111011",
  27110=>"111000100",
  27111=>"000011111",
  27112=>"000010000",
  27113=>"111111010",
  27114=>"000000000",
  27115=>"110111111",
  27116=>"111001111",
  27117=>"000000100",
  27118=>"111111111",
  27119=>"111000000",
  27120=>"000000111",
  27121=>"000000111",
  27122=>"100000100",
  27123=>"000000001",
  27124=>"000111111",
  27125=>"111111111",
  27126=>"000000111",
  27127=>"100000000",
  27128=>"000000111",
  27129=>"011000111",
  27130=>"111000011",
  27131=>"101000000",
  27132=>"000010111",
  27133=>"011001000",
  27134=>"000000001",
  27135=>"000000000",
  27136=>"110000000",
  27137=>"000000001",
  27138=>"000000000",
  27139=>"000000000",
  27140=>"111111111",
  27141=>"111111111",
  27142=>"000000000",
  27143=>"111111111",
  27144=>"101000111",
  27145=>"111111000",
  27146=>"000000000",
  27147=>"000000000",
  27148=>"110111111",
  27149=>"111111111",
  27150=>"010110011",
  27151=>"111111111",
  27152=>"000111011",
  27153=>"011001001",
  27154=>"111111111",
  27155=>"001001001",
  27156=>"000000000",
  27157=>"110111111",
  27158=>"000000011",
  27159=>"101111011",
  27160=>"000000100",
  27161=>"000000000",
  27162=>"111100100",
  27163=>"100000000",
  27164=>"000000000",
  27165=>"000000110",
  27166=>"111111111",
  27167=>"000111110",
  27168=>"111111111",
  27169=>"000000000",
  27170=>"110000000",
  27171=>"111111111",
  27172=>"000000000",
  27173=>"111000111",
  27174=>"011011010",
  27175=>"001010000",
  27176=>"011011010",
  27177=>"000000000",
  27178=>"111111111",
  27179=>"000100010",
  27180=>"111101000",
  27181=>"110110000",
  27182=>"010110100",
  27183=>"000101111",
  27184=>"111111111",
  27185=>"111111110",
  27186=>"111001001",
  27187=>"000011001",
  27188=>"101100100",
  27189=>"001011000",
  27190=>"111110111",
  27191=>"000010000",
  27192=>"000000000",
  27193=>"000000100",
  27194=>"111111111",
  27195=>"110110111",
  27196=>"000000000",
  27197=>"111111000",
  27198=>"110001011",
  27199=>"000000111",
  27200=>"000000000",
  27201=>"000000000",
  27202=>"000000000",
  27203=>"111111010",
  27204=>"100000000",
  27205=>"000000000",
  27206=>"110101001",
  27207=>"000000000",
  27208=>"000001001",
  27209=>"111111111",
  27210=>"111111111",
  27211=>"110110111",
  27212=>"100111111",
  27213=>"111111000",
  27214=>"000000000",
  27215=>"000000000",
  27216=>"000000000",
  27217=>"111111111",
  27218=>"001111001",
  27219=>"000001000",
  27220=>"111111000",
  27221=>"000000001",
  27222=>"111011000",
  27223=>"011001000",
  27224=>"000000000",
  27225=>"000000000",
  27226=>"000000000",
  27227=>"111011001",
  27228=>"000000000",
  27229=>"111111111",
  27230=>"000000000",
  27231=>"000011001",
  27232=>"111111111",
  27233=>"100111111",
  27234=>"000000000",
  27235=>"000000101",
  27236=>"111010000",
  27237=>"011000000",
  27238=>"000100110",
  27239=>"100011011",
  27240=>"111111101",
  27241=>"000000100",
  27242=>"000000111",
  27243=>"111111110",
  27244=>"111110010",
  27245=>"111000111",
  27246=>"111111111",
  27247=>"111111111",
  27248=>"001111111",
  27249=>"001000000",
  27250=>"101110110",
  27251=>"111111111",
  27252=>"110000000",
  27253=>"111011000",
  27254=>"000000111",
  27255=>"111111111",
  27256=>"000000111",
  27257=>"000000100",
  27258=>"111000000",
  27259=>"111111111",
  27260=>"000010010",
  27261=>"111111001",
  27262=>"111111101",
  27263=>"100000000",
  27264=>"000000111",
  27265=>"111111111",
  27266=>"000001111",
  27267=>"001111011",
  27268=>"111001001",
  27269=>"000000100",
  27270=>"110110000",
  27271=>"111111111",
  27272=>"110000000",
  27273=>"111100000",
  27274=>"111111111",
  27275=>"111110000",
  27276=>"000000000",
  27277=>"000010000",
  27278=>"000010111",
  27279=>"111111001",
  27280=>"100000111",
  27281=>"111101000",
  27282=>"000000000",
  27283=>"100000000",
  27284=>"001111111",
  27285=>"000000000",
  27286=>"000111111",
  27287=>"110100111",
  27288=>"001000100",
  27289=>"011111100",
  27290=>"111001111",
  27291=>"100111111",
  27292=>"111100100",
  27293=>"111000101",
  27294=>"000000000",
  27295=>"111111111",
  27296=>"001001000",
  27297=>"000000001",
  27298=>"000000000",
  27299=>"111011001",
  27300=>"100000001",
  27301=>"000000000",
  27302=>"111111001",
  27303=>"110110110",
  27304=>"000110110",
  27305=>"111111111",
  27306=>"111111111",
  27307=>"101111111",
  27308=>"000000000",
  27309=>"000110110",
  27310=>"011001111",
  27311=>"111100000",
  27312=>"111111010",
  27313=>"000000000",
  27314=>"101111111",
  27315=>"111111111",
  27316=>"111111111",
  27317=>"001000000",
  27318=>"011001001",
  27319=>"001001001",
  27320=>"111000100",
  27321=>"000000000",
  27322=>"111110010",
  27323=>"011110110",
  27324=>"001000011",
  27325=>"111111111",
  27326=>"111100100",
  27327=>"111000000",
  27328=>"111110000",
  27329=>"000001000",
  27330=>"111111111",
  27331=>"000110010",
  27332=>"111111111",
  27333=>"000000000",
  27334=>"110111111",
  27335=>"000111000",
  27336=>"011000000",
  27337=>"000101111",
  27338=>"001001001",
  27339=>"111111111",
  27340=>"001011111",
  27341=>"000001000",
  27342=>"011000100",
  27343=>"000000110",
  27344=>"111000011",
  27345=>"100001111",
  27346=>"110111111",
  27347=>"111001111",
  27348=>"000011011",
  27349=>"111111110",
  27350=>"100000000",
  27351=>"111111111",
  27352=>"000001001",
  27353=>"111111111",
  27354=>"100100110",
  27355=>"000011111",
  27356=>"000000000",
  27357=>"010110110",
  27358=>"101111111",
  27359=>"000100100",
  27360=>"000111010",
  27361=>"000000000",
  27362=>"111000000",
  27363=>"111111011",
  27364=>"000011011",
  27365=>"111100110",
  27366=>"000001000",
  27367=>"000000000",
  27368=>"010111111",
  27369=>"101000111",
  27370=>"000000111",
  27371=>"111111111",
  27372=>"111111100",
  27373=>"000000010",
  27374=>"011110111",
  27375=>"110000111",
  27376=>"000000111",
  27377=>"000000111",
  27378=>"000001111",
  27379=>"010111111",
  27380=>"110000000",
  27381=>"000110110",
  27382=>"111111000",
  27383=>"000000101",
  27384=>"111100000",
  27385=>"111111111",
  27386=>"000000000",
  27387=>"000000000",
  27388=>"111101001",
  27389=>"000000001",
  27390=>"000011011",
  27391=>"111000000",
  27392=>"111101101",
  27393=>"011010010",
  27394=>"111000011",
  27395=>"111111111",
  27396=>"000101101",
  27397=>"111101111",
  27398=>"111000111",
  27399=>"000000100",
  27400=>"101000001",
  27401=>"111000000",
  27402=>"011111111",
  27403=>"000000100",
  27404=>"101111111",
  27405=>"110111001",
  27406=>"010010000",
  27407=>"000000000",
  27408=>"000010111",
  27409=>"011111111",
  27410=>"111111111",
  27411=>"111111111",
  27412=>"111111111",
  27413=>"110000011",
  27414=>"011111000",
  27415=>"000000000",
  27416=>"100001000",
  27417=>"000000001",
  27418=>"000000000",
  27419=>"111111001",
  27420=>"110110111",
  27421=>"110110111",
  27422=>"111111111",
  27423=>"011111001",
  27424=>"010010000",
  27425=>"100111111",
  27426=>"000000111",
  27427=>"111111011",
  27428=>"101111111",
  27429=>"111111111",
  27430=>"111100110",
  27431=>"111111011",
  27432=>"011011001",
  27433=>"000001001",
  27434=>"000000000",
  27435=>"100111111",
  27436=>"111111111",
  27437=>"010000000",
  27438=>"111111111",
  27439=>"111111111",
  27440=>"001011111",
  27441=>"011000000",
  27442=>"100001111",
  27443=>"000111111",
  27444=>"110000001",
  27445=>"111111000",
  27446=>"111111111",
  27447=>"100100101",
  27448=>"111111111",
  27449=>"111111111",
  27450=>"011011011",
  27451=>"000000100",
  27452=>"011000000",
  27453=>"000111100",
  27454=>"111011011",
  27455=>"101000111",
  27456=>"101000011",
  27457=>"011111011",
  27458=>"100111111",
  27459=>"000100000",
  27460=>"000000011",
  27461=>"111000000",
  27462=>"011010000",
  27463=>"100010111",
  27464=>"111111111",
  27465=>"000110111",
  27466=>"010111111",
  27467=>"011111111",
  27468=>"011111011",
  27469=>"000011000",
  27470=>"110010111",
  27471=>"111111001",
  27472=>"011011000",
  27473=>"111111111",
  27474=>"111111111",
  27475=>"111111111",
  27476=>"111001101",
  27477=>"011011011",
  27478=>"000000111",
  27479=>"000101111",
  27480=>"000000000",
  27481=>"001101111",
  27482=>"010000111",
  27483=>"110111101",
  27484=>"111111111",
  27485=>"000000000",
  27486=>"000100101",
  27487=>"000000000",
  27488=>"110000000",
  27489=>"000000000",
  27490=>"111111111",
  27491=>"111000110",
  27492=>"110111000",
  27493=>"111001000",
  27494=>"101101101",
  27495=>"000111110",
  27496=>"110111111",
  27497=>"000000000",
  27498=>"111111011",
  27499=>"100110100",
  27500=>"000000000",
  27501=>"111111111",
  27502=>"000000000",
  27503=>"111111111",
  27504=>"011111111",
  27505=>"111111001",
  27506=>"000000101",
  27507=>"011011001",
  27508=>"111011001",
  27509=>"111001101",
  27510=>"011111100",
  27511=>"000011110",
  27512=>"111011000",
  27513=>"000111001",
  27514=>"000000111",
  27515=>"111111000",
  27516=>"101111111",
  27517=>"111111111",
  27518=>"111111000",
  27519=>"111111111",
  27520=>"110111110",
  27521=>"000001011",
  27522=>"010000000",
  27523=>"111111111",
  27524=>"000100110",
  27525=>"000110000",
  27526=>"100100111",
  27527=>"110000100",
  27528=>"110000111",
  27529=>"011011111",
  27530=>"100000000",
  27531=>"000000000",
  27532=>"110110111",
  27533=>"000010000",
  27534=>"000000000",
  27535=>"101000000",
  27536=>"111111111",
  27537=>"111111111",
  27538=>"100101100",
  27539=>"000000000",
  27540=>"000000000",
  27541=>"111111011",
  27542=>"111111110",
  27543=>"010010111",
  27544=>"111111000",
  27545=>"000111111",
  27546=>"000000111",
  27547=>"001011000",
  27548=>"000000000",
  27549=>"000001111",
  27550=>"000000000",
  27551=>"110111000",
  27552=>"001000000",
  27553=>"000000011",
  27554=>"001100000",
  27555=>"100111111",
  27556=>"101100111",
  27557=>"111111111",
  27558=>"000000111",
  27559=>"000100111",
  27560=>"111111110",
  27561=>"000111111",
  27562=>"000100101",
  27563=>"000000000",
  27564=>"111111000",
  27565=>"111100110",
  27566=>"000000100",
  27567=>"111010010",
  27568=>"000000000",
  27569=>"011111010",
  27570=>"111111111",
  27571=>"001000000",
  27572=>"000111111",
  27573=>"100000101",
  27574=>"011111111",
  27575=>"101001001",
  27576=>"111111111",
  27577=>"111111111",
  27578=>"010000100",
  27579=>"110111011",
  27580=>"110111111",
  27581=>"000001011",
  27582=>"111101100",
  27583=>"010010010",
  27584=>"000000111",
  27585=>"111001101",
  27586=>"000000000",
  27587=>"111111111",
  27588=>"111110111",
  27589=>"110000001",
  27590=>"101101111",
  27591=>"000000000",
  27592=>"011101111",
  27593=>"000011000",
  27594=>"111111111",
  27595=>"100100100",
  27596=>"100000000",
  27597=>"000100000",
  27598=>"100001011",
  27599=>"000111111",
  27600=>"000000001",
  27601=>"000100101",
  27602=>"111111111",
  27603=>"000011000",
  27604=>"000000000",
  27605=>"000111111",
  27606=>"000000000",
  27607=>"111101001",
  27608=>"000000011",
  27609=>"000000000",
  27610=>"000000001",
  27611=>"001000000",
  27612=>"110111111",
  27613=>"110111110",
  27614=>"001001111",
  27615=>"110011010",
  27616=>"000000000",
  27617=>"111111000",
  27618=>"000000100",
  27619=>"111111111",
  27620=>"001011111",
  27621=>"111111000",
  27622=>"101100111",
  27623=>"000000000",
  27624=>"010111011",
  27625=>"111111111",
  27626=>"000001011",
  27627=>"001000000",
  27628=>"000000111",
  27629=>"111111110",
  27630=>"000101111",
  27631=>"000000000",
  27632=>"000000000",
  27633=>"111111111",
  27634=>"000000000",
  27635=>"001000100",
  27636=>"100001011",
  27637=>"000000000",
  27638=>"000000000",
  27639=>"000000110",
  27640=>"100100111",
  27641=>"111011011",
  27642=>"111111001",
  27643=>"110111111",
  27644=>"101111111",
  27645=>"011111110",
  27646=>"000000000",
  27647=>"000100111",
  27648=>"001001000",
  27649=>"111111100",
  27650=>"000000111",
  27651=>"000000000",
  27652=>"111001100",
  27653=>"000000000",
  27654=>"000000000",
  27655=>"001000111",
  27656=>"001000011",
  27657=>"000000000",
  27658=>"111110000",
  27659=>"000000100",
  27660=>"111111000",
  27661=>"001000000",
  27662=>"001101000",
  27663=>"000000000",
  27664=>"000000000",
  27665=>"000000101",
  27666=>"111111111",
  27667=>"110111111",
  27668=>"000001111",
  27669=>"111111111",
  27670=>"111101001",
  27671=>"000000000",
  27672=>"000000000",
  27673=>"000000000",
  27674=>"000000000",
  27675=>"000110101",
  27676=>"111110000",
  27677=>"000000110",
  27678=>"011111111",
  27679=>"110000001",
  27680=>"111111111",
  27681=>"111111010",
  27682=>"111111110",
  27683=>"100000000",
  27684=>"000000110",
  27685=>"000000000",
  27686=>"110101000",
  27687=>"111111001",
  27688=>"101000000",
  27689=>"000000000",
  27690=>"000000101",
  27691=>"101000001",
  27692=>"111111000",
  27693=>"111111011",
  27694=>"000000101",
  27695=>"111110000",
  27696=>"111111111",
  27697=>"000000000",
  27698=>"101000100",
  27699=>"000100110",
  27700=>"111110110",
  27701=>"111000000",
  27702=>"111000001",
  27703=>"000000000",
  27704=>"110100000",
  27705=>"000011000",
  27706=>"011111111",
  27707=>"001000111",
  27708=>"101111111",
  27709=>"000100111",
  27710=>"000000000",
  27711=>"000000000",
  27712=>"111001000",
  27713=>"111111111",
  27714=>"111000000",
  27715=>"000110111",
  27716=>"111111111",
  27717=>"111111111",
  27718=>"000000001",
  27719=>"100100100",
  27720=>"100100110",
  27721=>"000111111",
  27722=>"000000101",
  27723=>"000011111",
  27724=>"011011010",
  27725=>"111001011",
  27726=>"000000000",
  27727=>"000000000",
  27728=>"111111111",
  27729=>"000111111",
  27730=>"111111111",
  27731=>"000000000",
  27732=>"000001001",
  27733=>"000111000",
  27734=>"111001011",
  27735=>"111111111",
  27736=>"111111111",
  27737=>"000000111",
  27738=>"111111011",
  27739=>"100000000",
  27740=>"001000001",
  27741=>"111111111",
  27742=>"000010000",
  27743=>"001000000",
  27744=>"111111111",
  27745=>"010000000",
  27746=>"000001001",
  27747=>"111110000",
  27748=>"000000000",
  27749=>"111111111",
  27750=>"000000111",
  27751=>"111111111",
  27752=>"111010010",
  27753=>"111111000",
  27754=>"100000000",
  27755=>"111111000",
  27756=>"000000000",
  27757=>"001000000",
  27758=>"000001111",
  27759=>"000000000",
  27760=>"110110100",
  27761=>"111111111",
  27762=>"010010110",
  27763=>"111111111",
  27764=>"000000000",
  27765=>"101011011",
  27766=>"111010000",
  27767=>"000000111",
  27768=>"011001111",
  27769=>"000000001",
  27770=>"000000000",
  27771=>"000000000",
  27772=>"000111111",
  27773=>"000000000",
  27774=>"000000000",
  27775=>"011111111",
  27776=>"101101111",
  27777=>"000111111",
  27778=>"111100000",
  27779=>"000000000",
  27780=>"000000000",
  27781=>"101000111",
  27782=>"100110110",
  27783=>"111111101",
  27784=>"001000010",
  27785=>"111111111",
  27786=>"111111011",
  27787=>"111111111",
  27788=>"111101111",
  27789=>"111111110",
  27790=>"111111000",
  27791=>"111111111",
  27792=>"000001001",
  27793=>"000000000",
  27794=>"110110000",
  27795=>"000000000",
  27796=>"000000001",
  27797=>"110110111",
  27798=>"111111111",
  27799=>"000000000",
  27800=>"000000100",
  27801=>"011101101",
  27802=>"000000111",
  27803=>"100110110",
  27804=>"000000000",
  27805=>"001100000",
  27806=>"111111101",
  27807=>"000001111",
  27808=>"100110000",
  27809=>"100111111",
  27810=>"111000000",
  27811=>"011010110",
  27812=>"000100111",
  27813=>"110111111",
  27814=>"111111011",
  27815=>"110000000",
  27816=>"000000000",
  27817=>"011000100",
  27818=>"001011111",
  27819=>"000000000",
  27820=>"011001110",
  27821=>"001110110",
  27822=>"111111111",
  27823=>"101100001",
  27824=>"111111000",
  27825=>"000000000",
  27826=>"111111111",
  27827=>"000000000",
  27828=>"000000000",
  27829=>"000000000",
  27830=>"111111111",
  27831=>"111111111",
  27832=>"100001011",
  27833=>"111001000",
  27834=>"101000000",
  27835=>"000000000",
  27836=>"110000000",
  27837=>"100101111",
  27838=>"101111111",
  27839=>"000000000",
  27840=>"100110011",
  27841=>"111011011",
  27842=>"000101001",
  27843=>"000000000",
  27844=>"011011001",
  27845=>"111111001",
  27846=>"000000001",
  27847=>"111111111",
  27848=>"000000001",
  27849=>"000000000",
  27850=>"000000000",
  27851=>"000000000",
  27852=>"000100000",
  27853=>"110110111",
  27854=>"111111000",
  27855=>"000000100",
  27856=>"001011111",
  27857=>"001001011",
  27858=>"100100110",
  27859=>"000000000",
  27860=>"000000111",
  27861=>"111111111",
  27862=>"000000000",
  27863=>"111110100",
  27864=>"111000000",
  27865=>"111111000",
  27866=>"111100000",
  27867=>"111111111",
  27868=>"111111111",
  27869=>"110110110",
  27870=>"000000000",
  27871=>"000000000",
  27872=>"000000111",
  27873=>"111011000",
  27874=>"100000000",
  27875=>"000111000",
  27876=>"000000000",
  27877=>"000000000",
  27878=>"111111111",
  27879=>"111110111",
  27880=>"000111111",
  27881=>"001111100",
  27882=>"000000111",
  27883=>"011000000",
  27884=>"000010000",
  27885=>"111111111",
  27886=>"111111111",
  27887=>"001000000",
  27888=>"111000000",
  27889=>"111100001",
  27890=>"000000000",
  27891=>"000000000",
  27892=>"000000000",
  27893=>"111000100",
  27894=>"100100000",
  27895=>"000010110",
  27896=>"000000100",
  27897=>"001001000",
  27898=>"111111010",
  27899=>"000000000",
  27900=>"111100000",
  27901=>"000100000",
  27902=>"000000000",
  27903=>"111101110",
  27904=>"000000111",
  27905=>"010000000",
  27906=>"000011010",
  27907=>"001000100",
  27908=>"111111111",
  27909=>"000000000",
  27910=>"001111111",
  27911=>"001001001",
  27912=>"000001111",
  27913=>"000100110",
  27914=>"111111111",
  27915=>"111111100",
  27916=>"000000000",
  27917=>"011111111",
  27918=>"111000001",
  27919=>"000000111",
  27920=>"011000111",
  27921=>"101000000",
  27922=>"000000000",
  27923=>"111111000",
  27924=>"000100000",
  27925=>"111011001",
  27926=>"111110100",
  27927=>"011111000",
  27928=>"100110110",
  27929=>"000000000",
  27930=>"110100010",
  27931=>"111000100",
  27932=>"100101111",
  27933=>"000111000",
  27934=>"000000110",
  27935=>"111111100",
  27936=>"101100000",
  27937=>"011111111",
  27938=>"111111000",
  27939=>"000000000",
  27940=>"000000001",
  27941=>"000000000",
  27942=>"011110110",
  27943=>"000101001",
  27944=>"000000000",
  27945=>"110110111",
  27946=>"001111000",
  27947=>"010111000",
  27948=>"000100111",
  27949=>"000000000",
  27950=>"100000111",
  27951=>"000001001",
  27952=>"000001000",
  27953=>"101100000",
  27954=>"000000000",
  27955=>"000000000",
  27956=>"000000010",
  27957=>"100000000",
  27958=>"010010101",
  27959=>"110100001",
  27960=>"000000000",
  27961=>"000000000",
  27962=>"000000000",
  27963=>"011111111",
  27964=>"111111111",
  27965=>"110111110",
  27966=>"100001001",
  27967=>"111111010",
  27968=>"000001000",
  27969=>"001111000",
  27970=>"000000001",
  27971=>"011011111",
  27972=>"111111111",
  27973=>"000110110",
  27974=>"011111000",
  27975=>"111111111",
  27976=>"000000010",
  27977=>"101001111",
  27978=>"101101000",
  27979=>"110100101",
  27980=>"000000000",
  27981=>"111111011",
  27982=>"000000011",
  27983=>"000001111",
  27984=>"111101111",
  27985=>"001111010",
  27986=>"000110111",
  27987=>"111111111",
  27988=>"111001111",
  27989=>"011011111",
  27990=>"000000000",
  27991=>"110000000",
  27992=>"000000000",
  27993=>"000000100",
  27994=>"100111001",
  27995=>"001001111",
  27996=>"111111000",
  27997=>"110111111",
  27998=>"000110110",
  27999=>"111111010",
  28000=>"100111111",
  28001=>"000000000",
  28002=>"100111111",
  28003=>"000000100",
  28004=>"001001001",
  28005=>"100110000",
  28006=>"111100111",
  28007=>"011001001",
  28008=>"011110000",
  28009=>"110010011",
  28010=>"000010010",
  28011=>"000000000",
  28012=>"011001000",
  28013=>"000000000",
  28014=>"111111010",
  28015=>"111111001",
  28016=>"111111111",
  28017=>"001011111",
  28018=>"011011111",
  28019=>"110110000",
  28020=>"000000000",
  28021=>"100100000",
  28022=>"111111111",
  28023=>"000110110",
  28024=>"111111111",
  28025=>"000000000",
  28026=>"111100111",
  28027=>"011000000",
  28028=>"101100000",
  28029=>"001000000",
  28030=>"000011000",
  28031=>"111101000",
  28032=>"111111110",
  28033=>"111111101",
  28034=>"000000011",
  28035=>"000000000",
  28036=>"011100110",
  28037=>"000001000",
  28038=>"111111111",
  28039=>"111100000",
  28040=>"000010110",
  28041=>"000000000",
  28042=>"011011011",
  28043=>"111111111",
  28044=>"111111111",
  28045=>"011001100",
  28046=>"000100111",
  28047=>"111111111",
  28048=>"000000000",
  28049=>"101000000",
  28050=>"101100111",
  28051=>"111111110",
  28052=>"111111111",
  28053=>"111000000",
  28054=>"000011111",
  28055=>"101001000",
  28056=>"001000000",
  28057=>"111111111",
  28058=>"000000111",
  28059=>"001001001",
  28060=>"000110100",
  28061=>"000000000",
  28062=>"000000000",
  28063=>"000010000",
  28064=>"111111111",
  28065=>"000000100",
  28066=>"010110110",
  28067=>"111011011",
  28068=>"000101111",
  28069=>"111011011",
  28070=>"111111111",
  28071=>"000001101",
  28072=>"000000000",
  28073=>"011111111",
  28074=>"111111100",
  28075=>"110111111",
  28076=>"110000000",
  28077=>"111011111",
  28078=>"111111111",
  28079=>"111110100",
  28080=>"100110111",
  28081=>"111111111",
  28082=>"000000000",
  28083=>"000000000",
  28084=>"111111111",
  28085=>"001001001",
  28086=>"000110111",
  28087=>"000100000",
  28088=>"111100110",
  28089=>"011111101",
  28090=>"100100000",
  28091=>"000001111",
  28092=>"000000000",
  28093=>"000000000",
  28094=>"100110000",
  28095=>"000000111",
  28096=>"000010000",
  28097=>"110000000",
  28098=>"000000000",
  28099=>"000100111",
  28100=>"111111111",
  28101=>"001001001",
  28102=>"111111010",
  28103=>"111000010",
  28104=>"110000000",
  28105=>"011000001",
  28106=>"000000000",
  28107=>"000000000",
  28108=>"101000000",
  28109=>"000000000",
  28110=>"100111111",
  28111=>"111011011",
  28112=>"111111111",
  28113=>"000000011",
  28114=>"011010010",
  28115=>"000000000",
  28116=>"011011001",
  28117=>"001001111",
  28118=>"000000000",
  28119=>"010011011",
  28120=>"110100100",
  28121=>"111101111",
  28122=>"000000000",
  28123=>"000000000",
  28124=>"011000000",
  28125=>"111101001",
  28126=>"000000000",
  28127=>"000000001",
  28128=>"111111000",
  28129=>"110000000",
  28130=>"000000000",
  28131=>"001100100",
  28132=>"111110000",
  28133=>"001000000",
  28134=>"101111000",
  28135=>"111011000",
  28136=>"111101101",
  28137=>"010011011",
  28138=>"100110111",
  28139=>"100100111",
  28140=>"000110111",
  28141=>"110110000",
  28142=>"111111111",
  28143=>"111111111",
  28144=>"100000000",
  28145=>"100100100",
  28146=>"000000000",
  28147=>"110111111",
  28148=>"000001000",
  28149=>"111100000",
  28150=>"001001000",
  28151=>"001100100",
  28152=>"000000000",
  28153=>"110111111",
  28154=>"011001001",
  28155=>"000000000",
  28156=>"111111111",
  28157=>"000001111",
  28158=>"111111100",
  28159=>"000000111",
  28160=>"111111111",
  28161=>"110000000",
  28162=>"000000111",
  28163=>"011111110",
  28164=>"001001000",
  28165=>"110010000",
  28166=>"011000001",
  28167=>"000100111",
  28168=>"111111000",
  28169=>"011111000",
  28170=>"001000000",
  28171=>"100111101",
  28172=>"000001001",
  28173=>"111101111",
  28174=>"001011100",
  28175=>"111110100",
  28176=>"110110110",
  28177=>"000000010",
  28178=>"000000000",
  28179=>"000010000",
  28180=>"111011000",
  28181=>"000101111",
  28182=>"111111111",
  28183=>"111111111",
  28184=>"110111111",
  28185=>"001000000",
  28186=>"111110111",
  28187=>"111011001",
  28188=>"000000000",
  28189=>"110011001",
  28190=>"000010000",
  28191=>"111111111",
  28192=>"000000000",
  28193=>"111111111",
  28194=>"111111111",
  28195=>"000000000",
  28196=>"000000000",
  28197=>"000000000",
  28198=>"000000000",
  28199=>"111101111",
  28200=>"001111111",
  28201=>"000000000",
  28202=>"011111111",
  28203=>"001000000",
  28204=>"111111000",
  28205=>"000000111",
  28206=>"111111111",
  28207=>"111010000",
  28208=>"000000000",
  28209=>"000000000",
  28210=>"001001111",
  28211=>"011001111",
  28212=>"000110110",
  28213=>"111111111",
  28214=>"000100111",
  28215=>"111111111",
  28216=>"111110110",
  28217=>"000000101",
  28218=>"100000000",
  28219=>"000000000",
  28220=>"111101000",
  28221=>"111111111",
  28222=>"000001000",
  28223=>"101100110",
  28224=>"111111111",
  28225=>"001001001",
  28226=>"001000000",
  28227=>"111100000",
  28228=>"100101101",
  28229=>"111110000",
  28230=>"000000111",
  28231=>"001111111",
  28232=>"001101101",
  28233=>"111001001",
  28234=>"000000000",
  28235=>"111110110",
  28236=>"111111110",
  28237=>"000000000",
  28238=>"101000000",
  28239=>"011000000",
  28240=>"000000100",
  28241=>"101101111",
  28242=>"001010000",
  28243=>"001000001",
  28244=>"000000000",
  28245=>"101100000",
  28246=>"101100110",
  28247=>"111100000",
  28248=>"100000000",
  28249=>"111000000",
  28250=>"101000000",
  28251=>"100000000",
  28252=>"000000111",
  28253=>"100000110",
  28254=>"111111111",
  28255=>"001000000",
  28256=>"000000000",
  28257=>"111001010",
  28258=>"000111111",
  28259=>"011011011",
  28260=>"000111111",
  28261=>"000011011",
  28262=>"001001000",
  28263=>"000000010",
  28264=>"000000000",
  28265=>"110110111",
  28266=>"100000111",
  28267=>"110000000",
  28268=>"110001001",
  28269=>"000000000",
  28270=>"111000000",
  28271=>"111110110",
  28272=>"000010110",
  28273=>"110110000",
  28274=>"000100100",
  28275=>"011000000",
  28276=>"000001000",
  28277=>"000110111",
  28278=>"000000000",
  28279=>"000000000",
  28280=>"000011011",
  28281=>"001111111",
  28282=>"000000101",
  28283=>"111000001",
  28284=>"111111111",
  28285=>"100100110",
  28286=>"000010000",
  28287=>"111111010",
  28288=>"000111111",
  28289=>"111000000",
  28290=>"111110010",
  28291=>"001011011",
  28292=>"000000000",
  28293=>"000000000",
  28294=>"100100001",
  28295=>"000000110",
  28296=>"000000000",
  28297=>"111111000",
  28298=>"000010111",
  28299=>"100111111",
  28300=>"111111110",
  28301=>"101111111",
  28302=>"110111000",
  28303=>"001001000",
  28304=>"111111011",
  28305=>"111110000",
  28306=>"111011000",
  28307=>"011001000",
  28308=>"000100111",
  28309=>"000000000",
  28310=>"111000000",
  28311=>"111111111",
  28312=>"000000000",
  28313=>"011111111",
  28314=>"001011111",
  28315=>"000111111",
  28316=>"111101101",
  28317=>"000000000",
  28318=>"111111000",
  28319=>"111111100",
  28320=>"110110111",
  28321=>"000000000",
  28322=>"000000000",
  28323=>"000100000",
  28324=>"000000111",
  28325=>"000000000",
  28326=>"010000111",
  28327=>"110111111",
  28328=>"101100001",
  28329=>"000000000",
  28330=>"000000000",
  28331=>"000000000",
  28332=>"000000000",
  28333=>"111111101",
  28334=>"100111111",
  28335=>"110110111",
  28336=>"000000000",
  28337=>"000000000",
  28338=>"111110111",
  28339=>"000000001",
  28340=>"000000000",
  28341=>"100110001",
  28342=>"000000000",
  28343=>"000000000",
  28344=>"101100100",
  28345=>"111111111",
  28346=>"000000000",
  28347=>"100000000",
  28348=>"000000000",
  28349=>"111101111",
  28350=>"000000000",
  28351=>"000111111",
  28352=>"111111111",
  28353=>"111111001",
  28354=>"100100111",
  28355=>"110110111",
  28356=>"000000000",
  28357=>"000111111",
  28358=>"001111111",
  28359=>"111110100",
  28360=>"000000000",
  28361=>"111100000",
  28362=>"001100101",
  28363=>"111111100",
  28364=>"100100101",
  28365=>"010101000",
  28366=>"000111111",
  28367=>"011000000",
  28368=>"000000000",
  28369=>"000000000",
  28370=>"001011001",
  28371=>"000000000",
  28372=>"100101111",
  28373=>"001111000",
  28374=>"101100000",
  28375=>"000000111",
  28376=>"000100101",
  28377=>"000110110",
  28378=>"101101111",
  28379=>"000111111",
  28380=>"100000100",
  28381=>"000000000",
  28382=>"000110000",
  28383=>"110110100",
  28384=>"111111111",
  28385=>"111111111",
  28386=>"000001111",
  28387=>"111111011",
  28388=>"001001111",
  28389=>"000001000",
  28390=>"111111111",
  28391=>"001000000",
  28392=>"111000000",
  28393=>"000010111",
  28394=>"111111111",
  28395=>"111111110",
  28396=>"000000000",
  28397=>"111111000",
  28398=>"010001000",
  28399=>"001000000",
  28400=>"100000111",
  28401=>"000000000",
  28402=>"111001101",
  28403=>"000000111",
  28404=>"111111111",
  28405=>"000110000",
  28406=>"111111000",
  28407=>"000000100",
  28408=>"001111111",
  28409=>"100100000",
  28410=>"111111111",
  28411=>"000000000",
  28412=>"000001001",
  28413=>"111111001",
  28414=>"111111111",
  28415=>"000000011",
  28416=>"100101001",
  28417=>"100100100",
  28418=>"000000111",
  28419=>"000010000",
  28420=>"000100111",
  28421=>"000110100",
  28422=>"110110000",
  28423=>"110110111",
  28424=>"000000111",
  28425=>"000000010",
  28426=>"011100100",
  28427=>"111010000",
  28428=>"111101100",
  28429=>"100000010",
  28430=>"000000000",
  28431=>"000000000",
  28432=>"111101111",
  28433=>"111111111",
  28434=>"000000110",
  28435=>"111011001",
  28436=>"000000011",
  28437=>"001000111",
  28438=>"111110101",
  28439=>"111111111",
  28440=>"000011111",
  28441=>"111111111",
  28442=>"111111110",
  28443=>"111111111",
  28444=>"000000001",
  28445=>"100000001",
  28446=>"111111000",
  28447=>"111111110",
  28448=>"111000100",
  28449=>"000111111",
  28450=>"000101101",
  28451=>"111110111",
  28452=>"111110100",
  28453=>"101111101",
  28454=>"100110110",
  28455=>"010010010",
  28456=>"011011011",
  28457=>"000111111",
  28458=>"111110110",
  28459=>"000000111",
  28460=>"111111100",
  28461=>"000001001",
  28462=>"111111100",
  28463=>"000000000",
  28464=>"010000000",
  28465=>"100110000",
  28466=>"000000110",
  28467=>"010111100",
  28468=>"110101001",
  28469=>"000000000",
  28470=>"000110100",
  28471=>"100000001",
  28472=>"000000000",
  28473=>"111111111",
  28474=>"000111111",
  28475=>"000000000",
  28476=>"001001000",
  28477=>"111000111",
  28478=>"000000000",
  28479=>"101111000",
  28480=>"000000000",
  28481=>"100100100",
  28482=>"101111111",
  28483=>"111111000",
  28484=>"111111000",
  28485=>"111100100",
  28486=>"000000001",
  28487=>"111001100",
  28488=>"000010000",
  28489=>"000000011",
  28490=>"000100100",
  28491=>"110010000",
  28492=>"000010111",
  28493=>"110111000",
  28494=>"100000000",
  28495=>"001011001",
  28496=>"001111111",
  28497=>"111101111",
  28498=>"000000000",
  28499=>"111111111",
  28500=>"000011011",
  28501=>"111111111",
  28502=>"000000000",
  28503=>"111110111",
  28504=>"100110111",
  28505=>"000000101",
  28506=>"111110000",
  28507=>"000110111",
  28508=>"111111001",
  28509=>"011111111",
  28510=>"000000110",
  28511=>"110100000",
  28512=>"111111111",
  28513=>"111110111",
  28514=>"000001100",
  28515=>"111101000",
  28516=>"111111111",
  28517=>"101001000",
  28518=>"000000000",
  28519=>"000000000",
  28520=>"001001000",
  28521=>"000110000",
  28522=>"000001111",
  28523=>"000000000",
  28524=>"111111000",
  28525=>"100100111",
  28526=>"111111100",
  28527=>"000000000",
  28528=>"000000000",
  28529=>"111011011",
  28530=>"111111011",
  28531=>"101111101",
  28532=>"001011001",
  28533=>"101111100",
  28534=>"000000000",
  28535=>"001000000",
  28536=>"111001000",
  28537=>"111110010",
  28538=>"111111000",
  28539=>"001001111",
  28540=>"001000001",
  28541=>"011011111",
  28542=>"110111111",
  28543=>"011111111",
  28544=>"101111000",
  28545=>"111111110",
  28546=>"111111111",
  28547=>"000000000",
  28548=>"111111111",
  28549=>"111101111",
  28550=>"110011000",
  28551=>"101100110",
  28552=>"111011111",
  28553=>"011001000",
  28554=>"111011010",
  28555=>"000000000",
  28556=>"111111111",
  28557=>"111111110",
  28558=>"111111100",
  28559=>"000000010",
  28560=>"111111111",
  28561=>"111110000",
  28562=>"111010010",
  28563=>"000000110",
  28564=>"100000000",
  28565=>"011111010",
  28566=>"011101100",
  28567=>"111111001",
  28568=>"111011111",
  28569=>"000000000",
  28570=>"101110111",
  28571=>"011111000",
  28572=>"111111000",
  28573=>"111111000",
  28574=>"000100100",
  28575=>"000000100",
  28576=>"111011001",
  28577=>"101111100",
  28578=>"100110001",
  28579=>"000001011",
  28580=>"001111111",
  28581=>"000000000",
  28582=>"111111111",
  28583=>"111001000",
  28584=>"100001000",
  28585=>"000010000",
  28586=>"000111111",
  28587=>"000110111",
  28588=>"000000000",
  28589=>"100100000",
  28590=>"000011111",
  28591=>"000000000",
  28592=>"000000000",
  28593=>"110010110",
  28594=>"000110111",
  28595=>"000000000",
  28596=>"000000100",
  28597=>"000100110",
  28598=>"111111101",
  28599=>"010110111",
  28600=>"110000000",
  28601=>"111001001",
  28602=>"111111111",
  28603=>"000000000",
  28604=>"110111111",
  28605=>"001001000",
  28606=>"000000111",
  28607=>"111100100",
  28608=>"000000000",
  28609=>"111111111",
  28610=>"000000000",
  28611=>"000000000",
  28612=>"101100111",
  28613=>"111111111",
  28614=>"000110111",
  28615=>"100000111",
  28616=>"000001111",
  28617=>"111001111",
  28618=>"111010000",
  28619=>"111111101",
  28620=>"110000110",
  28621=>"111100110",
  28622=>"000010000",
  28623=>"111100000",
  28624=>"000000000",
  28625=>"100111111",
  28626=>"110100111",
  28627=>"111111111",
  28628=>"001100101",
  28629=>"101101001",
  28630=>"000000000",
  28631=>"000011011",
  28632=>"000100100",
  28633=>"111011111",
  28634=>"111111111",
  28635=>"111111111",
  28636=>"111111111",
  28637=>"100110111",
  28638=>"010011011",
  28639=>"100100001",
  28640=>"111111111",
  28641=>"000000000",
  28642=>"000000000",
  28643=>"001000000",
  28644=>"011111111",
  28645=>"111111111",
  28646=>"001111111",
  28647=>"111001000",
  28648=>"000000000",
  28649=>"000100101",
  28650=>"000000000",
  28651=>"110111110",
  28652=>"000000000",
  28653=>"111111011",
  28654=>"000000100",
  28655=>"101011111",
  28656=>"000000000",
  28657=>"111001000",
  28658=>"100101110",
  28659=>"011001000",
  28660=>"111111100",
  28661=>"111111111",
  28662=>"001001001",
  28663=>"111111000",
  28664=>"000000111",
  28665=>"100101001",
  28666=>"000000010",
  28667=>"111110111",
  28668=>"011010110",
  28669=>"000100101",
  28670=>"111101111",
  28671=>"100100101",
  28672=>"110110010",
  28673=>"111101111",
  28674=>"111000000",
  28675=>"111111000",
  28676=>"111110010",
  28677=>"001101111",
  28678=>"111101000",
  28679=>"001111111",
  28680=>"000000110",
  28681=>"000001111",
  28682=>"111110001",
  28683=>"111111111",
  28684=>"001001001",
  28685=>"111111111",
  28686=>"111111011",
  28687=>"101101111",
  28688=>"000000110",
  28689=>"111111111",
  28690=>"000000000",
  28691=>"110110110",
  28692=>"111011001",
  28693=>"011001111",
  28694=>"000000000",
  28695=>"000110110",
  28696=>"100100101",
  28697=>"100100000",
  28698=>"000001111",
  28699=>"100000111",
  28700=>"100100000",
  28701=>"011011001",
  28702=>"000000000",
  28703=>"111110110",
  28704=>"000000001",
  28705=>"110111111",
  28706=>"111100000",
  28707=>"000000000",
  28708=>"111001000",
  28709=>"111111110",
  28710=>"111111100",
  28711=>"001011000",
  28712=>"000000001",
  28713=>"000000000",
  28714=>"100000000",
  28715=>"111110111",
  28716=>"111110111",
  28717=>"001001000",
  28718=>"001000101",
  28719=>"111111001",
  28720=>"111111110",
  28721=>"000000000",
  28722=>"010011001",
  28723=>"111111010",
  28724=>"111111001",
  28725=>"001111011",
  28726=>"111010011",
  28727=>"001000000",
  28728=>"110100000",
  28729=>"000000000",
  28730=>"111001111",
  28731=>"011111111",
  28732=>"001000111",
  28733=>"110000111",
  28734=>"111001001",
  28735=>"001000000",
  28736=>"000010110",
  28737=>"011001111",
  28738=>"110110000",
  28739=>"000001011",
  28740=>"011111111",
  28741=>"100000000",
  28742=>"111100000",
  28743=>"111111111",
  28744=>"011011001",
  28745=>"111001001",
  28746=>"111111111",
  28747=>"101001111",
  28748=>"001011111",
  28749=>"010010111",
  28750=>"011010010",
  28751=>"110110110",
  28752=>"100111111",
  28753=>"010111111",
  28754=>"101000110",
  28755=>"110110111",
  28756=>"000100100",
  28757=>"111100111",
  28758=>"000001001",
  28759=>"000000111",
  28760=>"000000000",
  28761=>"111111111",
  28762=>"000000000",
  28763=>"111001001",
  28764=>"000000000",
  28765=>"111111011",
  28766=>"111110111",
  28767=>"111111011",
  28768=>"000000000",
  28769=>"000000100",
  28770=>"110111111",
  28771=>"000111111",
  28772=>"000001011",
  28773=>"111111111",
  28774=>"001111111",
  28775=>"111001101",
  28776=>"111000000",
  28777=>"000000000",
  28778=>"000100111",
  28779=>"111111111",
  28780=>"111111000",
  28781=>"111111111",
  28782=>"000000000",
  28783=>"000111011",
  28784=>"100111111",
  28785=>"111111001",
  28786=>"100100111",
  28787=>"000010111",
  28788=>"000000000",
  28789=>"111111111",
  28790=>"001000000",
  28791=>"100100101",
  28792=>"000001000",
  28793=>"000000000",
  28794=>"001001001",
  28795=>"000000001",
  28796=>"100111100",
  28797=>"111011111",
  28798=>"101001000",
  28799=>"111111111",
  28800=>"001001001",
  28801=>"111111111",
  28802=>"010010100",
  28803=>"000000001",
  28804=>"000100111",
  28805=>"000111111",
  28806=>"110110010",
  28807=>"000001000",
  28808=>"000000000",
  28809=>"000000001",
  28810=>"111100101",
  28811=>"111111001",
  28812=>"111111111",
  28813=>"110110111",
  28814=>"110111010",
  28815=>"111111111",
  28816=>"110111000",
  28817=>"110110000",
  28818=>"000011111",
  28819=>"110110111",
  28820=>"000000111",
  28821=>"000001101",
  28822=>"011111010",
  28823=>"000001111",
  28824=>"001000100",
  28825=>"110111100",
  28826=>"111111101",
  28827=>"111100100",
  28828=>"111111110",
  28829=>"001111111",
  28830=>"111111111",
  28831=>"001001001",
  28832=>"000000110",
  28833=>"000110001",
  28834=>"111111001",
  28835=>"000000000",
  28836=>"001001001",
  28837=>"101001001",
  28838=>"000000000",
  28839=>"111111111",
  28840=>"111011001",
  28841=>"100111111",
  28842=>"111100100",
  28843=>"000001001",
  28844=>"111111000",
  28845=>"001001011",
  28846=>"001000111",
  28847=>"001111101",
  28848=>"111111111",
  28849=>"011011000",
  28850=>"011111011",
  28851=>"000000000",
  28852=>"000000001",
  28853=>"011111111",
  28854=>"000101111",
  28855=>"000011111",
  28856=>"101111111",
  28857=>"000011000",
  28858=>"000111111",
  28859=>"000000100",
  28860=>"111111111",
  28861=>"110000000",
  28862=>"000111111",
  28863=>"001000001",
  28864=>"111111111",
  28865=>"000001111",
  28866=>"001000000",
  28867=>"111101111",
  28868=>"011111111",
  28869=>"111000000",
  28870=>"000000111",
  28871=>"111011111",
  28872=>"000011111",
  28873=>"110111111",
  28874=>"000000000",
  28875=>"000001011",
  28876=>"111111101",
  28877=>"100101101",
  28878=>"000000110",
  28879=>"110010011",
  28880=>"111100000",
  28881=>"001001011",
  28882=>"000000000",
  28883=>"110111111",
  28884=>"111110000",
  28885=>"110110110",
  28886=>"000000000",
  28887=>"001000000",
  28888=>"000000011",
  28889=>"110010000",
  28890=>"111111111",
  28891=>"100100101",
  28892=>"111111110",
  28893=>"111111101",
  28894=>"001101111",
  28895=>"101111111",
  28896=>"011000010",
  28897=>"001000000",
  28898=>"000000000",
  28899=>"001000001",
  28900=>"000000000",
  28901=>"100000100",
  28902=>"111111111",
  28903=>"100001001",
  28904=>"000000001",
  28905=>"000101101",
  28906=>"111111111",
  28907=>"001001000",
  28908=>"000000000",
  28909=>"000000111",
  28910=>"111000000",
  28911=>"000011111",
  28912=>"000000001",
  28913=>"000001000",
  28914=>"000111111",
  28915=>"110011000",
  28916=>"111001000",
  28917=>"101001011",
  28918=>"110000000",
  28919=>"001111111",
  28920=>"000111111",
  28921=>"000000111",
  28922=>"110111011",
  28923=>"110000000",
  28924=>"111110100",
  28925=>"110110010",
  28926=>"100111000",
  28927=>"101100111",
  28928=>"011111111",
  28929=>"000100001",
  28930=>"111101111",
  28931=>"000000001",
  28932=>"111001111",
  28933=>"100101001",
  28934=>"000111111",
  28935=>"110000001",
  28936=>"011011011",
  28937=>"000000000",
  28938=>"000001101",
  28939=>"100000000",
  28940=>"001000001",
  28941=>"111110000",
  28942=>"111111001",
  28943=>"001001111",
  28944=>"111000000",
  28945=>"110011010",
  28946=>"000100111",
  28947=>"000000000",
  28948=>"101000011",
  28949=>"000000110",
  28950=>"100100110",
  28951=>"000000000",
  28952=>"111110010",
  28953=>"111111000",
  28954=>"001001111",
  28955=>"111001000",
  28956=>"111100000",
  28957=>"000000000",
  28958=>"000000000",
  28959=>"000000011",
  28960=>"010000000",
  28961=>"000000000",
  28962=>"111010001",
  28963=>"000000100",
  28964=>"110000000",
  28965=>"111111111",
  28966=>"000001001",
  28967=>"111111111",
  28968=>"101100110",
  28969=>"111111010",
  28970=>"000101101",
  28971=>"011011000",
  28972=>"111111111",
  28973=>"000010011",
  28974=>"111111111",
  28975=>"110000011",
  28976=>"001001111",
  28977=>"111111000",
  28978=>"111111010",
  28979=>"111111111",
  28980=>"001101111",
  28981=>"000100010",
  28982=>"100000000",
  28983=>"111111111",
  28984=>"000000111",
  28985=>"101111111",
  28986=>"000000000",
  28987=>"000000000",
  28988=>"111011011",
  28989=>"111111011",
  28990=>"000000000",
  28991=>"000100110",
  28992=>"000111111",
  28993=>"000110000",
  28994=>"110000011",
  28995=>"111111111",
  28996=>"101011111",
  28997=>"010000001",
  28998=>"000000000",
  28999=>"011110110",
  29000=>"100111000",
  29001=>"111000111",
  29002=>"100000011",
  29003=>"000000111",
  29004=>"000001111",
  29005=>"001000111",
  29006=>"000000111",
  29007=>"000110111",
  29008=>"110111110",
  29009=>"000000110",
  29010=>"110110111",
  29011=>"000001111",
  29012=>"111111111",
  29013=>"011000000",
  29014=>"000000011",
  29015=>"000000001",
  29016=>"000000000",
  29017=>"000000000",
  29018=>"011111110",
  29019=>"000001001",
  29020=>"001000000",
  29021=>"000001001",
  29022=>"100000000",
  29023=>"000010011",
  29024=>"110110000",
  29025=>"000000001",
  29026=>"000100100",
  29027=>"001000000",
  29028=>"111111011",
  29029=>"000000011",
  29030=>"000000111",
  29031=>"001010111",
  29032=>"110000000",
  29033=>"101111111",
  29034=>"000100000",
  29035=>"000110110",
  29036=>"000000101",
  29037=>"011111111",
  29038=>"000000111",
  29039=>"110110000",
  29040=>"000000001",
  29041=>"000000000",
  29042=>"000001011",
  29043=>"001000011",
  29044=>"000010011",
  29045=>"101111111",
  29046=>"110000111",
  29047=>"101111111",
  29048=>"111001101",
  29049=>"111000111",
  29050=>"111111111",
  29051=>"100110010",
  29052=>"010000000",
  29053=>"000000000",
  29054=>"101101111",
  29055=>"000011001",
  29056=>"000000110",
  29057=>"000111011",
  29058=>"000000000",
  29059=>"000000001",
  29060=>"111101101",
  29061=>"011111001",
  29062=>"001001001",
  29063=>"101001001",
  29064=>"111001100",
  29065=>"111111111",
  29066=>"101111111",
  29067=>"111111111",
  29068=>"111111111",
  29069=>"000110110",
  29070=>"000000001",
  29071=>"111111111",
  29072=>"000000000",
  29073=>"110000000",
  29074=>"000000001",
  29075=>"001100000",
  29076=>"000110000",
  29077=>"000100111",
  29078=>"110110000",
  29079=>"111111011",
  29080=>"001000100",
  29081=>"111000110",
  29082=>"011111110",
  29083=>"111000000",
  29084=>"000011000",
  29085=>"111111000",
  29086=>"000001001",
  29087=>"111111111",
  29088=>"001001000",
  29089=>"011011011",
  29090=>"000000001",
  29091=>"101101000",
  29092=>"111111000",
  29093=>"000101010",
  29094=>"001001001",
  29095=>"000001011",
  29096=>"110110111",
  29097=>"111001000",
  29098=>"000000000",
  29099=>"000100101",
  29100=>"000001111",
  29101=>"100001100",
  29102=>"000000110",
  29103=>"000000100",
  29104=>"000000000",
  29105=>"001101101",
  29106=>"100000000",
  29107=>"111111111",
  29108=>"001011111",
  29109=>"000000101",
  29110=>"101111111",
  29111=>"111111111",
  29112=>"111010000",
  29113=>"000000000",
  29114=>"110000000",
  29115=>"000000000",
  29116=>"110100000",
  29117=>"111111111",
  29118=>"000000110",
  29119=>"010111110",
  29120=>"110110000",
  29121=>"111111111",
  29122=>"000000000",
  29123=>"001001111",
  29124=>"000000011",
  29125=>"100001001",
  29126=>"000000000",
  29127=>"111111111",
  29128=>"000001000",
  29129=>"100100010",
  29130=>"001000000",
  29131=>"101101111",
  29132=>"110110000",
  29133=>"110110110",
  29134=>"100000000",
  29135=>"010111111",
  29136=>"110110111",
  29137=>"000000001",
  29138=>"111111111",
  29139=>"000000000",
  29140=>"111111000",
  29141=>"010000000",
  29142=>"000000000",
  29143=>"100100100",
  29144=>"110110110",
  29145=>"000000011",
  29146=>"000000000",
  29147=>"000011111",
  29148=>"000011011",
  29149=>"011101111",
  29150=>"111111101",
  29151=>"000000111",
  29152=>"000100110",
  29153=>"101000110",
  29154=>"111010000",
  29155=>"000111111",
  29156=>"000010011",
  29157=>"000000000",
  29158=>"011001001",
  29159=>"110000000",
  29160=>"111111111",
  29161=>"000110111",
  29162=>"111001100",
  29163=>"110111011",
  29164=>"000001111",
  29165=>"110100100",
  29166=>"100000111",
  29167=>"111111111",
  29168=>"000000000",
  29169=>"000000000",
  29170=>"000011011",
  29171=>"000001011",
  29172=>"000000111",
  29173=>"001001001",
  29174=>"111111111",
  29175=>"110110110",
  29176=>"011111000",
  29177=>"000000010",
  29178=>"000000000",
  29179=>"000000001",
  29180=>"111110000",
  29181=>"011011011",
  29182=>"100100000",
  29183=>"111111000",
  29184=>"000000000",
  29185=>"000001011",
  29186=>"001111111",
  29187=>"000111111",
  29188=>"000000100",
  29189=>"001000000",
  29190=>"110111111",
  29191=>"001001111",
  29192=>"000100100",
  29193=>"111000000",
  29194=>"111111111",
  29195=>"001001001",
  29196=>"000000100",
  29197=>"010000000",
  29198=>"111011011",
  29199=>"110111111",
  29200=>"000000110",
  29201=>"000110111",
  29202=>"000000000",
  29203=>"100000000",
  29204=>"111111000",
  29205=>"111111111",
  29206=>"111111111",
  29207=>"000000000",
  29208=>"110110000",
  29209=>"110100011",
  29210=>"111111111",
  29211=>"000000011",
  29212=>"111111111",
  29213=>"000000000",
  29214=>"110110111",
  29215=>"111111111",
  29216=>"000010010",
  29217=>"111111101",
  29218=>"110111111",
  29219=>"111000111",
  29220=>"111111101",
  29221=>"111111111",
  29222=>"111000000",
  29223=>"000111100",
  29224=>"111111111",
  29225=>"111111111",
  29226=>"111111110",
  29227=>"110101111",
  29228=>"100110000",
  29229=>"111111000",
  29230=>"111111100",
  29231=>"001111000",
  29232=>"100000000",
  29233=>"010011011",
  29234=>"001011111",
  29235=>"110111111",
  29236=>"000000000",
  29237=>"000000000",
  29238=>"000110110",
  29239=>"100000010",
  29240=>"011000000",
  29241=>"111110000",
  29242=>"000000000",
  29243=>"000000000",
  29244=>"000000100",
  29245=>"110000000",
  29246=>"000000000",
  29247=>"000000000",
  29248=>"000010111",
  29249=>"011011000",
  29250=>"010111111",
  29251=>"100000100",
  29252=>"000000000",
  29253=>"100110100",
  29254=>"111000000",
  29255=>"111111111",
  29256=>"111111101",
  29257=>"000000111",
  29258=>"111111111",
  29259=>"111111111",
  29260=>"000100000",
  29261=>"001111001",
  29262=>"000000000",
  29263=>"111111111",
  29264=>"111110110",
  29265=>"000000000",
  29266=>"111111111",
  29267=>"110110110",
  29268=>"000000000",
  29269=>"000011001",
  29270=>"110100100",
  29271=>"000000000",
  29272=>"111111111",
  29273=>"000000000",
  29274=>"111111111",
  29275=>"000010110",
  29276=>"001000000",
  29277=>"000001000",
  29278=>"111111101",
  29279=>"000000001",
  29280=>"111111111",
  29281=>"000000000",
  29282=>"010000000",
  29283=>"110001011",
  29284=>"111111111",
  29285=>"100100111",
  29286=>"000000011",
  29287=>"111101110",
  29288=>"111111110",
  29289=>"111101111",
  29290=>"100000111",
  29291=>"000000000",
  29292=>"000000000",
  29293=>"111111111",
  29294=>"000000000",
  29295=>"000000000",
  29296=>"000000000",
  29297=>"000000000",
  29298=>"000000010",
  29299=>"110101000",
  29300=>"000000000",
  29301=>"000000000",
  29302=>"000001000",
  29303=>"001111111",
  29304=>"101000000",
  29305=>"101111111",
  29306=>"110010000",
  29307=>"000000000",
  29308=>"000001000",
  29309=>"111111111",
  29310=>"000000111",
  29311=>"011011011",
  29312=>"111111111",
  29313=>"111111000",
  29314=>"000000000",
  29315=>"010000000",
  29316=>"011000000",
  29317=>"111111111",
  29318=>"011011010",
  29319=>"000111111",
  29320=>"111111110",
  29321=>"111111111",
  29322=>"111111111",
  29323=>"111110110",
  29324=>"111111111",
  29325=>"111111111",
  29326=>"111011111",
  29327=>"011001010",
  29328=>"111111111",
  29329=>"000000111",
  29330=>"011011111",
  29331=>"111111101",
  29332=>"000111111",
  29333=>"111111111",
  29334=>"000000000",
  29335=>"000000111",
  29336=>"000000111",
  29337=>"001011011",
  29338=>"010000000",
  29339=>"001001000",
  29340=>"001000000",
  29341=>"010000111",
  29342=>"111001000",
  29343=>"000010010",
  29344=>"111111111",
  29345=>"001001001",
  29346=>"000111111",
  29347=>"111011111",
  29348=>"000000000",
  29349=>"001111011",
  29350=>"111111111",
  29351=>"000000000",
  29352=>"000001111",
  29353=>"000000001",
  29354=>"100100100",
  29355=>"000001001",
  29356=>"000000000",
  29357=>"000000000",
  29358=>"000000000",
  29359=>"000000000",
  29360=>"111111111",
  29361=>"111111111",
  29362=>"111111000",
  29363=>"000111000",
  29364=>"111011111",
  29365=>"000000000",
  29366=>"110111100",
  29367=>"111111111",
  29368=>"100000010",
  29369=>"111111110",
  29370=>"000000000",
  29371=>"000000001",
  29372=>"111001001",
  29373=>"000010000",
  29374=>"000000000",
  29375=>"000000101",
  29376=>"100000000",
  29377=>"111111111",
  29378=>"010111111",
  29379=>"111111111",
  29380=>"000000000",
  29381=>"000111001",
  29382=>"110111000",
  29383=>"000000000",
  29384=>"111111111",
  29385=>"000110000",
  29386=>"110100100",
  29387=>"111111111",
  29388=>"100100000",
  29389=>"000000000",
  29390=>"111111000",
  29391=>"010010110",
  29392=>"111111111",
  29393=>"110111110",
  29394=>"001000000",
  29395=>"000000000",
  29396=>"001001001",
  29397=>"001000101",
  29398=>"110000100",
  29399=>"000000000",
  29400=>"001011011",
  29401=>"000100100",
  29402=>"000010111",
  29403=>"000111111",
  29404=>"111111011",
  29405=>"111101001",
  29406=>"111001001",
  29407=>"000000000",
  29408=>"111111100",
  29409=>"101111100",
  29410=>"111111011",
  29411=>"100111111",
  29412=>"101111111",
  29413=>"011011111",
  29414=>"000111111",
  29415=>"111111111",
  29416=>"101000000",
  29417=>"000000111",
  29418=>"110000111",
  29419=>"001111111",
  29420=>"000000100",
  29421=>"000100000",
  29422=>"110000011",
  29423=>"111111111",
  29424=>"110111111",
  29425=>"000000000",
  29426=>"000000100",
  29427=>"011111000",
  29428=>"111111111",
  29429=>"000000000",
  29430=>"000000011",
  29431=>"001001000",
  29432=>"000000000",
  29433=>"111111100",
  29434=>"111111111",
  29435=>"111101111",
  29436=>"000000000",
  29437=>"111111111",
  29438=>"110111101",
  29439=>"111111111",
  29440=>"110110010",
  29441=>"100100110",
  29442=>"111111111",
  29443=>"001011001",
  29444=>"000000111",
  29445=>"111101000",
  29446=>"000000111",
  29447=>"100000111",
  29448=>"110111110",
  29449=>"011011111",
  29450=>"000000000",
  29451=>"000000001",
  29452=>"001000111",
  29453=>"101101111",
  29454=>"011111111",
  29455=>"111000000",
  29456=>"011000001",
  29457=>"111000000",
  29458=>"000000000",
  29459=>"111101111",
  29460=>"000000000",
  29461=>"110000000",
  29462=>"000010000",
  29463=>"111111111",
  29464=>"000000010",
  29465=>"100001000",
  29466=>"011011011",
  29467=>"111111000",
  29468=>"111111111",
  29469=>"000001000",
  29470=>"111111110",
  29471=>"001001000",
  29472=>"010100011",
  29473=>"000000000",
  29474=>"000000000",
  29475=>"000000110",
  29476=>"000000000",
  29477=>"111110111",
  29478=>"000010010",
  29479=>"000001011",
  29480=>"100111111",
  29481=>"000000000",
  29482=>"111101111",
  29483=>"111111111",
  29484=>"000010000",
  29485=>"100000000",
  29486=>"111011111",
  29487=>"000000111",
  29488=>"000000000",
  29489=>"000000000",
  29490=>"111111111",
  29491=>"100100010",
  29492=>"111011000",
  29493=>"110000000",
  29494=>"000000000",
  29495=>"111111111",
  29496=>"100100000",
  29497=>"000000000",
  29498=>"010000000",
  29499=>"000000000",
  29500=>"111111111",
  29501=>"101000000",
  29502=>"111100000",
  29503=>"000000110",
  29504=>"111111111",
  29505=>"000000000",
  29506=>"110110110",
  29507=>"100110111",
  29508=>"000000011",
  29509=>"110111111",
  29510=>"111111011",
  29511=>"000000000",
  29512=>"011111111",
  29513=>"111111111",
  29514=>"100110010",
  29515=>"000000000",
  29516=>"111001001",
  29517=>"111000000",
  29518=>"100111111",
  29519=>"000000000",
  29520=>"110110110",
  29521=>"000001101",
  29522=>"000000111",
  29523=>"000000000",
  29524=>"000000000",
  29525=>"111111011",
  29526=>"001000111",
  29527=>"111111111",
  29528=>"111111111",
  29529=>"111111111",
  29530=>"111111111",
  29531=>"000000000",
  29532=>"000111111",
  29533=>"000000000",
  29534=>"100100000",
  29535=>"111111010",
  29536=>"000000000",
  29537=>"111111111",
  29538=>"001001000",
  29539=>"001101111",
  29540=>"111111010",
  29541=>"010100111",
  29542=>"111111011",
  29543=>"001001000",
  29544=>"111101000",
  29545=>"000000000",
  29546=>"000000000",
  29547=>"110111111",
  29548=>"001000000",
  29549=>"111111111",
  29550=>"111111111",
  29551=>"000100100",
  29552=>"111111111",
  29553=>"111011001",
  29554=>"000111001",
  29555=>"100111111",
  29556=>"111011000",
  29557=>"111111110",
  29558=>"111111111",
  29559=>"111111000",
  29560=>"111111111",
  29561=>"000000000",
  29562=>"111100111",
  29563=>"111011000",
  29564=>"000001101",
  29565=>"011000100",
  29566=>"000000000",
  29567=>"111111111",
  29568=>"101001001",
  29569=>"110111111",
  29570=>"000000001",
  29571=>"000100111",
  29572=>"000000111",
  29573=>"000000001",
  29574=>"111111111",
  29575=>"011011000",
  29576=>"000000000",
  29577=>"001000000",
  29578=>"111111111",
  29579=>"000000101",
  29580=>"111000000",
  29581=>"100100000",
  29582=>"000000000",
  29583=>"000110110",
  29584=>"001001011",
  29585=>"000000000",
  29586=>"000000000",
  29587=>"100000000",
  29588=>"011001101",
  29589=>"000110011",
  29590=>"100000000",
  29591=>"001000000",
  29592=>"000000110",
  29593=>"010111111",
  29594=>"110000010",
  29595=>"011111110",
  29596=>"111111011",
  29597=>"111110111",
  29598=>"111101001",
  29599=>"111000000",
  29600=>"000000001",
  29601=>"001000000",
  29602=>"111100100",
  29603=>"000000000",
  29604=>"111111111",
  29605=>"111100000",
  29606=>"111111111",
  29607=>"000000000",
  29608=>"110111100",
  29609=>"111011011",
  29610=>"110110111",
  29611=>"100100000",
  29612=>"000000000",
  29613=>"001010110",
  29614=>"110110000",
  29615=>"000100111",
  29616=>"100000111",
  29617=>"111111111",
  29618=>"111111111",
  29619=>"000000000",
  29620=>"111111111",
  29621=>"011000000",
  29622=>"000000000",
  29623=>"111010000",
  29624=>"001000000",
  29625=>"010010111",
  29626=>"000011000",
  29627=>"100000000",
  29628=>"111111111",
  29629=>"111111111",
  29630=>"111000000",
  29631=>"110110111",
  29632=>"100000000",
  29633=>"000000000",
  29634=>"000000000",
  29635=>"000000000",
  29636=>"110110111",
  29637=>"011111111",
  29638=>"111111111",
  29639=>"111100000",
  29640=>"000000000",
  29641=>"010111111",
  29642=>"110111111",
  29643=>"000000000",
  29644=>"000010000",
  29645=>"110110110",
  29646=>"000100000",
  29647=>"111110111",
  29648=>"100100111",
  29649=>"101101000",
  29650=>"000000000",
  29651=>"111111111",
  29652=>"000000000",
  29653=>"000000100",
  29654=>"111111111",
  29655=>"100000000",
  29656=>"111111000",
  29657=>"111100100",
  29658=>"011010000",
  29659=>"110100100",
  29660=>"111111111",
  29661=>"101111111",
  29662=>"000000000",
  29663=>"110000100",
  29664=>"001000000",
  29665=>"101110110",
  29666=>"111111111",
  29667=>"000000000",
  29668=>"111111111",
  29669=>"000000000",
  29670=>"000100101",
  29671=>"111011001",
  29672=>"010001011",
  29673=>"000000000",
  29674=>"000011000",
  29675=>"011001011",
  29676=>"001000000",
  29677=>"000000000",
  29678=>"001000000",
  29679=>"000000100",
  29680=>"111111111",
  29681=>"110111111",
  29682=>"111111111",
  29683=>"111111100",
  29684=>"111111111",
  29685=>"000100000",
  29686=>"000000000",
  29687=>"010001000",
  29688=>"111111011",
  29689=>"001000001",
  29690=>"100110110",
  29691=>"000000000",
  29692=>"111111111",
  29693=>"011000000",
  29694=>"100000001",
  29695=>"000000001",
  29696=>"111111111",
  29697=>"111111111",
  29698=>"000001111",
  29699=>"011111111",
  29700=>"101111111",
  29701=>"000000001",
  29702=>"000000011",
  29703=>"111111111",
  29704=>"111111111",
  29705=>"111111111",
  29706=>"111111111",
  29707=>"111001000",
  29708=>"111101111",
  29709=>"111101111",
  29710=>"110110000",
  29711=>"001001001",
  29712=>"111111111",
  29713=>"010110111",
  29714=>"000000010",
  29715=>"000010001",
  29716=>"011000110",
  29717=>"001101000",
  29718=>"111111010",
  29719=>"111100000",
  29720=>"001011111",
  29721=>"111110000",
  29722=>"011000000",
  29723=>"011111111",
  29724=>"001011010",
  29725=>"011000000",
  29726=>"111110010",
  29727=>"111100000",
  29728=>"001111111",
  29729=>"111111000",
  29730=>"001000111",
  29731=>"111011000",
  29732=>"001111111",
  29733=>"000000011",
  29734=>"000000000",
  29735=>"111110000",
  29736=>"011111100",
  29737=>"000111000",
  29738=>"111111111",
  29739=>"000000000",
  29740=>"111001000",
  29741=>"011011000",
  29742=>"111000000",
  29743=>"111111111",
  29744=>"001111110",
  29745=>"000111111",
  29746=>"010110111",
  29747=>"111111111",
  29748=>"111111000",
  29749=>"111101100",
  29750=>"000000000",
  29751=>"000000000",
  29752=>"110110000",
  29753=>"111111110",
  29754=>"111000000",
  29755=>"001000001",
  29756=>"000000000",
  29757=>"100000000",
  29758=>"111110111",
  29759=>"000000000",
  29760=>"001000000",
  29761=>"110111100",
  29762=>"101001000",
  29763=>"101000000",
  29764=>"100100111",
  29765=>"111000101",
  29766=>"000000001",
  29767=>"000000000",
  29768=>"111110111",
  29769=>"000000000",
  29770=>"111111111",
  29771=>"000000011",
  29772=>"101111000",
  29773=>"000111111",
  29774=>"001000000",
  29775=>"111101000",
  29776=>"110001000",
  29777=>"011111111",
  29778=>"101111111",
  29779=>"000000000",
  29780=>"011111111",
  29781=>"111000010",
  29782=>"000111110",
  29783=>"011001111",
  29784=>"000111111",
  29785=>"111000000",
  29786=>"011111111",
  29787=>"011000100",
  29788=>"000110111",
  29789=>"110111001",
  29790=>"000001111",
  29791=>"111100111",
  29792=>"100100000",
  29793=>"000000000",
  29794=>"011111111",
  29795=>"111111111",
  29796=>"000000000",
  29797=>"111111111",
  29798=>"111111000",
  29799=>"111111111",
  29800=>"000000000",
  29801=>"011110110",
  29802=>"111111000",
  29803=>"000111111",
  29804=>"101101111",
  29805=>"000000111",
  29806=>"001000001",
  29807=>"000000111",
  29808=>"100000000",
  29809=>"000000000",
  29810=>"110111111",
  29811=>"001001001",
  29812=>"000000001",
  29813=>"000000000",
  29814=>"000000011",
  29815=>"000100100",
  29816=>"111111111",
  29817=>"000011000",
  29818=>"111111111",
  29819=>"000000111",
  29820=>"111011001",
  29821=>"111111111",
  29822=>"111111111",
  29823=>"111111111",
  29824=>"000000000",
  29825=>"000000000",
  29826=>"110000000",
  29827=>"000000101",
  29828=>"000000000",
  29829=>"000000001",
  29830=>"101111111",
  29831=>"001000000",
  29832=>"000000000",
  29833=>"000000111",
  29834=>"100111111",
  29835=>"010000110",
  29836=>"111111110",
  29837=>"000000111",
  29838=>"001000000",
  29839=>"011000000",
  29840=>"111111000",
  29841=>"000111111",
  29842=>"111111000",
  29843=>"111111000",
  29844=>"110010111",
  29845=>"011001011",
  29846=>"111011011",
  29847=>"111110000",
  29848=>"111111111",
  29849=>"000011011",
  29850=>"111111111",
  29851=>"011001000",
  29852=>"100000000",
  29853=>"101001000",
  29854=>"111111111",
  29855=>"111111001",
  29856=>"111110100",
  29857=>"001000000",
  29858=>"000000111",
  29859=>"000000111",
  29860=>"000001101",
  29861=>"000000000",
  29862=>"110010110",
  29863=>"111110010",
  29864=>"111011011",
  29865=>"111111000",
  29866=>"000000101",
  29867=>"111111111",
  29868=>"111011111",
  29869=>"000000000",
  29870=>"000000000",
  29871=>"111010000",
  29872=>"111110000",
  29873=>"111101101",
  29874=>"010110110",
  29875=>"110110000",
  29876=>"111110100",
  29877=>"001100100",
  29878=>"000101111",
  29879=>"110110111",
  29880=>"111111111",
  29881=>"111010000",
  29882=>"000000001",
  29883=>"011001110",
  29884=>"111000011",
  29885=>"000010000",
  29886=>"000111111",
  29887=>"001001001",
  29888=>"000000111",
  29889=>"100000111",
  29890=>"111111111",
  29891=>"000000000",
  29892=>"001000000",
  29893=>"000101111",
  29894=>"100111111",
  29895=>"000000010",
  29896=>"011011000",
  29897=>"000000000",
  29898=>"000000000",
  29899=>"000000011",
  29900=>"000000001",
  29901=>"000000000",
  29902=>"011001000",
  29903=>"000000000",
  29904=>"000000001",
  29905=>"010011111",
  29906=>"001011011",
  29907=>"000000000",
  29908=>"001001001",
  29909=>"000000000",
  29910=>"000011111",
  29911=>"110000100",
  29912=>"110110010",
  29913=>"100000111",
  29914=>"000000000",
  29915=>"111111000",
  29916=>"111000001",
  29917=>"111000000",
  29918=>"000111011",
  29919=>"100111001",
  29920=>"010111000",
  29921=>"001111100",
  29922=>"011111111",
  29923=>"010110111",
  29924=>"100001011",
  29925=>"110000000",
  29926=>"111111000",
  29927=>"111000010",
  29928=>"000000101",
  29929=>"100101110",
  29930=>"110001111",
  29931=>"000000111",
  29932=>"000000111",
  29933=>"111110010",
  29934=>"111000011",
  29935=>"000000111",
  29936=>"000000000",
  29937=>"000110111",
  29938=>"111100100",
  29939=>"100111111",
  29940=>"111011111",
  29941=>"001111111",
  29942=>"111111111",
  29943=>"011000100",
  29944=>"000000011",
  29945=>"000000000",
  29946=>"000000000",
  29947=>"010000000",
  29948=>"111111111",
  29949=>"001001000",
  29950=>"111001000",
  29951=>"011000000",
  29952=>"111001001",
  29953=>"001000000",
  29954=>"111111000",
  29955=>"000000000",
  29956=>"111111110",
  29957=>"000000000",
  29958=>"111000000",
  29959=>"000000001",
  29960=>"111111111",
  29961=>"111000000",
  29962=>"000000111",
  29963=>"111111011",
  29964=>"000000110",
  29965=>"111111111",
  29966=>"001111111",
  29967=>"001001011",
  29968=>"000000000",
  29969=>"000000100",
  29970=>"001000000",
  29971=>"100111111",
  29972=>"001010111",
  29973=>"101111111",
  29974=>"111010000",
  29975=>"000010111",
  29976=>"111010000",
  29977=>"000000000",
  29978=>"111111001",
  29979=>"010000000",
  29980=>"111110000",
  29981=>"000000111",
  29982=>"000000000",
  29983=>"001100111",
  29984=>"010110111",
  29985=>"010010001",
  29986=>"000111111",
  29987=>"101111111",
  29988=>"001000010",
  29989=>"001000000",
  29990=>"110111101",
  29991=>"000000110",
  29992=>"011000111",
  29993=>"111111110",
  29994=>"111000000",
  29995=>"010111111",
  29996=>"111011000",
  29997=>"110110100",
  29998=>"000010111",
  29999=>"111000000",
  30000=>"111001000",
  30001=>"000000000",
  30002=>"101001000",
  30003=>"000110111",
  30004=>"111000000",
  30005=>"011000111",
  30006=>"000000000",
  30007=>"000000011",
  30008=>"011111111",
  30009=>"111111111",
  30010=>"000000111",
  30011=>"001001100",
  30012=>"111011011",
  30013=>"000000111",
  30014=>"111111111",
  30015=>"100111001",
  30016=>"010000100",
  30017=>"111000000",
  30018=>"000000111",
  30019=>"111011111",
  30020=>"000000000",
  30021=>"100010110",
  30022=>"011111111",
  30023=>"010111111",
  30024=>"111111111",
  30025=>"000000000",
  30026=>"111000000",
  30027=>"010011000",
  30028=>"001000000",
  30029=>"001000111",
  30030=>"000000110",
  30031=>"111001100",
  30032=>"111000000",
  30033=>"111111111",
  30034=>"101000000",
  30035=>"010000111",
  30036=>"000000000",
  30037=>"111111110",
  30038=>"111111000",
  30039=>"000000001",
  30040=>"110100000",
  30041=>"111111110",
  30042=>"000000000",
  30043=>"101000111",
  30044=>"000111101",
  30045=>"111111011",
  30046=>"000000111",
  30047=>"111100000",
  30048=>"111111111",
  30049=>"001001111",
  30050=>"111111111",
  30051=>"111011000",
  30052=>"000000111",
  30053=>"111111111",
  30054=>"110110110",
  30055=>"000001000",
  30056=>"010001001",
  30057=>"000000100",
  30058=>"011000000",
  30059=>"101001000",
  30060=>"000110100",
  30061=>"000100000",
  30062=>"000000000",
  30063=>"000000111",
  30064=>"101000001",
  30065=>"111111110",
  30066=>"101000001",
  30067=>"000000000",
  30068=>"101000111",
  30069=>"100000000",
  30070=>"010000000",
  30071=>"011111011",
  30072=>"111111000",
  30073=>"000000101",
  30074=>"111011000",
  30075=>"001110110",
  30076=>"111101100",
  30077=>"110110110",
  30078=>"000011111",
  30079=>"000000111",
  30080=>"101111111",
  30081=>"000111001",
  30082=>"001001001",
  30083=>"111011011",
  30084=>"111000000",
  30085=>"111111000",
  30086=>"111101000",
  30087=>"000000111",
  30088=>"111001000",
  30089=>"111111000",
  30090=>"111111001",
  30091=>"111000111",
  30092=>"000001001",
  30093=>"011000000",
  30094=>"110010110",
  30095=>"000111111",
  30096=>"111001000",
  30097=>"001100111",
  30098=>"000010010",
  30099=>"011011100",
  30100=>"001001001",
  30101=>"001101011",
  30102=>"001011001",
  30103=>"100111100",
  30104=>"111111111",
  30105=>"000001000",
  30106=>"010111111",
  30107=>"000000000",
  30108=>"111111111",
  30109=>"111111000",
  30110=>"001001000",
  30111=>"000000110",
  30112=>"000000000",
  30113=>"111111111",
  30114=>"000010011",
  30115=>"000011000",
  30116=>"100000000",
  30117=>"000000000",
  30118=>"000111010",
  30119=>"111011011",
  30120=>"111010000",
  30121=>"000000000",
  30122=>"000000001",
  30123=>"000000000",
  30124=>"000000111",
  30125=>"101111111",
  30126=>"011111000",
  30127=>"000110010",
  30128=>"001111000",
  30129=>"000000010",
  30130=>"111010000",
  30131=>"010111111",
  30132=>"000000000",
  30133=>"111000000",
  30134=>"100100000",
  30135=>"000000111",
  30136=>"000000100",
  30137=>"000001011",
  30138=>"000101111",
  30139=>"001000000",
  30140=>"111111011",
  30141=>"101000011",
  30142=>"000011110",
  30143=>"111011010",
  30144=>"110100100",
  30145=>"000000000",
  30146=>"111010010",
  30147=>"000000000",
  30148=>"100111111",
  30149=>"110111111",
  30150=>"110111000",
  30151=>"000000111",
  30152=>"000001111",
  30153=>"000000111",
  30154=>"111011001",
  30155=>"111101000",
  30156=>"111110111",
  30157=>"000111111",
  30158=>"000111111",
  30159=>"000110000",
  30160=>"000000110",
  30161=>"110111111",
  30162=>"111011000",
  30163=>"000100110",
  30164=>"001001101",
  30165=>"111111011",
  30166=>"000011111",
  30167=>"100000111",
  30168=>"111111000",
  30169=>"100100111",
  30170=>"111111111",
  30171=>"110111111",
  30172=>"111011000",
  30173=>"001100000",
  30174=>"111111000",
  30175=>"011011000",
  30176=>"111011000",
  30177=>"111000011",
  30178=>"011111111",
  30179=>"000100111",
  30180=>"101101111",
  30181=>"000000111",
  30182=>"000000001",
  30183=>"000000111",
  30184=>"111111011",
  30185=>"000100111",
  30186=>"000110111",
  30187=>"000110111",
  30188=>"111010000",
  30189=>"000000100",
  30190=>"000100110",
  30191=>"101100000",
  30192=>"000000110",
  30193=>"110111001",
  30194=>"000000111",
  30195=>"010000000",
  30196=>"111000101",
  30197=>"011001000",
  30198=>"000110111",
  30199=>"111111100",
  30200=>"000001111",
  30201=>"111110110",
  30202=>"111111111",
  30203=>"111111110",
  30204=>"000000000",
  30205=>"001111111",
  30206=>"111111001",
  30207=>"101000000",
  30208=>"001001001",
  30209=>"111000111",
  30210=>"111000001",
  30211=>"000000000",
  30212=>"001000000",
  30213=>"111000000",
  30214=>"000010000",
  30215=>"000000001",
  30216=>"001000010",
  30217=>"000000000",
  30218=>"111000000",
  30219=>"000111111",
  30220=>"100110000",
  30221=>"111111111",
  30222=>"000111111",
  30223=>"000000111",
  30224=>"110100110",
  30225=>"010111111",
  30226=>"000000101",
  30227=>"000111111",
  30228=>"011011011",
  30229=>"000101111",
  30230=>"111111011",
  30231=>"111111001",
  30232=>"110111110",
  30233=>"100000000",
  30234=>"000111111",
  30235=>"111100100",
  30236=>"101101111",
  30237=>"111111111",
  30238=>"000000000",
  30239=>"000000010",
  30240=>"100000000",
  30241=>"000000111",
  30242=>"000000100",
  30243=>"111100110",
  30244=>"000111111",
  30245=>"000000001",
  30246=>"110111110",
  30247=>"100111000",
  30248=>"001000000",
  30249=>"000000000",
  30250=>"100000000",
  30251=>"011000011",
  30252=>"101111111",
  30253=>"000000000",
  30254=>"000000001",
  30255=>"000000000",
  30256=>"100111110",
  30257=>"001001111",
  30258=>"111111001",
  30259=>"011100100",
  30260=>"000000000",
  30261=>"000001111",
  30262=>"001000001",
  30263=>"001000011",
  30264=>"000000000",
  30265=>"000001001",
  30266=>"111111111",
  30267=>"111110000",
  30268=>"000000001",
  30269=>"000000000",
  30270=>"011000000",
  30271=>"111111111",
  30272=>"111111111",
  30273=>"110111111",
  30274=>"000010111",
  30275=>"000011000",
  30276=>"000001001",
  30277=>"000000100",
  30278=>"001111111",
  30279=>"111111110",
  30280=>"011011001",
  30281=>"011011010",
  30282=>"000000011",
  30283=>"000000101",
  30284=>"111110100",
  30285=>"100100110",
  30286=>"100100111",
  30287=>"111111111",
  30288=>"111111111",
  30289=>"110110000",
  30290=>"100001000",
  30291=>"000000000",
  30292=>"110110110",
  30293=>"010111111",
  30294=>"100000100",
  30295=>"000101111",
  30296=>"111000000",
  30297=>"000000111",
  30298=>"111011000",
  30299=>"000110110",
  30300=>"001001101",
  30301=>"000000000",
  30302=>"011010010",
  30303=>"111111011",
  30304=>"111000000",
  30305=>"000000011",
  30306=>"111111111",
  30307=>"110000010",
  30308=>"001001011",
  30309=>"000000000",
  30310=>"000000001",
  30311=>"000000110",
  30312=>"000011000",
  30313=>"000000011",
  30314=>"011000000",
  30315=>"111000100",
  30316=>"000001000",
  30317=>"000000000",
  30318=>"101001001",
  30319=>"000111000",
  30320=>"011000011",
  30321=>"011011111",
  30322=>"000000011",
  30323=>"111111010",
  30324=>"111111010",
  30325=>"010111011",
  30326=>"111111000",
  30327=>"000000000",
  30328=>"000000001",
  30329=>"101001011",
  30330=>"101001001",
  30331=>"000011111",
  30332=>"100000000",
  30333=>"000001001",
  30334=>"101000000",
  30335=>"000010000",
  30336=>"000100000",
  30337=>"111111110",
  30338=>"000001001",
  30339=>"001111000",
  30340=>"110111110",
  30341=>"000001000",
  30342=>"000000000",
  30343=>"000000000",
  30344=>"111110000",
  30345=>"011111111",
  30346=>"111111111",
  30347=>"111111111",
  30348=>"110111011",
  30349=>"000000000",
  30350=>"000010000",
  30351=>"110110110",
  30352=>"101101111",
  30353=>"011000000",
  30354=>"111111101",
  30355=>"010111111",
  30356=>"011111010",
  30357=>"111010111",
  30358=>"111111111",
  30359=>"000001001",
  30360=>"001001101",
  30361=>"100110110",
  30362=>"111111111",
  30363=>"111111111",
  30364=>"101000000",
  30365=>"111001011",
  30366=>"001011111",
  30367=>"000000000",
  30368=>"000000000",
  30369=>"100111001",
  30370=>"111111111",
  30371=>"000101111",
  30372=>"000000001",
  30373=>"111100100",
  30374=>"001111111",
  30375=>"000000000",
  30376=>"000000000",
  30377=>"000000011",
  30378=>"000000101",
  30379=>"100000000",
  30380=>"111111111",
  30381=>"111111001",
  30382=>"111111010",
  30383=>"000111110",
  30384=>"010001000",
  30385=>"001011000",
  30386=>"111111010",
  30387=>"010111011",
  30388=>"000000110",
  30389=>"000111110",
  30390=>"110111110",
  30391=>"001000001",
  30392=>"000000001",
  30393=>"000001001",
  30394=>"001011111",
  30395=>"111010011",
  30396=>"000000001",
  30397=>"111001111",
  30398=>"101001111",
  30399=>"000000001",
  30400=>"001000000",
  30401=>"000000000",
  30402=>"101000011",
  30403=>"000000010",
  30404=>"001001111",
  30405=>"000000000",
  30406=>"110110000",
  30407=>"110111110",
  30408=>"011111111",
  30409=>"111111111",
  30410=>"000000000",
  30411=>"000000001",
  30412=>"000100101",
  30413=>"000000000",
  30414=>"111001101",
  30415=>"000000111",
  30416=>"000000000",
  30417=>"000000110",
  30418=>"111111111",
  30419=>"111111111",
  30420=>"101111111",
  30421=>"000110010",
  30422=>"000000010",
  30423=>"111000000",
  30424=>"100110100",
  30425=>"110110000",
  30426=>"101000000",
  30427=>"000111111",
  30428=>"011011000",
  30429=>"111111010",
  30430=>"000000000",
  30431=>"001000111",
  30432=>"111011001",
  30433=>"111111111",
  30434=>"111111111",
  30435=>"000000000",
  30436=>"100100001",
  30437=>"011011011",
  30438=>"000010001",
  30439=>"011000000",
  30440=>"000001100",
  30441=>"000000110",
  30442=>"000000111",
  30443=>"011000100",
  30444=>"111100100",
  30445=>"111001000",
  30446=>"111000000",
  30447=>"000000000",
  30448=>"001000000",
  30449=>"111000000",
  30450=>"000111111",
  30451=>"001000111",
  30452=>"010001000",
  30453=>"110100100",
  30454=>"101001110",
  30455=>"000000000",
  30456=>"111111110",
  30457=>"111000000",
  30458=>"110111110",
  30459=>"110010010",
  30460=>"001100000",
  30461=>"110111110",
  30462=>"111111001",
  30463=>"000000000",
  30464=>"101000001",
  30465=>"100100100",
  30466=>"000000001",
  30467=>"111111000",
  30468=>"000000000",
  30469=>"110000000",
  30470=>"001111111",
  30471=>"110110110",
  30472=>"111111001",
  30473=>"000000001",
  30474=>"111111111",
  30475=>"011000000",
  30476=>"100000000",
  30477=>"100100111",
  30478=>"000000111",
  30479=>"111011011",
  30480=>"100111011",
  30481=>"111111111",
  30482=>"010110111",
  30483=>"000000000",
  30484=>"010111111",
  30485=>"000111111",
  30486=>"100110110",
  30487=>"000000000",
  30488=>"011011001",
  30489=>"111111001",
  30490=>"000000000",
  30491=>"111000000",
  30492=>"101001001",
  30493=>"101100000",
  30494=>"000000000",
  30495=>"111101111",
  30496=>"000000000",
  30497=>"111111000",
  30498=>"111111100",
  30499=>"000000010",
  30500=>"000001111",
  30501=>"011011111",
  30502=>"001111111",
  30503=>"111111011",
  30504=>"001110000",
  30505=>"000111111",
  30506=>"010010111",
  30507=>"110101000",
  30508=>"000000000",
  30509=>"111000110",
  30510=>"111111111",
  30511=>"000000100",
  30512=>"101000000",
  30513=>"000001101",
  30514=>"011000111",
  30515=>"000000001",
  30516=>"111010000",
  30517=>"101100100",
  30518=>"000000000",
  30519=>"001001000",
  30520=>"000000000",
  30521=>"000111000",
  30522=>"011001000",
  30523=>"111111111",
  30524=>"111001000",
  30525=>"000000000",
  30526=>"101000000",
  30527=>"100100000",
  30528=>"000000111",
  30529=>"111011000",
  30530=>"100111000",
  30531=>"110010000",
  30532=>"000010000",
  30533=>"001001000",
  30534=>"000111111",
  30535=>"000011011",
  30536=>"000000000",
  30537=>"010010111",
  30538=>"000000000",
  30539=>"000001001",
  30540=>"111011111",
  30541=>"000110111",
  30542=>"111111000",
  30543=>"000000000",
  30544=>"001000000",
  30545=>"000000111",
  30546=>"010000000",
  30547=>"000100111",
  30548=>"111111111",
  30549=>"001011000",
  30550=>"000000001",
  30551=>"111110110",
  30552=>"110111000",
  30553=>"000000111",
  30554=>"001000000",
  30555=>"111110100",
  30556=>"111011011",
  30557=>"111001001",
  30558=>"001001001",
  30559=>"111111111",
  30560=>"000000000",
  30561=>"111111111",
  30562=>"100010100",
  30563=>"100111010",
  30564=>"000011001",
  30565=>"101000001",
  30566=>"000100111",
  30567=>"111111011",
  30568=>"011001000",
  30569=>"000000000",
  30570=>"000000000",
  30571=>"000000100",
  30572=>"000000000",
  30573=>"110111101",
  30574=>"010111111",
  30575=>"111010000",
  30576=>"010001011",
  30577=>"111001001",
  30578=>"000000000",
  30579=>"001111110",
  30580=>"011111111",
  30581=>"011000000",
  30582=>"111100000",
  30583=>"110100100",
  30584=>"000000000",
  30585=>"111111011",
  30586=>"110111111",
  30587=>"111111000",
  30588=>"000001111",
  30589=>"001000000",
  30590=>"111111010",
  30591=>"000000001",
  30592=>"001001011",
  30593=>"011110111",
  30594=>"000001001",
  30595=>"100101011",
  30596=>"011000111",
  30597=>"010111010",
  30598=>"111111111",
  30599=>"000011000",
  30600=>"111111101",
  30601=>"111111011",
  30602=>"111111111",
  30603=>"000000111",
  30604=>"000000001",
  30605=>"110111110",
  30606=>"000000111",
  30607=>"000000000",
  30608=>"000111110",
  30609=>"000000000",
  30610=>"000001011",
  30611=>"001000000",
  30612=>"000000111",
  30613=>"010111111",
  30614=>"111101100",
  30615=>"000011111",
  30616=>"110111111",
  30617=>"111101001",
  30618=>"000000000",
  30619=>"000000000",
  30620=>"111111010",
  30621=>"101000000",
  30622=>"000000000",
  30623=>"000000111",
  30624=>"111111001",
  30625=>"110100100",
  30626=>"110111111",
  30627=>"000000000",
  30628=>"000111111",
  30629=>"000011111",
  30630=>"111111111",
  30631=>"111111111",
  30632=>"010000000",
  30633=>"000000000",
  30634=>"110000000",
  30635=>"011011111",
  30636=>"000100110",
  30637=>"110100111",
  30638=>"001001111",
  30639=>"000000001",
  30640=>"000000001",
  30641=>"111111111",
  30642=>"101001111",
  30643=>"000100100",
  30644=>"001001000",
  30645=>"000001101",
  30646=>"110111110",
  30647=>"000000000",
  30648=>"000000001",
  30649=>"111111111",
  30650=>"000000111",
  30651=>"001000000",
  30652=>"110110000",
  30653=>"000100111",
  30654=>"000000001",
  30655=>"011000000",
  30656=>"110111101",
  30657=>"111111111",
  30658=>"111111111",
  30659=>"111111011",
  30660=>"111111111",
  30661=>"011111001",
  30662=>"000100110",
  30663=>"000000000",
  30664=>"111111111",
  30665=>"100111111",
  30666=>"000000000",
  30667=>"110001011",
  30668=>"000000111",
  30669=>"001111000",
  30670=>"110110110",
  30671=>"000000000",
  30672=>"110000110",
  30673=>"000000000",
  30674=>"111000000",
  30675=>"000000001",
  30676=>"100100100",
  30677=>"101001101",
  30678=>"000010110",
  30679=>"011000000",
  30680=>"000000000",
  30681=>"000110000",
  30682=>"000001111",
  30683=>"111111010",
  30684=>"000000001",
  30685=>"000011011",
  30686=>"111000000",
  30687=>"000000100",
  30688=>"111111111",
  30689=>"111111100",
  30690=>"111110000",
  30691=>"000110000",
  30692=>"000000010",
  30693=>"111111011",
  30694=>"111011010",
  30695=>"000000000",
  30696=>"110110110",
  30697=>"111111111",
  30698=>"111110100",
  30699=>"110110010",
  30700=>"000000111",
  30701=>"010111111",
  30702=>"000001111",
  30703=>"111111111",
  30704=>"000000000",
  30705=>"010000000",
  30706=>"010111011",
  30707=>"101111000",
  30708=>"000000111",
  30709=>"000000000",
  30710=>"111111000",
  30711=>"011011011",
  30712=>"110111010",
  30713=>"101100000",
  30714=>"000111110",
  30715=>"000010111",
  30716=>"111111000",
  30717=>"110110011",
  30718=>"111111111",
  30719=>"000111111",
  30720=>"000000000",
  30721=>"000000101",
  30722=>"000000000",
  30723=>"011010100",
  30724=>"111110000",
  30725=>"100000100",
  30726=>"011111011",
  30727=>"111111111",
  30728=>"111111010",
  30729=>"101001000",
  30730=>"110000000",
  30731=>"111110010",
  30732=>"000000110",
  30733=>"111111111",
  30734=>"111111111",
  30735=>"111111111",
  30736=>"111111101",
  30737=>"000000000",
  30738=>"111111011",
  30739=>"111100100",
  30740=>"000000000",
  30741=>"000000000",
  30742=>"001001001",
  30743=>"011011011",
  30744=>"000000111",
  30745=>"010111111",
  30746=>"101000101",
  30747=>"000000100",
  30748=>"110111010",
  30749=>"111111000",
  30750=>"011001011",
  30751=>"111001001",
  30752=>"000100111",
  30753=>"111011000",
  30754=>"110110100",
  30755=>"111111101",
  30756=>"001000000",
  30757=>"111110110",
  30758=>"000001000",
  30759=>"000100111",
  30760=>"000000110",
  30761=>"100110111",
  30762=>"101101001",
  30763=>"100111111",
  30764=>"101111111",
  30765=>"000010111",
  30766=>"001111111",
  30767=>"000000000",
  30768=>"100100100",
  30769=>"001000000",
  30770=>"011000011",
  30771=>"110110100",
  30772=>"101101000",
  30773=>"111110100",
  30774=>"111111001",
  30775=>"010010000",
  30776=>"000000000",
  30777=>"000100100",
  30778=>"000110010",
  30779=>"111110110",
  30780=>"001101111",
  30781=>"000000000",
  30782=>"000000000",
  30783=>"000000000",
  30784=>"000000111",
  30785=>"000101100",
  30786=>"111111111",
  30787=>"100100000",
  30788=>"000000110",
  30789=>"001001111",
  30790=>"011111000",
  30791=>"110000000",
  30792=>"001001011",
  30793=>"000111111",
  30794=>"000000000",
  30795=>"111111111",
  30796=>"000010111",
  30797=>"101101001",
  30798=>"101011111",
  30799=>"111111011",
  30800=>"000000000",
  30801=>"000001000",
  30802=>"000111111",
  30803=>"011001000",
  30804=>"101100000",
  30805=>"000001111",
  30806=>"110111001",
  30807=>"000000000",
  30808=>"111111110",
  30809=>"000000111",
  30810=>"101000000",
  30811=>"110001001",
  30812=>"010000000",
  30813=>"000000000",
  30814=>"101000000",
  30815=>"111100100",
  30816=>"000001111",
  30817=>"101111111",
  30818=>"000010100",
  30819=>"111101111",
  30820=>"111111110",
  30821=>"111111111",
  30822=>"111111110",
  30823=>"111101101",
  30824=>"000000000",
  30825=>"000000000",
  30826=>"000000000",
  30827=>"011010000",
  30828=>"000000110",
  30829=>"000000100",
  30830=>"001000000",
  30831=>"000000001",
  30832=>"110110110",
  30833=>"100111111",
  30834=>"110111010",
  30835=>"111111101",
  30836=>"000000000",
  30837=>"100111010",
  30838=>"000000110",
  30839=>"000000000",
  30840=>"111000110",
  30841=>"111100000",
  30842=>"111101101",
  30843=>"100001001",
  30844=>"001001011",
  30845=>"110110110",
  30846=>"111111011",
  30847=>"011111111",
  30848=>"010000000",
  30849=>"000000000",
  30850=>"111111111",
  30851=>"111111111",
  30852=>"111111000",
  30853=>"000010111",
  30854=>"000000000",
  30855=>"011000000",
  30856=>"111111010",
  30857=>"000100000",
  30858=>"010010010",
  30859=>"111111111",
  30860=>"000000100",
  30861=>"100111111",
  30862=>"001010000",
  30863=>"000000000",
  30864=>"111111111",
  30865=>"111111111",
  30866=>"100100000",
  30867=>"111000000",
  30868=>"000110110",
  30869=>"111111111",
  30870=>"111111101",
  30871=>"000000000",
  30872=>"100000000",
  30873=>"111111111",
  30874=>"111111110",
  30875=>"111111111",
  30876=>"000110001",
  30877=>"101001111",
  30878=>"010010000",
  30879=>"000111010",
  30880=>"000010000",
  30881=>"001100111",
  30882=>"011000010",
  30883=>"101100100",
  30884=>"110000011",
  30885=>"011111111",
  30886=>"000010111",
  30887=>"010011010",
  30888=>"000000000",
  30889=>"000101111",
  30890=>"000010010",
  30891=>"111111111",
  30892=>"111111000",
  30893=>"111011011",
  30894=>"111111111",
  30895=>"000000000",
  30896=>"000100100",
  30897=>"111110111",
  30898=>"000010010",
  30899=>"100111111",
  30900=>"000000000",
  30901=>"110110000",
  30902=>"011111111",
  30903=>"100110000",
  30904=>"111111110",
  30905=>"000110000",
  30906=>"111000001",
  30907=>"011000101",
  30908=>"100100000",
  30909=>"110110110",
  30910=>"110000000",
  30911=>"111110110",
  30912=>"111110000",
  30913=>"000000000",
  30914=>"010110110",
  30915=>"101101011",
  30916=>"000000010",
  30917=>"110110010",
  30918=>"111111111",
  30919=>"000100111",
  30920=>"000000000",
  30921=>"000000000",
  30922=>"100001101",
  30923=>"011000000",
  30924=>"010010000",
  30925=>"011111111",
  30926=>"001111111",
  30927=>"010010000",
  30928=>"000000110",
  30929=>"000000100",
  30930=>"111000100",
  30931=>"100100000",
  30932=>"111111110",
  30933=>"111110110",
  30934=>"111100111",
  30935=>"000000110",
  30936=>"000000000",
  30937=>"111111011",
  30938=>"000000000",
  30939=>"010000111",
  30940=>"111110100",
  30941=>"000000011",
  30942=>"000100110",
  30943=>"010010000",
  30944=>"000000111",
  30945=>"100111011",
  30946=>"111110111",
  30947=>"000000000",
  30948=>"110111101",
  30949=>"011000000",
  30950=>"110111111",
  30951=>"111111111",
  30952=>"100100000",
  30953=>"111111011",
  30954=>"111101101",
  30955=>"000000000",
  30956=>"000010111",
  30957=>"111111111",
  30958=>"011001111",
  30959=>"011000100",
  30960=>"011011001",
  30961=>"011111111",
  30962=>"000111111",
  30963=>"010011011",
  30964=>"101100001",
  30965=>"110000000",
  30966=>"101100111",
  30967=>"101101111",
  30968=>"000000001",
  30969=>"000000101",
  30970=>"000001000",
  30971=>"111111110",
  30972=>"000000000",
  30973=>"000001111",
  30974=>"001111001",
  30975=>"000000000",
  30976=>"010101111",
  30977=>"110100100",
  30978=>"111111111",
  30979=>"100100111",
  30980=>"000001001",
  30981=>"000000000",
  30982=>"111111011",
  30983=>"000000011",
  30984=>"111111000",
  30985=>"111111110",
  30986=>"001101101",
  30987=>"111101011",
  30988=>"000100100",
  30989=>"000111011",
  30990=>"010110110",
  30991=>"111111000",
  30992=>"111111001",
  30993=>"000111111",
  30994=>"100100111",
  30995=>"111111111",
  30996=>"010000000",
  30997=>"011111111",
  30998=>"111111001",
  30999=>"011100000",
  31000=>"111111111",
  31001=>"000000000",
  31002=>"111111000",
  31003=>"000000000",
  31004=>"111110110",
  31005=>"111111111",
  31006=>"000000000",
  31007=>"111111111",
  31008=>"000000011",
  31009=>"111110111",
  31010=>"000000001",
  31011=>"111111111",
  31012=>"111001000",
  31013=>"000001000",
  31014=>"000011000",
  31015=>"100100000",
  31016=>"111000000",
  31017=>"000000000",
  31018=>"000000000",
  31019=>"000000001",
  31020=>"010001000",
  31021=>"100000000",
  31022=>"111111111",
  31023=>"111100000",
  31024=>"011001001",
  31025=>"111111001",
  31026=>"000000000",
  31027=>"000000000",
  31028=>"000101100",
  31029=>"110100110",
  31030=>"100111111",
  31031=>"110111111",
  31032=>"001000111",
  31033=>"110111011",
  31034=>"111111011",
  31035=>"101001111",
  31036=>"000001001",
  31037=>"000000000",
  31038=>"011011111",
  31039=>"011000111",
  31040=>"001001111",
  31041=>"110111111",
  31042=>"111101100",
  31043=>"000001001",
  31044=>"111011000",
  31045=>"111111010",
  31046=>"000000000",
  31047=>"111011000",
  31048=>"111111111",
  31049=>"001110110",
  31050=>"000000010",
  31051=>"111110100",
  31052=>"000000000",
  31053=>"000000111",
  31054=>"111001000",
  31055=>"011011001",
  31056=>"001110111",
  31057=>"110110000",
  31058=>"000000110",
  31059=>"111111111",
  31060=>"000000001",
  31061=>"001000111",
  31062=>"000111100",
  31063=>"111111111",
  31064=>"011111111",
  31065=>"110000001",
  31066=>"100100100",
  31067=>"000101111",
  31068=>"100000100",
  31069=>"100000101",
  31070=>"111011111",
  31071=>"000000110",
  31072=>"100011111",
  31073=>"111101001",
  31074=>"111111111",
  31075=>"101001011",
  31076=>"110110110",
  31077=>"111001101",
  31078=>"100000000",
  31079=>"100000001",
  31080=>"110011000",
  31081=>"000111111",
  31082=>"001000011",
  31083=>"101101111",
  31084=>"011011001",
  31085=>"110101001",
  31086=>"000000000",
  31087=>"000000001",
  31088=>"011000101",
  31089=>"101000000",
  31090=>"110110000",
  31091=>"011011001",
  31092=>"000000001",
  31093=>"111111111",
  31094=>"011001011",
  31095=>"001011111",
  31096=>"001001001",
  31097=>"000000000",
  31098=>"110110111",
  31099=>"000000000",
  31100=>"011101111",
  31101=>"010111111",
  31102=>"101111101",
  31103=>"111111111",
  31104=>"000000001",
  31105=>"111111111",
  31106=>"000000000",
  31107=>"101000000",
  31108=>"000000100",
  31109=>"000000100",
  31110=>"111011011",
  31111=>"100100100",
  31112=>"111011111",
  31113=>"000010110",
  31114=>"111111101",
  31115=>"000001101",
  31116=>"111111111",
  31117=>"000010010",
  31118=>"111111000",
  31119=>"010011010",
  31120=>"101101111",
  31121=>"000000000",
  31122=>"101000000",
  31123=>"000000000",
  31124=>"101000000",
  31125=>"001000000",
  31126=>"000000100",
  31127=>"110110110",
  31128=>"000000100",
  31129=>"101001001",
  31130=>"011111111",
  31131=>"110111010",
  31132=>"111110100",
  31133=>"110000111",
  31134=>"111000000",
  31135=>"100110110",
  31136=>"001001001",
  31137=>"110100110",
  31138=>"000111011",
  31139=>"000000000",
  31140=>"000000011",
  31141=>"111111111",
  31142=>"000000101",
  31143=>"111111111",
  31144=>"000110000",
  31145=>"000000111",
  31146=>"010110110",
  31147=>"111111110",
  31148=>"111101101",
  31149=>"000100101",
  31150=>"011011101",
  31151=>"000000011",
  31152=>"111111100",
  31153=>"100001111",
  31154=>"000111000",
  31155=>"000001000",
  31156=>"000000000",
  31157=>"110000101",
  31158=>"111111111",
  31159=>"000000000",
  31160=>"000000110",
  31161=>"111101011",
  31162=>"000000000",
  31163=>"110010000",
  31164=>"000000111",
  31165=>"111111000",
  31166=>"111111010",
  31167=>"010010010",
  31168=>"101111111",
  31169=>"100111111",
  31170=>"000000000",
  31171=>"110000000",
  31172=>"000001000",
  31173=>"001011011",
  31174=>"100000000",
  31175=>"100000000",
  31176=>"110101111",
  31177=>"000000111",
  31178=>"110100100",
  31179=>"111111111",
  31180=>"000111110",
  31181=>"010010000",
  31182=>"000000001",
  31183=>"111011111",
  31184=>"001111111",
  31185=>"001011100",
  31186=>"011011111",
  31187=>"011111111",
  31188=>"000000010",
  31189=>"100100100",
  31190=>"101100100",
  31191=>"011111011",
  31192=>"000100100",
  31193=>"101101111",
  31194=>"111111111",
  31195=>"010000010",
  31196=>"111000000",
  31197=>"000011111",
  31198=>"111101111",
  31199=>"000000011",
  31200=>"000100110",
  31201=>"010000000",
  31202=>"001111111",
  31203=>"011000000",
  31204=>"000000111",
  31205=>"001001101",
  31206=>"111111110",
  31207=>"100100101",
  31208=>"000000000",
  31209=>"001101111",
  31210=>"000001101",
  31211=>"000000011",
  31212=>"110111111",
  31213=>"011001011",
  31214=>"000000000",
  31215=>"000000000",
  31216=>"001000000",
  31217=>"001111111",
  31218=>"100000000",
  31219=>"000000000",
  31220=>"111011000",
  31221=>"111111111",
  31222=>"000101001",
  31223=>"011000001",
  31224=>"000100111",
  31225=>"010010110",
  31226=>"111001101",
  31227=>"000000000",
  31228=>"000000000",
  31229=>"110110110",
  31230=>"110111000",
  31231=>"110100110",
  31232=>"000000000",
  31233=>"000000000",
  31234=>"111111111",
  31235=>"100000001",
  31236=>"001000000",
  31237=>"110000010",
  31238=>"001111111",
  31239=>"111111111",
  31240=>"111111111",
  31241=>"000000000",
  31242=>"111111111",
  31243=>"111111111",
  31244=>"000100000",
  31245=>"000000000",
  31246=>"011011000",
  31247=>"001111111",
  31248=>"111111001",
  31249=>"001000000",
  31250=>"101111111",
  31251=>"001001001",
  31252=>"111101111",
  31253=>"000000000",
  31254=>"111110000",
  31255=>"011111111",
  31256=>"011111111",
  31257=>"110111101",
  31258=>"011011110",
  31259=>"100000000",
  31260=>"000000000",
  31261=>"110111111",
  31262=>"001001001",
  31263=>"111111011",
  31264=>"011001011",
  31265=>"000011011",
  31266=>"011011011",
  31267=>"000000111",
  31268=>"111111111",
  31269=>"111111111",
  31270=>"011011000",
  31271=>"000100000",
  31272=>"111111010",
  31273=>"000000000",
  31274=>"000011111",
  31275=>"001000000",
  31276=>"110111111",
  31277=>"000000101",
  31278=>"100001010",
  31279=>"000111111",
  31280=>"000110111",
  31281=>"100100000",
  31282=>"000000000",
  31283=>"011101110",
  31284=>"000000011",
  31285=>"111111111",
  31286=>"000111111",
  31287=>"011011111",
  31288=>"111111000",
  31289=>"011000000",
  31290=>"000010000",
  31291=>"111011011",
  31292=>"111111111",
  31293=>"001000000",
  31294=>"010111011",
  31295=>"000000000",
  31296=>"101001000",
  31297=>"100100100",
  31298=>"000100110",
  31299=>"000000000",
  31300=>"000000000",
  31301=>"110111111",
  31302=>"000000000",
  31303=>"111110110",
  31304=>"010001001",
  31305=>"111111111",
  31306=>"000000101",
  31307=>"111111111",
  31308=>"000000000",
  31309=>"001000000",
  31310=>"100000000",
  31311=>"101111000",
  31312=>"001111011",
  31313=>"100110110",
  31314=>"111001000",
  31315=>"110100000",
  31316=>"111000110",
  31317=>"111111001",
  31318=>"000000000",
  31319=>"110111111",
  31320=>"011001101",
  31321=>"110100000",
  31322=>"000000111",
  31323=>"111001001",
  31324=>"101000000",
  31325=>"111110111",
  31326=>"001001001",
  31327=>"000110111",
  31328=>"111111111",
  31329=>"000000000",
  31330=>"001001000",
  31331=>"101111111",
  31332=>"111000000",
  31333=>"001001101",
  31334=>"010110001",
  31335=>"011000101",
  31336=>"111101001",
  31337=>"010000000",
  31338=>"110010000",
  31339=>"000000001",
  31340=>"000000000",
  31341=>"011000111",
  31342=>"111111000",
  31343=>"111111111",
  31344=>"000000000",
  31345=>"111111111",
  31346=>"100000000",
  31347=>"001011011",
  31348=>"111110110",
  31349=>"111111111",
  31350=>"111111000",
  31351=>"100101011",
  31352=>"111111101",
  31353=>"000000000",
  31354=>"111111111",
  31355=>"111111111",
  31356=>"000100111",
  31357=>"001000000",
  31358=>"111111111",
  31359=>"111111111",
  31360=>"000000111",
  31361=>"000000000",
  31362=>"000000000",
  31363=>"000000000",
  31364=>"110000100",
  31365=>"000000000",
  31366=>"111111111",
  31367=>"010111111",
  31368=>"000000100",
  31369=>"111111111",
  31370=>"111110100",
  31371=>"111000001",
  31372=>"000100110",
  31373=>"111111111",
  31374=>"000000110",
  31375=>"000000000",
  31376=>"000000000",
  31377=>"111111111",
  31378=>"000000001",
  31379=>"111111011",
  31380=>"000111111",
  31381=>"110000000",
  31382=>"111111111",
  31383=>"000000000",
  31384=>"111111011",
  31385=>"111111111",
  31386=>"000000000",
  31387=>"100111111",
  31388=>"111111111",
  31389=>"000000000",
  31390=>"000010111",
  31391=>"000000000",
  31392=>"101101000",
  31393=>"000000000",
  31394=>"111111111",
  31395=>"000001000",
  31396=>"000000110",
  31397=>"111101001",
  31398=>"110111110",
  31399=>"110000000",
  31400=>"001111100",
  31401=>"111111111",
  31402=>"000000000",
  31403=>"111111111",
  31404=>"011010000",
  31405=>"011011001",
  31406=>"110111111",
  31407=>"111111111",
  31408=>"110111000",
  31409=>"111111101",
  31410=>"000100000",
  31411=>"010111110",
  31412=>"001000110",
  31413=>"101000001",
  31414=>"000000000",
  31415=>"000101101",
  31416=>"000000000",
  31417=>"000111111",
  31418=>"000011011",
  31419=>"011111011",
  31420=>"000100000",
  31421=>"000000000",
  31422=>"111000111",
  31423=>"001000001",
  31424=>"110110110",
  31425=>"000000001",
  31426=>"101111111",
  31427=>"111111000",
  31428=>"000000000",
  31429=>"111111111",
  31430=>"110111011",
  31431=>"010111111",
  31432=>"111110010",
  31433=>"000000000",
  31434=>"000000000",
  31435=>"000110110",
  31436=>"010000000",
  31437=>"110110100",
  31438=>"100100000",
  31439=>"111100000",
  31440=>"111111111",
  31441=>"001111010",
  31442=>"111111111",
  31443=>"001001000",
  31444=>"111111000",
  31445=>"011111110",
  31446=>"111111111",
  31447=>"111100000",
  31448=>"111111111",
  31449=>"001001000",
  31450=>"000000000",
  31451=>"010010000",
  31452=>"111100101",
  31453=>"010000000",
  31454=>"000000100",
  31455=>"000000000",
  31456=>"000000000",
  31457=>"000101101",
  31458=>"111101101",
  31459=>"000011001",
  31460=>"111111100",
  31461=>"111001000",
  31462=>"000000000",
  31463=>"011010000",
  31464=>"110000000",
  31465=>"000000000",
  31466=>"111000000",
  31467=>"000000011",
  31468=>"000000010",
  31469=>"101000111",
  31470=>"000100100",
  31471=>"111111000",
  31472=>"011011110",
  31473=>"001001100",
  31474=>"000110111",
  31475=>"001011000",
  31476=>"001000000",
  31477=>"111111100",
  31478=>"111100110",
  31479=>"111110010",
  31480=>"010000000",
  31481=>"110110110",
  31482=>"111111111",
  31483=>"110000000",
  31484=>"111111110",
  31485=>"000000000",
  31486=>"111111000",
  31487=>"111000000",
  31488=>"010111111",
  31489=>"011010010",
  31490=>"000110000",
  31491=>"111111111",
  31492=>"011111011",
  31493=>"011001111",
  31494=>"000000000",
  31495=>"000111111",
  31496=>"001011010",
  31497=>"000000000",
  31498=>"000010000",
  31499=>"111111010",
  31500=>"100110110",
  31501=>"000010000",
  31502=>"111111111",
  31503=>"110100000",
  31504=>"111000000",
  31505=>"000111111",
  31506=>"111111111",
  31507=>"110000000",
  31508=>"011001011",
  31509=>"000111111",
  31510=>"010010000",
  31511=>"001000000",
  31512=>"000000000",
  31513=>"111011111",
  31514=>"000000111",
  31515=>"000000000",
  31516=>"110110000",
  31517=>"000001111",
  31518=>"111111111",
  31519=>"100100111",
  31520=>"000100111",
  31521=>"000000000",
  31522=>"000111100",
  31523=>"110100110",
  31524=>"001011111",
  31525=>"000000100",
  31526=>"000011011",
  31527=>"001001000",
  31528=>"000010111",
  31529=>"011111111",
  31530=>"011000000",
  31531=>"011001011",
  31532=>"111111111",
  31533=>"011111110",
  31534=>"111111111",
  31535=>"000000000",
  31536=>"111111111",
  31537=>"000000001",
  31538=>"011111111",
  31539=>"111111111",
  31540=>"111100100",
  31541=>"000000011",
  31542=>"110111110",
  31543=>"101111111",
  31544=>"000111111",
  31545=>"011011000",
  31546=>"000000010",
  31547=>"110111011",
  31548=>"000111110",
  31549=>"000000000",
  31550=>"111011011",
  31551=>"000000111",
  31552=>"011011001",
  31553=>"000000000",
  31554=>"111111111",
  31555=>"111000000",
  31556=>"000000000",
  31557=>"111010000",
  31558=>"000000000",
  31559=>"111111111",
  31560=>"111100100",
  31561=>"101101101",
  31562=>"111000000",
  31563=>"100100100",
  31564=>"000001000",
  31565=>"110110100",
  31566=>"000000000",
  31567=>"111110110",
  31568=>"111110000",
  31569=>"000000000",
  31570=>"000000000",
  31571=>"000001001",
  31572=>"000000000",
  31573=>"000011111",
  31574=>"100111001",
  31575=>"000001001",
  31576=>"100111000",
  31577=>"001111111",
  31578=>"111111111",
  31579=>"000000000",
  31580=>"011111001",
  31581=>"001001111",
  31582=>"111001000",
  31583=>"111111111",
  31584=>"111111111",
  31585=>"000010000",
  31586=>"100100101",
  31587=>"000000000",
  31588=>"000000110",
  31589=>"000000000",
  31590=>"111111111",
  31591=>"000010000",
  31592=>"011000000",
  31593=>"010000000",
  31594=>"011111010",
  31595=>"000000111",
  31596=>"101001111",
  31597=>"000000000",
  31598=>"110111111",
  31599=>"011111001",
  31600=>"000001011",
  31601=>"111001101",
  31602=>"000000110",
  31603=>"010011111",
  31604=>"000100000",
  31605=>"010011111",
  31606=>"111111001",
  31607=>"111101111",
  31608=>"000000001",
  31609=>"111111100",
  31610=>"111111111",
  31611=>"000010011",
  31612=>"101111101",
  31613=>"111111111",
  31614=>"111111111",
  31615=>"000000111",
  31616=>"000000000",
  31617=>"111111111",
  31618=>"011111111",
  31619=>"111111101",
  31620=>"111111000",
  31621=>"000000000",
  31622=>"000000010",
  31623=>"100100100",
  31624=>"111000000",
  31625=>"001011111",
  31626=>"100110000",
  31627=>"111111111",
  31628=>"101000111",
  31629=>"011000000",
  31630=>"000011000",
  31631=>"000000001",
  31632=>"100100100",
  31633=>"000000000",
  31634=>"110100110",
  31635=>"000110100",
  31636=>"000000001",
  31637=>"111110101",
  31638=>"111011001",
  31639=>"000000000",
  31640=>"111111111",
  31641=>"000000001",
  31642=>"001011000",
  31643=>"000110111",
  31644=>"010010011",
  31645=>"111000000",
  31646=>"111111111",
  31647=>"111100000",
  31648=>"000001111",
  31649=>"011011001",
  31650=>"000000100",
  31651=>"011010000",
  31652=>"011111111",
  31653=>"111111111",
  31654=>"111100101",
  31655=>"000000000",
  31656=>"000100111",
  31657=>"000001001",
  31658=>"000000000",
  31659=>"000000010",
  31660=>"111111111",
  31661=>"111000000",
  31662=>"000000000",
  31663=>"000001101",
  31664=>"111011011",
  31665=>"111111111",
  31666=>"001000000",
  31667=>"111111111",
  31668=>"001011111",
  31669=>"111111110",
  31670=>"111011001",
  31671=>"101100001",
  31672=>"111111100",
  31673=>"111111111",
  31674=>"100110111",
  31675=>"001000011",
  31676=>"000000000",
  31677=>"101000001",
  31678=>"010010010",
  31679=>"011011011",
  31680=>"000000001",
  31681=>"011001000",
  31682=>"000000000",
  31683=>"000000000",
  31684=>"001011111",
  31685=>"000000000",
  31686=>"000100110",
  31687=>"000010000",
  31688=>"001011010",
  31689=>"110110111",
  31690=>"111101111",
  31691=>"000000000",
  31692=>"111111111",
  31693=>"000000000",
  31694=>"000000000",
  31695=>"111111111",
  31696=>"000001101",
  31697=>"010011001",
  31698=>"000000110",
  31699=>"000000000",
  31700=>"001011011",
  31701=>"110110111",
  31702=>"111101101",
  31703=>"000000000",
  31704=>"111111111",
  31705=>"111001001",
  31706=>"000100100",
  31707=>"010011111",
  31708=>"111111011",
  31709=>"000000000",
  31710=>"111110111",
  31711=>"011111011",
  31712=>"000000000",
  31713=>"111111011",
  31714=>"000000000",
  31715=>"111111001",
  31716=>"000000110",
  31717=>"111101111",
  31718=>"111111011",
  31719=>"111111111",
  31720=>"000000010",
  31721=>"000000010",
  31722=>"001000000",
  31723=>"111011000",
  31724=>"011100101",
  31725=>"100100100",
  31726=>"000111111",
  31727=>"000000000",
  31728=>"000000000",
  31729=>"000101111",
  31730=>"111011111",
  31731=>"000000000",
  31732=>"000000100",
  31733=>"111111111",
  31734=>"000011011",
  31735=>"111111111",
  31736=>"010010001",
  31737=>"000110110",
  31738=>"111001011",
  31739=>"000000000",
  31740=>"111111111",
  31741=>"100111111",
  31742=>"110111111",
  31743=>"110111111",
  31744=>"111111111",
  31745=>"000000111",
  31746=>"111000001",
  31747=>"000000000",
  31748=>"000000000",
  31749=>"101101101",
  31750=>"110111010",
  31751=>"111111111",
  31752=>"001000111",
  31753=>"100110110",
  31754=>"100000000",
  31755=>"111110101",
  31756=>"110110110",
  31757=>"000000000",
  31758=>"001011011",
  31759=>"000000000",
  31760=>"000111111",
  31761=>"000111101",
  31762=>"000000000",
  31763=>"111000000",
  31764=>"111000000",
  31765=>"011011001",
  31766=>"110000001",
  31767=>"111111000",
  31768=>"000000100",
  31769=>"110010000",
  31770=>"001001000",
  31771=>"100100110",
  31772=>"111111111",
  31773=>"000101111",
  31774=>"100100110",
  31775=>"100100000",
  31776=>"000101111",
  31777=>"110000000",
  31778=>"000000000",
  31779=>"111111111",
  31780=>"111111111",
  31781=>"111110110",
  31782=>"000000000",
  31783=>"000000000",
  31784=>"000010111",
  31785=>"111111000",
  31786=>"000001000",
  31787=>"000000000",
  31788=>"100111111",
  31789=>"000111111",
  31790=>"101100000",
  31791=>"100000000",
  31792=>"001100000",
  31793=>"000000000",
  31794=>"011000000",
  31795=>"000000100",
  31796=>"000110111",
  31797=>"001001011",
  31798=>"111111111",
  31799=>"000100110",
  31800=>"011011100",
  31801=>"000000001",
  31802=>"000010010",
  31803=>"000101111",
  31804=>"101000000",
  31805=>"111011001",
  31806=>"110111110",
  31807=>"001001111",
  31808=>"000000011",
  31809=>"100000000",
  31810=>"010010010",
  31811=>"000111111",
  31812=>"111001000",
  31813=>"111111000",
  31814=>"011011111",
  31815=>"000000000",
  31816=>"011111111",
  31817=>"111111111",
  31818=>"000000000",
  31819=>"001000001",
  31820=>"001101111",
  31821=>"101000000",
  31822=>"011011111",
  31823=>"010010010",
  31824=>"011001111",
  31825=>"010000000",
  31826=>"111011000",
  31827=>"010110110",
  31828=>"001000000",
  31829=>"111111110",
  31830=>"000000000",
  31831=>"111111110",
  31832=>"000000100",
  31833=>"101000101",
  31834=>"111111111",
  31835=>"111000110",
  31836=>"111111111",
  31837=>"101000000",
  31838=>"011111111",
  31839=>"111011011",
  31840=>"000000111",
  31841=>"000000000",
  31842=>"000000000",
  31843=>"111111111",
  31844=>"111011000",
  31845=>"101111111",
  31846=>"011111111",
  31847=>"111110000",
  31848=>"111110000",
  31849=>"000001001",
  31850=>"000000000",
  31851=>"101101111",
  31852=>"010111111",
  31853=>"001000101",
  31854=>"001000111",
  31855=>"111110111",
  31856=>"111001011",
  31857=>"111110101",
  31858=>"111110000",
  31859=>"111111010",
  31860=>"111011010",
  31861=>"110111110",
  31862=>"000000000",
  31863=>"010111100",
  31864=>"101101100",
  31865=>"101001011",
  31866=>"111100100",
  31867=>"011000000",
  31868=>"001000101",
  31869=>"111001000",
  31870=>"110000000",
  31871=>"111111101",
  31872=>"000111010",
  31873=>"011011000",
  31874=>"111111111",
  31875=>"001101000",
  31876=>"000100100",
  31877=>"101101111",
  31878=>"111111001",
  31879=>"000000000",
  31880=>"000110111",
  31881=>"001000000",
  31882=>"100000000",
  31883=>"111111010",
  31884=>"000000101",
  31885=>"001001001",
  31886=>"010000000",
  31887=>"111111111",
  31888=>"101001001",
  31889=>"110011010",
  31890=>"011110010",
  31891=>"111111111",
  31892=>"000000000",
  31893=>"011111111",
  31894=>"110111010",
  31895=>"000000111",
  31896=>"000000000",
  31897=>"010000111",
  31898=>"011011101",
  31899=>"000000000",
  31900=>"000000000",
  31901=>"101000000",
  31902=>"001001111",
  31903=>"000000000",
  31904=>"111011000",
  31905=>"000001000",
  31906=>"110000110",
  31907=>"111111111",
  31908=>"100000101",
  31909=>"000110111",
  31910=>"101101101",
  31911=>"111100000",
  31912=>"000000000",
  31913=>"101000000",
  31914=>"010011000",
  31915=>"111110000",
  31916=>"011000000",
  31917=>"100101111",
  31918=>"101101111",
  31919=>"000000001",
  31920=>"000010000",
  31921=>"111111011",
  31922=>"111111110",
  31923=>"111111000",
  31924=>"111110000",
  31925=>"111111111",
  31926=>"000111111",
  31927=>"010111111",
  31928=>"110111110",
  31929=>"011011111",
  31930=>"101000000",
  31931=>"100010110",
  31932=>"110111011",
  31933=>"000000000",
  31934=>"000010111",
  31935=>"000000000",
  31936=>"101000000",
  31937=>"001000000",
  31938=>"111111111",
  31939=>"111111111",
  31940=>"000011001",
  31941=>"000000111",
  31942=>"000000100",
  31943=>"111101101",
  31944=>"100111001",
  31945=>"000000001",
  31946=>"000000100",
  31947=>"001000000",
  31948=>"000000111",
  31949=>"111001001",
  31950=>"000111111",
  31951=>"000000010",
  31952=>"000001111",
  31953=>"101000001",
  31954=>"000100110",
  31955=>"110111110",
  31956=>"011101111",
  31957=>"111111111",
  31958=>"101000000",
  31959=>"111011011",
  31960=>"101101000",
  31961=>"110111110",
  31962=>"000000110",
  31963=>"001000000",
  31964=>"001001000",
  31965=>"111000000",
  31966=>"111101101",
  31967=>"010010000",
  31968=>"000000000",
  31969=>"000000000",
  31970=>"101101001",
  31971=>"000000001",
  31972=>"110111100",
  31973=>"110000110",
  31974=>"010010010",
  31975=>"111110110",
  31976=>"111111111",
  31977=>"101001001",
  31978=>"000000000",
  31979=>"000011110",
  31980=>"101000000",
  31981=>"001001001",
  31982=>"111100000",
  31983=>"111111111",
  31984=>"011001100",
  31985=>"111000000",
  31986=>"110000110",
  31987=>"111010000",
  31988=>"010000000",
  31989=>"111100100",
  31990=>"111110010",
  31991=>"000000000",
  31992=>"111111111",
  31993=>"000000000",
  31994=>"000000000",
  31995=>"111111111",
  31996=>"011111011",
  31997=>"110110110",
  31998=>"011000000",
  31999=>"111111110",
  32000=>"100000000",
  32001=>"111101101",
  32002=>"001000000",
  32003=>"111111110",
  32004=>"011000000",
  32005=>"101110000",
  32006=>"111111111",
  32007=>"000000111",
  32008=>"011111111",
  32009=>"111110111",
  32010=>"111110101",
  32011=>"111111110",
  32012=>"001000000",
  32013=>"111110000",
  32014=>"011000000",
  32015=>"100000000",
  32016=>"111111111",
  32017=>"000000000",
  32018=>"000000000",
  32019=>"101100100",
  32020=>"011111111",
  32021=>"111111111",
  32022=>"111111100",
  32023=>"111111111",
  32024=>"111101111",
  32025=>"101000000",
  32026=>"000000000",
  32027=>"010000000",
  32028=>"100100111",
  32029=>"000001000",
  32030=>"010000000",
  32031=>"111011001",
  32032=>"011011000",
  32033=>"100110111",
  32034=>"010000010",
  32035=>"000100110",
  32036=>"011001011",
  32037=>"000000111",
  32038=>"010111111",
  32039=>"100000000",
  32040=>"000100100",
  32041=>"000000100",
  32042=>"000000101",
  32043=>"111001000",
  32044=>"000010110",
  32045=>"001111111",
  32046=>"111100101",
  32047=>"000000000",
  32048=>"100100111",
  32049=>"011000000",
  32050=>"111111111",
  32051=>"000100000",
  32052=>"111101001",
  32053=>"100111111",
  32054=>"001100000",
  32055=>"111001001",
  32056=>"000000000",
  32057=>"111111111",
  32058=>"110110110",
  32059=>"000000000",
  32060=>"000111111",
  32061=>"000000000",
  32062=>"110110110",
  32063=>"110110110",
  32064=>"111111001",
  32065=>"100000101",
  32066=>"111111111",
  32067=>"001111111",
  32068=>"000001001",
  32069=>"011111111",
  32070=>"110110000",
  32071=>"110000000",
  32072=>"111000001",
  32073=>"101100111",
  32074=>"000110110",
  32075=>"111111110",
  32076=>"111000111",
  32077=>"000100111",
  32078=>"000101111",
  32079=>"000110110",
  32080=>"000000000",
  32081=>"000110111",
  32082=>"110111110",
  32083=>"011111111",
  32084=>"000111111",
  32085=>"011011011",
  32086=>"000110000",
  32087=>"100100100",
  32088=>"000010000",
  32089=>"011111111",
  32090=>"000000000",
  32091=>"000000000",
  32092=>"001011011",
  32093=>"000000100",
  32094=>"000110110",
  32095=>"111110111",
  32096=>"111111101",
  32097=>"111001001",
  32098=>"110011011",
  32099=>"111001000",
  32100=>"000000000",
  32101=>"010110000",
  32102=>"000000111",
  32103=>"111111111",
  32104=>"100111111",
  32105=>"111001001",
  32106=>"011001111",
  32107=>"000000000",
  32108=>"100111111",
  32109=>"111111111",
  32110=>"111000000",
  32111=>"001010111",
  32112=>"111000111",
  32113=>"111111011",
  32114=>"111010111",
  32115=>"111101000",
  32116=>"010110010",
  32117=>"111111111",
  32118=>"000000000",
  32119=>"111110110",
  32120=>"111111011",
  32121=>"000011011",
  32122=>"110100000",
  32123=>"001001000",
  32124=>"110000000",
  32125=>"011110111",
  32126=>"000000000",
  32127=>"000000000",
  32128=>"000000110",
  32129=>"001111111",
  32130=>"111110110",
  32131=>"000000000",
  32132=>"011000011",
  32133=>"010000100",
  32134=>"011011000",
  32135=>"100000001",
  32136=>"101100000",
  32137=>"111100011",
  32138=>"000100100",
  32139=>"001000000",
  32140=>"111111111",
  32141=>"011000000",
  32142=>"000000000",
  32143=>"000000000",
  32144=>"111001000",
  32145=>"000000111",
  32146=>"001000001",
  32147=>"011111111",
  32148=>"111111000",
  32149=>"010000000",
  32150=>"000000000",
  32151=>"111100000",
  32152=>"110111111",
  32153=>"011011111",
  32154=>"000000000",
  32155=>"111101110",
  32156=>"001000000",
  32157=>"011000001",
  32158=>"111101000",
  32159=>"111010000",
  32160=>"111100100",
  32161=>"111111001",
  32162=>"000100110",
  32163=>"000000111",
  32164=>"000000111",
  32165=>"000010111",
  32166=>"100100111",
  32167=>"111101111",
  32168=>"110110000",
  32169=>"111111100",
  32170=>"001000111",
  32171=>"001010000",
  32172=>"101111000",
  32173=>"000000000",
  32174=>"000000000",
  32175=>"000000000",
  32176=>"001001111",
  32177=>"001101101",
  32178=>"000000010",
  32179=>"111011000",
  32180=>"111111111",
  32181=>"010011111",
  32182=>"001001000",
  32183=>"111111110",
  32184=>"111111000",
  32185=>"111111111",
  32186=>"100010000",
  32187=>"000110110",
  32188=>"000000000",
  32189=>"000000000",
  32190=>"001001011",
  32191=>"101100100",
  32192=>"000000001",
  32193=>"101100101",
  32194=>"010011000",
  32195=>"001111111",
  32196=>"110110110",
  32197=>"100110000",
  32198=>"111100000",
  32199=>"111111111",
  32200=>"111000000",
  32201=>"000000000",
  32202=>"000000000",
  32203=>"111110111",
  32204=>"000000000",
  32205=>"000000001",
  32206=>"011101101",
  32207=>"000100111",
  32208=>"111111111",
  32209=>"001000000",
  32210=>"111111111",
  32211=>"110110111",
  32212=>"110111111",
  32213=>"000000000",
  32214=>"000000000",
  32215=>"001011000",
  32216=>"000101111",
  32217=>"111000010",
  32218=>"000000111",
  32219=>"100110000",
  32220=>"111101111",
  32221=>"111111111",
  32222=>"000100111",
  32223=>"101111111",
  32224=>"111111111",
  32225=>"111111111",
  32226=>"110011001",
  32227=>"111111111",
  32228=>"011000000",
  32229=>"000000000",
  32230=>"010010000",
  32231=>"000000000",
  32232=>"110111111",
  32233=>"111111000",
  32234=>"001001011",
  32235=>"111111111",
  32236=>"000110111",
  32237=>"111111110",
  32238=>"111111000",
  32239=>"100001011",
  32240=>"111111000",
  32241=>"011001000",
  32242=>"111111111",
  32243=>"000000111",
  32244=>"000000000",
  32245=>"111111011",
  32246=>"111111111",
  32247=>"101001000",
  32248=>"010011111",
  32249=>"111111000",
  32250=>"000001101",
  32251=>"000000000",
  32252=>"000100111",
  32253=>"111001011",
  32254=>"111111100",
  32255=>"111111111",
  32256=>"111000110",
  32257=>"001011010",
  32258=>"111000000",
  32259=>"000000111",
  32260=>"000111110",
  32261=>"111000000",
  32262=>"000111111",
  32263=>"111100000",
  32264=>"111111000",
  32265=>"111000010",
  32266=>"000000010",
  32267=>"111111000",
  32268=>"100111011",
  32269=>"100000010",
  32270=>"000001111",
  32271=>"000111111",
  32272=>"000000001",
  32273=>"000111110",
  32274=>"000110100",
  32275=>"110110111",
  32276=>"101001111",
  32277=>"111000100",
  32278=>"101111111",
  32279=>"000101111",
  32280=>"000000111",
  32281=>"001000011",
  32282=>"000000110",
  32283=>"011110110",
  32284=>"000010111",
  32285=>"110111111",
  32286=>"100000110",
  32287=>"000000101",
  32288=>"111111001",
  32289=>"111111010",
  32290=>"111111100",
  32291=>"110110111",
  32292=>"000111111",
  32293=>"000000001",
  32294=>"111111111",
  32295=>"101000111",
  32296=>"000100110",
  32297=>"111111111",
  32298=>"111111111",
  32299=>"100000100",
  32300=>"000000011",
  32301=>"110000000",
  32302=>"001000000",
  32303=>"101000000",
  32304=>"111111000",
  32305=>"000001111",
  32306=>"111111111",
  32307=>"000000000",
  32308=>"000001001",
  32309=>"001111101",
  32310=>"000000000",
  32311=>"101111011",
  32312=>"111111000",
  32313=>"111110111",
  32314=>"111111010",
  32315=>"000000000",
  32316=>"111100000",
  32317=>"010111111",
  32318=>"011101111",
  32319=>"111001000",
  32320=>"111001001",
  32321=>"110110000",
  32322=>"001000000",
  32323=>"111000000",
  32324=>"000000001",
  32325=>"000000100",
  32326=>"011011010",
  32327=>"011011000",
  32328=>"111110000",
  32329=>"000000011",
  32330=>"100100101",
  32331=>"110100111",
  32332=>"000000111",
  32333=>"100000000",
  32334=>"000111000",
  32335=>"111001111",
  32336=>"110111110",
  32337=>"101110000",
  32338=>"111110000",
  32339=>"001000000",
  32340=>"000000100",
  32341=>"111100100",
  32342=>"111001111",
  32343=>"000000000",
  32344=>"110111110",
  32345=>"000000000",
  32346=>"111100110",
  32347=>"111111101",
  32348=>"000111111",
  32349=>"001000100",
  32350=>"111000000",
  32351=>"111101000",
  32352=>"101000000",
  32353=>"110110001",
  32354=>"011011001",
  32355=>"000000000",
  32356=>"111111011",
  32357=>"111000000",
  32358=>"111011000",
  32359=>"111010111",
  32360=>"101100111",
  32361=>"111111101",
  32362=>"111011000",
  32363=>"011111111",
  32364=>"110111111",
  32365=>"000000111",
  32366=>"111111111",
  32367=>"000000000",
  32368=>"111000111",
  32369=>"101110100",
  32370=>"000000111",
  32371=>"011001011",
  32372=>"000111111",
  32373=>"111111111",
  32374=>"110111101",
  32375=>"000000111",
  32376=>"111011001",
  32377=>"111111111",
  32378=>"000000110",
  32379=>"001000100",
  32380=>"111011111",
  32381=>"000110110",
  32382=>"000000111",
  32383=>"000000011",
  32384=>"100000000",
  32385=>"111111111",
  32386=>"000000011",
  32387=>"111100100",
  32388=>"111111111",
  32389=>"111101011",
  32390=>"111111000",
  32391=>"000000001",
  32392=>"000000000",
  32393=>"111000000",
  32394=>"011000011",
  32395=>"111111000",
  32396=>"100110111",
  32397=>"000000111",
  32398=>"100111111",
  32399=>"000100111",
  32400=>"101000111",
  32401=>"111011000",
  32402=>"110000000",
  32403=>"101100001",
  32404=>"111001101",
  32405=>"000101111",
  32406=>"111000000",
  32407=>"111100000",
  32408=>"110100101",
  32409=>"111011000",
  32410=>"100111011",
  32411=>"000000011",
  32412=>"111101100",
  32413=>"111110101",
  32414=>"111111110",
  32415=>"000000000",
  32416=>"111101111",
  32417=>"110000000",
  32418=>"000000000",
  32419=>"111111111",
  32420=>"000100110",
  32421=>"000111110",
  32422=>"101000000",
  32423=>"100101100",
  32424=>"100000000",
  32425=>"011011000",
  32426=>"000010010",
  32427=>"111001000",
  32428=>"111000100",
  32429=>"110010110",
  32430=>"111010110",
  32431=>"010011101",
  32432=>"111000000",
  32433=>"000101101",
  32434=>"111111010",
  32435=>"000000000",
  32436=>"111111111",
  32437=>"100100110",
  32438=>"111001111",
  32439=>"111111111",
  32440=>"111111111",
  32441=>"000000111",
  32442=>"000110111",
  32443=>"100100111",
  32444=>"100000000",
  32445=>"111110111",
  32446=>"100000011",
  32447=>"100110111",
  32448=>"000000000",
  32449=>"000000000",
  32450=>"000000000",
  32451=>"111011000",
  32452=>"000000100",
  32453=>"000000000",
  32454=>"000110111",
  32455=>"111111000",
  32456=>"111000001",
  32457=>"111011011",
  32458=>"000000001",
  32459=>"000111111",
  32460=>"000000000",
  32461=>"000100010",
  32462=>"000101001",
  32463=>"111001001",
  32464=>"110100000",
  32465=>"000001000",
  32466=>"100000010",
  32467=>"000000000",
  32468=>"110000000",
  32469=>"110110111",
  32470=>"111100100",
  32471=>"000000000",
  32472=>"000000011",
  32473=>"000000001",
  32474=>"111111111",
  32475=>"100100010",
  32476=>"111111111",
  32477=>"000000000",
  32478=>"000000000",
  32479=>"100100000",
  32480=>"111110110",
  32481=>"110111000",
  32482=>"111101000",
  32483=>"100000000",
  32484=>"001111111",
  32485=>"000111111",
  32486=>"100101111",
  32487=>"100000110",
  32488=>"111111001",
  32489=>"100010111",
  32490=>"111010111",
  32491=>"111010011",
  32492=>"000111111",
  32493=>"111111100",
  32494=>"111000111",
  32495=>"111000000",
  32496=>"100011011",
  32497=>"000111111",
  32498=>"000001111",
  32499=>"111000010",
  32500=>"111111011",
  32501=>"001111110",
  32502=>"111101001",
  32503=>"111110000",
  32504=>"110010010",
  32505=>"101111010",
  32506=>"101000111",
  32507=>"111000000",
  32508=>"000000110",
  32509=>"001111110",
  32510=>"100100000",
  32511=>"000000001",
  32512=>"110110000",
  32513=>"000100110",
  32514=>"111000000",
  32515=>"110011011",
  32516=>"000110000",
  32517=>"010110000",
  32518=>"010000000",
  32519=>"000000010",
  32520=>"101011111",
  32521=>"000000011",
  32522=>"100100000",
  32523=>"111111000",
  32524=>"001001111",
  32525=>"111011010",
  32526=>"010110111",
  32527=>"000100101",
  32528=>"101111111",
  32529=>"110100000",
  32530=>"111001111",
  32531=>"100000000",
  32532=>"000110110",
  32533=>"000000000",
  32534=>"001111111",
  32535=>"000000111",
  32536=>"000001111",
  32537=>"111000001",
  32538=>"111111111",
  32539=>"100111111",
  32540=>"111111110",
  32541=>"111110000",
  32542=>"011111000",
  32543=>"011011011",
  32544=>"110111000",
  32545=>"000000000",
  32546=>"100100111",
  32547=>"111011010",
  32548=>"110110011",
  32549=>"011111111",
  32550=>"110000000",
  32551=>"000000000",
  32552=>"000110111",
  32553=>"100000000",
  32554=>"111010000",
  32555=>"111100000",
  32556=>"001111111",
  32557=>"000110110",
  32558=>"000000110",
  32559=>"000000000",
  32560=>"111111110",
  32561=>"110000110",
  32562=>"100000000",
  32563=>"111111000",
  32564=>"110000000",
  32565=>"010000000",
  32566=>"001000110",
  32567=>"110000000",
  32568=>"100000000",
  32569=>"111000000",
  32570=>"100100101",
  32571=>"101001001",
  32572=>"111000101",
  32573=>"100000000",
  32574=>"111001001",
  32575=>"100000000",
  32576=>"111101000",
  32577=>"111011111",
  32578=>"111110000",
  32579=>"000111111",
  32580=>"000000001",
  32581=>"100100100",
  32582=>"011111111",
  32583=>"111111111",
  32584=>"111101111",
  32585=>"000000000",
  32586=>"001011111",
  32587=>"000001011",
  32588=>"000111011",
  32589=>"010110111",
  32590=>"100000000",
  32591=>"100100011",
  32592=>"000111111",
  32593=>"111001000",
  32594=>"001000111",
  32595=>"100010000",
  32596=>"011111111",
  32597=>"011001001",
  32598=>"000000111",
  32599=>"111111111",
  32600=>"111011011",
  32601=>"001000000",
  32602=>"111111111",
  32603=>"111111111",
  32604=>"110000000",
  32605=>"111111111",
  32606=>"111011111",
  32607=>"001000000",
  32608=>"111000000",
  32609=>"110101111",
  32610=>"001100100",
  32611=>"111111111",
  32612=>"111111111",
  32613=>"111000000",
  32614=>"111111111",
  32615=>"100000001",
  32616=>"101100110",
  32617=>"100011011",
  32618=>"000011111",
  32619=>"111011011",
  32620=>"110011000",
  32621=>"111111111",
  32622=>"000110010",
  32623=>"100000111",
  32624=>"001000000",
  32625=>"000000011",
  32626=>"000000011",
  32627=>"100100111",
  32628=>"111111011",
  32629=>"000001111",
  32630=>"111000000",
  32631=>"111111000",
  32632=>"111001101",
  32633=>"100000100",
  32634=>"000000000",
  32635=>"101111111",
  32636=>"000000011",
  32637=>"100000101",
  32638=>"110110000",
  32639=>"000111111",
  32640=>"110000000",
  32641=>"000000111",
  32642=>"000000111",
  32643=>"000110110",
  32644=>"111111000",
  32645=>"111111111",
  32646=>"111010000",
  32647=>"011111011",
  32648=>"001111011",
  32649=>"101000000",
  32650=>"000110000",
  32651=>"111111000",
  32652=>"111000000",
  32653=>"111111111",
  32654=>"111111111",
  32655=>"000000000",
  32656=>"000001001",
  32657=>"001000001",
  32658=>"110110111",
  32659=>"111001000",
  32660=>"000111100",
  32661=>"000011000",
  32662=>"000110111",
  32663=>"111101000",
  32664=>"001101111",
  32665=>"100100000",
  32666=>"110111011",
  32667=>"110110001",
  32668=>"111111001",
  32669=>"000011010",
  32670=>"101111111",
  32671=>"000001001",
  32672=>"000000000",
  32673=>"101001111",
  32674=>"100000000",
  32675=>"111100001",
  32676=>"110000101",
  32677=>"111111000",
  32678=>"000000000",
  32679=>"000000110",
  32680=>"010000000",
  32681=>"011010000",
  32682=>"111111010",
  32683=>"011001101",
  32684=>"011001000",
  32685=>"111000000",
  32686=>"110000011",
  32687=>"000000011",
  32688=>"000000000",
  32689=>"111101000",
  32690=>"000000010",
  32691=>"111000000",
  32692=>"111011011",
  32693=>"001001111",
  32694=>"000000100",
  32695=>"010111011",
  32696=>"111110000",
  32697=>"111110111",
  32698=>"111111000",
  32699=>"100100000",
  32700=>"000000000",
  32701=>"000011011",
  32702=>"111011100",
  32703=>"101101100",
  32704=>"111111001",
  32705=>"000000000",
  32706=>"000000000",
  32707=>"000000000",
  32708=>"000000000",
  32709=>"001000101",
  32710=>"101000001",
  32711=>"111100100",
  32712=>"100110111",
  32713=>"111111111",
  32714=>"101000001",
  32715=>"000000011",
  32716=>"000000000",
  32717=>"111111111",
  32718=>"100000000",
  32719=>"101111101",
  32720=>"111111000",
  32721=>"000100100",
  32722=>"000000000",
  32723=>"001001111",
  32724=>"100100110",
  32725=>"111110000",
  32726=>"110000000",
  32727=>"011111000",
  32728=>"101000000",
  32729=>"111111100",
  32730=>"000000001",
  32731=>"111111111",
  32732=>"110110111",
  32733=>"111001111",
  32734=>"000010011",
  32735=>"100100110",
  32736=>"000011001",
  32737=>"101111111",
  32738=>"111000000",
  32739=>"001011011",
  32740=>"111001000",
  32741=>"000111000",
  32742=>"000000001",
  32743=>"111000000",
  32744=>"101100111",
  32745=>"111010000",
  32746=>"001000000",
  32747=>"111111000",
  32748=>"000000000",
  32749=>"100100000",
  32750=>"111101111",
  32751=>"000000111",
  32752=>"000000111",
  32753=>"111110111",
  32754=>"100000000",
  32755=>"111100111",
  32756=>"011111111",
  32757=>"100000000",
  32758=>"111111011",
  32759=>"001000010",
  32760=>"010000000",
  32761=>"010011000",
  32762=>"000000000",
  32763=>"111000000",
  32764=>"111101001",
  32765=>"000000000",
  32766=>"111100000",
  32767=>"111001011",
  32768=>"000011011",
  32769=>"011011110",
  32770=>"111111111",
  32771=>"000000000",
  32772=>"001001111",
  32773=>"001100100",
  32774=>"111011111",
  32775=>"111000011",
  32776=>"111100000",
  32777=>"111111111",
  32778=>"111111111",
  32779=>"111111110",
  32780=>"111101101",
  32781=>"100000000",
  32782=>"101100111",
  32783=>"000000000",
  32784=>"000100111",
  32785=>"000111111",
  32786=>"110100110",
  32787=>"000000101",
  32788=>"111111111",
  32789=>"000000111",
  32790=>"000000000",
  32791=>"000011111",
  32792=>"100100100",
  32793=>"000111111",
  32794=>"011000111",
  32795=>"000111111",
  32796=>"011011111",
  32797=>"101001000",
  32798=>"000110111",
  32799=>"111001000",
  32800=>"000000000",
  32801=>"000000110",
  32802=>"111101000",
  32803=>"000000100",
  32804=>"111101000",
  32805=>"111111111",
  32806=>"001000000",
  32807=>"111100000",
  32808=>"101000000",
  32809=>"000000111",
  32810=>"000001001",
  32811=>"011001000",
  32812=>"000111111",
  32813=>"000111011",
  32814=>"111101000",
  32815=>"010000000",
  32816=>"000001110",
  32817=>"000001000",
  32818=>"100111100",
  32819=>"000100111",
  32820=>"111111111",
  32821=>"111111111",
  32822=>"100011111",
  32823=>"000000000",
  32824=>"101000001",
  32825=>"000011111",
  32826=>"000000000",
  32827=>"111000000",
  32828=>"111011000",
  32829=>"111111111",
  32830=>"111111000",
  32831=>"111111100",
  32832=>"111111111",
  32833=>"111111000",
  32834=>"011011011",
  32835=>"000000111",
  32836=>"010001000",
  32837=>"011000000",
  32838=>"000000000",
  32839=>"111111011",
  32840=>"110011000",
  32841=>"011001000",
  32842=>"111000100",
  32843=>"111111110",
  32844=>"101111000",
  32845=>"111101111",
  32846=>"000000101",
  32847=>"111111111",
  32848=>"011011000",
  32849=>"111111111",
  32850=>"000000111",
  32851=>"000011111",
  32852=>"100100111",
  32853=>"001011000",
  32854=>"011000000",
  32855=>"111111111",
  32856=>"011001111",
  32857=>"111000000",
  32858=>"000000100",
  32859=>"101111111",
  32860=>"111111111",
  32861=>"100110111",
  32862=>"111101100",
  32863=>"110100000",
  32864=>"000000000",
  32865=>"011011111",
  32866=>"000000000",
  32867=>"111000010",
  32868=>"101100000",
  32869=>"110111010",
  32870=>"000000001",
  32871=>"111111111",
  32872=>"000000000",
  32873=>"111111111",
  32874=>"010000110",
  32875=>"111110100",
  32876=>"111110000",
  32877=>"111111111",
  32878=>"011000000",
  32879=>"000000111",
  32880=>"111111111",
  32881=>"101001011",
  32882=>"000001111",
  32883=>"111101000",
  32884=>"000000000",
  32885=>"000101101",
  32886=>"000000000",
  32887=>"000001001",
  32888=>"111111000",
  32889=>"000000000",
  32890=>"000000000",
  32891=>"111000000",
  32892=>"111001001",
  32893=>"000000001",
  32894=>"000111111",
  32895=>"111000000",
  32896=>"100000000",
  32897=>"000111111",
  32898=>"011011111",
  32899=>"111111111",
  32900=>"000010000",
  32901=>"100000000",
  32902=>"011000000",
  32903=>"110011111",
  32904=>"000010111",
  32905=>"000000100",
  32906=>"001000000",
  32907=>"000100001",
  32908=>"000000000",
  32909=>"111111110",
  32910=>"111101011",
  32911=>"100100100",
  32912=>"011111111",
  32913=>"111111111",
  32914=>"000000000",
  32915=>"001001000",
  32916=>"111011111",
  32917=>"000101101",
  32918=>"111111111",
  32919=>"111000000",
  32920=>"000000100",
  32921=>"111000100",
  32922=>"000011011",
  32923=>"010111000",
  32924=>"111001100",
  32925=>"110110000",
  32926=>"101001001",
  32927=>"000000000",
  32928=>"000000111",
  32929=>"000010011",
  32930=>"110110000",
  32931=>"111111111",
  32932=>"010011001",
  32933=>"111001000",
  32934=>"000000000",
  32935=>"111101100",
  32936=>"000000111",
  32937=>"000000000",
  32938=>"001000000",
  32939=>"100100111",
  32940=>"011001000",
  32941=>"000111111",
  32942=>"011001000",
  32943=>"111111111",
  32944=>"110000000",
  32945=>"100100000",
  32946=>"111101111",
  32947=>"111000000",
  32948=>"000110110",
  32949=>"000111100",
  32950=>"111000000",
  32951=>"111111001",
  32952=>"111111001",
  32953=>"000000000",
  32954=>"001000000",
  32955=>"000000001",
  32956=>"000000000",
  32957=>"111101000",
  32958=>"101111000",
  32959=>"001000000",
  32960=>"111001000",
  32961=>"001000000",
  32962=>"000001111",
  32963=>"000000000",
  32964=>"100100000",
  32965=>"000010111",
  32966=>"100111001",
  32967=>"111110000",
  32968=>"000000000",
  32969=>"111111001",
  32970=>"000100111",
  32971=>"110000100",
  32972=>"000000110",
  32973=>"000000000",
  32974=>"001000000",
  32975=>"000111100",
  32976=>"000010000",
  32977=>"000000000",
  32978=>"000000000",
  32979=>"000000100",
  32980=>"001000000",
  32981=>"000000100",
  32982=>"010000010",
  32983=>"000000111",
  32984=>"010111111",
  32985=>"111111111",
  32986=>"011000000",
  32987=>"111000000",
  32988=>"111000000",
  32989=>"111000000",
  32990=>"000001111",
  32991=>"000100100",
  32992=>"000000111",
  32993=>"001011111",
  32994=>"111111111",
  32995=>"000000111",
  32996=>"100111011",
  32997=>"100111111",
  32998=>"000000000",
  32999=>"000100101",
  33000=>"000011011",
  33001=>"100100000",
  33002=>"111000110",
  33003=>"000010010",
  33004=>"111111000",
  33005=>"000000111",
  33006=>"101000000",
  33007=>"111111000",
  33008=>"111111000",
  33009=>"000111111",
  33010=>"000000000",
  33011=>"111000101",
  33012=>"000100100",
  33013=>"111001000",
  33014=>"000100110",
  33015=>"110111111",
  33016=>"000111111",
  33017=>"000000000",
  33018=>"111000000",
  33019=>"000000000",
  33020=>"000001001",
  33021=>"001001110",
  33022=>"000000000",
  33023=>"000000000",
  33024=>"111111111",
  33025=>"011000000",
  33026=>"111010111",
  33027=>"000100100",
  33028=>"001111000",
  33029=>"100000000",
  33030=>"111000100",
  33031=>"000000000",
  33032=>"011000000",
  33033=>"111011000",
  33034=>"110100000",
  33035=>"111110110",
  33036=>"000001101",
  33037=>"111111111",
  33038=>"001000000",
  33039=>"000000000",
  33040=>"101100001",
  33041=>"111111101",
  33042=>"111110000",
  33043=>"000000000",
  33044=>"111111001",
  33045=>"000000110",
  33046=>"000001011",
  33047=>"111101000",
  33048=>"001001111",
  33049=>"110110000",
  33050=>"000000000",
  33051=>"000100111",
  33052=>"000100110",
  33053=>"110000000",
  33054=>"000000000",
  33055=>"111111111",
  33056=>"110000001",
  33057=>"000100110",
  33058=>"111111111",
  33059=>"110111111",
  33060=>"000010111",
  33061=>"011011101",
  33062=>"111111111",
  33063=>"111100000",
  33064=>"000111111",
  33065=>"111111110",
  33066=>"000000111",
  33067=>"111100000",
  33068=>"111111001",
  33069=>"011000000",
  33070=>"000111111",
  33071=>"000001000",
  33072=>"111001000",
  33073=>"000100111",
  33074=>"000000000",
  33075=>"100111111",
  33076=>"011001000",
  33077=>"111111000",
  33078=>"100010000",
  33079=>"001011001",
  33080=>"000110111",
  33081=>"111010000",
  33082=>"000011111",
  33083=>"000000000",
  33084=>"000011111",
  33085=>"111111000",
  33086=>"111011000",
  33087=>"111111001",
  33088=>"100000000",
  33089=>"000011011",
  33090=>"111111011",
  33091=>"000010111",
  33092=>"111011000",
  33093=>"100000000",
  33094=>"000000111",
  33095=>"111111111",
  33096=>"000000000",
  33097=>"000000000",
  33098=>"000111001",
  33099=>"100000000",
  33100=>"001001111",
  33101=>"111111000",
  33102=>"011011100",
  33103=>"000000110",
  33104=>"110100111",
  33105=>"111100100",
  33106=>"111111110",
  33107=>"010001000",
  33108=>"011000010",
  33109=>"011011010",
  33110=>"111111111",
  33111=>"111101000",
  33112=>"011000000",
  33113=>"000000000",
  33114=>"011111111",
  33115=>"011101111",
  33116=>"111100100",
  33117=>"111111111",
  33118=>"111000000",
  33119=>"111100111",
  33120=>"110111111",
  33121=>"000111111",
  33122=>"000001111",
  33123=>"110011000",
  33124=>"001001001",
  33125=>"111000000",
  33126=>"000010111",
  33127=>"111111000",
  33128=>"111110110",
  33129=>"000111111",
  33130=>"001001001",
  33131=>"011000111",
  33132=>"000000000",
  33133=>"000000100",
  33134=>"111111011",
  33135=>"111111111",
  33136=>"010110111",
  33137=>"111111000",
  33138=>"000010000",
  33139=>"011100100",
  33140=>"000000000",
  33141=>"000111111",
  33142=>"000100111",
  33143=>"111010000",
  33144=>"000111000",
  33145=>"000111111",
  33146=>"100110111",
  33147=>"000010000",
  33148=>"000001001",
  33149=>"001011000",
  33150=>"100100001",
  33151=>"110111111",
  33152=>"000000000",
  33153=>"000011010",
  33154=>"000000001",
  33155=>"100000000",
  33156=>"110000000",
  33157=>"111111110",
  33158=>"101000010",
  33159=>"000000000",
  33160=>"111111111",
  33161=>"001000110",
  33162=>"111110100",
  33163=>"111111111",
  33164=>"000000000",
  33165=>"111111111",
  33166=>"111111000",
  33167=>"000000000",
  33168=>"000000110",
  33169=>"100000000",
  33170=>"001001001",
  33171=>"000110111",
  33172=>"111000000",
  33173=>"010010010",
  33174=>"000001011",
  33175=>"111101111",
  33176=>"000111111",
  33177=>"101001000",
  33178=>"110110111",
  33179=>"111111001",
  33180=>"100000000",
  33181=>"000000000",
  33182=>"111011001",
  33183=>"000000000",
  33184=>"000000000",
  33185=>"100110110",
  33186=>"011000101",
  33187=>"110000000",
  33188=>"111111000",
  33189=>"111111000",
  33190=>"111100000",
  33191=>"111111111",
  33192=>"110000000",
  33193=>"000000100",
  33194=>"111100111",
  33195=>"111111011",
  33196=>"000000111",
  33197=>"111111110",
  33198=>"111000000",
  33199=>"101000000",
  33200=>"111000000",
  33201=>"111111000",
  33202=>"000000111",
  33203=>"000000000",
  33204=>"111011011",
  33205=>"000000101",
  33206=>"000000111",
  33207=>"011111000",
  33208=>"001000000",
  33209=>"101111111",
  33210=>"000000000",
  33211=>"111011100",
  33212=>"011111111",
  33213=>"000111000",
  33214=>"101111111",
  33215=>"011001001",
  33216=>"100000000",
  33217=>"111111110",
  33218=>"000000111",
  33219=>"000000000",
  33220=>"011001000",
  33221=>"001000000",
  33222=>"100000000",
  33223=>"000001001",
  33224=>"001101111",
  33225=>"000000111",
  33226=>"111000000",
  33227=>"000001101",
  33228=>"000000000",
  33229=>"001000000",
  33230=>"000000010",
  33231=>"001011111",
  33232=>"110111111",
  33233=>"111111110",
  33234=>"000111011",
  33235=>"000000011",
  33236=>"100100100",
  33237=>"001000111",
  33238=>"101100111",
  33239=>"001111110",
  33240=>"111001000",
  33241=>"111101001",
  33242=>"111000000",
  33243=>"001000000",
  33244=>"011001011",
  33245=>"000000000",
  33246=>"100100000",
  33247=>"111100000",
  33248=>"010110111",
  33249=>"111111110",
  33250=>"111101000",
  33251=>"000000011",
  33252=>"111111111",
  33253=>"111000000",
  33254=>"000001001",
  33255=>"000000110",
  33256=>"111111110",
  33257=>"110111101",
  33258=>"111011000",
  33259=>"010110011",
  33260=>"110111011",
  33261=>"111110110",
  33262=>"111111000",
  33263=>"111000111",
  33264=>"001000101",
  33265=>"110000001",
  33266=>"011011000",
  33267=>"000000110",
  33268=>"111111000",
  33269=>"110110000",
  33270=>"111111000",
  33271=>"001111111",
  33272=>"000000010",
  33273=>"000000110",
  33274=>"000000111",
  33275=>"000000111",
  33276=>"110000100",
  33277=>"010000100",
  33278=>"000000011",
  33279=>"111111000",
  33280=>"111111101",
  33281=>"110110111",
  33282=>"101101000",
  33283=>"111001000",
  33284=>"111001000",
  33285=>"000000111",
  33286=>"010000001",
  33287=>"000000011",
  33288=>"100111011",
  33289=>"111111101",
  33290=>"111111011",
  33291=>"010001000",
  33292=>"110110100",
  33293=>"010000000",
  33294=>"101111110",
  33295=>"111011011",
  33296=>"000000101",
  33297=>"000000000",
  33298=>"011111111",
  33299=>"000000000",
  33300=>"111111111",
  33301=>"111111110",
  33302=>"110000000",
  33303=>"111111011",
  33304=>"111110110",
  33305=>"000001111",
  33306=>"111110000",
  33307=>"111000000",
  33308=>"111000000",
  33309=>"111111111",
  33310=>"111000000",
  33311=>"111110000",
  33312=>"000000010",
  33313=>"111110000",
  33314=>"000111111",
  33315=>"100100111",
  33316=>"111111111",
  33317=>"111111111",
  33318=>"111000000",
  33319=>"111101000",
  33320=>"111111111",
  33321=>"001011111",
  33322=>"000000000",
  33323=>"000101111",
  33324=>"110111111",
  33325=>"000000000",
  33326=>"111111111",
  33327=>"000000110",
  33328=>"000101001",
  33329=>"000110111",
  33330=>"100000001",
  33331=>"100100000",
  33332=>"111111101",
  33333=>"110110110",
  33334=>"111111111",
  33335=>"110111011",
  33336=>"000101111",
  33337=>"001001111",
  33338=>"111111111",
  33339=>"000000000",
  33340=>"001000000",
  33341=>"111111111",
  33342=>"001010111",
  33343=>"000101111",
  33344=>"000111111",
  33345=>"110110010",
  33346=>"000000000",
  33347=>"000011000",
  33348=>"100100111",
  33349=>"011111011",
  33350=>"111111111",
  33351=>"100111111",
  33352=>"000000000",
  33353=>"111111110",
  33354=>"001001000",
  33355=>"110000111",
  33356=>"000000000",
  33357=>"000000100",
  33358=>"000000111",
  33359=>"111101100",
  33360=>"111111111",
  33361=>"100000000",
  33362=>"001111111",
  33363=>"000000100",
  33364=>"000000000",
  33365=>"110111100",
  33366=>"111000000",
  33367=>"000001011",
  33368=>"111111111",
  33369=>"111111111",
  33370=>"110000000",
  33371=>"111000010",
  33372=>"111111111",
  33373=>"111111101",
  33374=>"111111000",
  33375=>"111111111",
  33376=>"111111111",
  33377=>"001000000",
  33378=>"111111011",
  33379=>"000000100",
  33380=>"000000000",
  33381=>"000000000",
  33382=>"000000000",
  33383=>"000111111",
  33384=>"111111111",
  33385=>"111100100",
  33386=>"111000000",
  33387=>"010111111",
  33388=>"000000000",
  33389=>"000000001",
  33390=>"111111000",
  33391=>"000000000",
  33392=>"111100000",
  33393=>"111111111",
  33394=>"000011011",
  33395=>"101000000",
  33396=>"011001010",
  33397=>"000000000",
  33398=>"011110110",
  33399=>"111111001",
  33400=>"000110010",
  33401=>"000000000",
  33402=>"111111111",
  33403=>"010000000",
  33404=>"110110111",
  33405=>"111001111",
  33406=>"111111111",
  33407=>"000000000",
  33408=>"111111000",
  33409=>"010000000",
  33410=>"000000100",
  33411=>"011001001",
  33412=>"100100100",
  33413=>"000001000",
  33414=>"111111111",
  33415=>"111111001",
  33416=>"000000000",
  33417=>"111111111",
  33418=>"111100111",
  33419=>"111111000",
  33420=>"100001011",
  33421=>"101000110",
  33422=>"111011001",
  33423=>"110100000",
  33424=>"000000000",
  33425=>"000000000",
  33426=>"111111111",
  33427=>"111111111",
  33428=>"101000000",
  33429=>"111110000",
  33430=>"110111111",
  33431=>"100000000",
  33432=>"111111111",
  33433=>"000000000",
  33434=>"011000001",
  33435=>"000000000",
  33436=>"011000010",
  33437=>"011011000",
  33438=>"000000111",
  33439=>"000000110",
  33440=>"111111111",
  33441=>"000100111",
  33442=>"111111101",
  33443=>"010011000",
  33444=>"111011011",
  33445=>"000000101",
  33446=>"000000000",
  33447=>"001000000",
  33448=>"111111111",
  33449=>"111111111",
  33450=>"000000111",
  33451=>"000000000",
  33452=>"110000000",
  33453=>"111000000",
  33454=>"111111111",
  33455=>"011101111",
  33456=>"111111111",
  33457=>"011111111",
  33458=>"000000000",
  33459=>"111111111",
  33460=>"111111111",
  33461=>"000000001",
  33462=>"101101111",
  33463=>"000100111",
  33464=>"111111000",
  33465=>"111111000",
  33466=>"111110110",
  33467=>"111000111",
  33468=>"111111111",
  33469=>"000000111",
  33470=>"000000110",
  33471=>"111000111",
  33472=>"001000000",
  33473=>"001001001",
  33474=>"011011111",
  33475=>"111010000",
  33476=>"110111000",
  33477=>"111111111",
  33478=>"110110111",
  33479=>"111111111",
  33480=>"000000000",
  33481=>"111110111",
  33482=>"111111110",
  33483=>"111011111",
  33484=>"111111101",
  33485=>"000000000",
  33486=>"111111111",
  33487=>"111111110",
  33488=>"111111100",
  33489=>"111111110",
  33490=>"000000011",
  33491=>"111111111",
  33492=>"101111101",
  33493=>"110111111",
  33494=>"111111010",
  33495=>"111101111",
  33496=>"111111101",
  33497=>"011001111",
  33498=>"000000000",
  33499=>"111000111",
  33500=>"111111000",
  33501=>"111111111",
  33502=>"001111111",
  33503=>"111010110",
  33504=>"110111111",
  33505=>"111111111",
  33506=>"111111111",
  33507=>"111111111",
  33508=>"111010000",
  33509=>"000000001",
  33510=>"111100000",
  33511=>"001001111",
  33512=>"000011001",
  33513=>"111111000",
  33514=>"011011111",
  33515=>"000000011",
  33516=>"101000000",
  33517=>"110111110",
  33518=>"000011111",
  33519=>"001111111",
  33520=>"000011111",
  33521=>"000000100",
  33522=>"001111000",
  33523=>"111111111",
  33524=>"110111111",
  33525=>"111111110",
  33526=>"000110000",
  33527=>"000000111",
  33528=>"110111111",
  33529=>"100010111",
  33530=>"111000111",
  33531=>"100000000",
  33532=>"011000100",
  33533=>"000000100",
  33534=>"010000000",
  33535=>"000000000",
  33536=>"111111111",
  33537=>"001001000",
  33538=>"110000000",
  33539=>"111111100",
  33540=>"000000010",
  33541=>"111111001",
  33542=>"101100111",
  33543=>"111000000",
  33544=>"111000111",
  33545=>"111111111",
  33546=>"100100000",
  33547=>"110000000",
  33548=>"000000000",
  33549=>"110000000",
  33550=>"100000000",
  33551=>"111001001",
  33552=>"111111110",
  33553=>"111101111",
  33554=>"100111111",
  33555=>"111011111",
  33556=>"011001011",
  33557=>"000110101",
  33558=>"110110100",
  33559=>"111111011",
  33560=>"111101111",
  33561=>"111001100",
  33562=>"111111001",
  33563=>"010000010",
  33564=>"000000100",
  33565=>"111111111",
  33566=>"000000000",
  33567=>"000100111",
  33568=>"001001111",
  33569=>"111111111",
  33570=>"111000000",
  33571=>"111111111",
  33572=>"011111110",
  33573=>"101111111",
  33574=>"001001101",
  33575=>"000000000",
  33576=>"101111111",
  33577=>"000000000",
  33578=>"001111111",
  33579=>"111111111",
  33580=>"111011000",
  33581=>"111011001",
  33582=>"000000111",
  33583=>"111111111",
  33584=>"000000001",
  33585=>"010011001",
  33586=>"000010000",
  33587=>"000100111",
  33588=>"111100100",
  33589=>"011000101",
  33590=>"101111111",
  33591=>"111000000",
  33592=>"111111110",
  33593=>"000000111",
  33594=>"000000000",
  33595=>"000000000",
  33596=>"000000011",
  33597=>"111111001",
  33598=>"001100111",
  33599=>"000000000",
  33600=>"000111110",
  33601=>"110111111",
  33602=>"000001000",
  33603=>"111111111",
  33604=>"001101111",
  33605=>"111111111",
  33606=>"000111111",
  33607=>"111111011",
  33608=>"000000111",
  33609=>"000000111",
  33610=>"100111111",
  33611=>"010101101",
  33612=>"010000000",
  33613=>"000000000",
  33614=>"111101101",
  33615=>"001000000",
  33616=>"111111111",
  33617=>"000100110",
  33618=>"011001111",
  33619=>"000000000",
  33620=>"111111111",
  33621=>"011111001",
  33622=>"100011111",
  33623=>"111111110",
  33624=>"111000011",
  33625=>"111000000",
  33626=>"000001000",
  33627=>"111111111",
  33628=>"000000010",
  33629=>"111111111",
  33630=>"111010011",
  33631=>"011111101",
  33632=>"111110110",
  33633=>"110111111",
  33634=>"100000000",
  33635=>"111011000",
  33636=>"010010010",
  33637=>"110110111",
  33638=>"100100101",
  33639=>"111001001",
  33640=>"111011011",
  33641=>"110111000",
  33642=>"000010000",
  33643=>"000000100",
  33644=>"100000000",
  33645=>"111111111",
  33646=>"111111111",
  33647=>"000000111",
  33648=>"000001001",
  33649=>"000000110",
  33650=>"010000011",
  33651=>"111111111",
  33652=>"000010110",
  33653=>"011000010",
  33654=>"011011010",
  33655=>"000010000",
  33656=>"001000111",
  33657=>"111000001",
  33658=>"110110010",
  33659=>"000000000",
  33660=>"100110111",
  33661=>"111111111",
  33662=>"000000001",
  33663=>"000000000",
  33664=>"100101110",
  33665=>"100111111",
  33666=>"111111110",
  33667=>"110111111",
  33668=>"101111000",
  33669=>"111110000",
  33670=>"111011000",
  33671=>"011000000",
  33672=>"000011111",
  33673=>"000000000",
  33674=>"000000000",
  33675=>"111111111",
  33676=>"000000001",
  33677=>"011111111",
  33678=>"001000111",
  33679=>"101000000",
  33680=>"000000011",
  33681=>"101101111",
  33682=>"111101101",
  33683=>"001000110",
  33684=>"111111000",
  33685=>"110110000",
  33686=>"111111000",
  33687=>"010011100",
  33688=>"111000000",
  33689=>"000000000",
  33690=>"111111000",
  33691=>"011001111",
  33692=>"111111110",
  33693=>"110110111",
  33694=>"110111011",
  33695=>"101101100",
  33696=>"011011000",
  33697=>"000000001",
  33698=>"111000000",
  33699=>"000011000",
  33700=>"100000000",
  33701=>"000000000",
  33702=>"000000011",
  33703=>"000000000",
  33704=>"111111110",
  33705=>"111011011",
  33706=>"111111111",
  33707=>"110011011",
  33708=>"000000000",
  33709=>"000110011",
  33710=>"000000000",
  33711=>"100000011",
  33712=>"011011000",
  33713=>"111111111",
  33714=>"110010111",
  33715=>"111111111",
  33716=>"000000111",
  33717=>"111001000",
  33718=>"000000000",
  33719=>"111000000",
  33720=>"111111111",
  33721=>"111111011",
  33722=>"111111111",
  33723=>"000111111",
  33724=>"110111111",
  33725=>"101000011",
  33726=>"111111111",
  33727=>"111100000",
  33728=>"111111111",
  33729=>"000001000",
  33730=>"000000000",
  33731=>"000011001",
  33732=>"111111111",
  33733=>"000000000",
  33734=>"111111111",
  33735=>"000110111",
  33736=>"111111111",
  33737=>"100101111",
  33738=>"111011011",
  33739=>"111111101",
  33740=>"111111000",
  33741=>"000000110",
  33742=>"111111101",
  33743=>"110000000",
  33744=>"110000101",
  33745=>"110111111",
  33746=>"000000000",
  33747=>"101101111",
  33748=>"100000100",
  33749=>"000000000",
  33750=>"000000000",
  33751=>"111100101",
  33752=>"101000000",
  33753=>"111110110",
  33754=>"000000100",
  33755=>"001111000",
  33756=>"101000000",
  33757=>"110111111",
  33758=>"000000011",
  33759=>"111111100",
  33760=>"010000110",
  33761=>"000100000",
  33762=>"111111111",
  33763=>"111000011",
  33764=>"111100111",
  33765=>"000010000",
  33766=>"111111101",
  33767=>"010000000",
  33768=>"110101111",
  33769=>"010111111",
  33770=>"011000000",
  33771=>"100001011",
  33772=>"111011011",
  33773=>"011010011",
  33774=>"000001111",
  33775=>"011010010",
  33776=>"111111111",
  33777=>"010011111",
  33778=>"001001011",
  33779=>"111111111",
  33780=>"111111111",
  33781=>"111100000",
  33782=>"111111111",
  33783=>"111111111",
  33784=>"001111111",
  33785=>"111001001",
  33786=>"110011011",
  33787=>"111111000",
  33788=>"100110100",
  33789=>"111000000",
  33790=>"000000000",
  33791=>"110111111",
  33792=>"000000110",
  33793=>"011011111",
  33794=>"100100000",
  33795=>"111111111",
  33796=>"000000101",
  33797=>"111111111",
  33798=>"111111111",
  33799=>"001101111",
  33800=>"000111111",
  33801=>"111110000",
  33802=>"010000100",
  33803=>"100000000",
  33804=>"111111110",
  33805=>"000101111",
  33806=>"100000000",
  33807=>"000000000",
  33808=>"010111011",
  33809=>"111111111",
  33810=>"000000000",
  33811=>"000000000",
  33812=>"001001111",
  33813=>"000000000",
  33814=>"111111010",
  33815=>"111011111",
  33816=>"111111111",
  33817=>"001000000",
  33818=>"111111111",
  33819=>"100100110",
  33820=>"000000000",
  33821=>"000001100",
  33822=>"110110100",
  33823=>"111111111",
  33824=>"111111111",
  33825=>"110110100",
  33826=>"000001100",
  33827=>"000000000",
  33828=>"000101111",
  33829=>"000000011",
  33830=>"100110000",
  33831=>"111000000",
  33832=>"111101110",
  33833=>"111111111",
  33834=>"000000000",
  33835=>"110111111",
  33836=>"111111111",
  33837=>"000000000",
  33838=>"111111111",
  33839=>"111001000",
  33840=>"000000011",
  33841=>"010000000",
  33842=>"100111111",
  33843=>"101000000",
  33844=>"111111110",
  33845=>"110110100",
  33846=>"110110000",
  33847=>"110000000",
  33848=>"011110110",
  33849=>"111011111",
  33850=>"000000000",
  33851=>"111111111",
  33852=>"101000000",
  33853=>"111111111",
  33854=>"001000011",
  33855=>"111111111",
  33856=>"001001000",
  33857=>"000100000",
  33858=>"000000000",
  33859=>"111000100",
  33860=>"101100110",
  33861=>"000000100",
  33862=>"000111011",
  33863=>"111111000",
  33864=>"111111111",
  33865=>"101101111",
  33866=>"111111111",
  33867=>"111111001",
  33868=>"000000101",
  33869=>"111111111",
  33870=>"000000000",
  33871=>"000000000",
  33872=>"111111000",
  33873=>"100000000",
  33874=>"001000000",
  33875=>"010010000",
  33876=>"100111111",
  33877=>"000010010",
  33878=>"011000110",
  33879=>"111111111",
  33880=>"110110110",
  33881=>"111101111",
  33882=>"111111000",
  33883=>"111111111",
  33884=>"011011011",
  33885=>"111111111",
  33886=>"000000111",
  33887=>"111111111",
  33888=>"101111111",
  33889=>"000000000",
  33890=>"111001111",
  33891=>"000000000",
  33892=>"000111111",
  33893=>"011011111",
  33894=>"000001000",
  33895=>"001101111",
  33896=>"111111111",
  33897=>"111111110",
  33898=>"000000000",
  33899=>"000000000",
  33900=>"000000100",
  33901=>"000000000",
  33902=>"000000000",
  33903=>"001001000",
  33904=>"100111111",
  33905=>"111111001",
  33906=>"001000000",
  33907=>"000000011",
  33908=>"001101111",
  33909=>"000111110",
  33910=>"000010000",
  33911=>"000000000",
  33912=>"000001111",
  33913=>"111110010",
  33914=>"000000000",
  33915=>"111111111",
  33916=>"110110100",
  33917=>"000000000",
  33918=>"001000000",
  33919=>"001001111",
  33920=>"000000000",
  33921=>"111101101",
  33922=>"111011111",
  33923=>"001001001",
  33924=>"111111101",
  33925=>"100000000",
  33926=>"111111100",
  33927=>"111100000",
  33928=>"000111111",
  33929=>"110111000",
  33930=>"011011001",
  33931=>"100111111",
  33932=>"111101110",
  33933=>"011111111",
  33934=>"111101001",
  33935=>"111111111",
  33936=>"000000000",
  33937=>"010011011",
  33938=>"111111111",
  33939=>"000011000",
  33940=>"001001000",
  33941=>"100001011",
  33942=>"111111111",
  33943=>"111000000",
  33944=>"000000000",
  33945=>"000001111",
  33946=>"000000000",
  33947=>"111111111",
  33948=>"000000111",
  33949=>"111111010",
  33950=>"111111111",
  33951=>"000001000",
  33952=>"110100111",
  33953=>"011111111",
  33954=>"000000010",
  33955=>"111111111",
  33956=>"001111110",
  33957=>"000000111",
  33958=>"000000000",
  33959=>"000000000",
  33960=>"000000000",
  33961=>"011000000",
  33962=>"000011111",
  33963=>"011000001",
  33964=>"100111111",
  33965=>"100110110",
  33966=>"011010000",
  33967=>"111111111",
  33968=>"111111111",
  33969=>"000011001",
  33970=>"010110010",
  33971=>"111111000",
  33972=>"111111111",
  33973=>"000111100",
  33974=>"111111111",
  33975=>"000111111",
  33976=>"011111111",
  33977=>"000000000",
  33978=>"001111111",
  33979=>"011001111",
  33980=>"101100111",
  33981=>"000001001",
  33982=>"111111111",
  33983=>"000010110",
  33984=>"111111111",
  33985=>"011000000",
  33986=>"011011111",
  33987=>"000001111",
  33988=>"010010000",
  33989=>"001100100",
  33990=>"010010010",
  33991=>"010000110",
  33992=>"000000010",
  33993=>"111111111",
  33994=>"011111111",
  33995=>"000000000",
  33996=>"111011111",
  33997=>"000000000",
  33998=>"111111111",
  33999=>"000000001",
  34000=>"110010000",
  34001=>"111111111",
  34002=>"000000000",
  34003=>"111111111",
  34004=>"100111111",
  34005=>"110000111",
  34006=>"000000000",
  34007=>"011010111",
  34008=>"111001111",
  34009=>"010110001",
  34010=>"111111000",
  34011=>"110011011",
  34012=>"100000001",
  34013=>"011000111",
  34014=>"000000000",
  34015=>"111011000",
  34016=>"111111111",
  34017=>"111111111",
  34018=>"000111111",
  34019=>"000000000",
  34020=>"000010000",
  34021=>"111111111",
  34022=>"000001000",
  34023=>"001001001",
  34024=>"000010001",
  34025=>"111000000",
  34026=>"000011111",
  34027=>"111101111",
  34028=>"011011000",
  34029=>"000000000",
  34030=>"000101111",
  34031=>"000111110",
  34032=>"000000000",
  34033=>"001000100",
  34034=>"000111111",
  34035=>"100000000",
  34036=>"010010000",
  34037=>"111111111",
  34038=>"001000000",
  34039=>"000000000",
  34040=>"001001111",
  34041=>"000000000",
  34042=>"000000000",
  34043=>"111111110",
  34044=>"000000001",
  34045=>"001111111",
  34046=>"000001011",
  34047=>"100110000",
  34048=>"110111000",
  34049=>"111111111",
  34050=>"000011011",
  34051=>"000011100",
  34052=>"110111111",
  34053=>"000010000",
  34054=>"101101110",
  34055=>"111011110",
  34056=>"000000000",
  34057=>"000000000",
  34058=>"110110000",
  34059=>"000000000",
  34060=>"000101111",
  34061=>"110100010",
  34062=>"111101110",
  34063=>"111011011",
  34064=>"111111111",
  34065=>"111111111",
  34066=>"000000000",
  34067=>"111111111",
  34068=>"100111111",
  34069=>"001001011",
  34070=>"111111111",
  34071=>"011111111",
  34072=>"000000000",
  34073=>"111110000",
  34074=>"110000000",
  34075=>"111000000",
  34076=>"100111111",
  34077=>"000000000",
  34078=>"001000001",
  34079=>"000001011",
  34080=>"111000000",
  34081=>"110010000",
  34082=>"011000000",
  34083=>"000000000",
  34084=>"000000010",
  34085=>"000000000",
  34086=>"101010011",
  34087=>"111011000",
  34088=>"101111101",
  34089=>"000000010",
  34090=>"001111111",
  34091=>"101110000",
  34092=>"111111111",
  34093=>"110111110",
  34094=>"000000000",
  34095=>"101000000",
  34096=>"110110110",
  34097=>"000000000",
  34098=>"110100000",
  34099=>"000000011",
  34100=>"111101000",
  34101=>"000000000",
  34102=>"101111111",
  34103=>"000000000",
  34104=>"000101000",
  34105=>"110111111",
  34106=>"000000001",
  34107=>"010010111",
  34108=>"000000000",
  34109=>"110111111",
  34110=>"000011001",
  34111=>"000000000",
  34112=>"100111111",
  34113=>"000000000",
  34114=>"011010000",
  34115=>"111111111",
  34116=>"111111110",
  34117=>"111111111",
  34118=>"111001001",
  34119=>"000000001",
  34120=>"000000000",
  34121=>"111111111",
  34122=>"011011111",
  34123=>"111101101",
  34124=>"111111000",
  34125=>"110110111",
  34126=>"000000110",
  34127=>"001000000",
  34128=>"100101101",
  34129=>"001000001",
  34130=>"111101111",
  34131=>"011001111",
  34132=>"111111111",
  34133=>"011011011",
  34134=>"110100101",
  34135=>"000000000",
  34136=>"000000000",
  34137=>"111111110",
  34138=>"001000000",
  34139=>"111000101",
  34140=>"111100000",
  34141=>"010000000",
  34142=>"111111001",
  34143=>"111111000",
  34144=>"111111111",
  34145=>"000111111",
  34146=>"000000011",
  34147=>"111111111",
  34148=>"100111111",
  34149=>"111001000",
  34150=>"000000001",
  34151=>"100000000",
  34152=>"111111111",
  34153=>"000000101",
  34154=>"011111111",
  34155=>"000000110",
  34156=>"100110100",
  34157=>"000000000",
  34158=>"101000111",
  34159=>"000000000",
  34160=>"111111111",
  34161=>"000000000",
  34162=>"000000001",
  34163=>"000000000",
  34164=>"000000000",
  34165=>"000000000",
  34166=>"111111111",
  34167=>"000110111",
  34168=>"111111111",
  34169=>"000111111",
  34170=>"000000000",
  34171=>"111111111",
  34172=>"011111111",
  34173=>"000110100",
  34174=>"000000000",
  34175=>"000000010",
  34176=>"100100100",
  34177=>"000000000",
  34178=>"000000000",
  34179=>"000000000",
  34180=>"000000111",
  34181=>"111111100",
  34182=>"011010000",
  34183=>"000100111",
  34184=>"000000000",
  34185=>"000000100",
  34186=>"000000000",
  34187=>"111111111",
  34188=>"111111111",
  34189=>"111111111",
  34190=>"000000000",
  34191=>"011011011",
  34192=>"000000000",
  34193=>"111111001",
  34194=>"000000000",
  34195=>"000000000",
  34196=>"000000000",
  34197=>"000000000",
  34198=>"011110110",
  34199=>"000000000",
  34200=>"011000100",
  34201=>"000011111",
  34202=>"001000111",
  34203=>"111111111",
  34204=>"101101011",
  34205=>"110110110",
  34206=>"000000000",
  34207=>"111111110",
  34208=>"111111011",
  34209=>"001001000",
  34210=>"111100000",
  34211=>"000000011",
  34212=>"111111111",
  34213=>"111111011",
  34214=>"000100000",
  34215=>"000000000",
  34216=>"111111101",
  34217=>"011000100",
  34218=>"110010000",
  34219=>"000110111",
  34220=>"000000000",
  34221=>"011111111",
  34222=>"000000111",
  34223=>"000100111",
  34224=>"000000000",
  34225=>"001010000",
  34226=>"000010000",
  34227=>"000000101",
  34228=>"000000000",
  34229=>"011000111",
  34230=>"111100100",
  34231=>"111111001",
  34232=>"000000000",
  34233=>"111000000",
  34234=>"010001001",
  34235=>"111000000",
  34236=>"111111110",
  34237=>"100001000",
  34238=>"111101111",
  34239=>"110111011",
  34240=>"011111111",
  34241=>"000000001",
  34242=>"111111010",
  34243=>"111111010",
  34244=>"111000000",
  34245=>"011000000",
  34246=>"111111111",
  34247=>"110100100",
  34248=>"000001000",
  34249=>"100000000",
  34250=>"001000000",
  34251=>"111111111",
  34252=>"111111010",
  34253=>"011001011",
  34254=>"111111111",
  34255=>"000000101",
  34256=>"000000000",
  34257=>"111111111",
  34258=>"111111111",
  34259=>"000001111",
  34260=>"000000000",
  34261=>"111101000",
  34262=>"000000011",
  34263=>"001001011",
  34264=>"111001000",
  34265=>"111011011",
  34266=>"011111000",
  34267=>"111111111",
  34268=>"011111111",
  34269=>"111011000",
  34270=>"111111111",
  34271=>"111110111",
  34272=>"110110000",
  34273=>"111111111",
  34274=>"001001111",
  34275=>"011000000",
  34276=>"100100111",
  34277=>"111010000",
  34278=>"110110111",
  34279=>"000000000",
  34280=>"111011000",
  34281=>"000000000",
  34282=>"001011011",
  34283=>"001101100",
  34284=>"011000000",
  34285=>"001001101",
  34286=>"000000000",
  34287=>"110010000",
  34288=>"000000000",
  34289=>"011101100",
  34290=>"101100100",
  34291=>"000000000",
  34292=>"000000010",
  34293=>"110000000",
  34294=>"000000000",
  34295=>"110110000",
  34296=>"011000000",
  34297=>"111111101",
  34298=>"110110000",
  34299=>"010010000",
  34300=>"111111111",
  34301=>"111000100",
  34302=>"100111111",
  34303=>"111111111",
  34304=>"111111111",
  34305=>"110111000",
  34306=>"000000000",
  34307=>"111111111",
  34308=>"000101111",
  34309=>"000101100",
  34310=>"111101001",
  34311=>"111111111",
  34312=>"111111111",
  34313=>"111111101",
  34314=>"100111111",
  34315=>"010111010",
  34316=>"001111111",
  34317=>"011011000",
  34318=>"000000000",
  34319=>"011000000",
  34320=>"110111111",
  34321=>"000111110",
  34322=>"111111110",
  34323=>"000001111",
  34324=>"111111111",
  34325=>"000000000",
  34326=>"011001011",
  34327=>"111010010",
  34328=>"010000000",
  34329=>"000000000",
  34330=>"101101000",
  34331=>"000000000",
  34332=>"000000000",
  34333=>"111000000",
  34334=>"001000000",
  34335=>"111110110",
  34336=>"111111111",
  34337=>"000000001",
  34338=>"011111111",
  34339=>"011011011",
  34340=>"111111111",
  34341=>"000000000",
  34342=>"111000000",
  34343=>"000000000",
  34344=>"000000000",
  34345=>"000001110",
  34346=>"111111111",
  34347=>"111111001",
  34348=>"111100101",
  34349=>"110111000",
  34350=>"101011000",
  34351=>"111111010",
  34352=>"001100110",
  34353=>"111101111",
  34354=>"011111111",
  34355=>"101000000",
  34356=>"111111111",
  34357=>"011011011",
  34358=>"111100000",
  34359=>"100100111",
  34360=>"010000000",
  34361=>"011011011",
  34362=>"000001011",
  34363=>"100000000",
  34364=>"000000001",
  34365=>"000000100",
  34366=>"000000000",
  34367=>"000000000",
  34368=>"111100100",
  34369=>"101111011",
  34370=>"000111111",
  34371=>"111011010",
  34372=>"000001001",
  34373=>"000000000",
  34374=>"111010111",
  34375=>"111111111",
  34376=>"011011011",
  34377=>"000000000",
  34378=>"010010010",
  34379=>"111111111",
  34380=>"111111111",
  34381=>"111111111",
  34382=>"111111101",
  34383=>"000000000",
  34384=>"000000000",
  34385=>"000000100",
  34386=>"010000000",
  34387=>"010011000",
  34388=>"000000100",
  34389=>"000000000",
  34390=>"011001100",
  34391=>"111101111",
  34392=>"111001001",
  34393=>"000000000",
  34394=>"110100000",
  34395=>"111011111",
  34396=>"111111111",
  34397=>"000000000",
  34398=>"111111111",
  34399=>"111100000",
  34400=>"000000000",
  34401=>"111111111",
  34402=>"011011000",
  34403=>"111111111",
  34404=>"111110100",
  34405=>"001000100",
  34406=>"001000000",
  34407=>"111110110",
  34408=>"110100000",
  34409=>"111111111",
  34410=>"000000000",
  34411=>"000000001",
  34412=>"000000000",
  34413=>"111111111",
  34414=>"000000000",
  34415=>"000100100",
  34416=>"111111111",
  34417=>"000000110",
  34418=>"101110111",
  34419=>"111101111",
  34420=>"000100111",
  34421=>"111111010",
  34422=>"000110110",
  34423=>"000000000",
  34424=>"111111111",
  34425=>"011001000",
  34426=>"000000000",
  34427=>"000000000",
  34428=>"001000000",
  34429=>"000000000",
  34430=>"001001001",
  34431=>"000000000",
  34432=>"111111111",
  34433=>"111100110",
  34434=>"111100000",
  34435=>"111111110",
  34436=>"000000000",
  34437=>"111001000",
  34438=>"000000100",
  34439=>"011110100",
  34440=>"111111110",
  34441=>"100100000",
  34442=>"111111111",
  34443=>"000000000",
  34444=>"011011011",
  34445=>"000000000",
  34446=>"000000011",
  34447=>"001011111",
  34448=>"000000000",
  34449=>"111111111",
  34450=>"110000000",
  34451=>"000000000",
  34452=>"001000000",
  34453=>"111110110",
  34454=>"000000000",
  34455=>"011111111",
  34456=>"000000000",
  34457=>"010110110",
  34458=>"111111001",
  34459=>"000000100",
  34460=>"000110110",
  34461=>"100000000",
  34462=>"111111111",
  34463=>"011000000",
  34464=>"001000000",
  34465=>"111000000",
  34466=>"111111110",
  34467=>"010111111",
  34468=>"000000011",
  34469=>"111110110",
  34470=>"000000001",
  34471=>"111110111",
  34472=>"011000110",
  34473=>"111111111",
  34474=>"000000011",
  34475=>"111111111",
  34476=>"011011010",
  34477=>"000001000",
  34478=>"011000000",
  34479=>"000011011",
  34480=>"000001000",
  34481=>"001001000",
  34482=>"111111111",
  34483=>"000000000",
  34484=>"001011001",
  34485=>"000110111",
  34486=>"010111111",
  34487=>"000000000",
  34488=>"111011001",
  34489=>"000000001",
  34490=>"010000000",
  34491=>"000000000",
  34492=>"011110000",
  34493=>"000000000",
  34494=>"111010000",
  34495=>"111111001",
  34496=>"001000000",
  34497=>"111111001",
  34498=>"000000000",
  34499=>"000000000",
  34500=>"000001000",
  34501=>"010011011",
  34502=>"000111111",
  34503=>"000000000",
  34504=>"101101101",
  34505=>"001000100",
  34506=>"001011111",
  34507=>"000000000",
  34508=>"111010111",
  34509=>"000000000",
  34510=>"000111110",
  34511=>"000000000",
  34512=>"001111111",
  34513=>"111011011",
  34514=>"111111000",
  34515=>"000010110",
  34516=>"111000000",
  34517=>"111001010",
  34518=>"111110100",
  34519=>"101000000",
  34520=>"111000000",
  34521=>"111111111",
  34522=>"011111111",
  34523=>"000000011",
  34524=>"111110111",
  34525=>"000100111",
  34526=>"000000000",
  34527=>"000000110",
  34528=>"000000000",
  34529=>"000111110",
  34530=>"011011010",
  34531=>"111111111",
  34532=>"111111001",
  34533=>"100100011",
  34534=>"000000001",
  34535=>"011111111",
  34536=>"000000100",
  34537=>"111111110",
  34538=>"001000000",
  34539=>"110111111",
  34540=>"000001111",
  34541=>"000000000",
  34542=>"000000100",
  34543=>"000000000",
  34544=>"111111111",
  34545=>"000000001",
  34546=>"111111000",
  34547=>"111011011",
  34548=>"111111111",
  34549=>"111001000",
  34550=>"100110000",
  34551=>"000111111",
  34552=>"000000000",
  34553=>"100100100",
  34554=>"111101111",
  34555=>"000000000",
  34556=>"111111010",
  34557=>"000001111",
  34558=>"011000110",
  34559=>"111111100",
  34560=>"001011111",
  34561=>"001001001",
  34562=>"111111111",
  34563=>"000000000",
  34564=>"111111111",
  34565=>"111101000",
  34566=>"000000000",
  34567=>"000000111",
  34568=>"111111010",
  34569=>"000000000",
  34570=>"000000000",
  34571=>"111111011",
  34572=>"111111111",
  34573=>"000000110",
  34574=>"000000000",
  34575=>"000000010",
  34576=>"011011111",
  34577=>"100100000",
  34578=>"001001001",
  34579=>"010111111",
  34580=>"010000011",
  34581=>"000111111",
  34582=>"011001001",
  34583=>"111110000",
  34584=>"111001101",
  34585=>"111111111",
  34586=>"001000000",
  34587=>"000000000",
  34588=>"000111111",
  34589=>"000000000",
  34590=>"000010000",
  34591=>"111111111",
  34592=>"011000000",
  34593=>"111101000",
  34594=>"000000000",
  34595=>"111000110",
  34596=>"110100000",
  34597=>"111001000",
  34598=>"111011111",
  34599=>"111011110",
  34600=>"010110011",
  34601=>"111111111",
  34602=>"000110110",
  34603=>"110111000",
  34604=>"111100111",
  34605=>"110000001",
  34606=>"100000000",
  34607=>"111000000",
  34608=>"111111001",
  34609=>"000000111",
  34610=>"111111111",
  34611=>"111111111",
  34612=>"000100000",
  34613=>"111111111",
  34614=>"111101000",
  34615=>"000111011",
  34616=>"111111111",
  34617=>"000000010",
  34618=>"001000100",
  34619=>"110010000",
  34620=>"000000000",
  34621=>"111000110",
  34622=>"110100111",
  34623=>"111111111",
  34624=>"000000000",
  34625=>"111111110",
  34626=>"000000000",
  34627=>"000000000",
  34628=>"000000000",
  34629=>"111111000",
  34630=>"000000010",
  34631=>"011111111",
  34632=>"111000000",
  34633=>"111111000",
  34634=>"011011000",
  34635=>"111111000",
  34636=>"111011000",
  34637=>"000000000",
  34638=>"011000000",
  34639=>"010010010",
  34640=>"010000000",
  34641=>"000000000",
  34642=>"000000000",
  34643=>"101111110",
  34644=>"010000011",
  34645=>"011111111",
  34646=>"111000010",
  34647=>"111000000",
  34648=>"111111111",
  34649=>"011001001",
  34650=>"000011111",
  34651=>"000000000",
  34652=>"100100100",
  34653=>"000000000",
  34654=>"000011000",
  34655=>"111111111",
  34656=>"011000000",
  34657=>"111000000",
  34658=>"001011100",
  34659=>"111011000",
  34660=>"011011011",
  34661=>"000000000",
  34662=>"000000011",
  34663=>"011000010",
  34664=>"001000000",
  34665=>"000000000",
  34666=>"000000111",
  34667=>"100100000",
  34668=>"111111001",
  34669=>"000000011",
  34670=>"100100000",
  34671=>"000000000",
  34672=>"111111110",
  34673=>"000000000",
  34674=>"001111110",
  34675=>"100110111",
  34676=>"000000000",
  34677=>"111111111",
  34678=>"100110111",
  34679=>"111100100",
  34680=>"001000000",
  34681=>"110111000",
  34682=>"111111111",
  34683=>"000000000",
  34684=>"010111111",
  34685=>"000010111",
  34686=>"000000011",
  34687=>"000000000",
  34688=>"100000000",
  34689=>"000110001",
  34690=>"110100100",
  34691=>"111111111",
  34692=>"000000010",
  34693=>"111111111",
  34694=>"111110111",
  34695=>"110110011",
  34696=>"001001001",
  34697=>"111100111",
  34698=>"001011000",
  34699=>"000000111",
  34700=>"011010110",
  34701=>"111101101",
  34702=>"111011000",
  34703=>"111111111",
  34704=>"101000100",
  34705=>"000000000",
  34706=>"111111000",
  34707=>"000000000",
  34708=>"000000000",
  34709=>"000001000",
  34710=>"010001001",
  34711=>"011111110",
  34712=>"110100000",
  34713=>"111110100",
  34714=>"111111111",
  34715=>"111111011",
  34716=>"000000110",
  34717=>"111111111",
  34718=>"110110111",
  34719=>"000100111",
  34720=>"000000000",
  34721=>"011000010",
  34722=>"000000000",
  34723=>"111111111",
  34724=>"111111011",
  34725=>"110111111",
  34726=>"111111111",
  34727=>"111000000",
  34728=>"111111001",
  34729=>"000110110",
  34730=>"111000111",
  34731=>"101000000",
  34732=>"111111111",
  34733=>"111101111",
  34734=>"111111111",
  34735=>"111001011",
  34736=>"000110111",
  34737=>"000000000",
  34738=>"011000110",
  34739=>"000000000",
  34740=>"000001001",
  34741=>"111111110",
  34742=>"111111001",
  34743=>"111111111",
  34744=>"011000000",
  34745=>"001111101",
  34746=>"111100000",
  34747=>"111111011",
  34748=>"101101101",
  34749=>"000000000",
  34750=>"111101000",
  34751=>"011011101",
  34752=>"001000000",
  34753=>"100000000",
  34754=>"000000000",
  34755=>"110111010",
  34756=>"101000110",
  34757=>"001001010",
  34758=>"111111111",
  34759=>"100100100",
  34760=>"000000111",
  34761=>"111100110",
  34762=>"001001000",
  34763=>"111000000",
  34764=>"111000000",
  34765=>"001000001",
  34766=>"110110000",
  34767=>"110000000",
  34768=>"111000000",
  34769=>"001000000",
  34770=>"011101111",
  34771=>"000000000",
  34772=>"110111110",
  34773=>"111111111",
  34774=>"111000000",
  34775=>"111111000",
  34776=>"001101001",
  34777=>"001111111",
  34778=>"110111111",
  34779=>"011101100",
  34780=>"000000000",
  34781=>"000000000",
  34782=>"111111111",
  34783=>"011011110",
  34784=>"111111111",
  34785=>"000000000",
  34786=>"111111011",
  34787=>"111111100",
  34788=>"000000010",
  34789=>"100000110",
  34790=>"111001111",
  34791=>"101000000",
  34792=>"000110111",
  34793=>"111011001",
  34794=>"010010000",
  34795=>"000000000",
  34796=>"000000000",
  34797=>"000110111",
  34798=>"111111111",
  34799=>"000000000",
  34800=>"000110111",
  34801=>"111111111",
  34802=>"000000011",
  34803=>"000000001",
  34804=>"111011111",
  34805=>"010111000",
  34806=>"011011111",
  34807=>"110110110",
  34808=>"000000001",
  34809=>"110111111",
  34810=>"111111111",
  34811=>"110000001",
  34812=>"000000000",
  34813=>"000000000",
  34814=>"000000000",
  34815=>"111111001",
  34816=>"111111111",
  34817=>"111111100",
  34818=>"000000000",
  34819=>"000000000",
  34820=>"111000000",
  34821=>"100000000",
  34822=>"111111111",
  34823=>"011001001",
  34824=>"011000000",
  34825=>"110111111",
  34826=>"000000000",
  34827=>"001000010",
  34828=>"011001000",
  34829=>"001000100",
  34830=>"111111111",
  34831=>"111111111",
  34832=>"110111011",
  34833=>"111110111",
  34834=>"000000000",
  34835=>"100110100",
  34836=>"000000111",
  34837=>"111011000",
  34838=>"000111111",
  34839=>"001011111",
  34840=>"111111111",
  34841=>"110101101",
  34842=>"011111110",
  34843=>"110111111",
  34844=>"111111001",
  34845=>"111111111",
  34846=>"110111100",
  34847=>"000000000",
  34848=>"101111111",
  34849=>"111011000",
  34850=>"111001001",
  34851=>"100100000",
  34852=>"111101101",
  34853=>"111111111",
  34854=>"001100100",
  34855=>"000000000",
  34856=>"111011011",
  34857=>"111101111",
  34858=>"111011001",
  34859=>"111111111",
  34860=>"111110111",
  34861=>"000000000",
  34862=>"111100111",
  34863=>"111101110",
  34864=>"000100100",
  34865=>"111101101",
  34866=>"101110111",
  34867=>"000000000",
  34868=>"000000001",
  34869=>"000100000",
  34870=>"001000101",
  34871=>"110000000",
  34872=>"000000000",
  34873=>"011111111",
  34874=>"000000000",
  34875=>"000000000",
  34876=>"000000000",
  34877=>"000111111",
  34878=>"110110111",
  34879=>"000001000",
  34880=>"001001111",
  34881=>"110000010",
  34882=>"111111111",
  34883=>"111110111",
  34884=>"111111111",
  34885=>"001001011",
  34886=>"111111000",
  34887=>"111111111",
  34888=>"001011001",
  34889=>"111110110",
  34890=>"000000000",
  34891=>"011011111",
  34892=>"000000000",
  34893=>"000000000",
  34894=>"000000000",
  34895=>"010011011",
  34896=>"010110000",
  34897=>"110110111",
  34898=>"111111111",
  34899=>"000000001",
  34900=>"001000000",
  34901=>"111111111",
  34902=>"110110000",
  34903=>"111111111",
  34904=>"110110111",
  34905=>"111111111",
  34906=>"111111111",
  34907=>"010000000",
  34908=>"101101001",
  34909=>"000000000",
  34910=>"000100100",
  34911=>"111111111",
  34912=>"011000000",
  34913=>"110111110",
  34914=>"111001011",
  34915=>"111111111",
  34916=>"010000000",
  34917=>"001011111",
  34918=>"111111000",
  34919=>"011011110",
  34920=>"100111111",
  34921=>"111111111",
  34922=>"001001000",
  34923=>"010110010",
  34924=>"001001100",
  34925=>"111100111",
  34926=>"111111010",
  34927=>"111111111",
  34928=>"000000000",
  34929=>"110111000",
  34930=>"110011011",
  34931=>"000000000",
  34932=>"111101101",
  34933=>"111111011",
  34934=>"111111010",
  34935=>"001000000",
  34936=>"111111111",
  34937=>"000001001",
  34938=>"111001000",
  34939=>"000000100",
  34940=>"110110000",
  34941=>"000001000",
  34942=>"000000000",
  34943=>"111111111",
  34944=>"110100100",
  34945=>"110001001",
  34946=>"000001100",
  34947=>"000000011",
  34948=>"111000111",
  34949=>"111110010",
  34950=>"110100000",
  34951=>"000000000",
  34952=>"000000011",
  34953=>"100110010",
  34954=>"000000000",
  34955=>"011111111",
  34956=>"111101111",
  34957=>"111111111",
  34958=>"111110000",
  34959=>"001000000",
  34960=>"000000000",
  34961=>"000011011",
  34962=>"100000001",
  34963=>"111111111",
  34964=>"001000100",
  34965=>"111010000",
  34966=>"000000000",
  34967=>"000000000",
  34968=>"001001101",
  34969=>"000100101",
  34970=>"000000111",
  34971=>"010110010",
  34972=>"111111001",
  34973=>"000000000",
  34974=>"111111111",
  34975=>"111011000",
  34976=>"111101111",
  34977=>"100000000",
  34978=>"010011111",
  34979=>"000000100",
  34980=>"000000000",
  34981=>"011011011",
  34982=>"000000000",
  34983=>"001000000",
  34984=>"100111111",
  34985=>"011111110",
  34986=>"000111111",
  34987=>"000000000",
  34988=>"100101111",
  34989=>"111111110",
  34990=>"111111111",
  34991=>"111111111",
  34992=>"111111111",
  34993=>"111111101",
  34994=>"000000000",
  34995=>"110000000",
  34996=>"000011110",
  34997=>"111111001",
  34998=>"011011000",
  34999=>"000011111",
  35000=>"100100000",
  35001=>"111111000",
  35002=>"000000111",
  35003=>"000111001",
  35004=>"011011001",
  35005=>"001010001",
  35006=>"111110100",
  35007=>"000000011",
  35008=>"011001000",
  35009=>"101101001",
  35010=>"100111011",
  35011=>"011000000",
  35012=>"110010000",
  35013=>"011011000",
  35014=>"111111101",
  35015=>"111110111",
  35016=>"011001111",
  35017=>"110110100",
  35018=>"000010111",
  35019=>"011111111",
  35020=>"000000010",
  35021=>"111111000",
  35022=>"000000000",
  35023=>"000010110",
  35024=>"000010010",
  35025=>"110100000",
  35026=>"111110010",
  35027=>"001000000",
  35028=>"001001001",
  35029=>"011011001",
  35030=>"000000000",
  35031=>"000000111",
  35032=>"000000000",
  35033=>"010010000",
  35034=>"111111111",
  35035=>"011111000",
  35036=>"111000000",
  35037=>"000000000",
  35038=>"011011111",
  35039=>"011001000",
  35040=>"110000000",
  35041=>"110110110",
  35042=>"000000000",
  35043=>"011111110",
  35044=>"000000000",
  35045=>"101100101",
  35046=>"001000000",
  35047=>"001001001",
  35048=>"111111111",
  35049=>"001011111",
  35050=>"111111111",
  35051=>"001000111",
  35052=>"001011011",
  35053=>"111001001",
  35054=>"011111111",
  35055=>"011111010",
  35056=>"111111001",
  35057=>"111111100",
  35058=>"111111111",
  35059=>"100000000",
  35060=>"111111111",
  35061=>"011110000",
  35062=>"001011111",
  35063=>"111111111",
  35064=>"101111111",
  35065=>"000000000",
  35066=>"000000000",
  35067=>"110111111",
  35068=>"001000001",
  35069=>"000110100",
  35070=>"001011110",
  35071=>"001000000",
  35072=>"001001000",
  35073=>"010010010",
  35074=>"000000000",
  35075=>"011111011",
  35076=>"111111111",
  35077=>"111000000",
  35078=>"111111111",
  35079=>"111011011",
  35080=>"111111111",
  35081=>"111111111",
  35082=>"000000000",
  35083=>"000000000",
  35084=>"110100000",
  35085=>"011111111",
  35086=>"111111100",
  35087=>"001111111",
  35088=>"000000100",
  35089=>"001000000",
  35090=>"000000000",
  35091=>"010000000",
  35092=>"001001111",
  35093=>"111111110",
  35094=>"000000011",
  35095=>"101001011",
  35096=>"111111111",
  35097=>"000000100",
  35098=>"000000000",
  35099=>"001001001",
  35100=>"111111111",
  35101=>"000000000",
  35102=>"111111111",
  35103=>"001011011",
  35104=>"000000000",
  35105=>"110010010",
  35106=>"111111111",
  35107=>"011001100",
  35108=>"000000100",
  35109=>"111111111",
  35110=>"000100100",
  35111=>"011011111",
  35112=>"111111111",
  35113=>"111111111",
  35114=>"110111111",
  35115=>"111111101",
  35116=>"111111110",
  35117=>"110110111",
  35118=>"001000000",
  35119=>"000000001",
  35120=>"011010000",
  35121=>"000000000",
  35122=>"001001000",
  35123=>"000000011",
  35124=>"111110000",
  35125=>"010000001",
  35126=>"011111111",
  35127=>"100000000",
  35128=>"111000000",
  35129=>"111110111",
  35130=>"000001001",
  35131=>"001111111",
  35132=>"000000011",
  35133=>"000000000",
  35134=>"000000000",
  35135=>"111111000",
  35136=>"000110110",
  35137=>"100100000",
  35138=>"000000000",
  35139=>"001000000",
  35140=>"111111111",
  35141=>"111111100",
  35142=>"111111111",
  35143=>"001000001",
  35144=>"000000000",
  35145=>"111111000",
  35146=>"111111100",
  35147=>"110100111",
  35148=>"000000000",
  35149=>"111111001",
  35150=>"111111111",
  35151=>"001111111",
  35152=>"001001011",
  35153=>"000000011",
  35154=>"111111111",
  35155=>"111111111",
  35156=>"111111110",
  35157=>"011011011",
  35158=>"111111100",
  35159=>"010011000",
  35160=>"001000100",
  35161=>"000010000",
  35162=>"111111011",
  35163=>"000010110",
  35164=>"111111111",
  35165=>"000000000",
  35166=>"000000000",
  35167=>"111111110",
  35168=>"110111000",
  35169=>"011111111",
  35170=>"011000111",
  35171=>"000000000",
  35172=>"111001111",
  35173=>"001011111",
  35174=>"010000100",
  35175=>"001001001",
  35176=>"011001001",
  35177=>"111000000",
  35178=>"111111000",
  35179=>"000000111",
  35180=>"000000000",
  35181=>"000111001",
  35182=>"011001000",
  35183=>"000000000",
  35184=>"000000000",
  35185=>"000011011",
  35186=>"000000000",
  35187=>"010100001",
  35188=>"000000011",
  35189=>"101011000",
  35190=>"001011001",
  35191=>"100100100",
  35192=>"111111111",
  35193=>"111111111",
  35194=>"000011111",
  35195=>"001011011",
  35196=>"111111110",
  35197=>"000000000",
  35198=>"111111000",
  35199=>"000001000",
  35200=>"111111000",
  35201=>"000110110",
  35202=>"010111111",
  35203=>"100100100",
  35204=>"111111111",
  35205=>"000000000",
  35206=>"010111111",
  35207=>"011111111",
  35208=>"100000000",
  35209=>"011011011",
  35210=>"001100100",
  35211=>"111110000",
  35212=>"111111111",
  35213=>"010010000",
  35214=>"011011001",
  35215=>"100000110",
  35216=>"010110110",
  35217=>"111111111",
  35218=>"111011010",
  35219=>"000000000",
  35220=>"111111010",
  35221=>"000000000",
  35222=>"000000000",
  35223=>"000000100",
  35224=>"000000000",
  35225=>"110111111",
  35226=>"111110110",
  35227=>"110111111",
  35228=>"111111111",
  35229=>"000000000",
  35230=>"011011111",
  35231=>"111111111",
  35232=>"111111001",
  35233=>"011011011",
  35234=>"000010010",
  35235=>"000100100",
  35236=>"111111111",
  35237=>"010111000",
  35238=>"100110110",
  35239=>"000000111",
  35240=>"100110100",
  35241=>"011001101",
  35242=>"000110111",
  35243=>"000000011",
  35244=>"110000110",
  35245=>"111111110",
  35246=>"000000100",
  35247=>"111111111",
  35248=>"011000000",
  35249=>"011001001",
  35250=>"000000000",
  35251=>"001111111",
  35252=>"000000100",
  35253=>"111111111",
  35254=>"111111111",
  35255=>"111001001",
  35256=>"111001000",
  35257=>"110111111",
  35258=>"001000001",
  35259=>"101101100",
  35260=>"000000000",
  35261=>"111101111",
  35262=>"110110110",
  35263=>"000000000",
  35264=>"000000000",
  35265=>"011011001",
  35266=>"000000000",
  35267=>"000000000",
  35268=>"100110000",
  35269=>"100100000",
  35270=>"010110100",
  35271=>"100111000",
  35272=>"000000000",
  35273=>"001111111",
  35274=>"110110100",
  35275=>"100111100",
  35276=>"001111000",
  35277=>"000001000",
  35278=>"111111000",
  35279=>"111111111",
  35280=>"110100000",
  35281=>"100100100",
  35282=>"110110000",
  35283=>"111111111",
  35284=>"110110111",
  35285=>"000000000",
  35286=>"111110100",
  35287=>"000000100",
  35288=>"000000000",
  35289=>"000110010",
  35290=>"111010000",
  35291=>"111111100",
  35292=>"111011011",
  35293=>"111111011",
  35294=>"100000000",
  35295=>"000000000",
  35296=>"010000000",
  35297=>"111111111",
  35298=>"001001011",
  35299=>"111000001",
  35300=>"000000000",
  35301=>"000001001",
  35302=>"110110000",
  35303=>"110010110",
  35304=>"111111111",
  35305=>"011111101",
  35306=>"111000101",
  35307=>"111101001",
  35308=>"000000000",
  35309=>"111111111",
  35310=>"000100100",
  35311=>"110110101",
  35312=>"000001001",
  35313=>"111111111",
  35314=>"110110111",
  35315=>"111010000",
  35316=>"000001111",
  35317=>"000000000",
  35318=>"000000000",
  35319=>"011011000",
  35320=>"000000000",
  35321=>"001101101",
  35322=>"111001111",
  35323=>"000000111",
  35324=>"111111000",
  35325=>"111111111",
  35326=>"000110111",
  35327=>"111111011",
  35328=>"000001001",
  35329=>"110111110",
  35330=>"111111111",
  35331=>"000000000",
  35332=>"110111111",
  35333=>"011011000",
  35334=>"100000000",
  35335=>"000000000",
  35336=>"100100000",
  35337=>"111111011",
  35338=>"001111111",
  35339=>"100000111",
  35340=>"000110110",
  35341=>"001001001",
  35342=>"000011011",
  35343=>"110111110",
  35344=>"110010110",
  35345=>"000000000",
  35346=>"000000000",
  35347=>"110111111",
  35348=>"111011001",
  35349=>"111111101",
  35350=>"111111110",
  35351=>"011111110",
  35352=>"000000100",
  35353=>"111111111",
  35354=>"000000000",
  35355=>"000100111",
  35356=>"111111111",
  35357=>"111111100",
  35358=>"100100100",
  35359=>"110110110",
  35360=>"000000000",
  35361=>"010111111",
  35362=>"001001000",
  35363=>"000000000",
  35364=>"000000000",
  35365=>"000000000",
  35366=>"000110111",
  35367=>"111100100",
  35368=>"000000000",
  35369=>"001011001",
  35370=>"000000000",
  35371=>"111100110",
  35372=>"001000100",
  35373=>"000000000",
  35374=>"000000000",
  35375=>"000110110",
  35376=>"000000111",
  35377=>"000000000",
  35378=>"011011011",
  35379=>"000000000",
  35380=>"100110111",
  35381=>"111111111",
  35382=>"110111111",
  35383=>"000010011",
  35384=>"111111111",
  35385=>"110010111",
  35386=>"111111111",
  35387=>"011111111",
  35388=>"000000000",
  35389=>"000001111",
  35390=>"000010100",
  35391=>"111110000",
  35392=>"000000000",
  35393=>"100000000",
  35394=>"100111111",
  35395=>"000000000",
  35396=>"110110110",
  35397=>"000001001",
  35398=>"000000000",
  35399=>"000001001",
  35400=>"011111011",
  35401=>"111001100",
  35402=>"010110111",
  35403=>"010111111",
  35404=>"000000111",
  35405=>"001100111",
  35406=>"111111101",
  35407=>"000110111",
  35408=>"011010000",
  35409=>"011011011",
  35410=>"000000000",
  35411=>"000000000",
  35412=>"111111111",
  35413=>"011011010",
  35414=>"000111111",
  35415=>"110110010",
  35416=>"000101111",
  35417=>"111001000",
  35418=>"111111110",
  35419=>"111110110",
  35420=>"000000000",
  35421=>"110111111",
  35422=>"000000000",
  35423=>"011000000",
  35424=>"000000000",
  35425=>"011111101",
  35426=>"000010000",
  35427=>"110111111",
  35428=>"111111100",
  35429=>"111111101",
  35430=>"001100100",
  35431=>"110100100",
  35432=>"000000000",
  35433=>"111111111",
  35434=>"111001011",
  35435=>"010110111",
  35436=>"000000100",
  35437=>"110101011",
  35438=>"010010110",
  35439=>"000000000",
  35440=>"111111000",
  35441=>"000001011",
  35442=>"111111111",
  35443=>"000011011",
  35444=>"011010011",
  35445=>"111111111",
  35446=>"000000000",
  35447=>"000000000",
  35448=>"011001001",
  35449=>"000010111",
  35450=>"101000000",
  35451=>"111111101",
  35452=>"100110100",
  35453=>"001001000",
  35454=>"110100000",
  35455=>"000110100",
  35456=>"011001000",
  35457=>"111110110",
  35458=>"000111111",
  35459=>"000000100",
  35460=>"000100111",
  35461=>"000000011",
  35462=>"001001000",
  35463=>"000000000",
  35464=>"011111111",
  35465=>"111111111",
  35466=>"000000000",
  35467=>"111111111",
  35468=>"101101111",
  35469=>"111111110",
  35470=>"111111101",
  35471=>"100100000",
  35472=>"001101101",
  35473=>"101101101",
  35474=>"011001000",
  35475=>"000000100",
  35476=>"000000000",
  35477=>"000100111",
  35478=>"001000000",
  35479=>"110111101",
  35480=>"000000000",
  35481=>"100110110",
  35482=>"000000010",
  35483=>"100000000",
  35484=>"111011000",
  35485=>"011111111",
  35486=>"001111111",
  35487=>"000000000",
  35488=>"111100000",
  35489=>"111111111",
  35490=>"111111111",
  35491=>"111110010",
  35492=>"000111111",
  35493=>"011000100",
  35494=>"111111111",
  35495=>"100100100",
  35496=>"011000000",
  35497=>"000000000",
  35498=>"110000000",
  35499=>"111111111",
  35500=>"001000000",
  35501=>"100111101",
  35502=>"000110111",
  35503=>"000011111",
  35504=>"000001001",
  35505=>"111110111",
  35506=>"010011011",
  35507=>"000000110",
  35508=>"000000100",
  35509=>"000000000",
  35510=>"001000000",
  35511=>"000000000",
  35512=>"000000011",
  35513=>"101101000",
  35514=>"000111111",
  35515=>"011110000",
  35516=>"111010011",
  35517=>"011111111",
  35518=>"111011011",
  35519=>"110100000",
  35520=>"000000000",
  35521=>"000001111",
  35522=>"011011001",
  35523=>"000010011",
  35524=>"011111111",
  35525=>"010011111",
  35526=>"001001001",
  35527=>"110110110",
  35528=>"111100111",
  35529=>"000001001",
  35530=>"100000000",
  35531=>"000010000",
  35532=>"111111111",
  35533=>"011010111",
  35534=>"000110110",
  35535=>"111000000",
  35536=>"011111111",
  35537=>"000000000",
  35538=>"000111101",
  35539=>"111110010",
  35540=>"000001001",
  35541=>"000000100",
  35542=>"111010000",
  35543=>"011000100",
  35544=>"011011001",
  35545=>"001001001",
  35546=>"011001100",
  35547=>"111011001",
  35548=>"001100110",
  35549=>"001001111",
  35550=>"111111111",
  35551=>"000011011",
  35552=>"000001111",
  35553=>"000000000",
  35554=>"010010111",
  35555=>"110010000",
  35556=>"111111111",
  35557=>"111111111",
  35558=>"110110110",
  35559=>"100110111",
  35560=>"111111110",
  35561=>"000101111",
  35562=>"101111111",
  35563=>"000111111",
  35564=>"000111111",
  35565=>"000010011",
  35566=>"000000011",
  35567=>"000000011",
  35568=>"111111111",
  35569=>"000000000",
  35570=>"011000000",
  35571=>"000001111",
  35572=>"111111111",
  35573=>"111000000",
  35574=>"100000100",
  35575=>"111110000",
  35576=>"000000010",
  35577=>"000000000",
  35578=>"000000001",
  35579=>"011001111",
  35580=>"110110100",
  35581=>"001100000",
  35582=>"111110111",
  35583=>"100000110",
  35584=>"000011001",
  35585=>"100000000",
  35586=>"111100100",
  35587=>"111011010",
  35588=>"111111001",
  35589=>"001001111",
  35590=>"000110111",
  35591=>"111111111",
  35592=>"000110111",
  35593=>"111111010",
  35594=>"000000000",
  35595=>"111111111",
  35596=>"101111111",
  35597=>"001000000",
  35598=>"000000001",
  35599=>"000010111",
  35600=>"110100100",
  35601=>"000000001",
  35602=>"101100101",
  35603=>"111111100",
  35604=>"100001000",
  35605=>"111111011",
  35606=>"111111111",
  35607=>"000000001",
  35608=>"000000001",
  35609=>"110101110",
  35610=>"010011011",
  35611=>"000000001",
  35612=>"111111110",
  35613=>"000011100",
  35614=>"001001000",
  35615=>"010110100",
  35616=>"001001000",
  35617=>"101111110",
  35618=>"000000011",
  35619=>"011111011",
  35620=>"011011011",
  35621=>"000000000",
  35622=>"000111101",
  35623=>"010110000",
  35624=>"111011110",
  35625=>"110100110",
  35626=>"011100000",
  35627=>"111111111",
  35628=>"011110111",
  35629=>"001001000",
  35630=>"000111001",
  35631=>"000000010",
  35632=>"111011011",
  35633=>"000110110",
  35634=>"000000000",
  35635=>"010010100",
  35636=>"011001011",
  35637=>"000000000",
  35638=>"011011000",
  35639=>"111111011",
  35640=>"000001001",
  35641=>"111111111",
  35642=>"011111000",
  35643=>"000100101",
  35644=>"110010010",
  35645=>"111111111",
  35646=>"010000100",
  35647=>"110111111",
  35648=>"001111101",
  35649=>"110110110",
  35650=>"111111011",
  35651=>"111100000",
  35652=>"000011110",
  35653=>"111011001",
  35654=>"000000000",
  35655=>"000000100",
  35656=>"000000000",
  35657=>"000000010",
  35658=>"011000000",
  35659=>"011110000",
  35660=>"111011111",
  35661=>"111111111",
  35662=>"000100101",
  35663=>"111111111",
  35664=>"011011001",
  35665=>"110111111",
  35666=>"100010000",
  35667=>"000000101",
  35668=>"000000000",
  35669=>"011011001",
  35670=>"000000000",
  35671=>"111111111",
  35672=>"000000001",
  35673=>"000000111",
  35674=>"000000000",
  35675=>"000000111",
  35676=>"011111111",
  35677=>"000000000",
  35678=>"011001001",
  35679=>"111011010",
  35680=>"000000000",
  35681=>"111111111",
  35682=>"000000001",
  35683=>"000000000",
  35684=>"000001001",
  35685=>"000000000",
  35686=>"010000010",
  35687=>"001011000",
  35688=>"110110111",
  35689=>"000010111",
  35690=>"000000000",
  35691=>"111111000",
  35692=>"001001001",
  35693=>"000000110",
  35694=>"111111110",
  35695=>"001011000",
  35696=>"000000000",
  35697=>"000000101",
  35698=>"001001111",
  35699=>"000000000",
  35700=>"001000000",
  35701=>"000100100",
  35702=>"111100110",
  35703=>"111111111",
  35704=>"011000000",
  35705=>"111111010",
  35706=>"111001001",
  35707=>"111111010",
  35708=>"000000000",
  35709=>"111111111",
  35710=>"000000000",
  35711=>"111111111",
  35712=>"000000110",
  35713=>"111111001",
  35714=>"000000000",
  35715=>"111101000",
  35716=>"000011111",
  35717=>"011111111",
  35718=>"111011111",
  35719=>"000000000",
  35720=>"111101101",
  35721=>"000000110",
  35722=>"000110111",
  35723=>"111111111",
  35724=>"011000000",
  35725=>"100111111",
  35726=>"110111111",
  35727=>"000000000",
  35728=>"000000000",
  35729=>"110110110",
  35730=>"000000011",
  35731=>"111110110",
  35732=>"001000000",
  35733=>"000000000",
  35734=>"000000110",
  35735=>"001001001",
  35736=>"000000111",
  35737=>"001000000",
  35738=>"000000000",
  35739=>"010111111",
  35740=>"011010110",
  35741=>"111111110",
  35742=>"001001101",
  35743=>"000000000",
  35744=>"100100100",
  35745=>"011011001",
  35746=>"000110100",
  35747=>"111111111",
  35748=>"010110000",
  35749=>"000000000",
  35750=>"001001001",
  35751=>"111111000",
  35752=>"000000000",
  35753=>"011111110",
  35754=>"000000001",
  35755=>"001001001",
  35756=>"000000000",
  35757=>"000000110",
  35758=>"110111111",
  35759=>"111111111",
  35760=>"100111111",
  35761=>"010010111",
  35762=>"011111111",
  35763=>"000111111",
  35764=>"000000000",
  35765=>"010010000",
  35766=>"111101001",
  35767=>"111000111",
  35768=>"111111111",
  35769=>"000110111",
  35770=>"001111110",
  35771=>"001001001",
  35772=>"000111111",
  35773=>"111100000",
  35774=>"001111111",
  35775=>"111000000",
  35776=>"000001000",
  35777=>"111011001",
  35778=>"110110010",
  35779=>"000111110",
  35780=>"001001111",
  35781=>"011110110",
  35782=>"000000000",
  35783=>"111011000",
  35784=>"000001011",
  35785=>"111111001",
  35786=>"101000001",
  35787=>"111111111",
  35788=>"010011000",
  35789=>"000000000",
  35790=>"000000000",
  35791=>"000000000",
  35792=>"001000001",
  35793=>"001000000",
  35794=>"111111111",
  35795=>"111111001",
  35796=>"111111111",
  35797=>"111111010",
  35798=>"001000000",
  35799=>"011011000",
  35800=>"111111111",
  35801=>"111111000",
  35802=>"100111000",
  35803=>"111111111",
  35804=>"010001000",
  35805=>"001111001",
  35806=>"000011111",
  35807=>"000100011",
  35808=>"011001111",
  35809=>"111111111",
  35810=>"000000000",
  35811=>"111111111",
  35812=>"110110111",
  35813=>"111111111",
  35814=>"000001011",
  35815=>"011011000",
  35816=>"111110100",
  35817=>"000000010",
  35818=>"000110111",
  35819=>"000010000",
  35820=>"111111111",
  35821=>"000000100",
  35822=>"110110111",
  35823=>"011011101",
  35824=>"001000100",
  35825=>"010111111",
  35826=>"000000111",
  35827=>"000011111",
  35828=>"000001001",
  35829=>"000000000",
  35830=>"110110000",
  35831=>"110110100",
  35832=>"001011010",
  35833=>"001101101",
  35834=>"000111111",
  35835=>"011010000",
  35836=>"010000000",
  35837=>"100000010",
  35838=>"000001010",
  35839=>"000001111",
  35840=>"011001001",
  35841=>"101111111",
  35842=>"000000111",
  35843=>"110111111",
  35844=>"001001001",
  35845=>"111111111",
  35846=>"010111000",
  35847=>"000000000",
  35848=>"000000001",
  35849=>"001111110",
  35850=>"111111111",
  35851=>"011111111",
  35852=>"110110110",
  35853=>"000000001",
  35854=>"000000111",
  35855=>"000000000",
  35856=>"000111111",
  35857=>"000010101",
  35858=>"010110111",
  35859=>"110100000",
  35860=>"001000000",
  35861=>"000111110",
  35862=>"101100100",
  35863=>"111111111",
  35864=>"111111101",
  35865=>"011011011",
  35866=>"001000000",
  35867=>"000100100",
  35868=>"001001011",
  35869=>"101000000",
  35870=>"011011011",
  35871=>"011011010",
  35872=>"100100110",
  35873=>"001111111",
  35874=>"010111000",
  35875=>"111111110",
  35876=>"000000000",
  35877=>"110110000",
  35878=>"111111000",
  35879=>"011111000",
  35880=>"011001000",
  35881=>"000100100",
  35882=>"100101111",
  35883=>"001000000",
  35884=>"000111111",
  35885=>"000010000",
  35886=>"010110111",
  35887=>"000000000",
  35888=>"001001101",
  35889=>"111111110",
  35890=>"111100000",
  35891=>"000000111",
  35892=>"010110100",
  35893=>"110011011",
  35894=>"110000000",
  35895=>"000000000",
  35896=>"100111111",
  35897=>"000011011",
  35898=>"000111011",
  35899=>"111111111",
  35900=>"111111111",
  35901=>"000000001",
  35902=>"100100000",
  35903=>"111101111",
  35904=>"111001000",
  35905=>"000000101",
  35906=>"000110111",
  35907=>"000011111",
  35908=>"111111111",
  35909=>"010010000",
  35910=>"011111011",
  35911=>"111111110",
  35912=>"001001000",
  35913=>"000010010",
  35914=>"100000000",
  35915=>"101000000",
  35916=>"000011111",
  35917=>"110110110",
  35918=>"001000000",
  35919=>"110111111",
  35920=>"111011010",
  35921=>"111011011",
  35922=>"001000111",
  35923=>"000111000",
  35924=>"000011001",
  35925=>"100111001",
  35926=>"111111111",
  35927=>"001111000",
  35928=>"110111000",
  35929=>"111001111",
  35930=>"000000000",
  35931=>"001000000",
  35932=>"111011111",
  35933=>"100000100",
  35934=>"000000001",
  35935=>"000000000",
  35936=>"000000000",
  35937=>"000000010",
  35938=>"111001001",
  35939=>"111111111",
  35940=>"111010001",
  35941=>"000000111",
  35942=>"100111111",
  35943=>"000000000",
  35944=>"000000000",
  35945=>"111111011",
  35946=>"011111111",
  35947=>"010011111",
  35948=>"100111111",
  35949=>"101000111",
  35950=>"111111111",
  35951=>"000110000",
  35952=>"011011011",
  35953=>"000111111",
  35954=>"000000000",
  35955=>"101001011",
  35956=>"000000000",
  35957=>"000000000",
  35958=>"110110010",
  35959=>"100100111",
  35960=>"001001011",
  35961=>"001000000",
  35962=>"000000000",
  35963=>"001001011",
  35964=>"111110110",
  35965=>"111100110",
  35966=>"010111111",
  35967=>"111001111",
  35968=>"010011000",
  35969=>"111110010",
  35970=>"101000001",
  35971=>"100110000",
  35972=>"000000011",
  35973=>"111001001",
  35974=>"111111101",
  35975=>"101101110",
  35976=>"111111110",
  35977=>"000001001",
  35978=>"111111000",
  35979=>"010010010",
  35980=>"000000000",
  35981=>"101011000",
  35982=>"101101111",
  35983=>"000110110",
  35984=>"101001111",
  35985=>"111111111",
  35986=>"100000000",
  35987=>"110111110",
  35988=>"011010000",
  35989=>"101001001",
  35990=>"000000000",
  35991=>"101000000",
  35992=>"101000100",
  35993=>"111111111",
  35994=>"000100111",
  35995=>"000110100",
  35996=>"111110111",
  35997=>"001000001",
  35998=>"000000011",
  35999=>"111010000",
  36000=>"110010111",
  36001=>"000111111",
  36002=>"110110111",
  36003=>"100001000",
  36004=>"110100001",
  36005=>"000010000",
  36006=>"101001000",
  36007=>"000000000",
  36008=>"101100111",
  36009=>"001001111",
  36010=>"000000000",
  36011=>"001000000",
  36012=>"000100100",
  36013=>"000000000",
  36014=>"000000100",
  36015=>"100111111",
  36016=>"111111111",
  36017=>"111111001",
  36018=>"111111010",
  36019=>"000001111",
  36020=>"100000000",
  36021=>"001001000",
  36022=>"000010000",
  36023=>"000000000",
  36024=>"000000111",
  36025=>"001011111",
  36026=>"000000000",
  36027=>"110000101",
  36028=>"111100100",
  36029=>"111111001",
  36030=>"001000000",
  36031=>"110110110",
  36032=>"011101000",
  36033=>"101111111",
  36034=>"111111110",
  36035=>"111011011",
  36036=>"111110000",
  36037=>"000100100",
  36038=>"001111111",
  36039=>"111001000",
  36040=>"000000000",
  36041=>"111111111",
  36042=>"000000000",
  36043=>"111111111",
  36044=>"000001000",
  36045=>"111111111",
  36046=>"110110010",
  36047=>"110010111",
  36048=>"110100010",
  36049=>"000000000",
  36050=>"100100101",
  36051=>"000010000",
  36052=>"110100000",
  36053=>"101001111",
  36054=>"111111111",
  36055=>"111111000",
  36056=>"000000000",
  36057=>"111111111",
  36058=>"000111000",
  36059=>"001111111",
  36060=>"000000000",
  36061=>"001001001",
  36062=>"000000000",
  36063=>"111111001",
  36064=>"000000000",
  36065=>"000000000",
  36066=>"111010000",
  36067=>"111111100",
  36068=>"111011111",
  36069=>"000000000",
  36070=>"101111100",
  36071=>"000000001",
  36072=>"101100000",
  36073=>"001000000",
  36074=>"010111111",
  36075=>"100001000",
  36076=>"111111111",
  36077=>"000011111",
  36078=>"111000011",
  36079=>"111100000",
  36080=>"100000000",
  36081=>"011011011",
  36082=>"011011000",
  36083=>"010000000",
  36084=>"111111111",
  36085=>"101001000",
  36086=>"011011111",
  36087=>"111101111",
  36088=>"000000000",
  36089=>"111000010",
  36090=>"000000001",
  36091=>"111111111",
  36092=>"110110110",
  36093=>"111000100",
  36094=>"000000000",
  36095=>"000111111",
  36096=>"000000000",
  36097=>"101100100",
  36098=>"111111110",
  36099=>"111111111",
  36100=>"000111000",
  36101=>"001111111",
  36102=>"001001000",
  36103=>"000000100",
  36104=>"001111111",
  36105=>"001000000",
  36106=>"110100101",
  36107=>"110110010",
  36108=>"001111101",
  36109=>"000000000",
  36110=>"000111111",
  36111=>"111100000",
  36112=>"000000000",
  36113=>"110111111",
  36114=>"000001011",
  36115=>"001000110",
  36116=>"000101010",
  36117=>"000110110",
  36118=>"000000000",
  36119=>"111111000",
  36120=>"000000000",
  36121=>"101100000",
  36122=>"001000000",
  36123=>"000000110",
  36124=>"001101000",
  36125=>"110111111",
  36126=>"111111010",
  36127=>"111011111",
  36128=>"100000000",
  36129=>"111111010",
  36130=>"111111001",
  36131=>"100100000",
  36132=>"100100111",
  36133=>"101001001",
  36134=>"011111000",
  36135=>"000000100",
  36136=>"001000000",
  36137=>"000000000",
  36138=>"000110110",
  36139=>"000000000",
  36140=>"110111111",
  36141=>"000110000",
  36142=>"000000000",
  36143=>"000010000",
  36144=>"111111111",
  36145=>"000000100",
  36146=>"111011001",
  36147=>"000000110",
  36148=>"000111111",
  36149=>"111111011",
  36150=>"111111000",
  36151=>"010110010",
  36152=>"000010011",
  36153=>"110110000",
  36154=>"000000100",
  36155=>"000101111",
  36156=>"111111111",
  36157=>"010111111",
  36158=>"111111000",
  36159=>"000001111",
  36160=>"011000000",
  36161=>"001001001",
  36162=>"000101101",
  36163=>"001000000",
  36164=>"111111000",
  36165=>"000010011",
  36166=>"111111111",
  36167=>"110110110",
  36168=>"111111111",
  36169=>"000000110",
  36170=>"000110000",
  36171=>"101011011",
  36172=>"000000000",
  36173=>"000000100",
  36174=>"000000110",
  36175=>"111111111",
  36176=>"111001000",
  36177=>"000000010",
  36178=>"000000001",
  36179=>"110111111",
  36180=>"010010000",
  36181=>"001011011",
  36182=>"111111111",
  36183=>"000011111",
  36184=>"101111111",
  36185=>"000000001",
  36186=>"011011000",
  36187=>"011000000",
  36188=>"000000111",
  36189=>"000110100",
  36190=>"111111110",
  36191=>"111111011",
  36192=>"111111111",
  36193=>"111001000",
  36194=>"100000001",
  36195=>"000100000",
  36196=>"110110110",
  36197=>"111000011",
  36198=>"100000110",
  36199=>"110100000",
  36200=>"100110111",
  36201=>"111111011",
  36202=>"011000000",
  36203=>"001001000",
  36204=>"000001010",
  36205=>"001000110",
  36206=>"000000000",
  36207=>"111111000",
  36208=>"111111111",
  36209=>"111111111",
  36210=>"111111111",
  36211=>"001011000",
  36212=>"100101100",
  36213=>"000000000",
  36214=>"111111111",
  36215=>"100110000",
  36216=>"000000000",
  36217=>"000000000",
  36218=>"111011111",
  36219=>"001001000",
  36220=>"000000001",
  36221=>"000000001",
  36222=>"111011011",
  36223=>"111111111",
  36224=>"000000001",
  36225=>"001111001",
  36226=>"111111110",
  36227=>"111101000",
  36228=>"111100000",
  36229=>"111011001",
  36230=>"000000111",
  36231=>"000000000",
  36232=>"000000000",
  36233=>"111111110",
  36234=>"111001111",
  36235=>"000010111",
  36236=>"111110111",
  36237=>"111111001",
  36238=>"000000000",
  36239=>"000000000",
  36240=>"000000111",
  36241=>"000000111",
  36242=>"101110000",
  36243=>"111001000",
  36244=>"010110111",
  36245=>"000000000",
  36246=>"000000000",
  36247=>"110110100",
  36248=>"000101111",
  36249=>"110111011",
  36250=>"000111111",
  36251=>"000000000",
  36252=>"111100000",
  36253=>"111000111",
  36254=>"110000000",
  36255=>"111111111",
  36256=>"111111101",
  36257=>"101000000",
  36258=>"111111001",
  36259=>"100100100",
  36260=>"001000001",
  36261=>"000000010",
  36262=>"101000111",
  36263=>"101111001",
  36264=>"000000100",
  36265=>"100110111",
  36266=>"110110110",
  36267=>"010000000",
  36268=>"111111111",
  36269=>"000001111",
  36270=>"100000111",
  36271=>"000000111",
  36272=>"011000111",
  36273=>"101100000",
  36274=>"110111111",
  36275=>"111111110",
  36276=>"000000000",
  36277=>"110110110",
  36278=>"110111110",
  36279=>"111110000",
  36280=>"110111101",
  36281=>"110110111",
  36282=>"110110110",
  36283=>"111100111",
  36284=>"010111111",
  36285=>"101101101",
  36286=>"010111111",
  36287=>"001011111",
  36288=>"000000001",
  36289=>"111001111",
  36290=>"010111011",
  36291=>"111111000",
  36292=>"000000111",
  36293=>"011001101",
  36294=>"001000110",
  36295=>"001000111",
  36296=>"010000000",
  36297=>"001011000",
  36298=>"111110110",
  36299=>"000100111",
  36300=>"111111000",
  36301=>"111111111",
  36302=>"000001001",
  36303=>"111111011",
  36304=>"000111111",
  36305=>"111011111",
  36306=>"111111111",
  36307=>"111111110",
  36308=>"100001000",
  36309=>"110111111",
  36310=>"001000011",
  36311=>"011111011",
  36312=>"011001000",
  36313=>"010111011",
  36314=>"111101100",
  36315=>"000001111",
  36316=>"110000000",
  36317=>"100000000",
  36318=>"111100110",
  36319=>"001000011",
  36320=>"111111111",
  36321=>"001001000",
  36322=>"000000111",
  36323=>"000000111",
  36324=>"001011111",
  36325=>"000000000",
  36326=>"100000000",
  36327=>"111100100",
  36328=>"011000000",
  36329=>"111001000",
  36330=>"101111111",
  36331=>"111100000",
  36332=>"111101101",
  36333=>"000001001",
  36334=>"111011000",
  36335=>"111000000",
  36336=>"010111011",
  36337=>"000110111",
  36338=>"111111111",
  36339=>"000000111",
  36340=>"000000010",
  36341=>"000110111",
  36342=>"001001000",
  36343=>"111111111",
  36344=>"110110111",
  36345=>"001001001",
  36346=>"000000000",
  36347=>"110111110",
  36348=>"100000000",
  36349=>"111101100",
  36350=>"011110000",
  36351=>"011000000",
  36352=>"000000000",
  36353=>"111111111",
  36354=>"111111111",
  36355=>"111111111",
  36356=>"000110111",
  36357=>"000000000",
  36358=>"001001000",
  36359=>"100111111",
  36360=>"110000000",
  36361=>"111101111",
  36362=>"001111111",
  36363=>"111111111",
  36364=>"101101101",
  36365=>"000000000",
  36366=>"110111111",
  36367=>"011011011",
  36368=>"011001111",
  36369=>"000001001",
  36370=>"000000000",
  36371=>"111111111",
  36372=>"111111000",
  36373=>"001000000",
  36374=>"010111111",
  36375=>"111111111",
  36376=>"101011111",
  36377=>"111011111",
  36378=>"101000100",
  36379=>"001000111",
  36380=>"000000000",
  36381=>"011001011",
  36382=>"111011100",
  36383=>"001111101",
  36384=>"000010000",
  36385=>"011111111",
  36386=>"001000000",
  36387=>"111111111",
  36388=>"100110111",
  36389=>"001000111",
  36390=>"000000001",
  36391=>"111111111",
  36392=>"111101101",
  36393=>"000000000",
  36394=>"111111111",
  36395=>"111111111",
  36396=>"111111100",
  36397=>"000000111",
  36398=>"001001000",
  36399=>"000000100",
  36400=>"000000000",
  36401=>"000100101",
  36402=>"000001001",
  36403=>"000000000",
  36404=>"010000000",
  36405=>"000000000",
  36406=>"000000000",
  36407=>"111001111",
  36408=>"000000000",
  36409=>"101000000",
  36410=>"000000011",
  36411=>"000000000",
  36412=>"000111111",
  36413=>"000111011",
  36414=>"111111011",
  36415=>"000000000",
  36416=>"111000000",
  36417=>"101111011",
  36418=>"111111111",
  36419=>"100000000",
  36420=>"110110110",
  36421=>"010011001",
  36422=>"000000000",
  36423=>"111111111",
  36424=>"011010111",
  36425=>"000000011",
  36426=>"111111111",
  36427=>"110110110",
  36428=>"110100111",
  36429=>"000010110",
  36430=>"101000001",
  36431=>"001000000",
  36432=>"001000000",
  36433=>"000000111",
  36434=>"001001111",
  36435=>"011000001",
  36436=>"111101111",
  36437=>"111111011",
  36438=>"111111111",
  36439=>"010111011",
  36440=>"110111111",
  36441=>"000000010",
  36442=>"000011111",
  36443=>"001011001",
  36444=>"011111111",
  36445=>"111111010",
  36446=>"001000000",
  36447=>"011000000",
  36448=>"111111111",
  36449=>"111110110",
  36450=>"110100100",
  36451=>"111111111",
  36452=>"110110010",
  36453=>"100110000",
  36454=>"001011000",
  36455=>"000000000",
  36456=>"000110111",
  36457=>"101100110",
  36458=>"010110001",
  36459=>"000000111",
  36460=>"111110000",
  36461=>"111111011",
  36462=>"110100111",
  36463=>"010110010",
  36464=>"111111111",
  36465=>"100110000",
  36466=>"100000000",
  36467=>"000000111",
  36468=>"001000000",
  36469=>"000010111",
  36470=>"000111111",
  36471=>"000000100",
  36472=>"110111100",
  36473=>"000011011",
  36474=>"011001000",
  36475=>"000000110",
  36476=>"100100100",
  36477=>"001000000",
  36478=>"011111011",
  36479=>"111111010",
  36480=>"000000000",
  36481=>"111011111",
  36482=>"111110111",
  36483=>"110110100",
  36484=>"100000001",
  36485=>"000000000",
  36486=>"000000000",
  36487=>"011000000",
  36488=>"000000001",
  36489=>"111111111",
  36490=>"111111111",
  36491=>"000001101",
  36492=>"110111011",
  36493=>"000000000",
  36494=>"100000000",
  36495=>"101110111",
  36496=>"111101111",
  36497=>"101101111",
  36498=>"100111111",
  36499=>"111001101",
  36500=>"100001001",
  36501=>"111100000",
  36502=>"111111000",
  36503=>"110100100",
  36504=>"000000000",
  36505=>"001111111",
  36506=>"000000101",
  36507=>"111111100",
  36508=>"011111111",
  36509=>"001000001",
  36510=>"101100000",
  36511=>"110111111",
  36512=>"111111010",
  36513=>"100000111",
  36514=>"000000001",
  36515=>"000100100",
  36516=>"110111110",
  36517=>"011100110",
  36518=>"111111111",
  36519=>"110000000",
  36520=>"000000111",
  36521=>"000101100",
  36522=>"000000000",
  36523=>"111111111",
  36524=>"001000000",
  36525=>"111111111",
  36526=>"000000100",
  36527=>"111000000",
  36528=>"000001111",
  36529=>"111100000",
  36530=>"101111101",
  36531=>"000000000",
  36532=>"011011111",
  36533=>"111001000",
  36534=>"111101111",
  36535=>"001000100",
  36536=>"111011011",
  36537=>"000000000",
  36538=>"111111100",
  36539=>"000000001",
  36540=>"111111010",
  36541=>"000000111",
  36542=>"000000111",
  36543=>"000000000",
  36544=>"100000000",
  36545=>"000010111",
  36546=>"011011000",
  36547=>"000000001",
  36548=>"000000000",
  36549=>"111011000",
  36550=>"110110000",
  36551=>"000100110",
  36552=>"000100110",
  36553=>"111111000",
  36554=>"100110101",
  36555=>"000000000",
  36556=>"001000000",
  36557=>"111011000",
  36558=>"000000000",
  36559=>"001100100",
  36560=>"010111111",
  36561=>"100000000",
  36562=>"000100000",
  36563=>"111111111",
  36564=>"100100000",
  36565=>"011111110",
  36566=>"111111010",
  36567=>"001000000",
  36568=>"111001011",
  36569=>"000000100",
  36570=>"011011111",
  36571=>"001000001",
  36572=>"111111111",
  36573=>"110111111",
  36574=>"000000000",
  36575=>"000000000",
  36576=>"100000000",
  36577=>"001111111",
  36578=>"111001001",
  36579=>"000000000",
  36580=>"111111111",
  36581=>"000000000",
  36582=>"110110111",
  36583=>"000011000",
  36584=>"100000100",
  36585=>"111110111",
  36586=>"000000000",
  36587=>"111001111",
  36588=>"111111011",
  36589=>"100000000",
  36590=>"111111111",
  36591=>"111111000",
  36592=>"110111111",
  36593=>"000000110",
  36594=>"000000111",
  36595=>"111101100",
  36596=>"000000000",
  36597=>"010110000",
  36598=>"000000000",
  36599=>"000010011",
  36600=>"000000000",
  36601=>"010011010",
  36602=>"001000000",
  36603=>"100000111",
  36604=>"111111111",
  36605=>"011000000",
  36606=>"111111111",
  36607=>"011010000",
  36608=>"110110111",
  36609=>"111111111",
  36610=>"110110111",
  36611=>"111111111",
  36612=>"000100111",
  36613=>"100000001",
  36614=>"000000000",
  36615=>"000110111",
  36616=>"000000000",
  36617=>"000000111",
  36618=>"000000000",
  36619=>"011111111",
  36620=>"000000000",
  36621=>"001000001",
  36622=>"100000000",
  36623=>"010000000",
  36624=>"000000000",
  36625=>"000000111",
  36626=>"111111111",
  36627=>"000111111",
  36628=>"100000000",
  36629=>"010010000",
  36630=>"111000000",
  36631=>"000111100",
  36632=>"111111111",
  36633=>"111000000",
  36634=>"000000000",
  36635=>"011000111",
  36636=>"110100110",
  36637=>"111001000",
  36638=>"111111111",
  36639=>"000000101",
  36640=>"010100111",
  36641=>"000000111",
  36642=>"111111111",
  36643=>"000000000",
  36644=>"000010111",
  36645=>"000000000",
  36646=>"000000100",
  36647=>"111111111",
  36648=>"000110110",
  36649=>"000000000",
  36650=>"111111111",
  36651=>"001111111",
  36652=>"000011000",
  36653=>"000000000",
  36654=>"000000111",
  36655=>"001111111",
  36656=>"001001001",
  36657=>"111000000",
  36658=>"111111111",
  36659=>"110100110",
  36660=>"000000000",
  36661=>"000000000",
  36662=>"000010111",
  36663=>"000000000",
  36664=>"000000111",
  36665=>"110010000",
  36666=>"000111111",
  36667=>"111111011",
  36668=>"111111111",
  36669=>"001111111",
  36670=>"011011111",
  36671=>"011011111",
  36672=>"000000000",
  36673=>"111101110",
  36674=>"111111111",
  36675=>"111011010",
  36676=>"110110000",
  36677=>"110100111",
  36678=>"001000000",
  36679=>"101001000",
  36680=>"001101111",
  36681=>"000000000",
  36682=>"010100000",
  36683=>"000001011",
  36684=>"110000000",
  36685=>"110100100",
  36686=>"111111110",
  36687=>"110010110",
  36688=>"100110000",
  36689=>"110110100",
  36690=>"111111111",
  36691=>"111111111",
  36692=>"110111011",
  36693=>"011011011",
  36694=>"011111111",
  36695=>"000000000",
  36696=>"101111111",
  36697=>"111111111",
  36698=>"000000000",
  36699=>"111110111",
  36700=>"100100100",
  36701=>"000000000",
  36702=>"000000101",
  36703=>"110111111",
  36704=>"000000001",
  36705=>"000000000",
  36706=>"100000011",
  36707=>"000000111",
  36708=>"000001000",
  36709=>"000000000",
  36710=>"000000011",
  36711=>"000000111",
  36712=>"000110101",
  36713=>"100101111",
  36714=>"011111110",
  36715=>"000000000",
  36716=>"000000011",
  36717=>"111111000",
  36718=>"000000000",
  36719=>"000000111",
  36720=>"000000000",
  36721=>"001000000",
  36722=>"111111111",
  36723=>"110100100",
  36724=>"101111100",
  36725=>"000111111",
  36726=>"000000000",
  36727=>"111111111",
  36728=>"111101001",
  36729=>"111111001",
  36730=>"000011110",
  36731=>"100100111",
  36732=>"000100111",
  36733=>"011011110",
  36734=>"000000000",
  36735=>"111111111",
  36736=>"111111111",
  36737=>"110110100",
  36738=>"111111111",
  36739=>"111111111",
  36740=>"011010111",
  36741=>"000000000",
  36742=>"100100111",
  36743=>"000000100",
  36744=>"111111111",
  36745=>"111111111",
  36746=>"000101100",
  36747=>"000111111",
  36748=>"110100111",
  36749=>"001100110",
  36750=>"000000111",
  36751=>"000000000",
  36752=>"111111111",
  36753=>"001000000",
  36754=>"001000000",
  36755=>"111111110",
  36756=>"111111111",
  36757=>"111000000",
  36758=>"110110111",
  36759=>"111111111",
  36760=>"001111111",
  36761=>"000010110",
  36762=>"000000000",
  36763=>"011111111",
  36764=>"001111111",
  36765=>"000000000",
  36766=>"001001101",
  36767=>"011011000",
  36768=>"011001000",
  36769=>"100100110",
  36770=>"110111111",
  36771=>"000111111",
  36772=>"111110110",
  36773=>"001000000",
  36774=>"000000000",
  36775=>"111111111",
  36776=>"000000000",
  36777=>"011110100",
  36778=>"111111000",
  36779=>"101111111",
  36780=>"011111000",
  36781=>"000001000",
  36782=>"001000000",
  36783=>"111111111",
  36784=>"101000110",
  36785=>"111111000",
  36786=>"101111111",
  36787=>"000000001",
  36788=>"000000000",
  36789=>"011001001",
  36790=>"110100100",
  36791=>"000000000",
  36792=>"000000110",
  36793=>"110110110",
  36794=>"000000111",
  36795=>"111000000",
  36796=>"111100000",
  36797=>"001001001",
  36798=>"000101101",
  36799=>"101101001",
  36800=>"111111001",
  36801=>"100000000",
  36802=>"000100000",
  36803=>"000000010",
  36804=>"000000000",
  36805=>"000000111",
  36806=>"010111111",
  36807=>"110110111",
  36808=>"110110000",
  36809=>"111111011",
  36810=>"011100100",
  36811=>"000000011",
  36812=>"100100100",
  36813=>"000000000",
  36814=>"110111111",
  36815=>"111110111",
  36816=>"110110101",
  36817=>"110111111",
  36818=>"010000110",
  36819=>"111000000",
  36820=>"110111111",
  36821=>"111110100",
  36822=>"000000000",
  36823=>"111111111",
  36824=>"000000101",
  36825=>"111111111",
  36826=>"000110101",
  36827=>"000110110",
  36828=>"000111110",
  36829=>"011011000",
  36830=>"011000000",
  36831=>"111111100",
  36832=>"000000000",
  36833=>"111111111",
  36834=>"000101111",
  36835=>"000000100",
  36836=>"000000001",
  36837=>"111111111",
  36838=>"101000111",
  36839=>"111111010",
  36840=>"000001001",
  36841=>"000000000",
  36842=>"000001001",
  36843=>"101100100",
  36844=>"000000000",
  36845=>"111111111",
  36846=>"100111111",
  36847=>"100000010",
  36848=>"000101111",
  36849=>"110111011",
  36850=>"010001100",
  36851=>"111111000",
  36852=>"111111111",
  36853=>"011000000",
  36854=>"111111010",
  36855=>"111111110",
  36856=>"010111001",
  36857=>"010110110",
  36858=>"100000000",
  36859=>"111111100",
  36860=>"111111111",
  36861=>"111110000",
  36862=>"111100100",
  36863=>"111001001",
  36864=>"111111111",
  36865=>"111111000",
  36866=>"111111111",
  36867=>"000000000",
  36868=>"011111111",
  36869=>"000101111",
  36870=>"000000000",
  36871=>"111111111",
  36872=>"111111001",
  36873=>"110110111",
  36874=>"111111111",
  36875=>"011011011",
  36876=>"011001000",
  36877=>"111111111",
  36878=>"000000100",
  36879=>"000000000",
  36880=>"000000000",
  36881=>"111111111",
  36882=>"000001111",
  36883=>"111111111",
  36884=>"000000000",
  36885=>"111010000",
  36886=>"000000000",
  36887=>"000000000",
  36888=>"011011100",
  36889=>"100000000",
  36890=>"110000010",
  36891=>"100001111",
  36892=>"110000000",
  36893=>"000011111",
  36894=>"111111110",
  36895=>"001000000",
  36896=>"000000000",
  36897=>"100000000",
  36898=>"100100001",
  36899=>"111011000",
  36900=>"111111110",
  36901=>"000000000",
  36902=>"111111111",
  36903=>"000000101",
  36904=>"100100000",
  36905=>"000000101",
  36906=>"111111111",
  36907=>"000110111",
  36908=>"000000000",
  36909=>"000000000",
  36910=>"111111111",
  36911=>"100101101",
  36912=>"000000000",
  36913=>"000000011",
  36914=>"000000000",
  36915=>"111111010",
  36916=>"111111001",
  36917=>"110000000",
  36918=>"111110100",
  36919=>"111101111",
  36920=>"000001000",
  36921=>"000010111",
  36922=>"000000001",
  36923=>"000000000",
  36924=>"000000000",
  36925=>"111000100",
  36926=>"111111111",
  36927=>"000000000",
  36928=>"100000001",
  36929=>"000101101",
  36930=>"000010011",
  36931=>"000000011",
  36932=>"001000001",
  36933=>"000111111",
  36934=>"111111011",
  36935=>"111111111",
  36936=>"100110000",
  36937=>"000000001",
  36938=>"101000000",
  36939=>"100000000",
  36940=>"111111111",
  36941=>"000000110",
  36942=>"000000000",
  36943=>"000000000",
  36944=>"000000000",
  36945=>"000000011",
  36946=>"111111000",
  36947=>"000000011",
  36948=>"000111111",
  36949=>"111011111",
  36950=>"011011001",
  36951=>"111111001",
  36952=>"111111110",
  36953=>"000000000",
  36954=>"100101100",
  36955=>"001001001",
  36956=>"000000000",
  36957=>"111101000",
  36958=>"111111001",
  36959=>"111011000",
  36960=>"000000000",
  36961=>"110110000",
  36962=>"111111011",
  36963=>"000000100",
  36964=>"000011111",
  36965=>"000000000",
  36966=>"001000000",
  36967=>"110110110",
  36968=>"111111111",
  36969=>"000010110",
  36970=>"111001011",
  36971=>"000000000",
  36972=>"101111111",
  36973=>"000000000",
  36974=>"000110111",
  36975=>"000000000",
  36976=>"000011111",
  36977=>"110111111",
  36978=>"111111111",
  36979=>"111111001",
  36980=>"111001011",
  36981=>"111111001",
  36982=>"000000000",
  36983=>"000000001",
  36984=>"000000000",
  36985=>"000000000",
  36986=>"001000000",
  36987=>"000000000",
  36988=>"000000000",
  36989=>"000000010",
  36990=>"000100000",
  36991=>"111111111",
  36992=>"000000000",
  36993=>"000000111",
  36994=>"000111111",
  36995=>"111111101",
  36996=>"000000000",
  36997=>"000000000",
  36998=>"000000100",
  36999=>"000000111",
  37000=>"000000000",
  37001=>"001000000",
  37002=>"000000111",
  37003=>"100111111",
  37004=>"100000001",
  37005=>"000010000",
  37006=>"100100101",
  37007=>"111111111",
  37008=>"000000000",
  37009=>"010111111",
  37010=>"000010110",
  37011=>"100000000",
  37012=>"001011011",
  37013=>"110110100",
  37014=>"011001000",
  37015=>"000000001",
  37016=>"001010010",
  37017=>"000011111",
  37018=>"111111110",
  37019=>"110110100",
  37020=>"111111111",
  37021=>"010011001",
  37022=>"000000000",
  37023=>"111111111",
  37024=>"000000000",
  37025=>"100011011",
  37026=>"000000001",
  37027=>"000000110",
  37028=>"111111111",
  37029=>"011000100",
  37030=>"100111111",
  37031=>"110000001",
  37032=>"000000001",
  37033=>"000000000",
  37034=>"100000000",
  37035=>"000111111",
  37036=>"111011011",
  37037=>"100110100",
  37038=>"111110111",
  37039=>"000000111",
  37040=>"000000000",
  37041=>"111110110",
  37042=>"100111111",
  37043=>"111101111",
  37044=>"111000000",
  37045=>"000001000",
  37046=>"000000000",
  37047=>"000001011",
  37048=>"010111111",
  37049=>"111101100",
  37050=>"000111001",
  37051=>"001000000",
  37052=>"000000000",
  37053=>"000101000",
  37054=>"101111111",
  37055=>"011000011",
  37056=>"000000000",
  37057=>"111000100",
  37058=>"101101111",
  37059=>"100000111",
  37060=>"000101111",
  37061=>"111000111",
  37062=>"011001001",
  37063=>"111110111",
  37064=>"111111000",
  37065=>"111111011",
  37066=>"110000111",
  37067=>"001000000",
  37068=>"101001111",
  37069=>"001111111",
  37070=>"000000111",
  37071=>"000001001",
  37072=>"100110111",
  37073=>"111111110",
  37074=>"000000000",
  37075=>"001111110",
  37076=>"000000000",
  37077=>"100010000",
  37078=>"111000000",
  37079=>"110000000",
  37080=>"010011111",
  37081=>"111000001",
  37082=>"011111111",
  37083=>"000000011",
  37084=>"110110110",
  37085=>"100100100",
  37086=>"111111111",
  37087=>"000000100",
  37088=>"000000000",
  37089=>"111111111",
  37090=>"000110000",
  37091=>"110100111",
  37092=>"000000000",
  37093=>"110110000",
  37094=>"000000000",
  37095=>"111111111",
  37096=>"001111111",
  37097=>"111111010",
  37098=>"000000000",
  37099=>"100100001",
  37100=>"010010000",
  37101=>"000001001",
  37102=>"111001100",
  37103=>"111111111",
  37104=>"111111001",
  37105=>"100100001",
  37106=>"000000000",
  37107=>"000000000",
  37108=>"000100101",
  37109=>"001011011",
  37110=>"000000011",
  37111=>"111000000",
  37112=>"000100111",
  37113=>"111000110",
  37114=>"000000000",
  37115=>"000000000",
  37116=>"111100000",
  37117=>"101000001",
  37118=>"111111111",
  37119=>"111111111",
  37120=>"001000000",
  37121=>"000000100",
  37122=>"111101000",
  37123=>"000000000",
  37124=>"111011011",
  37125=>"001111111",
  37126=>"010011000",
  37127=>"000100101",
  37128=>"000000000",
  37129=>"000000000",
  37130=>"101101000",
  37131=>"111111110",
  37132=>"101101100",
  37133=>"000000000",
  37134=>"111111111",
  37135=>"000111111",
  37136=>"000000111",
  37137=>"100100100",
  37138=>"110111011",
  37139=>"000000000",
  37140=>"110110110",
  37141=>"000000010",
  37142=>"111111101",
  37143=>"110100100",
  37144=>"001000001",
  37145=>"100100111",
  37146=>"111111111",
  37147=>"000000001",
  37148=>"001000110",
  37149=>"001101111",
  37150=>"000000000",
  37151=>"000100000",
  37152=>"010010111",
  37153=>"001000100",
  37154=>"101100000",
  37155=>"001001001",
  37156=>"100110110",
  37157=>"000000000",
  37158=>"111111111",
  37159=>"111111011",
  37160=>"111111111",
  37161=>"111111111",
  37162=>"111111111",
  37163=>"000111110",
  37164=>"111111111",
  37165=>"000000101",
  37166=>"111111111",
  37167=>"010000000",
  37168=>"000000011",
  37169=>"111111111",
  37170=>"011001001",
  37171=>"000001111",
  37172=>"000000000",
  37173=>"000010111",
  37174=>"010010000",
  37175=>"111111111",
  37176=>"000000000",
  37177=>"000000000",
  37178=>"011000000",
  37179=>"000000000",
  37180=>"110000000",
  37181=>"110011111",
  37182=>"111111111",
  37183=>"111111111",
  37184=>"001111000",
  37185=>"001000100",
  37186=>"000000000",
  37187=>"000000000",
  37188=>"000000000",
  37189=>"111000001",
  37190=>"111111111",
  37191=>"000000000",
  37192=>"000000000",
  37193=>"011011011",
  37194=>"011100000",
  37195=>"111001100",
  37196=>"000110111",
  37197=>"000011111",
  37198=>"111111101",
  37199=>"111111111",
  37200=>"000100110",
  37201=>"001001001",
  37202=>"000000000",
  37203=>"000001011",
  37204=>"001000000",
  37205=>"110110000",
  37206=>"111111111",
  37207=>"000000000",
  37208=>"111111111",
  37209=>"111000101",
  37210=>"100110101",
  37211=>"000000111",
  37212=>"111111111",
  37213=>"000000010",
  37214=>"111111111",
  37215=>"000000000",
  37216=>"111111111",
  37217=>"000000000",
  37218=>"111111111",
  37219=>"111000000",
  37220=>"010111111",
  37221=>"100110111",
  37222=>"111111111",
  37223=>"001000110",
  37224=>"100000100",
  37225=>"111111111",
  37226=>"111111111",
  37227=>"100111011",
  37228=>"001001000",
  37229=>"011111001",
  37230=>"000000000",
  37231=>"111110110",
  37232=>"100000100",
  37233=>"111000000",
  37234=>"000001111",
  37235=>"100100111",
  37236=>"111111111",
  37237=>"111111111",
  37238=>"011000110",
  37239=>"111111111",
  37240=>"111111111",
  37241=>"111111111",
  37242=>"000000100",
  37243=>"101000000",
  37244=>"111111001",
  37245=>"000000000",
  37246=>"000000010",
  37247=>"000000000",
  37248=>"110110111",
  37249=>"111100000",
  37250=>"111111111",
  37251=>"101100100",
  37252=>"111000000",
  37253=>"110000000",
  37254=>"111110101",
  37255=>"111000000",
  37256=>"000000001",
  37257=>"001010111",
  37258=>"111100000",
  37259=>"111000111",
  37260=>"001000000",
  37261=>"111111111",
  37262=>"001000000",
  37263=>"000000000",
  37264=>"111000000",
  37265=>"111101101",
  37266=>"000111111",
  37267=>"111110111",
  37268=>"101001001",
  37269=>"010010011",
  37270=>"111111111",
  37271=>"000000000",
  37272=>"111111100",
  37273=>"111111110",
  37274=>"011010011",
  37275=>"110111111",
  37276=>"000000000",
  37277=>"111000111",
  37278=>"000000000",
  37279=>"000000000",
  37280=>"100001000",
  37281=>"111111111",
  37282=>"011110110",
  37283=>"111111111",
  37284=>"100110111",
  37285=>"111111101",
  37286=>"001000001",
  37287=>"111111111",
  37288=>"111101101",
  37289=>"111111111",
  37290=>"100000101",
  37291=>"000000000",
  37292=>"001011111",
  37293=>"011011011",
  37294=>"001000100",
  37295=>"111111101",
  37296=>"110111111",
  37297=>"000010111",
  37298=>"111000000",
  37299=>"000000000",
  37300=>"111101111",
  37301=>"000001111",
  37302=>"111111111",
  37303=>"111001011",
  37304=>"000001001",
  37305=>"111000000",
  37306=>"111011011",
  37307=>"111111111",
  37308=>"100000000",
  37309=>"000000110",
  37310=>"000010010",
  37311=>"111110110",
  37312=>"000000111",
  37313=>"111111111",
  37314=>"111111111",
  37315=>"111111110",
  37316=>"000000111",
  37317=>"111011111",
  37318=>"000000000",
  37319=>"111001111",
  37320=>"111000000",
  37321=>"110111111",
  37322=>"000000000",
  37323=>"000000000",
  37324=>"000011111",
  37325=>"100111111",
  37326=>"111111111",
  37327=>"000001101",
  37328=>"111011101",
  37329=>"001111011",
  37330=>"000000001",
  37331=>"010000000",
  37332=>"111000000",
  37333=>"111111100",
  37334=>"110110100",
  37335=>"100000000",
  37336=>"000000110",
  37337=>"111100111",
  37338=>"111110010",
  37339=>"000001111",
  37340=>"001100111",
  37341=>"000000001",
  37342=>"000000111",
  37343=>"111111111",
  37344=>"000000111",
  37345=>"000000000",
  37346=>"100110111",
  37347=>"000000000",
  37348=>"101111110",
  37349=>"001000000",
  37350=>"000111101",
  37351=>"110100011",
  37352=>"001010010",
  37353=>"001000000",
  37354=>"111111111",
  37355=>"100001111",
  37356=>"000111000",
  37357=>"000000001",
  37358=>"111111000",
  37359=>"011000001",
  37360=>"000101000",
  37361=>"000111111",
  37362=>"111000111",
  37363=>"101100000",
  37364=>"100000001",
  37365=>"110000000",
  37366=>"111111111",
  37367=>"000000000",
  37368=>"000000000",
  37369=>"001111011",
  37370=>"001000111",
  37371=>"000000000",
  37372=>"111111100",
  37373=>"111111111",
  37374=>"100000110",
  37375=>"000000000",
  37376=>"000000111",
  37377=>"111100000",
  37378=>"111010100",
  37379=>"011110111",
  37380=>"010110110",
  37381=>"110000000",
  37382=>"000000001",
  37383=>"111111111",
  37384=>"110000100",
  37385=>"000000010",
  37386=>"000000000",
  37387=>"000011000",
  37388=>"000000110",
  37389=>"000111111",
  37390=>"000000010",
  37391=>"000101001",
  37392=>"111111001",
  37393=>"111111111",
  37394=>"111110000",
  37395=>"111101000",
  37396=>"111100000",
  37397=>"111010000",
  37398=>"000000000",
  37399=>"011011001",
  37400=>"000011010",
  37401=>"000000000",
  37402=>"000000000",
  37403=>"111111101",
  37404=>"000111111",
  37405=>"111111101",
  37406=>"000000010",
  37407=>"111111110",
  37408=>"000000000",
  37409=>"111111111",
  37410=>"001001001",
  37411=>"110000001",
  37412=>"000110010",
  37413=>"001000000",
  37414=>"111111111",
  37415=>"110111111",
  37416=>"111111111",
  37417=>"000000110",
  37418=>"100000000",
  37419=>"010000011",
  37420=>"000000000",
  37421=>"000000010",
  37422=>"101110111",
  37423=>"111000110",
  37424=>"111111111",
  37425=>"000001001",
  37426=>"100111110",
  37427=>"011111111",
  37428=>"111111111",
  37429=>"010111110",
  37430=>"101111110",
  37431=>"011111111",
  37432=>"011111000",
  37433=>"000000000",
  37434=>"001000000",
  37435=>"100110011",
  37436=>"111101111",
  37437=>"000010110",
  37438=>"100110100",
  37439=>"000001001",
  37440=>"000000000",
  37441=>"000111111",
  37442=>"000000000",
  37443=>"110111000",
  37444=>"011011111",
  37445=>"001000100",
  37446=>"111000111",
  37447=>"000000000",
  37448=>"000000001",
  37449=>"000000000",
  37450=>"101001101",
  37451=>"010010111",
  37452=>"000000010",
  37453=>"111110110",
  37454=>"000000000",
  37455=>"111111111",
  37456=>"110000000",
  37457=>"011111111",
  37458=>"111111001",
  37459=>"011100000",
  37460=>"000000000",
  37461=>"010010110",
  37462=>"001000011",
  37463=>"011000000",
  37464=>"000000000",
  37465=>"111000111",
  37466=>"111111111",
  37467=>"011011000",
  37468=>"000110110",
  37469=>"111111111",
  37470=>"000001111",
  37471=>"100111111",
  37472=>"100000000",
  37473=>"111111111",
  37474=>"111100101",
  37475=>"101000000",
  37476=>"010000111",
  37477=>"111001101",
  37478=>"011111111",
  37479=>"100100000",
  37480=>"010011111",
  37481=>"000011111",
  37482=>"110000111",
  37483=>"111111111",
  37484=>"010110111",
  37485=>"100101111",
  37486=>"000000000",
  37487=>"111011000",
  37488=>"000000111",
  37489=>"000001111",
  37490=>"101101111",
  37491=>"010110000",
  37492=>"001001111",
  37493=>"001000000",
  37494=>"111111111",
  37495=>"000000000",
  37496=>"000000000",
  37497=>"010000000",
  37498=>"000000110",
  37499=>"000000000",
  37500=>"000110110",
  37501=>"111101111",
  37502=>"000000000",
  37503=>"000010000",
  37504=>"000000000",
  37505=>"111111111",
  37506=>"111111011",
  37507=>"000001001",
  37508=>"000111111",
  37509=>"101000000",
  37510=>"000001000",
  37511=>"011000000",
  37512=>"001001001",
  37513=>"100100101",
  37514=>"000000000",
  37515=>"111111111",
  37516=>"111111101",
  37517=>"000000000",
  37518=>"000010110",
  37519=>"000000000",
  37520=>"101101111",
  37521=>"000000000",
  37522=>"000001111",
  37523=>"100110110",
  37524=>"111110010",
  37525=>"000000000",
  37526=>"100111000",
  37527=>"000000101",
  37528=>"111111111",
  37529=>"000000001",
  37530=>"111011011",
  37531=>"111111111",
  37532=>"100000000",
  37533=>"111111111",
  37534=>"011100111",
  37535=>"111111111",
  37536=>"000000000",
  37537=>"111000111",
  37538=>"000000100",
  37539=>"000001111",
  37540=>"001001110",
  37541=>"111011001",
  37542=>"110111010",
  37543=>"000001101",
  37544=>"000000001",
  37545=>"000000000",
  37546=>"000111111",
  37547=>"111111111",
  37548=>"000001001",
  37549=>"000110100",
  37550=>"111000100",
  37551=>"110110000",
  37552=>"110111000",
  37553=>"000011000",
  37554=>"000111010",
  37555=>"010111011",
  37556=>"111111111",
  37557=>"100001011",
  37558=>"001100100",
  37559=>"000100100",
  37560=>"011000000",
  37561=>"000000000",
  37562=>"000101111",
  37563=>"101001001",
  37564=>"111000000",
  37565=>"111111111",
  37566=>"000000000",
  37567=>"101000000",
  37568=>"000000000",
  37569=>"011001011",
  37570=>"000000111",
  37571=>"100111001",
  37572=>"010010110",
  37573=>"000111111",
  37574=>"010001111",
  37575=>"000110100",
  37576=>"111111100",
  37577=>"000000000",
  37578=>"110000100",
  37579=>"001000000",
  37580=>"111111111",
  37581=>"111111111",
  37582=>"000000000",
  37583=>"000000000",
  37584=>"110001011",
  37585=>"000111111",
  37586=>"000111111",
  37587=>"000000100",
  37588=>"000000011",
  37589=>"110001011",
  37590=>"110110111",
  37591=>"111110110",
  37592=>"000010000",
  37593=>"111110111",
  37594=>"000000000",
  37595=>"000011111",
  37596=>"111111001",
  37597=>"111111101",
  37598=>"111111111",
  37599=>"000000101",
  37600=>"000000111",
  37601=>"111111111",
  37602=>"100000001",
  37603=>"000000011",
  37604=>"000000000",
  37605=>"110110110",
  37606=>"000000000",
  37607=>"111000000",
  37608=>"000101001",
  37609=>"000000000",
  37610=>"111111111",
  37611=>"010000000",
  37612=>"111000000",
  37613=>"100110111",
  37614=>"111111111",
  37615=>"001000000",
  37616=>"001000111",
  37617=>"111111111",
  37618=>"111011011",
  37619=>"001111111",
  37620=>"000000000",
  37621=>"000111111",
  37622=>"001011001",
  37623=>"111101001",
  37624=>"000000000",
  37625=>"000000000",
  37626=>"000000011",
  37627=>"000010000",
  37628=>"011111110",
  37629=>"010111111",
  37630=>"111001001",
  37631=>"011111111",
  37632=>"000110010",
  37633=>"000100101",
  37634=>"000000010",
  37635=>"000000000",
  37636=>"001011000",
  37637=>"000000000",
  37638=>"000011111",
  37639=>"110111000",
  37640=>"011111111",
  37641=>"111100100",
  37642=>"111111111",
  37643=>"100000000",
  37644=>"000000000",
  37645=>"111111111",
  37646=>"111111111",
  37647=>"111111111",
  37648=>"011111111",
  37649=>"000000110",
  37650=>"000000001",
  37651=>"100000101",
  37652=>"000000000",
  37653=>"111000000",
  37654=>"100110110",
  37655=>"111111111",
  37656=>"100000000",
  37657=>"000000011",
  37658=>"110100000",
  37659=>"110100001",
  37660=>"011111111",
  37661=>"000000111",
  37662=>"111111111",
  37663=>"000000000",
  37664=>"011011011",
  37665=>"000100000",
  37666=>"001010000",
  37667=>"111111111",
  37668=>"111111111",
  37669=>"111111111",
  37670=>"000000000",
  37671=>"111101111",
  37672=>"111111111",
  37673=>"100000000",
  37674=>"001100111",
  37675=>"000100011",
  37676=>"101111101",
  37677=>"110000010",
  37678=>"101111111",
  37679=>"000100100",
  37680=>"110110100",
  37681=>"100100111",
  37682=>"011011011",
  37683=>"111111111",
  37684=>"010000000",
  37685=>"000000101",
  37686=>"000000010",
  37687=>"000100111",
  37688=>"000110000",
  37689=>"000000000",
  37690=>"111001001",
  37691=>"111111111",
  37692=>"111111000",
  37693=>"111110000",
  37694=>"000000000",
  37695=>"111110110",
  37696=>"111000000",
  37697=>"111110110",
  37698=>"111111111",
  37699=>"100000000",
  37700=>"000000000",
  37701=>"111111101",
  37702=>"000000000",
  37703=>"111111101",
  37704=>"111111111",
  37705=>"010000000",
  37706=>"111100100",
  37707=>"000011011",
  37708=>"111111111",
  37709=>"000000000",
  37710=>"111111111",
  37711=>"100000000",
  37712=>"001111001",
  37713=>"000001111",
  37714=>"000000110",
  37715=>"000000000",
  37716=>"000000000",
  37717=>"011011011",
  37718=>"111110000",
  37719=>"101111000",
  37720=>"000000011",
  37721=>"111111110",
  37722=>"111110110",
  37723=>"000000001",
  37724=>"111111111",
  37725=>"000000000",
  37726=>"000000001",
  37727=>"001001110",
  37728=>"100110110",
  37729=>"110110111",
  37730=>"000001111",
  37731=>"111111111",
  37732=>"000000110",
  37733=>"001000100",
  37734=>"000111111",
  37735=>"110111111",
  37736=>"000100100",
  37737=>"010011000",
  37738=>"000001111",
  37739=>"000000000",
  37740=>"111111111",
  37741=>"001000110",
  37742=>"000000000",
  37743=>"000000001",
  37744=>"011011111",
  37745=>"000001000",
  37746=>"111101100",
  37747=>"000001001",
  37748=>"000000001",
  37749=>"111111111",
  37750=>"111111110",
  37751=>"111111110",
  37752=>"111000000",
  37753=>"000111111",
  37754=>"000000000",
  37755=>"000000000",
  37756=>"000001111",
  37757=>"011000000",
  37758=>"111110110",
  37759=>"011000000",
  37760=>"000100100",
  37761=>"001101111",
  37762=>"000000001",
  37763=>"000101001",
  37764=>"011111111",
  37765=>"000100100",
  37766=>"111101000",
  37767=>"100000111",
  37768=>"000000111",
  37769=>"111111000",
  37770=>"110111111",
  37771=>"111110110",
  37772=>"111000111",
  37773=>"000110110",
  37774=>"111011001",
  37775=>"000100000",
  37776=>"000111111",
  37777=>"111111111",
  37778=>"111111000",
  37779=>"111011010",
  37780=>"011010010",
  37781=>"000000000",
  37782=>"011000110",
  37783=>"000110110",
  37784=>"010000000",
  37785=>"110110001",
  37786=>"000010010",
  37787=>"001100110",
  37788=>"000000010",
  37789=>"111010110",
  37790=>"001001000",
  37791=>"100111010",
  37792=>"101111111",
  37793=>"100100101",
  37794=>"000000000",
  37795=>"111111000",
  37796=>"010111111",
  37797=>"110111010",
  37798=>"000110000",
  37799=>"111111011",
  37800=>"100100000",
  37801=>"110000011",
  37802=>"101001101",
  37803=>"011011011",
  37804=>"111111000",
  37805=>"000000000",
  37806=>"111111111",
  37807=>"000011000",
  37808=>"111111111",
  37809=>"010111000",
  37810=>"001000000",
  37811=>"000011000",
  37812=>"000000111",
  37813=>"111111100",
  37814=>"100100000",
  37815=>"001000001",
  37816=>"111111100",
  37817=>"111111111",
  37818=>"001000001",
  37819=>"001100110",
  37820=>"111110000",
  37821=>"111111001",
  37822=>"100000000",
  37823=>"000100001",
  37824=>"000001111",
  37825=>"000000000",
  37826=>"111111111",
  37827=>"111111011",
  37828=>"100010011",
  37829=>"111111111",
  37830=>"111011000",
  37831=>"010000011",
  37832=>"110110000",
  37833=>"000000000",
  37834=>"000000101",
  37835=>"011111111",
  37836=>"011000000",
  37837=>"111001000",
  37838=>"110010110",
  37839=>"000110111",
  37840=>"000000000",
  37841=>"110111111",
  37842=>"111111111",
  37843=>"001001111",
  37844=>"111111111",
  37845=>"111000011",
  37846=>"110111111",
  37847=>"000011111",
  37848=>"000110111",
  37849=>"001111111",
  37850=>"110110100",
  37851=>"110100111",
  37852=>"000001101",
  37853=>"101101101",
  37854=>"111111011",
  37855=>"000001001",
  37856=>"000110110",
  37857=>"111111111",
  37858=>"111111000",
  37859=>"001000101",
  37860=>"111111111",
  37861=>"000000111",
  37862=>"111000000",
  37863=>"001000000",
  37864=>"000000000",
  37865=>"001001100",
  37866=>"000000100",
  37867=>"000001001",
  37868=>"111111001",
  37869=>"000000001",
  37870=>"111111000",
  37871=>"000000111",
  37872=>"001001000",
  37873=>"000000000",
  37874=>"011001001",
  37875=>"111111000",
  37876=>"000000000",
  37877=>"110000111",
  37878=>"110111110",
  37879=>"110111101",
  37880=>"000000000",
  37881=>"000111100",
  37882=>"000001000",
  37883=>"111111001",
  37884=>"000000000",
  37885=>"111011011",
  37886=>"110100000",
  37887=>"000000111",
  37888=>"100000000",
  37889=>"111111111",
  37890=>"111000111",
  37891=>"011000000",
  37892=>"001000001",
  37893=>"111011111",
  37894=>"111111110",
  37895=>"111111111",
  37896=>"111111011",
  37897=>"111011001",
  37898=>"111111000",
  37899=>"000000100",
  37900=>"000010100",
  37901=>"000000011",
  37902=>"011111111",
  37903=>"001000000",
  37904=>"111111000",
  37905=>"000000001",
  37906=>"000000000",
  37907=>"111101111",
  37908=>"111111111",
  37909=>"111111000",
  37910=>"010111110",
  37911=>"000000000",
  37912=>"000000000",
  37913=>"011100100",
  37914=>"000110000",
  37915=>"000000000",
  37916=>"000000000",
  37917=>"000010010",
  37918=>"000000111",
  37919=>"000000111",
  37920=>"000000000",
  37921=>"110111111",
  37922=>"100001111",
  37923=>"111111001",
  37924=>"101000111",
  37925=>"000000000",
  37926=>"000000000",
  37927=>"111111000",
  37928=>"000010110",
  37929=>"111101000",
  37930=>"111111101",
  37931=>"001010111",
  37932=>"010011011",
  37933=>"111110110",
  37934=>"000000110",
  37935=>"001111111",
  37936=>"000000000",
  37937=>"000000000",
  37938=>"111111111",
  37939=>"111011011",
  37940=>"000000000",
  37941=>"000000000",
  37942=>"111111101",
  37943=>"011011000",
  37944=>"100100000",
  37945=>"000001111",
  37946=>"000001111",
  37947=>"000001011",
  37948=>"111000000",
  37949=>"000000000",
  37950=>"111111111",
  37951=>"001000000",
  37952=>"011011111",
  37953=>"000000110",
  37954=>"111011000",
  37955=>"011111111",
  37956=>"011001011",
  37957=>"011011001",
  37958=>"111100000",
  37959=>"000000000",
  37960=>"111011001",
  37961=>"111010010",
  37962=>"011001001",
  37963=>"000000000",
  37964=>"000111111",
  37965=>"000000000",
  37966=>"001000011",
  37967=>"000000111",
  37968=>"000111111",
  37969=>"111111110",
  37970=>"000000000",
  37971=>"001001000",
  37972=>"000000000",
  37973=>"000000000",
  37974=>"100000001",
  37975=>"000000101",
  37976=>"111101111",
  37977=>"100000000",
  37978=>"111111011",
  37979=>"111101001",
  37980=>"100000001",
  37981=>"000000000",
  37982=>"000000000",
  37983=>"000000000",
  37984=>"110110111",
  37985=>"111111011",
  37986=>"101000001",
  37987=>"000000011",
  37988=>"000111000",
  37989=>"000000000",
  37990=>"111111000",
  37991=>"111111111",
  37992=>"000000100",
  37993=>"111001000",
  37994=>"111111111",
  37995=>"000110111",
  37996=>"111111111",
  37997=>"000000000",
  37998=>"001001111",
  37999=>"000000111",
  38000=>"000000000",
  38001=>"111111011",
  38002=>"000011111",
  38003=>"000001000",
  38004=>"110100100",
  38005=>"000001000",
  38006=>"111101000",
  38007=>"000000111",
  38008=>"000100111",
  38009=>"000000001",
  38010=>"111100000",
  38011=>"000000001",
  38012=>"000000010",
  38013=>"000000000",
  38014=>"000000000",
  38015=>"000010111",
  38016=>"000100110",
  38017=>"001000011",
  38018=>"110111000",
  38019=>"110100111",
  38020=>"000101111",
  38021=>"111000000",
  38022=>"100100000",
  38023=>"101011111",
  38024=>"110100010",
  38025=>"011111100",
  38026=>"111111111",
  38027=>"111111010",
  38028=>"110010110",
  38029=>"000000011",
  38030=>"110011110",
  38031=>"011011011",
  38032=>"000000101",
  38033=>"000000000",
  38034=>"111111001",
  38035=>"000000000",
  38036=>"111111000",
  38037=>"001001011",
  38038=>"000111111",
  38039=>"001000000",
  38040=>"100000001",
  38041=>"110111111",
  38042=>"000100111",
  38043=>"001001011",
  38044=>"111110000",
  38045=>"111111111",
  38046=>"111111000",
  38047=>"111111001",
  38048=>"000000000",
  38049=>"111011000",
  38050=>"011011111",
  38051=>"000100111",
  38052=>"001001000",
  38053=>"100000101",
  38054=>"001101101",
  38055=>"000001000",
  38056=>"000011000",
  38057=>"000000000",
  38058=>"111111111",
  38059=>"000000110",
  38060=>"011011111",
  38061=>"000001011",
  38062=>"000000011",
  38063=>"111111000",
  38064=>"111111111",
  38065=>"011011010",
  38066=>"000100000",
  38067=>"101000000",
  38068=>"000000000",
  38069=>"000000000",
  38070=>"000000000",
  38071=>"000000101",
  38072=>"000000000",
  38073=>"111111111",
  38074=>"111100100",
  38075=>"110110110",
  38076=>"000000011",
  38077=>"111111111",
  38078=>"000111001",
  38079=>"111011001",
  38080=>"000111110",
  38081=>"000111001",
  38082=>"000011011",
  38083=>"000000000",
  38084=>"000001111",
  38085=>"000000000",
  38086=>"001111111",
  38087=>"111111101",
  38088=>"011111010",
  38089=>"101101101",
  38090=>"001101101",
  38091=>"000000001",
  38092=>"000000011",
  38093=>"000011000",
  38094=>"000111111",
  38095=>"111111011",
  38096=>"000000001",
  38097=>"000001001",
  38098=>"011000000",
  38099=>"111111111",
  38100=>"001001111",
  38101=>"001011111",
  38102=>"000000000",
  38103=>"111111110",
  38104=>"111111000",
  38105=>"110111110",
  38106=>"001111111",
  38107=>"000000000",
  38108=>"111111111",
  38109=>"000000000",
  38110=>"111101000",
  38111=>"000000000",
  38112=>"000000000",
  38113=>"111111111",
  38114=>"111111110",
  38115=>"100000011",
  38116=>"001000001",
  38117=>"111111111",
  38118=>"000000100",
  38119=>"101101111",
  38120=>"111111111",
  38121=>"011010000",
  38122=>"000000001",
  38123=>"001001111",
  38124=>"111111000",
  38125=>"000000111",
  38126=>"111111111",
  38127=>"111001101",
  38128=>"000111111",
  38129=>"110000000",
  38130=>"001111111",
  38131=>"111110001",
  38132=>"111001001",
  38133=>"000000000",
  38134=>"111111111",
  38135=>"111111111",
  38136=>"000000110",
  38137=>"111111111",
  38138=>"100000000",
  38139=>"100000101",
  38140=>"000001111",
  38141=>"111011000",
  38142=>"111101111",
  38143=>"010110000",
  38144=>"111110000",
  38145=>"100100100",
  38146=>"111111011",
  38147=>"010111111",
  38148=>"111111111",
  38149=>"001010110",
  38150=>"110101111",
  38151=>"000000001",
  38152=>"111001001",
  38153=>"110110110",
  38154=>"011111111",
  38155=>"000110111",
  38156=>"110100100",
  38157=>"100100101",
  38158=>"100000000",
  38159=>"000111111",
  38160=>"000111000",
  38161=>"111000000",
  38162=>"000100110",
  38163=>"111111111",
  38164=>"001001111",
  38165=>"111111000",
  38166=>"001000000",
  38167=>"110111111",
  38168=>"001010010",
  38169=>"010000111",
  38170=>"001000111",
  38171=>"000000000",
  38172=>"100110111",
  38173=>"110000000",
  38174=>"111111111",
  38175=>"100000000",
  38176=>"011000000",
  38177=>"111111111",
  38178=>"000101111",
  38179=>"110011111",
  38180=>"011000110",
  38181=>"111111111",
  38182=>"110000000",
  38183=>"111111111",
  38184=>"011110111",
  38185=>"000000000",
  38186=>"110010111",
  38187=>"011001001",
  38188=>"000110100",
  38189=>"100110110",
  38190=>"000000111",
  38191=>"000000000",
  38192=>"111011001",
  38193=>"111111000",
  38194=>"000000000",
  38195=>"111111000",
  38196=>"000001000",
  38197=>"000000000",
  38198=>"111111101",
  38199=>"000111111",
  38200=>"011011000",
  38201=>"111111111",
  38202=>"111000000",
  38203=>"100100001",
  38204=>"000100111",
  38205=>"001001111",
  38206=>"101000000",
  38207=>"111010000",
  38208=>"111101111",
  38209=>"111111111",
  38210=>"111100111",
  38211=>"000110110",
  38212=>"000001101",
  38213=>"000000000",
  38214=>"010110100",
  38215=>"111111000",
  38216=>"111111011",
  38217=>"001000000",
  38218=>"110000111",
  38219=>"100100100",
  38220=>"001000100",
  38221=>"001001001",
  38222=>"111011011",
  38223=>"000000111",
  38224=>"111111001",
  38225=>"010000000",
  38226=>"000001000",
  38227=>"000000111",
  38228=>"100111111",
  38229=>"111011001",
  38230=>"111000000",
  38231=>"100000000",
  38232=>"011001111",
  38233=>"000000000",
  38234=>"101000000",
  38235=>"011000001",
  38236=>"111111111",
  38237=>"111001001",
  38238=>"111100000",
  38239=>"111011000",
  38240=>"111111101",
  38241=>"000000000",
  38242=>"100110111",
  38243=>"101001000",
  38244=>"000000111",
  38245=>"000000000",
  38246=>"011010000",
  38247=>"111111110",
  38248=>"001011001",
  38249=>"011110100",
  38250=>"000010000",
  38251=>"000111110",
  38252=>"000001111",
  38253=>"110111001",
  38254=>"000000000",
  38255=>"000000111",
  38256=>"111111111",
  38257=>"111110000",
  38258=>"111000000",
  38259=>"100000000",
  38260=>"000000000",
  38261=>"000000000",
  38262=>"111000111",
  38263=>"000001000",
  38264=>"111100000",
  38265=>"000111111",
  38266=>"111111111",
  38267=>"001110000",
  38268=>"010011111",
  38269=>"000111111",
  38270=>"000000000",
  38271=>"000000000",
  38272=>"010011000",
  38273=>"011111111",
  38274=>"110111111",
  38275=>"110111001",
  38276=>"000000000",
  38277=>"000000000",
  38278=>"001111111",
  38279=>"110110111",
  38280=>"000111111",
  38281=>"011111111",
  38282=>"011001011",
  38283=>"000111111",
  38284=>"000000101",
  38285=>"110110110",
  38286=>"010110110",
  38287=>"000000101",
  38288=>"000111111",
  38289=>"000000111",
  38290=>"011011111",
  38291=>"000000011",
  38292=>"000000000",
  38293=>"000000000",
  38294=>"111111111",
  38295=>"101100000",
  38296=>"101111111",
  38297=>"000001111",
  38298=>"010111110",
  38299=>"110111111",
  38300=>"111111111",
  38301=>"000000111",
  38302=>"111000000",
  38303=>"000011001",
  38304=>"000000100",
  38305=>"111111001",
  38306=>"110010011",
  38307=>"000100101",
  38308=>"000100111",
  38309=>"111111111",
  38310=>"000000000",
  38311=>"001111111",
  38312=>"000000011",
  38313=>"000000000",
  38314=>"111111111",
  38315=>"110100011",
  38316=>"111111111",
  38317=>"000000001",
  38318=>"111000000",
  38319=>"100100100",
  38320=>"000000111",
  38321=>"000000011",
  38322=>"000111111",
  38323=>"000000001",
  38324=>"001000000",
  38325=>"111111111",
  38326=>"110111110",
  38327=>"000111111",
  38328=>"111111110",
  38329=>"100111101",
  38330=>"000000001",
  38331=>"000000000",
  38332=>"111111111",
  38333=>"000010110",
  38334=>"111111011",
  38335=>"111001000",
  38336=>"000000001",
  38337=>"001000011",
  38338=>"111100000",
  38339=>"000000000",
  38340=>"100000001",
  38341=>"111110000",
  38342=>"111000000",
  38343=>"111111111",
  38344=>"110111111",
  38345=>"000000000",
  38346=>"111000000",
  38347=>"000000000",
  38348=>"001100000",
  38349=>"000001000",
  38350=>"011111101",
  38351=>"000011111",
  38352=>"100000011",
  38353=>"111110000",
  38354=>"111111111",
  38355=>"111000000",
  38356=>"100101111",
  38357=>"000000011",
  38358=>"000000000",
  38359=>"010110110",
  38360=>"001001011",
  38361=>"000000000",
  38362=>"000000001",
  38363=>"111111000",
  38364=>"111111111",
  38365=>"111011111",
  38366=>"111000000",
  38367=>"100111111",
  38368=>"111001000",
  38369=>"001000000",
  38370=>"000001000",
  38371=>"000001011",
  38372=>"111100000",
  38373=>"000000000",
  38374=>"000011011",
  38375=>"000000000",
  38376=>"110111110",
  38377=>"000100000",
  38378=>"111110000",
  38379=>"111100111",
  38380=>"001010111",
  38381=>"110011000",
  38382=>"101100111",
  38383=>"111111011",
  38384=>"000000000",
  38385=>"111000000",
  38386=>"101110110",
  38387=>"000000011",
  38388=>"000010000",
  38389=>"001000000",
  38390=>"000101111",
  38391=>"011011000",
  38392=>"011000000",
  38393=>"000000000",
  38394=>"111111111",
  38395=>"111111111",
  38396=>"000100111",
  38397=>"000001001",
  38398=>"011011001",
  38399=>"000000111",
  38400=>"111111110",
  38401=>"000000111",
  38402=>"000111111",
  38403=>"111111000",
  38404=>"000000000",
  38405=>"001000000",
  38406=>"111111111",
  38407=>"111111111",
  38408=>"000101111",
  38409=>"001001011",
  38410=>"100000111",
  38411=>"111011011",
  38412=>"101111111",
  38413=>"000001011",
  38414=>"100110110",
  38415=>"001001100",
  38416=>"000000100",
  38417=>"000101011",
  38418=>"001111011",
  38419=>"000111000",
  38420=>"111111001",
  38421=>"110111111",
  38422=>"010111111",
  38423=>"100110111",
  38424=>"100100000",
  38425=>"001000000",
  38426=>"000001011",
  38427=>"000000010",
  38428=>"000000011",
  38429=>"000001111",
  38430=>"000000000",
  38431=>"000000011",
  38432=>"111111111",
  38433=>"000000000",
  38434=>"111111101",
  38435=>"000000000",
  38436=>"000000000",
  38437=>"111000100",
  38438=>"111111000",
  38439=>"000000011",
  38440=>"001111111",
  38441=>"000000000",
  38442=>"111111111",
  38443=>"000000100",
  38444=>"011000100",
  38445=>"111111111",
  38446=>"111000000",
  38447=>"001111111",
  38448=>"100000000",
  38449=>"000000000",
  38450=>"000100100",
  38451=>"000001001",
  38452=>"000001001",
  38453=>"110111100",
  38454=>"000000000",
  38455=>"111111111",
  38456=>"111111010",
  38457=>"000000000",
  38458=>"111101101",
  38459=>"010110010",
  38460=>"000100000",
  38461=>"000000000",
  38462=>"011000100",
  38463=>"000000000",
  38464=>"011110000",
  38465=>"000000011",
  38466=>"000111111",
  38467=>"111111000",
  38468=>"000110110",
  38469=>"001000010",
  38470=>"111111011",
  38471=>"111111111",
  38472=>"111111110",
  38473=>"111111000",
  38474=>"000100101",
  38475=>"111001000",
  38476=>"000000000",
  38477=>"101000000",
  38478=>"100100111",
  38479=>"000000000",
  38480=>"111111011",
  38481=>"111111111",
  38482=>"000011111",
  38483=>"111111100",
  38484=>"111000000",
  38485=>"000001111",
  38486=>"111011000",
  38487=>"111111011",
  38488=>"110111111",
  38489=>"111001101",
  38490=>"111111111",
  38491=>"000000111",
  38492=>"111110000",
  38493=>"000000000",
  38494=>"000000000",
  38495=>"100000111",
  38496=>"110000000",
  38497=>"100111110",
  38498=>"000111111",
  38499=>"000000110",
  38500=>"110010000",
  38501=>"111111111",
  38502=>"000000010",
  38503=>"111111111",
  38504=>"111001000",
  38505=>"000111111",
  38506=>"000101111",
  38507=>"111111111",
  38508=>"100101101",
  38509=>"000001011",
  38510=>"101001111",
  38511=>"000000000",
  38512=>"111100000",
  38513=>"111010000",
  38514=>"010001011",
  38515=>"000000101",
  38516=>"000000000",
  38517=>"000000000",
  38518=>"000111111",
  38519=>"000000000",
  38520=>"111111111",
  38521=>"011000000",
  38522=>"000000000",
  38523=>"000000111",
  38524=>"110110110",
  38525=>"000111111",
  38526=>"000000000",
  38527=>"000110111",
  38528=>"000000111",
  38529=>"111111000",
  38530=>"111000000",
  38531=>"111011000",
  38532=>"111111111",
  38533=>"001001001",
  38534=>"100101000",
  38535=>"110010110",
  38536=>"000000111",
  38537=>"111111011",
  38538=>"000000000",
  38539=>"111111001",
  38540=>"000001001",
  38541=>"111000000",
  38542=>"000011111",
  38543=>"111111111",
  38544=>"000000000",
  38545=>"111000000",
  38546=>"000000000",
  38547=>"110000000",
  38548=>"111001011",
  38549=>"111111111",
  38550=>"111110000",
  38551=>"111000111",
  38552=>"101000111",
  38553=>"100000111",
  38554=>"000111111",
  38555=>"000000000",
  38556=>"111111000",
  38557=>"000000111",
  38558=>"111101000",
  38559=>"000011011",
  38560=>"111111111",
  38561=>"000000000",
  38562=>"111000001",
  38563=>"100000000",
  38564=>"000000000",
  38565=>"111111011",
  38566=>"001101111",
  38567=>"001111001",
  38568=>"111111111",
  38569=>"000000000",
  38570=>"111111111",
  38571=>"000000100",
  38572=>"000000000",
  38573=>"000010111",
  38574=>"111110111",
  38575=>"101100001",
  38576=>"111111000",
  38577=>"100000000",
  38578=>"111111111",
  38579=>"000101111",
  38580=>"000111110",
  38581=>"111111000",
  38582=>"001000000",
  38583=>"011011000",
  38584=>"111111111",
  38585=>"000111111",
  38586=>"001101001",
  38587=>"000000100",
  38588=>"000000001",
  38589=>"111111000",
  38590=>"111111111",
  38591=>"101111111",
  38592=>"011011111",
  38593=>"000011111",
  38594=>"000000001",
  38595=>"001000000",
  38596=>"000000111",
  38597=>"000110111",
  38598=>"000111111",
  38599=>"110111000",
  38600=>"011111110",
  38601=>"111111111",
  38602=>"100111111",
  38603=>"000000000",
  38604=>"011111111",
  38605=>"000111110",
  38606=>"111111000",
  38607=>"111001000",
  38608=>"110111001",
  38609=>"000000010",
  38610=>"000000000",
  38611=>"011001000",
  38612=>"010000000",
  38613=>"000000000",
  38614=>"111111000",
  38615=>"000000111",
  38616=>"000001111",
  38617=>"000000110",
  38618=>"000000000",
  38619=>"111000110",
  38620=>"111111111",
  38621=>"111011111",
  38622=>"011111111",
  38623=>"000111000",
  38624=>"111100111",
  38625=>"111111000",
  38626=>"110100100",
  38627=>"001011111",
  38628=>"001111000",
  38629=>"000000111",
  38630=>"111110111",
  38631=>"110000000",
  38632=>"010000000",
  38633=>"110100000",
  38634=>"001100001",
  38635=>"000000000",
  38636=>"000000000",
  38637=>"011000111",
  38638=>"000111111",
  38639=>"000000100",
  38640=>"111111111",
  38641=>"111111111",
  38642=>"001000000",
  38643=>"000000111",
  38644=>"111111000",
  38645=>"111000001",
  38646=>"000110010",
  38647=>"111001000",
  38648=>"111111011",
  38649=>"110111111",
  38650=>"111110000",
  38651=>"010111111",
  38652=>"000100000",
  38653=>"111111000",
  38654=>"001101111",
  38655=>"100101111",
  38656=>"001010000",
  38657=>"000000111",
  38658=>"000000000",
  38659=>"111111100",
  38660=>"001000000",
  38661=>"000001111",
  38662=>"000000000",
  38663=>"100110110",
  38664=>"001011111",
  38665=>"001000001",
  38666=>"111111111",
  38667=>"110110100",
  38668=>"011011111",
  38669=>"111111000",
  38670=>"110110000",
  38671=>"111111111",
  38672=>"101001011",
  38673=>"000000000",
  38674=>"000001001",
  38675=>"000000011",
  38676=>"000011000",
  38677=>"010010111",
  38678=>"110110110",
  38679=>"111111000",
  38680=>"101011011",
  38681=>"000000000",
  38682=>"111000000",
  38683=>"111111111",
  38684=>"011111001",
  38685=>"111111111",
  38686=>"000000110",
  38687=>"010000111",
  38688=>"100000000",
  38689=>"101000000",
  38690=>"000000000",
  38691=>"111111111",
  38692=>"010000111",
  38693=>"011111111",
  38694=>"111111001",
  38695=>"001001000",
  38696=>"010111111",
  38697=>"011001001",
  38698=>"000110111",
  38699=>"111111001",
  38700=>"000000000",
  38701=>"000000111",
  38702=>"101101011",
  38703=>"011011111",
  38704=>"111101100",
  38705=>"111101001",
  38706=>"100100111",
  38707=>"000011111",
  38708=>"111101111",
  38709=>"011110000",
  38710=>"111000001",
  38711=>"111011111",
  38712=>"110110000",
  38713=>"111000000",
  38714=>"111111111",
  38715=>"000001101",
  38716=>"000000000",
  38717=>"000101001",
  38718=>"111001000",
  38719=>"000000111",
  38720=>"000000111",
  38721=>"001001001",
  38722=>"111111000",
  38723=>"111001111",
  38724=>"000000000",
  38725=>"111111000",
  38726=>"000000000",
  38727=>"000000011",
  38728=>"000000000",
  38729=>"000000111",
  38730=>"000100111",
  38731=>"000000111",
  38732=>"011011000",
  38733=>"110000000",
  38734=>"111111111",
  38735=>"000100111",
  38736=>"011111011",
  38737=>"111111000",
  38738=>"111111101",
  38739=>"111100111",
  38740=>"000000000",
  38741=>"011011001",
  38742=>"001111111",
  38743=>"000000000",
  38744=>"111101111",
  38745=>"111111111",
  38746=>"010000111",
  38747=>"000000000",
  38748=>"000111111",
  38749=>"011011111",
  38750=>"001111111",
  38751=>"111111111",
  38752=>"100111100",
  38753=>"000000000",
  38754=>"001010010",
  38755=>"111100111",
  38756=>"100110111",
  38757=>"010111111",
  38758=>"111001001",
  38759=>"000011111",
  38760=>"000000110",
  38761=>"000011111",
  38762=>"111100111",
  38763=>"000111010",
  38764=>"000001111",
  38765=>"000000000",
  38766=>"111111111",
  38767=>"000000000",
  38768=>"001011011",
  38769=>"000001001",
  38770=>"000000101",
  38771=>"001111111",
  38772=>"000000000",
  38773=>"000000000",
  38774=>"000000111",
  38775=>"111010000",
  38776=>"000000000",
  38777=>"000000000",
  38778=>"001001111",
  38779=>"111111111",
  38780=>"100000011",
  38781=>"101001000",
  38782=>"111111001",
  38783=>"000011111",
  38784=>"000000000",
  38785=>"000000000",
  38786=>"110011000",
  38787=>"001001000",
  38788=>"111111001",
  38789=>"010111111",
  38790=>"100100001",
  38791=>"111111111",
  38792=>"000000111",
  38793=>"111000000",
  38794=>"001111111",
  38795=>"111111111",
  38796=>"111101111",
  38797=>"000001001",
  38798=>"111000111",
  38799=>"011001000",
  38800=>"000000000",
  38801=>"000000111",
  38802=>"101000000",
  38803=>"000000000",
  38804=>"111111000",
  38805=>"000110100",
  38806=>"111111111",
  38807=>"000100000",
  38808=>"111111000",
  38809=>"001000000",
  38810=>"000000000",
  38811=>"111111111",
  38812=>"000000000",
  38813=>"111000000",
  38814=>"000001001",
  38815=>"110000000",
  38816=>"011111111",
  38817=>"000110110",
  38818=>"111111100",
  38819=>"001100000",
  38820=>"111111111",
  38821=>"111111100",
  38822=>"000001001",
  38823=>"000000000",
  38824=>"010111000",
  38825=>"001000101",
  38826=>"111111111",
  38827=>"111111100",
  38828=>"000000000",
  38829=>"000001111",
  38830=>"000110111",
  38831=>"100000000",
  38832=>"110111111",
  38833=>"111111111",
  38834=>"101011111",
  38835=>"000001000",
  38836=>"001001011",
  38837=>"000000000",
  38838=>"001111000",
  38839=>"000011110",
  38840=>"111111100",
  38841=>"000000000",
  38842=>"111111000",
  38843=>"000000001",
  38844=>"111111000",
  38845=>"111111100",
  38846=>"100111111",
  38847=>"110111100",
  38848=>"000000101",
  38849=>"000000111",
  38850=>"111101111",
  38851=>"000000000",
  38852=>"000011111",
  38853=>"011011111",
  38854=>"000000000",
  38855=>"001000000",
  38856=>"000000000",
  38857=>"111111111",
  38858=>"111111111",
  38859=>"001111000",
  38860=>"000101000",
  38861=>"111111111",
  38862=>"100100101",
  38863=>"001111101",
  38864=>"000000111",
  38865=>"111000011",
  38866=>"000000000",
  38867=>"100000111",
  38868=>"001010110",
  38869=>"001001000",
  38870=>"000000000",
  38871=>"000000111",
  38872=>"001000000",
  38873=>"111100000",
  38874=>"000010111",
  38875=>"000010000",
  38876=>"111111001",
  38877=>"111111111",
  38878=>"000000011",
  38879=>"110111111",
  38880=>"110111111",
  38881=>"000000000",
  38882=>"111000111",
  38883=>"110111111",
  38884=>"110000010",
  38885=>"001001000",
  38886=>"101001101",
  38887=>"011111111",
  38888=>"111011111",
  38889=>"111111111",
  38890=>"011011111",
  38891=>"111111111",
  38892=>"110000001",
  38893=>"001000001",
  38894=>"000111111",
  38895=>"000111111",
  38896=>"000000110",
  38897=>"000100000",
  38898=>"111011001",
  38899=>"000100101",
  38900=>"111001011",
  38901=>"100000000",
  38902=>"000000111",
  38903=>"000111111",
  38904=>"000000111",
  38905=>"001001011",
  38906=>"000000000",
  38907=>"111111000",
  38908=>"000011011",
  38909=>"111111111",
  38910=>"111011000",
  38911=>"001000000",
  38912=>"111101101",
  38913=>"000000000",
  38914=>"000001000",
  38915=>"001111000",
  38916=>"100111111",
  38917=>"111111111",
  38918=>"000000000",
  38919=>"111001001",
  38920=>"000000000",
  38921=>"100100110",
  38922=>"101101011",
  38923=>"000000000",
  38924=>"010000000",
  38925=>"011101111",
  38926=>"000000011",
  38927=>"000000000",
  38928=>"111111111",
  38929=>"111111111",
  38930=>"111111100",
  38931=>"101001000",
  38932=>"111111111",
  38933=>"000000000",
  38934=>"100000000",
  38935=>"110110110",
  38936=>"000100000",
  38937=>"100000000",
  38938=>"000000111",
  38939=>"100000000",
  38940=>"000000000",
  38941=>"000110000",
  38942=>"000000100",
  38943=>"101111111",
  38944=>"010000000",
  38945=>"000100011",
  38946=>"111110111",
  38947=>"000000010",
  38948=>"111001001",
  38949=>"111111111",
  38950=>"001001000",
  38951=>"000100000",
  38952=>"111111111",
  38953=>"000000111",
  38954=>"111111111",
  38955=>"000100100",
  38956=>"110010010",
  38957=>"000000000",
  38958=>"111111001",
  38959=>"000000000",
  38960=>"111111111",
  38961=>"000000000",
  38962=>"100111111",
  38963=>"100100000",
  38964=>"111111111",
  38965=>"000011111",
  38966=>"111111111",
  38967=>"100111111",
  38968=>"000000111",
  38969=>"000000001",
  38970=>"000000000",
  38971=>"111001000",
  38972=>"111111111",
  38973=>"111110100",
  38974=>"111111110",
  38975=>"101111111",
  38976=>"111111111",
  38977=>"111111111",
  38978=>"100111111",
  38979=>"111111110",
  38980=>"111111110",
  38981=>"000000000",
  38982=>"000000000",
  38983=>"000000000",
  38984=>"111001001",
  38985=>"111111111",
  38986=>"000000111",
  38987=>"000000000",
  38988=>"111111000",
  38989=>"111110110",
  38990=>"000100111",
  38991=>"111010111",
  38992=>"000000000",
  38993=>"000000000",
  38994=>"111100000",
  38995=>"000000110",
  38996=>"111100100",
  38997=>"000000001",
  38998=>"000110011",
  38999=>"000000001",
  39000=>"000000000",
  39001=>"000000001",
  39002=>"000000111",
  39003=>"111111111",
  39004=>"000000000",
  39005=>"000110111",
  39006=>"001000000",
  39007=>"111111111",
  39008=>"011111111",
  39009=>"000000110",
  39010=>"000110111",
  39011=>"000000000",
  39012=>"100100000",
  39013=>"000000000",
  39014=>"100100110",
  39015=>"000000000",
  39016=>"000001111",
  39017=>"111111100",
  39018=>"000000000",
  39019=>"100000010",
  39020=>"101101101",
  39021=>"111111111",
  39022=>"100100000",
  39023=>"000100111",
  39024=>"000111111",
  39025=>"000100111",
  39026=>"000000100",
  39027=>"000000000",
  39028=>"111111000",
  39029=>"110110000",
  39030=>"111110110",
  39031=>"110001000",
  39032=>"100110110",
  39033=>"110111111",
  39034=>"111111111",
  39035=>"101100100",
  39036=>"100100100",
  39037=>"111001000",
  39038=>"111111111",
  39039=>"100111111",
  39040=>"000000000",
  39041=>"000100100",
  39042=>"111111111",
  39043=>"000100100",
  39044=>"001000000",
  39045=>"111111111",
  39046=>"000111100",
  39047=>"000000000",
  39048=>"001000000",
  39049=>"111111111",
  39050=>"111111000",
  39051=>"011001001",
  39052=>"000000100",
  39053=>"000100110",
  39054=>"111111111",
  39055=>"111111111",
  39056=>"111111111",
  39057=>"000010111",
  39058=>"111111111",
  39059=>"000001000",
  39060=>"000000000",
  39061=>"111111111",
  39062=>"000000111",
  39063=>"000000000",
  39064=>"000000110",
  39065=>"000000000",
  39066=>"000000000",
  39067=>"111111111",
  39068=>"100000000",
  39069=>"100000001",
  39070=>"111111111",
  39071=>"000000000",
  39072=>"000000000",
  39073=>"000000000",
  39074=>"111110000",
  39075=>"000000000",
  39076=>"011011100",
  39077=>"000000000",
  39078=>"000000000",
  39079=>"000000111",
  39080=>"111111111",
  39081=>"000000000",
  39082=>"000000011",
  39083=>"111110110",
  39084=>"111111100",
  39085=>"111111101",
  39086=>"101111111",
  39087=>"000000011",
  39088=>"111111000",
  39089=>"111011111",
  39090=>"110110110",
  39091=>"010000111",
  39092=>"101001111",
  39093=>"011000000",
  39094=>"111111111",
  39095=>"111110100",
  39096=>"111111111",
  39097=>"001000000",
  39098=>"111111000",
  39099=>"111111010",
  39100=>"000100111",
  39101=>"000000000",
  39102=>"111111111",
  39103=>"000000100",
  39104=>"111111110",
  39105=>"000000000",
  39106=>"001000000",
  39107=>"111111111",
  39108=>"001001000",
  39109=>"101111111",
  39110=>"001000000",
  39111=>"111111111",
  39112=>"111011000",
  39113=>"111000111",
  39114=>"000000000",
  39115=>"000000000",
  39116=>"000000000",
  39117=>"111011000",
  39118=>"111111111",
  39119=>"100100111",
  39120=>"001001011",
  39121=>"011011000",
  39122=>"000000000",
  39123=>"000000000",
  39124=>"001001111",
  39125=>"111111111",
  39126=>"111111111",
  39127=>"000000000",
  39128=>"111111111",
  39129=>"000100000",
  39130=>"000001000",
  39131=>"001111111",
  39132=>"000000000",
  39133=>"111111111",
  39134=>"000111110",
  39135=>"000100100",
  39136=>"111111111",
  39137=>"010110110",
  39138=>"000000100",
  39139=>"111111001",
  39140=>"000000000",
  39141=>"111111111",
  39142=>"111111110",
  39143=>"111111111",
  39144=>"110010100",
  39145=>"000000000",
  39146=>"111010000",
  39147=>"111111111",
  39148=>"000000000",
  39149=>"000111111",
  39150=>"000000000",
  39151=>"000000000",
  39152=>"100100000",
  39153=>"111010001",
  39154=>"111010000",
  39155=>"000000110",
  39156=>"000000000",
  39157=>"111111110",
  39158=>"001100111",
  39159=>"000000100",
  39160=>"100000101",
  39161=>"000000000",
  39162=>"111111111",
  39163=>"000001001",
  39164=>"101001001",
  39165=>"000000111",
  39166=>"001101101",
  39167=>"001000000",
  39168=>"000000000",
  39169=>"111111111",
  39170=>"000000111",
  39171=>"000110010",
  39172=>"100000000",
  39173=>"000011010",
  39174=>"001001111",
  39175=>"000000000",
  39176=>"000000000",
  39177=>"000000010",
  39178=>"111111110",
  39179=>"000000000",
  39180=>"111111111",
  39181=>"100000000",
  39182=>"111111000",
  39183=>"111101111",
  39184=>"001100000",
  39185=>"100100001",
  39186=>"100000111",
  39187=>"111011001",
  39188=>"000000000",
  39189=>"111111101",
  39190=>"011111111",
  39191=>"111000000",
  39192=>"111111111",
  39193=>"000000000",
  39194=>"101111100",
  39195=>"000100100",
  39196=>"000001101",
  39197=>"000100000",
  39198=>"000000000",
  39199=>"011010000",
  39200=>"000001001",
  39201=>"000000000",
  39202=>"000000111",
  39203=>"000000000",
  39204=>"110110000",
  39205=>"111111111",
  39206=>"110111111",
  39207=>"000010000",
  39208=>"000000000",
  39209=>"110100000",
  39210=>"000000000",
  39211=>"000000111",
  39212=>"110100111",
  39213=>"111011001",
  39214=>"000111111",
  39215=>"001000111",
  39216=>"101100110",
  39217=>"111110110",
  39218=>"101000000",
  39219=>"111110000",
  39220=>"011111111",
  39221=>"100000000",
  39222=>"011111111",
  39223=>"000000000",
  39224=>"111111111",
  39225=>"000000000",
  39226=>"111110000",
  39227=>"110111110",
  39228=>"000101111",
  39229=>"100111111",
  39230=>"000111111",
  39231=>"100110000",
  39232=>"000111111",
  39233=>"011111010",
  39234=>"111110111",
  39235=>"111111111",
  39236=>"000110000",
  39237=>"111011001",
  39238=>"111111111",
  39239=>"000000000",
  39240=>"101101111",
  39241=>"000000010",
  39242=>"000000000",
  39243=>"001011111",
  39244=>"111001011",
  39245=>"000111111",
  39246=>"000000000",
  39247=>"100110110",
  39248=>"111111111",
  39249=>"000001111",
  39250=>"000111111",
  39251=>"000000111",
  39252=>"000000000",
  39253=>"011011011",
  39254=>"000000000",
  39255=>"111000111",
  39256=>"111000000",
  39257=>"000010000",
  39258=>"000000000",
  39259=>"111111110",
  39260=>"000000000",
  39261=>"000000000",
  39262=>"001100100",
  39263=>"111111111",
  39264=>"001101101",
  39265=>"011000000",
  39266=>"001000001",
  39267=>"000000000",
  39268=>"000010111",
  39269=>"000000100",
  39270=>"000000000",
  39271=>"000110010",
  39272=>"001111100",
  39273=>"000000000",
  39274=>"000000000",
  39275=>"000000101",
  39276=>"001101100",
  39277=>"000000000",
  39278=>"000111111",
  39279=>"000111111",
  39280=>"000000111",
  39281=>"010000101",
  39282=>"001000000",
  39283=>"001000000",
  39284=>"000110000",
  39285=>"000000101",
  39286=>"111111111",
  39287=>"110111000",
  39288=>"000000000",
  39289=>"000000000",
  39290=>"000000000",
  39291=>"000010111",
  39292=>"100100001",
  39293=>"111111111",
  39294=>"111000000",
  39295=>"111111111",
  39296=>"111111111",
  39297=>"111111111",
  39298=>"010010110",
  39299=>"000000000",
  39300=>"101111111",
  39301=>"011011011",
  39302=>"111111011",
  39303=>"111111111",
  39304=>"000000111",
  39305=>"000000100",
  39306=>"000000000",
  39307=>"010010011",
  39308=>"111111111",
  39309=>"111111111",
  39310=>"111111100",
  39311=>"000000000",
  39312=>"111111111",
  39313=>"111000000",
  39314=>"111000000",
  39315=>"000000101",
  39316=>"111000000",
  39317=>"011011011",
  39318=>"000000100",
  39319=>"101000001",
  39320=>"010100110",
  39321=>"110110111",
  39322=>"000000000",
  39323=>"000000111",
  39324=>"110110100",
  39325=>"000000000",
  39326=>"000000000",
  39327=>"100000000",
  39328=>"110110111",
  39329=>"000000110",
  39330=>"000000000",
  39331=>"100111111",
  39332=>"100101101",
  39333=>"110000000",
  39334=>"111111101",
  39335=>"001001100",
  39336=>"111011000",
  39337=>"111111110",
  39338=>"000000000",
  39339=>"001001111",
  39340=>"000000000",
  39341=>"001000011",
  39342=>"000001101",
  39343=>"000100100",
  39344=>"000000000",
  39345=>"111110100",
  39346=>"000000000",
  39347=>"111111111",
  39348=>"000000000",
  39349=>"111111000",
  39350=>"111101101",
  39351=>"111111111",
  39352=>"110111000",
  39353=>"111111111",
  39354=>"111011010",
  39355=>"111111001",
  39356=>"000001111",
  39357=>"011101111",
  39358=>"110111111",
  39359=>"011011111",
  39360=>"111111011",
  39361=>"111111111",
  39362=>"111111011",
  39363=>"111111001",
  39364=>"000000101",
  39365=>"111111111",
  39366=>"001011011",
  39367=>"111111111",
  39368=>"001000111",
  39369=>"101111000",
  39370=>"101111011",
  39371=>"001011111",
  39372=>"110011111",
  39373=>"111000001",
  39374=>"011111111",
  39375=>"001101000",
  39376=>"000000011",
  39377=>"000100111",
  39378=>"111111011",
  39379=>"000010000",
  39380=>"111111011",
  39381=>"000000000",
  39382=>"000000000",
  39383=>"000111011",
  39384=>"101101111",
  39385=>"010111110",
  39386=>"111110000",
  39387=>"000000000",
  39388=>"000111110",
  39389=>"001000000",
  39390=>"000000000",
  39391=>"111000000",
  39392=>"001011110",
  39393=>"000000000",
  39394=>"000000110",
  39395=>"111111111",
  39396=>"001111111",
  39397=>"110010111",
  39398=>"011011010",
  39399=>"001001100",
  39400=>"000000000",
  39401=>"001011111",
  39402=>"000111111",
  39403=>"111111111",
  39404=>"100000000",
  39405=>"001110100",
  39406=>"000001011",
  39407=>"111111111",
  39408=>"011001001",
  39409=>"110111110",
  39410=>"000000111",
  39411=>"110111111",
  39412=>"111111111",
  39413=>"110111111",
  39414=>"000000100",
  39415=>"101111111",
  39416=>"110111111",
  39417=>"100101111",
  39418=>"100010000",
  39419=>"001001001",
  39420=>"000010110",
  39421=>"000000100",
  39422=>"111111111",
  39423=>"000000000",
  39424=>"110111110",
  39425=>"110100000",
  39426=>"101000100",
  39427=>"111111010",
  39428=>"100000010",
  39429=>"111111011",
  39430=>"111101111",
  39431=>"001000101",
  39432=>"111000000",
  39433=>"000000000",
  39434=>"001000111",
  39435=>"011111011",
  39436=>"001000100",
  39437=>"100000000",
  39438=>"000000010",
  39439=>"000000110",
  39440=>"111100000",
  39441=>"000000100",
  39442=>"110000000",
  39443=>"011111111",
  39444=>"111111111",
  39445=>"000000001",
  39446=>"100111111",
  39447=>"110110100",
  39448=>"000000000",
  39449=>"100110000",
  39450=>"000000101",
  39451=>"111111111",
  39452=>"100000000",
  39453=>"111011000",
  39454=>"000000000",
  39455=>"111111100",
  39456=>"110111110",
  39457=>"000000000",
  39458=>"111111111",
  39459=>"100000110",
  39460=>"000000000",
  39461=>"001000000",
  39462=>"100001000",
  39463=>"111111111",
  39464=>"100000111",
  39465=>"111000000",
  39466=>"001000010",
  39467=>"111111111",
  39468=>"000000111",
  39469=>"111111000",
  39470=>"000000000",
  39471=>"000010010",
  39472=>"000000000",
  39473=>"110111111",
  39474=>"100101011",
  39475=>"001000110",
  39476=>"110110110",
  39477=>"000100100",
  39478=>"110101100",
  39479=>"000000001",
  39480=>"000000111",
  39481=>"000000111",
  39482=>"000000000",
  39483=>"010000011",
  39484=>"101101100",
  39485=>"000000000",
  39486=>"000111111",
  39487=>"100100100",
  39488=>"000000000",
  39489=>"101010000",
  39490=>"111111111",
  39491=>"111111000",
  39492=>"000000000",
  39493=>"110110000",
  39494=>"000001000",
  39495=>"100101101",
  39496=>"111011011",
  39497=>"001000001",
  39498=>"111111000",
  39499=>"100000000",
  39500=>"110110000",
  39501=>"011001111",
  39502=>"001000010",
  39503=>"110000000",
  39504=>"000110110",
  39505=>"111001001",
  39506=>"111111010",
  39507=>"000000000",
  39508=>"110100101",
  39509=>"100000000",
  39510=>"000000011",
  39511=>"110110110",
  39512=>"110111111",
  39513=>"101001111",
  39514=>"000000001",
  39515=>"111111111",
  39516=>"111110010",
  39517=>"001001111",
  39518=>"011001000",
  39519=>"011011001",
  39520=>"111101111",
  39521=>"000000111",
  39522=>"111001111",
  39523=>"100111111",
  39524=>"000100110",
  39525=>"000000000",
  39526=>"111001000",
  39527=>"111011011",
  39528=>"011010001",
  39529=>"001001101",
  39530=>"111101111",
  39531=>"000000000",
  39532=>"100101001",
  39533=>"111111111",
  39534=>"000010000",
  39535=>"000000000",
  39536=>"000000000",
  39537=>"000000000",
  39538=>"111111111",
  39539=>"000000000",
  39540=>"000100111",
  39541=>"000000000",
  39542=>"000000000",
  39543=>"000000101",
  39544=>"000000000",
  39545=>"000000000",
  39546=>"000001000",
  39547=>"111111000",
  39548=>"100110110",
  39549=>"000000000",
  39550=>"000000000",
  39551=>"000000111",
  39552=>"000000110",
  39553=>"111111101",
  39554=>"111001011",
  39555=>"111011111",
  39556=>"111111111",
  39557=>"010010000",
  39558=>"110111000",
  39559=>"110110010",
  39560=>"111111100",
  39561=>"000000000",
  39562=>"000000000",
  39563=>"110110100",
  39564=>"100000000",
  39565=>"111111111",
  39566=>"101000000",
  39567=>"100100000",
  39568=>"000000000",
  39569=>"000000000",
  39570=>"111111000",
  39571=>"000000001",
  39572=>"000000000",
  39573=>"000000000",
  39574=>"101111111",
  39575=>"100100110",
  39576=>"000000011",
  39577=>"111111111",
  39578=>"100111111",
  39579=>"011000000",
  39580=>"001011001",
  39581=>"110000000",
  39582=>"110000000",
  39583=>"111000000",
  39584=>"000000101",
  39585=>"110110110",
  39586=>"000000011",
  39587=>"011111110",
  39588=>"000000100",
  39589=>"011011111",
  39590=>"111111111",
  39591=>"011111111",
  39592=>"111111011",
  39593=>"000000101",
  39594=>"111111111",
  39595=>"000000000",
  39596=>"011000001",
  39597=>"100100000",
  39598=>"000110000",
  39599=>"001001111",
  39600=>"111010000",
  39601=>"111111100",
  39602=>"111111111",
  39603=>"000000100",
  39604=>"111001100",
  39605=>"000000111",
  39606=>"000000100",
  39607=>"000000000",
  39608=>"110111111",
  39609=>"001001111",
  39610=>"000000000",
  39611=>"111111000",
  39612=>"111001001",
  39613=>"010110110",
  39614=>"111110000",
  39615=>"110111010",
  39616=>"000000100",
  39617=>"101101111",
  39618=>"001001111",
  39619=>"001000011",
  39620=>"001111101",
  39621=>"101111111",
  39622=>"000000000",
  39623=>"000000000",
  39624=>"000000000",
  39625=>"000100000",
  39626=>"000000001",
  39627=>"110110000",
  39628=>"001000001",
  39629=>"111111111",
  39630=>"111000000",
  39631=>"111111000",
  39632=>"000000000",
  39633=>"110111011",
  39634=>"110111111",
  39635=>"000000000",
  39636=>"110111001",
  39637=>"011011011",
  39638=>"111111000",
  39639=>"111011101",
  39640=>"001011011",
  39641=>"110110111",
  39642=>"111000000",
  39643=>"111001000",
  39644=>"111111110",
  39645=>"111111000",
  39646=>"101111001",
  39647=>"000000000",
  39648=>"111000001",
  39649=>"000000111",
  39650=>"111000110",
  39651=>"000000000",
  39652=>"000000000",
  39653=>"110110110",
  39654=>"000000000",
  39655=>"100100111",
  39656=>"001000000",
  39657=>"110111000",
  39658=>"001001011",
  39659=>"001001001",
  39660=>"010110110",
  39661=>"000011011",
  39662=>"011001000",
  39663=>"110111111",
  39664=>"000000100",
  39665=>"111111000",
  39666=>"000010110",
  39667=>"100000111",
  39668=>"000000000",
  39669=>"110010000",
  39670=>"011000000",
  39671=>"111001001",
  39672=>"000000000",
  39673=>"000000000",
  39674=>"100000000",
  39675=>"000000000",
  39676=>"100110000",
  39677=>"000000000",
  39678=>"000111111",
  39679=>"001000001",
  39680=>"110110111",
  39681=>"000010110",
  39682=>"111111111",
  39683=>"011110111",
  39684=>"100101011",
  39685=>"000000000",
  39686=>"000000000",
  39687=>"111000000",
  39688=>"000000001",
  39689=>"000000111",
  39690=>"111111010",
  39691=>"111011001",
  39692=>"001101111",
  39693=>"111110111",
  39694=>"111111111",
  39695=>"000001001",
  39696=>"000000000",
  39697=>"110111110",
  39698=>"101100111",
  39699=>"110000000",
  39700=>"100111111",
  39701=>"111111111",
  39702=>"001011001",
  39703=>"111111111",
  39704=>"110111111",
  39705=>"001000010",
  39706=>"000001000",
  39707=>"000100110",
  39708=>"111110100",
  39709=>"111000000",
  39710=>"010111100",
  39711=>"111111111",
  39712=>"000000000",
  39713=>"110111111",
  39714=>"111111000",
  39715=>"000000001",
  39716=>"000000000",
  39717=>"111011000",
  39718=>"000110110",
  39719=>"000000001",
  39720=>"111111011",
  39721=>"111111010",
  39722=>"100000110",
  39723=>"000000000",
  39724=>"000000000",
  39725=>"100001000",
  39726=>"000000000",
  39727=>"000000100",
  39728=>"000001000",
  39729=>"000000000",
  39730=>"000000001",
  39731=>"000000000",
  39732=>"011011001",
  39733=>"101111110",
  39734=>"001000000",
  39735=>"111100000",
  39736=>"000000100",
  39737=>"101101101",
  39738=>"011011111",
  39739=>"111111111",
  39740=>"000000011",
  39741=>"111111111",
  39742=>"000111111",
  39743=>"000100100",
  39744=>"010000000",
  39745=>"111111000",
  39746=>"000111111",
  39747=>"000000001",
  39748=>"000010011",
  39749=>"001000000",
  39750=>"000000000",
  39751=>"000000100",
  39752=>"000000001",
  39753=>"110110000",
  39754=>"001000000",
  39755=>"100001001",
  39756=>"011000000",
  39757=>"111101100",
  39758=>"001010011",
  39759=>"010010011",
  39760=>"100100100",
  39761=>"000000000",
  39762=>"000000110",
  39763=>"111111111",
  39764=>"000000000",
  39765=>"011011011",
  39766=>"111000000",
  39767=>"110111111",
  39768=>"111111000",
  39769=>"101000111",
  39770=>"000000000",
  39771=>"000000011",
  39772=>"000001011",
  39773=>"010010010",
  39774=>"000000000",
  39775=>"100000000",
  39776=>"000000101",
  39777=>"100000111",
  39778=>"000000100",
  39779=>"111111111",
  39780=>"100100000",
  39781=>"000000000",
  39782=>"111000000",
  39783=>"000110110",
  39784=>"000000000",
  39785=>"001000000",
  39786=>"111111010",
  39787=>"010111111",
  39788=>"000001000",
  39789=>"000110111",
  39790=>"000111111",
  39791=>"000000000",
  39792=>"000111000",
  39793=>"110100000",
  39794=>"110100111",
  39795=>"111111111",
  39796=>"000111011",
  39797=>"100100100",
  39798=>"111111000",
  39799=>"111111111",
  39800=>"000000111",
  39801=>"000000000",
  39802=>"000101111",
  39803=>"000000000",
  39804=>"000010010",
  39805=>"001001001",
  39806=>"001111111",
  39807=>"111111111",
  39808=>"000001000",
  39809=>"111011111",
  39810=>"111111111",
  39811=>"000111111",
  39812=>"111111111",
  39813=>"000001111",
  39814=>"100111111",
  39815=>"010011011",
  39816=>"111111000",
  39817=>"101001000",
  39818=>"111111111",
  39819=>"011011000",
  39820=>"001001111",
  39821=>"000111111",
  39822=>"111101101",
  39823=>"000000000",
  39824=>"000000100",
  39825=>"110111111",
  39826=>"111111111",
  39827=>"111111100",
  39828=>"000000000",
  39829=>"000010110",
  39830=>"110011011",
  39831=>"000101111",
  39832=>"111111111",
  39833=>"100111011",
  39834=>"100100101",
  39835=>"000000111",
  39836=>"111111011",
  39837=>"100100110",
  39838=>"111110010",
  39839=>"111000000",
  39840=>"001001001",
  39841=>"011111000",
  39842=>"010000000",
  39843=>"111111010",
  39844=>"000011000",
  39845=>"001101000",
  39846=>"111111001",
  39847=>"111111111",
  39848=>"000100100",
  39849=>"000000010",
  39850=>"011110110",
  39851=>"100100110",
  39852=>"100000110",
  39853=>"111110000",
  39854=>"100111000",
  39855=>"011011011",
  39856=>"100000000",
  39857=>"111000000",
  39858=>"111111111",
  39859=>"100100111",
  39860=>"100000000",
  39861=>"100100000",
  39862=>"111110100",
  39863=>"011011110",
  39864=>"111111111",
  39865=>"111010000",
  39866=>"000000000",
  39867=>"000000000",
  39868=>"111111111",
  39869=>"111111111",
  39870=>"100101111",
  39871=>"000011000",
  39872=>"001000000",
  39873=>"000000000",
  39874=>"000101101",
  39875=>"000000010",
  39876=>"111111111",
  39877=>"100100100",
  39878=>"111111111",
  39879=>"100000011",
  39880=>"000000000",
  39881=>"000100000",
  39882=>"101001001",
  39883=>"111111000",
  39884=>"000000000",
  39885=>"010111111",
  39886=>"111011011",
  39887=>"000111111",
  39888=>"011010000",
  39889=>"111000010",
  39890=>"111111111",
  39891=>"111110000",
  39892=>"000000000",
  39893=>"110111111",
  39894=>"111101000",
  39895=>"110110111",
  39896=>"110111111",
  39897=>"100100100",
  39898=>"000000010",
  39899=>"111111100",
  39900=>"111111111",
  39901=>"000000011",
  39902=>"000000011",
  39903=>"000100000",
  39904=>"110010010",
  39905=>"000000001",
  39906=>"000000110",
  39907=>"000000100",
  39908=>"111111011",
  39909=>"001111110",
  39910=>"100100110",
  39911=>"011011010",
  39912=>"111110110",
  39913=>"000100110",
  39914=>"000000000",
  39915=>"011111011",
  39916=>"100100000",
  39917=>"111100100",
  39918=>"000000110",
  39919=>"000010110",
  39920=>"111000111",
  39921=>"111111000",
  39922=>"000000111",
  39923=>"000000000",
  39924=>"100111011",
  39925=>"000000100",
  39926=>"000000000",
  39927=>"000000000",
  39928=>"111111111",
  39929=>"110111111",
  39930=>"000000001",
  39931=>"111001000",
  39932=>"111111000",
  39933=>"111111111",
  39934=>"000000000",
  39935=>"100110111",
  39936=>"000000000",
  39937=>"000000000",
  39938=>"001101111",
  39939=>"000000000",
  39940=>"001001111",
  39941=>"001000000",
  39942=>"000000000",
  39943=>"111111100",
  39944=>"111111101",
  39945=>"000000000",
  39946=>"100111111",
  39947=>"111111111",
  39948=>"000000000",
  39949=>"000000000",
  39950=>"100100100",
  39951=>"000100111",
  39952=>"111111111",
  39953=>"000000000",
  39954=>"111111111",
  39955=>"000001101",
  39956=>"000000111",
  39957=>"001000001",
  39958=>"000000000",
  39959=>"111100111",
  39960=>"111111111",
  39961=>"100101111",
  39962=>"001000000",
  39963=>"000000000",
  39964=>"111111111",
  39965=>"000000000",
  39966=>"001001001",
  39967=>"000100000",
  39968=>"111110000",
  39969=>"111111110",
  39970=>"001001111",
  39971=>"100100110",
  39972=>"000000000",
  39973=>"111000000",
  39974=>"000000000",
  39975=>"111101111",
  39976=>"100100110",
  39977=>"000000000",
  39978=>"111111111",
  39979=>"111111111",
  39980=>"100000101",
  39981=>"000000000",
  39982=>"111111000",
  39983=>"111111111",
  39984=>"100000000",
  39985=>"000000000",
  39986=>"000000100",
  39987=>"110100000",
  39988=>"110111111",
  39989=>"000100001",
  39990=>"000101101",
  39991=>"100100110",
  39992=>"000000000",
  39993=>"110100110",
  39994=>"000001111",
  39995=>"000111111",
  39996=>"000010011",
  39997=>"000000000",
  39998=>"011010000",
  39999=>"111000000",
  40000=>"111001000",
  40001=>"000000000",
  40002=>"111011111",
  40003=>"000000000",
  40004=>"111011000",
  40005=>"001001111",
  40006=>"111111010",
  40007=>"010000000",
  40008=>"001001011",
  40009=>"000000000",
  40010=>"111100111",
  40011=>"000000000",
  40012=>"000000000",
  40013=>"010000011",
  40014=>"111111111",
  40015=>"000000000",
  40016=>"000000000",
  40017=>"111111111",
  40018=>"110000000",
  40019=>"111011001",
  40020=>"000000001",
  40021=>"111111111",
  40022=>"100100000",
  40023=>"000111010",
  40024=>"000000000",
  40025=>"111110111",
  40026=>"000001011",
  40027=>"000110110",
  40028=>"000000000",
  40029=>"111111111",
  40030=>"000000100",
  40031=>"001000111",
  40032=>"000000000",
  40033=>"011000000",
  40034=>"000000000",
  40035=>"100000000",
  40036=>"111111000",
  40037=>"001000000",
  40038=>"000010000",
  40039=>"111111111",
  40040=>"000111001",
  40041=>"111101100",
  40042=>"000111111",
  40043=>"000000000",
  40044=>"000000000",
  40045=>"001111111",
  40046=>"111111111",
  40047=>"000000000",
  40048=>"000000001",
  40049=>"000000000",
  40050=>"011111111",
  40051=>"000000000",
  40052=>"111111111",
  40053=>"101101111",
  40054=>"111100100",
  40055=>"111111001",
  40056=>"001111111",
  40057=>"111111110",
  40058=>"010111010",
  40059=>"111111111",
  40060=>"110110110",
  40061=>"000000111",
  40062=>"110000000",
  40063=>"000000110",
  40064=>"111110101",
  40065=>"000000101",
  40066=>"001000000",
  40067=>"000000000",
  40068=>"111111011",
  40069=>"101111001",
  40070=>"000000000",
  40071=>"100000000",
  40072=>"001111000",
  40073=>"100000000",
  40074=>"000000000",
  40075=>"000000000",
  40076=>"100011111",
  40077=>"010100000",
  40078=>"000001000",
  40079=>"111111111",
  40080=>"111111000",
  40081=>"100000111",
  40082=>"000000011",
  40083=>"010111000",
  40084=>"011011000",
  40085=>"000000111",
  40086=>"111101111",
  40087=>"000000000",
  40088=>"001111111",
  40089=>"001001111",
  40090=>"000000110",
  40091=>"000000000",
  40092=>"000000000",
  40093=>"101111111",
  40094=>"100111011",
  40095=>"000111111",
  40096=>"000100111",
  40097=>"110110010",
  40098=>"111101111",
  40099=>"000000111",
  40100=>"000000000",
  40101=>"111111111",
  40102=>"110110000",
  40103=>"110011001",
  40104=>"100100111",
  40105=>"000001101",
  40106=>"111000000",
  40107=>"110110110",
  40108=>"101111111",
  40109=>"001000000",
  40110=>"111001000",
  40111=>"111111001",
  40112=>"010111111",
  40113=>"111111111",
  40114=>"111111111",
  40115=>"111111111",
  40116=>"111000000",
  40117=>"111111111",
  40118=>"000000000",
  40119=>"000110111",
  40120=>"110111111",
  40121=>"000110111",
  40122=>"000000000",
  40123=>"000000000",
  40124=>"111111111",
  40125=>"111111111",
  40126=>"111111111",
  40127=>"000000001",
  40128=>"110111111",
  40129=>"110111111",
  40130=>"011001000",
  40131=>"110110000",
  40132=>"101101111",
  40133=>"101110110",
  40134=>"010110111",
  40135=>"000000000",
  40136=>"000001111",
  40137=>"000111111",
  40138=>"000000110",
  40139=>"111111110",
  40140=>"001000000",
  40141=>"111100101",
  40142=>"111111001",
  40143=>"111111111",
  40144=>"000100100",
  40145=>"000000000",
  40146=>"101111111",
  40147=>"000000000",
  40148=>"000000001",
  40149=>"111111111",
  40150=>"000000000",
  40151=>"101000000",
  40152=>"100100100",
  40153=>"100100101",
  40154=>"000000000",
  40155=>"000110101",
  40156=>"000111010",
  40157=>"000001101",
  40158=>"010111110",
  40159=>"000010000",
  40160=>"000000000",
  40161=>"000000000",
  40162=>"111111111",
  40163=>"111111111",
  40164=>"001111110",
  40165=>"000000001",
  40166=>"000000000",
  40167=>"111111111",
  40168=>"000000111",
  40169=>"111111111",
  40170=>"111111111",
  40171=>"000000000",
  40172=>"000111100",
  40173=>"000010000",
  40174=>"111111111",
  40175=>"011111011",
  40176=>"111111111",
  40177=>"100100111",
  40178=>"000000010",
  40179=>"000000000",
  40180=>"101111010",
  40181=>"100110100",
  40182=>"000100011",
  40183=>"000000000",
  40184=>"111110100",
  40185=>"000000000",
  40186=>"000110111",
  40187=>"000001001",
  40188=>"010110111",
  40189=>"000001110",
  40190=>"000111111",
  40191=>"011001100",
  40192=>"000000111",
  40193=>"000001001",
  40194=>"111111111",
  40195=>"000011111",
  40196=>"101101111",
  40197=>"000000000",
  40198=>"100110111",
  40199=>"000100001",
  40200=>"000000110",
  40201=>"111111111",
  40202=>"000000000",
  40203=>"000000101",
  40204=>"000000011",
  40205=>"000000111",
  40206=>"101111111",
  40207=>"110111111",
  40208=>"110111000",
  40209=>"111111111",
  40210=>"000000000",
  40211=>"110000111",
  40212=>"101101000",
  40213=>"111111111",
  40214=>"100100100",
  40215=>"011011000",
  40216=>"000001111",
  40217=>"000000000",
  40218=>"000011011",
  40219=>"001000100",
  40220=>"110110110",
  40221=>"000000000",
  40222=>"111111111",
  40223=>"000000000",
  40224=>"100110111",
  40225=>"111011111",
  40226=>"000000011",
  40227=>"001001101",
  40228=>"000000000",
  40229=>"001011011",
  40230=>"000100000",
  40231=>"100000010",
  40232=>"100111100",
  40233=>"000001111",
  40234=>"000000000",
  40235=>"000000000",
  40236=>"000111111",
  40237=>"100111101",
  40238=>"111110000",
  40239=>"000000000",
  40240=>"110111011",
  40241=>"000111111",
  40242=>"111111111",
  40243=>"011000000",
  40244=>"100100000",
  40245=>"000000100",
  40246=>"001001000",
  40247=>"000000000",
  40248=>"000111111",
  40249=>"000000000",
  40250=>"101111111",
  40251=>"111111001",
  40252=>"000000001",
  40253=>"000001001",
  40254=>"101111000",
  40255=>"000000000",
  40256=>"000000000",
  40257=>"111111111",
  40258=>"000000000",
  40259=>"110110011",
  40260=>"111111101",
  40261=>"000000000",
  40262=>"111111111",
  40263=>"111111010",
  40264=>"111111110",
  40265=>"000000000",
  40266=>"001001101",
  40267=>"010000000",
  40268=>"000000000",
  40269=>"011010000",
  40270=>"010011001",
  40271=>"000000000",
  40272=>"000001011",
  40273=>"000101101",
  40274=>"000000111",
  40275=>"000000000",
  40276=>"000000001",
  40277=>"001001001",
  40278=>"111111111",
  40279=>"000000000",
  40280=>"000111111",
  40281=>"111000000",
  40282=>"111111111",
  40283=>"111000000",
  40284=>"000000000",
  40285=>"111111111",
  40286=>"111111001",
  40287=>"111110110",
  40288=>"111111111",
  40289=>"000001111",
  40290=>"111111100",
  40291=>"000000000",
  40292=>"010000000",
  40293=>"000111111",
  40294=>"000000000",
  40295=>"001100010",
  40296=>"011000000",
  40297=>"110000000",
  40298=>"110111011",
  40299=>"000000001",
  40300=>"011011001",
  40301=>"010111000",
  40302=>"000111111",
  40303=>"111011000",
  40304=>"100111000",
  40305=>"111111111",
  40306=>"110010111",
  40307=>"100110111",
  40308=>"000000000",
  40309=>"000000000",
  40310=>"000000001",
  40311=>"000000000",
  40312=>"110111111",
  40313=>"000000000",
  40314=>"111111111",
  40315=>"110110110",
  40316=>"110111111",
  40317=>"110111111",
  40318=>"111001000",
  40319=>"111111110",
  40320=>"011000000",
  40321=>"111111110",
  40322=>"100100111",
  40323=>"100101110",
  40324=>"101000111",
  40325=>"000000000",
  40326=>"000100111",
  40327=>"010110010",
  40328=>"000000000",
  40329=>"000000000",
  40330=>"000000111",
  40331=>"111111011",
  40332=>"000000100",
  40333=>"010000001",
  40334=>"100101101",
  40335=>"000100100",
  40336=>"000000000",
  40337=>"000000000",
  40338=>"111000111",
  40339=>"000000000",
  40340=>"111111111",
  40341=>"000010000",
  40342=>"000000111",
  40343=>"101111110",
  40344=>"101111111",
  40345=>"110111011",
  40346=>"111110110",
  40347=>"111111111",
  40348=>"111111111",
  40349=>"000000000",
  40350=>"111111111",
  40351=>"110110000",
  40352=>"000000000",
  40353=>"110100100",
  40354=>"110111110",
  40355=>"000001001",
  40356=>"111111101",
  40357=>"110100111",
  40358=>"000000000",
  40359=>"111111111",
  40360=>"110110000",
  40361=>"000000000",
  40362=>"000100111",
  40363=>"000111111",
  40364=>"000000000",
  40365=>"111111000",
  40366=>"000000000",
  40367=>"010111011",
  40368=>"000000001",
  40369=>"111110111",
  40370=>"001011011",
  40371=>"111101111",
  40372=>"100000100",
  40373=>"111111111",
  40374=>"000000000",
  40375=>"000100000",
  40376=>"011111111",
  40377=>"111000111",
  40378=>"110000000",
  40379=>"111111111",
  40380=>"111111000",
  40381=>"100000000",
  40382=>"111001000",
  40383=>"000000100",
  40384=>"100111000",
  40385=>"111111111",
  40386=>"111111111",
  40387=>"111100000",
  40388=>"101111111",
  40389=>"000001011",
  40390=>"000000110",
  40391=>"111111111",
  40392=>"010110011",
  40393=>"111010000",
  40394=>"000001001",
  40395=>"000000000",
  40396=>"000000000",
  40397=>"000011000",
  40398=>"000000000",
  40399=>"111000000",
  40400=>"111111111",
  40401=>"000000000",
  40402=>"100000011",
  40403=>"111111111",
  40404=>"000000000",
  40405=>"111000111",
  40406=>"000000001",
  40407=>"000100011",
  40408=>"000000000",
  40409=>"111111111",
  40410=>"111111000",
  40411=>"000000111",
  40412=>"000101101",
  40413=>"111100000",
  40414=>"100000000",
  40415=>"100100110",
  40416=>"111011000",
  40417=>"000000010",
  40418=>"000010000",
  40419=>"100000101",
  40420=>"111001000",
  40421=>"000111000",
  40422=>"111111111",
  40423=>"110000000",
  40424=>"111101111",
  40425=>"011111111",
  40426=>"111111011",
  40427=>"000101101",
  40428=>"101111111",
  40429=>"111111001",
  40430=>"111111111",
  40431=>"111111111",
  40432=>"000111110",
  40433=>"000110111",
  40434=>"010011111",
  40435=>"111111110",
  40436=>"000000000",
  40437=>"100100111",
  40438=>"100000000",
  40439=>"111001001",
  40440=>"111111110",
  40441=>"000000011",
  40442=>"000000000",
  40443=>"000000000",
  40444=>"000100000",
  40445=>"111111111",
  40446=>"000000000",
  40447=>"001001000",
  40448=>"111001011",
  40449=>"000000000",
  40450=>"000000000",
  40451=>"000100110",
  40452=>"011010001",
  40453=>"000101001",
  40454=>"000000000",
  40455=>"111111111",
  40456=>"100100001",
  40457=>"111111111",
  40458=>"000000111",
  40459=>"111111000",
  40460=>"000000001",
  40461=>"111111111",
  40462=>"000000000",
  40463=>"011001001",
  40464=>"011111111",
  40465=>"111100000",
  40466=>"111111111",
  40467=>"000000111",
  40468=>"000000000",
  40469=>"111111101",
  40470=>"011110000",
  40471=>"101000101",
  40472=>"111111011",
  40473=>"111001111",
  40474=>"000000111",
  40475=>"000110110",
  40476=>"111111111",
  40477=>"011011011",
  40478=>"011111101",
  40479=>"100100000",
  40480=>"011111111",
  40481=>"000110110",
  40482=>"001101111",
  40483=>"000111110",
  40484=>"000000000",
  40485=>"111111000",
  40486=>"000000000",
  40487=>"000000101",
  40488=>"100000000",
  40489=>"000000000",
  40490=>"111111111",
  40491=>"110111111",
  40492=>"000100001",
  40493=>"000001000",
  40494=>"111101101",
  40495=>"011000010",
  40496=>"111111111",
  40497=>"111111010",
  40498=>"100001001",
  40499=>"000000000",
  40500=>"111111101",
  40501=>"111111111",
  40502=>"111111110",
  40503=>"111111111",
  40504=>"001001111",
  40505=>"011111111",
  40506=>"001001111",
  40507=>"111111111",
  40508=>"101001111",
  40509=>"111000000",
  40510=>"011001001",
  40511=>"000000000",
  40512=>"000000000",
  40513=>"000000000",
  40514=>"000001011",
  40515=>"001111000",
  40516=>"000000000",
  40517=>"001001001",
  40518=>"111111111",
  40519=>"000010111",
  40520=>"000000001",
  40521=>"000000011",
  40522=>"111111111",
  40523=>"000000000",
  40524=>"010111111",
  40525=>"111111111",
  40526=>"000000100",
  40527=>"000000111",
  40528=>"000000000",
  40529=>"111111111",
  40530=>"000000000",
  40531=>"001001000",
  40532=>"111111001",
  40533=>"000000000",
  40534=>"000001111",
  40535=>"111110111",
  40536=>"000000111",
  40537=>"001000000",
  40538=>"000000000",
  40539=>"000000000",
  40540=>"000000101",
  40541=>"111111111",
  40542=>"000000000",
  40543=>"001001000",
  40544=>"000000000",
  40545=>"000000000",
  40546=>"000000000",
  40547=>"000000000",
  40548=>"000000100",
  40549=>"000000100",
  40550=>"000000000",
  40551=>"000110111",
  40552=>"001011111",
  40553=>"000001011",
  40554=>"001000000",
  40555=>"000000000",
  40556=>"011011110",
  40557=>"000000000",
  40558=>"101111111",
  40559=>"000000000",
  40560=>"110111111",
  40561=>"111111100",
  40562=>"010000000",
  40563=>"000000000",
  40564=>"111101001",
  40565=>"100111001",
  40566=>"100000111",
  40567=>"000000011",
  40568=>"000111111",
  40569=>"100100000",
  40570=>"000000010",
  40571=>"000000000",
  40572=>"110110110",
  40573=>"000000111",
  40574=>"111110110",
  40575=>"000000000",
  40576=>"000000000",
  40577=>"000000000",
  40578=>"111111000",
  40579=>"111111111",
  40580=>"001001111",
  40581=>"000000111",
  40582=>"110111100",
  40583=>"000000000",
  40584=>"000000011",
  40585=>"000000001",
  40586=>"000000000",
  40587=>"011001111",
  40588=>"000000000",
  40589=>"000111111",
  40590=>"111001000",
  40591=>"000000100",
  40592=>"100000000",
  40593=>"100000101",
  40594=>"000000010",
  40595=>"011111000",
  40596=>"011111111",
  40597=>"000101101",
  40598=>"001000000",
  40599=>"111101111",
  40600=>"001000001",
  40601=>"111101100",
  40602=>"100111111",
  40603=>"111000100",
  40604=>"111111011",
  40605=>"000000101",
  40606=>"111111111",
  40607=>"111111110",
  40608=>"000000000",
  40609=>"000000000",
  40610=>"110110111",
  40611=>"001000000",
  40612=>"000000000",
  40613=>"111111111",
  40614=>"010011000",
  40615=>"001001111",
  40616=>"000100000",
  40617=>"111111000",
  40618=>"110111010",
  40619=>"100001111",
  40620=>"100000111",
  40621=>"110110110",
  40622=>"111111111",
  40623=>"000001111",
  40624=>"111111111",
  40625=>"111100110",
  40626=>"010111111",
  40627=>"001111101",
  40628=>"111110111",
  40629=>"010111111",
  40630=>"011001001",
  40631=>"001111010",
  40632=>"101000000",
  40633=>"111111011",
  40634=>"000000111",
  40635=>"011010000",
  40636=>"000000000",
  40637=>"111111111",
  40638=>"111111111",
  40639=>"100100110",
  40640=>"111101100",
  40641=>"111100000",
  40642=>"111111000",
  40643=>"111111111",
  40644=>"001000000",
  40645=>"000000000",
  40646=>"111111110",
  40647=>"111111000",
  40648=>"011011111",
  40649=>"100000000",
  40650=>"000000000",
  40651=>"000000000",
  40652=>"111101111",
  40653=>"011001000",
  40654=>"001001111",
  40655=>"000010100",
  40656=>"000100111",
  40657=>"111111111",
  40658=>"000111111",
  40659=>"011011001",
  40660=>"111111001",
  40661=>"111011001",
  40662=>"000000000",
  40663=>"001001000",
  40664=>"111111111",
  40665=>"111111111",
  40666=>"000000000",
  40667=>"100000111",
  40668=>"111111111",
  40669=>"011111111",
  40670=>"000000000",
  40671=>"001001111",
  40672=>"000000011",
  40673=>"000000011",
  40674=>"111111111",
  40675=>"011001000",
  40676=>"100110111",
  40677=>"000000000",
  40678=>"100110110",
  40679=>"111111111",
  40680=>"111100100",
  40681=>"000000100",
  40682=>"111011111",
  40683=>"100000000",
  40684=>"011111111",
  40685=>"000000000",
  40686=>"000000101",
  40687=>"011000000",
  40688=>"000000011",
  40689=>"001101101",
  40690=>"111110000",
  40691=>"000100111",
  40692=>"011010011",
  40693=>"000100100",
  40694=>"000011000",
  40695=>"000000000",
  40696=>"000000000",
  40697=>"111111111",
  40698=>"000000000",
  40699=>"000001111",
  40700=>"110110110",
  40701=>"000000000",
  40702=>"111110111",
  40703=>"100100000",
  40704=>"000000000",
  40705=>"001001000",
  40706=>"111111011",
  40707=>"011111111",
  40708=>"000000000",
  40709=>"111111111",
  40710=>"000000101",
  40711=>"011011000",
  40712=>"000000000",
  40713=>"000000000",
  40714=>"000100000",
  40715=>"001001111",
  40716=>"110100110",
  40717=>"110100000",
  40718=>"100100000",
  40719=>"011111000",
  40720=>"000100000",
  40721=>"000000001",
  40722=>"000000111",
  40723=>"000001011",
  40724=>"000000000",
  40725=>"000000010",
  40726=>"110110110",
  40727=>"001000000",
  40728=>"110111101",
  40729=>"110001000",
  40730=>"001101111",
  40731=>"001001000",
  40732=>"000000000",
  40733=>"000110111",
  40734=>"111111011",
  40735=>"010010000",
  40736=>"000000000",
  40737=>"000010111",
  40738=>"000000111",
  40739=>"011111111",
  40740=>"000000110",
  40741=>"001101001",
  40742=>"000000000",
  40743=>"000000001",
  40744=>"111111111",
  40745=>"011001001",
  40746=>"111111000",
  40747=>"111011000",
  40748=>"000001111",
  40749=>"000000100",
  40750=>"111110000",
  40751=>"011111111",
  40752=>"011011111",
  40753=>"001000000",
  40754=>"111111111",
  40755=>"011010000",
  40756=>"111101110",
  40757=>"111111111",
  40758=>"000001000",
  40759=>"000000001",
  40760=>"000010011",
  40761=>"010011111",
  40762=>"000010111",
  40763=>"000000111",
  40764=>"001001011",
  40765=>"111110111",
  40766=>"010111000",
  40767=>"111111111",
  40768=>"000000100",
  40769=>"000000000",
  40770=>"111101111",
  40771=>"000000100",
  40772=>"001100100",
  40773=>"111111111",
  40774=>"111111000",
  40775=>"111111111",
  40776=>"000111101",
  40777=>"010110001",
  40778=>"110000000",
  40779=>"011111111",
  40780=>"000000001",
  40781=>"000100110",
  40782=>"001011000",
  40783=>"110000000",
  40784=>"011011011",
  40785=>"000000111",
  40786=>"011111111",
  40787=>"111111111",
  40788=>"000100000",
  40789=>"001011001",
  40790=>"111011010",
  40791=>"111111111",
  40792=>"111111111",
  40793=>"010000000",
  40794=>"111010111",
  40795=>"111111100",
  40796=>"001100000",
  40797=>"000000101",
  40798=>"100101001",
  40799=>"111111111",
  40800=>"000000000",
  40801=>"000000000",
  40802=>"111111011",
  40803=>"001111111",
  40804=>"111111111",
  40805=>"000000000",
  40806=>"000000111",
  40807=>"000000110",
  40808=>"110110110",
  40809=>"000000000",
  40810=>"000111111",
  40811=>"100100000",
  40812=>"100111001",
  40813=>"000111111",
  40814=>"000000000",
  40815=>"000000001",
  40816=>"010111111",
  40817=>"011000111",
  40818=>"111111111",
  40819=>"111111111",
  40820=>"000000000",
  40821=>"101000100",
  40822=>"000000111",
  40823=>"111111011",
  40824=>"000000000",
  40825=>"100110011",
  40826=>"111111111",
  40827=>"100111111",
  40828=>"110111111",
  40829=>"000000111",
  40830=>"000000000",
  40831=>"000111111",
  40832=>"111111110",
  40833=>"111110110",
  40834=>"000000111",
  40835=>"110000010",
  40836=>"111111111",
  40837=>"111111000",
  40838=>"000000000",
  40839=>"111000000",
  40840=>"000000000",
  40841=>"111011001",
  40842=>"000000000",
  40843=>"000000000",
  40844=>"111001001",
  40845=>"111110100",
  40846=>"111100111",
  40847=>"000000001",
  40848=>"111111110",
  40849=>"001000100",
  40850=>"100000100",
  40851=>"000100100",
  40852=>"110010010",
  40853=>"000010000",
  40854=>"010010000",
  40855=>"000001001",
  40856=>"000001001",
  40857=>"011110111",
  40858=>"111111010",
  40859=>"101111101",
  40860=>"001111111",
  40861=>"111111111",
  40862=>"000000000",
  40863=>"111111111",
  40864=>"011100110",
  40865=>"001000000",
  40866=>"011111100",
  40867=>"000001000",
  40868=>"000000111",
  40869=>"000111011",
  40870=>"111111110",
  40871=>"101111111",
  40872=>"001001000",
  40873=>"111111001",
  40874=>"000000100",
  40875=>"000001001",
  40876=>"100000000",
  40877=>"110111000",
  40878=>"000100111",
  40879=>"010011111",
  40880=>"000010111",
  40881=>"000000000",
  40882=>"011001000",
  40883=>"000000000",
  40884=>"001000111",
  40885=>"110010111",
  40886=>"111111111",
  40887=>"000001111",
  40888=>"011011111",
  40889=>"111111111",
  40890=>"111111000",
  40891=>"001001111",
  40892=>"111111111",
  40893=>"000000000",
  40894=>"100100000",
  40895=>"000110100",
  40896=>"100000000",
  40897=>"100111110",
  40898=>"111111111",
  40899=>"011011010",
  40900=>"000001001",
  40901=>"010011011",
  40902=>"001000000",
  40903=>"000000000",
  40904=>"000100100",
  40905=>"000000000",
  40906=>"000000000",
  40907=>"111111111",
  40908=>"000011000",
  40909=>"111111111",
  40910=>"000000010",
  40911=>"000000000",
  40912=>"111111001",
  40913=>"111111111",
  40914=>"111111111",
  40915=>"111111111",
  40916=>"111111011",
  40917=>"111111111",
  40918=>"000000000",
  40919=>"000000000",
  40920=>"001101111",
  40921=>"110111101",
  40922=>"111111000",
  40923=>"001011000",
  40924=>"000101100",
  40925=>"111111000",
  40926=>"000011111",
  40927=>"111111111",
  40928=>"001000000",
  40929=>"111111111",
  40930=>"110000000",
  40931=>"111111111",
  40932=>"011111111",
  40933=>"111101111",
  40934=>"000000111",
  40935=>"000000000",
  40936=>"111111111",
  40937=>"111010011",
  40938=>"000000011",
  40939=>"001100100",
  40940=>"000000000",
  40941=>"001001001",
  40942=>"011011111",
  40943=>"001001001",
  40944=>"001101111",
  40945=>"111111111",
  40946=>"110000011",
  40947=>"000000000",
  40948=>"110000000",
  40949=>"111111111",
  40950=>"000000000",
  40951=>"000000100",
  40952=>"000000000",
  40953=>"111011001",
  40954=>"101101101",
  40955=>"111111100",
  40956=>"111111111",
  40957=>"100000000",
  40958=>"111111111",
  40959=>"000001000",
  40960=>"011110111",
  40961=>"111110000",
  40962=>"111111101",
  40963=>"111111000",
  40964=>"001011111",
  40965=>"111111100",
  40966=>"000000000",
  40967=>"111111111",
  40968=>"000000111",
  40969=>"111001000",
  40970=>"000010000",
  40971=>"000000000",
  40972=>"000001000",
  40973=>"010000000",
  40974=>"000101000",
  40975=>"000000100",
  40976=>"111111111",
  40977=>"100101111",
  40978=>"000111111",
  40979=>"111111111",
  40980=>"000000001",
  40981=>"111110111",
  40982=>"111000010",
  40983=>"000001111",
  40984=>"111110100",
  40985=>"000111110",
  40986=>"111101111",
  40987=>"000101111",
  40988=>"111111111",
  40989=>"101001000",
  40990=>"111111111",
  40991=>"110100000",
  40992=>"110110110",
  40993=>"111111111",
  40994=>"100000100",
  40995=>"000000000",
  40996=>"111111111",
  40997=>"001001000",
  40998=>"000000000",
  40999=>"111111101",
  41000=>"111111111",
  41001=>"010010011",
  41002=>"111101101",
  41003=>"010110000",
  41004=>"000000000",
  41005=>"000100111",
  41006=>"001000100",
  41007=>"011111111",
  41008=>"000000000",
  41009=>"000000100",
  41010=>"000001001",
  41011=>"011111111",
  41012=>"000000100",
  41013=>"001111111",
  41014=>"101101111",
  41015=>"111111111",
  41016=>"000000011",
  41017=>"110111011",
  41018=>"001000000",
  41019=>"000001111",
  41020=>"111111111",
  41021=>"101111111",
  41022=>"111101110",
  41023=>"111111111",
  41024=>"101110100",
  41025=>"111111111",
  41026=>"111000100",
  41027=>"101110111",
  41028=>"000000100",
  41029=>"111111011",
  41030=>"000000111",
  41031=>"000000000",
  41032=>"011011001",
  41033=>"000000001",
  41034=>"000000000",
  41035=>"111111001",
  41036=>"101000111",
  41037=>"000000111",
  41038=>"000001000",
  41039=>"111111111",
  41040=>"000000000",
  41041=>"000000001",
  41042=>"000000000",
  41043=>"000000000",
  41044=>"000101111",
  41045=>"100111111",
  41046=>"100000000",
  41047=>"001111111",
  41048=>"111111111",
  41049=>"101000000",
  41050=>"111111111",
  41051=>"010010000",
  41052=>"111111011",
  41053=>"000000100",
  41054=>"111111111",
  41055=>"110111111",
  41056=>"000000011",
  41057=>"001001001",
  41058=>"000000000",
  41059=>"110111100",
  41060=>"111111000",
  41061=>"000000111",
  41062=>"111111111",
  41063=>"000000000",
  41064=>"000000100",
  41065=>"111100000",
  41066=>"011111000",
  41067=>"000000001",
  41068=>"111111111",
  41069=>"111111111",
  41070=>"101100111",
  41071=>"000000110",
  41072=>"000000000",
  41073=>"000011000",
  41074=>"000100111",
  41075=>"111010000",
  41076=>"101111011",
  41077=>"110110000",
  41078=>"000000000",
  41079=>"000111111",
  41080=>"000000000",
  41081=>"011111011",
  41082=>"000000000",
  41083=>"000000000",
  41084=>"000000000",
  41085=>"111111111",
  41086=>"000000000",
  41087=>"000000000",
  41088=>"110000000",
  41089=>"000001111",
  41090=>"011111111",
  41091=>"000000000",
  41092=>"111111000",
  41093=>"111100111",
  41094=>"111111111",
  41095=>"000000000",
  41096=>"000000000",
  41097=>"000011010",
  41098=>"111100000",
  41099=>"111111011",
  41100=>"000000000",
  41101=>"000000000",
  41102=>"111111111",
  41103=>"000000000",
  41104=>"111101101",
  41105=>"000000101",
  41106=>"000111011",
  41107=>"010110110",
  41108=>"010010010",
  41109=>"111111111",
  41110=>"010000000",
  41111=>"000000000",
  41112=>"001001001",
  41113=>"000000000",
  41114=>"000000000",
  41115=>"111111111",
  41116=>"111110111",
  41117=>"000000111",
  41118=>"100000000",
  41119=>"000000000",
  41120=>"010010010",
  41121=>"000011011",
  41122=>"000000000",
  41123=>"000110010",
  41124=>"100000000",
  41125=>"000000000",
  41126=>"000111111",
  41127=>"000111000",
  41128=>"000110111",
  41129=>"000000000",
  41130=>"000000110",
  41131=>"000000100",
  41132=>"111110110",
  41133=>"101111111",
  41134=>"000000010",
  41135=>"011011101",
  41136=>"111001111",
  41137=>"000000000",
  41138=>"100101100",
  41139=>"000011100",
  41140=>"010010010",
  41141=>"101000110",
  41142=>"000001001",
  41143=>"011001110",
  41144=>"001001111",
  41145=>"011001111",
  41146=>"111100000",
  41147=>"100000111",
  41148=>"111111101",
  41149=>"111111100",
  41150=>"000100101",
  41151=>"000000100",
  41152=>"000000000",
  41153=>"000000000",
  41154=>"111111111",
  41155=>"110110111",
  41156=>"100111111",
  41157=>"011111111",
  41158=>"000010111",
  41159=>"000011111",
  41160=>"000000000",
  41161=>"000000000",
  41162=>"000000001",
  41163=>"000000000",
  41164=>"100101111",
  41165=>"000001000",
  41166=>"000000000",
  41167=>"001001111",
  41168=>"000000100",
  41169=>"111111110",
  41170=>"111111111",
  41171=>"000000000",
  41172=>"000000001",
  41173=>"000000000",
  41174=>"111111111",
  41175=>"011011110",
  41176=>"110110000",
  41177=>"111111111",
  41178=>"000000000",
  41179=>"111111111",
  41180=>"011001111",
  41181=>"111111011",
  41182=>"010111111",
  41183=>"000000001",
  41184=>"101001111",
  41185=>"110110011",
  41186=>"000000000",
  41187=>"111111111",
  41188=>"110111111",
  41189=>"110110110",
  41190=>"000000000",
  41191=>"111111111",
  41192=>"101101000",
  41193=>"011011000",
  41194=>"011011110",
  41195=>"111100111",
  41196=>"111001100",
  41197=>"100111111",
  41198=>"110111111",
  41199=>"011000000",
  41200=>"000000000",
  41201=>"000000000",
  41202=>"111110111",
  41203=>"000000000",
  41204=>"000001100",
  41205=>"010011111",
  41206=>"001011111",
  41207=>"111110010",
  41208=>"111111111",
  41209=>"000000010",
  41210=>"001011101",
  41211=>"000000000",
  41212=>"010011111",
  41213=>"010000000",
  41214=>"110000000",
  41215=>"010000100",
  41216=>"111111110",
  41217=>"111111100",
  41218=>"111101100",
  41219=>"111111111",
  41220=>"111000000",
  41221=>"000111111",
  41222=>"111111100",
  41223=>"011010110",
  41224=>"100101111",
  41225=>"111111000",
  41226=>"101111101",
  41227=>"000100110",
  41228=>"111111101",
  41229=>"001101111",
  41230=>"111111111",
  41231=>"000000000",
  41232=>"000000011",
  41233=>"011011111",
  41234=>"000000000",
  41235=>"100000001",
  41236=>"000000000",
  41237=>"000000000",
  41238=>"000111100",
  41239=>"000000100",
  41240=>"000000000",
  41241=>"111111010",
  41242=>"000000000",
  41243=>"010000111",
  41244=>"100111111",
  41245=>"111111111",
  41246=>"111111111",
  41247=>"000000000",
  41248=>"000000000",
  41249=>"000000000",
  41250=>"000000101",
  41251=>"000000000",
  41252=>"000000000",
  41253=>"000000000",
  41254=>"111101111",
  41255=>"100000000",
  41256=>"000000000",
  41257=>"001000000",
  41258=>"111111100",
  41259=>"111111111",
  41260=>"000000000",
  41261=>"110110110",
  41262=>"110100100",
  41263=>"111111110",
  41264=>"000110110",
  41265=>"011111111",
  41266=>"111101001",
  41267=>"000110110",
  41268=>"001001001",
  41269=>"100110111",
  41270=>"111011011",
  41271=>"000000111",
  41272=>"011111111",
  41273=>"001000000",
  41274=>"001000000",
  41275=>"111111101",
  41276=>"111111111",
  41277=>"001001000",
  41278=>"000100100",
  41279=>"011100100",
  41280=>"011000000",
  41281=>"011011000",
  41282=>"111011111",
  41283=>"100000001",
  41284=>"101000100",
  41285=>"111111111",
  41286=>"000000000",
  41287=>"110110110",
  41288=>"111111111",
  41289=>"000000100",
  41290=>"111111111",
  41291=>"110110110",
  41292=>"000000000",
  41293=>"000111111",
  41294=>"001000100",
  41295=>"110110110",
  41296=>"000000100",
  41297=>"000000000",
  41298=>"001001000",
  41299=>"001001000",
  41300=>"000000100",
  41301=>"011010000",
  41302=>"111000000",
  41303=>"001001001",
  41304=>"111111111",
  41305=>"111111111",
  41306=>"101001000",
  41307=>"000101100",
  41308=>"000000000",
  41309=>"111000100",
  41310=>"000001001",
  41311=>"000000001",
  41312=>"001000000",
  41313=>"000000000",
  41314=>"111111111",
  41315=>"111111111",
  41316=>"100100100",
  41317=>"001000000",
  41318=>"110111111",
  41319=>"001000001",
  41320=>"001001001",
  41321=>"010110110",
  41322=>"100101111",
  41323=>"111111111",
  41324=>"001001000",
  41325=>"000000000",
  41326=>"000000000",
  41327=>"000000000",
  41328=>"110111111",
  41329=>"000000000",
  41330=>"011011000",
  41331=>"111111111",
  41332=>"111110110",
  41333=>"111111000",
  41334=>"111111011",
  41335=>"010000000",
  41336=>"011111111",
  41337=>"111111111",
  41338=>"000011010",
  41339=>"110110110",
  41340=>"000000000",
  41341=>"000010111",
  41342=>"111011011",
  41343=>"111100100",
  41344=>"000000000",
  41345=>"000000010",
  41346=>"100100100",
  41347=>"111111111",
  41348=>"111111111",
  41349=>"000000000",
  41350=>"000000000",
  41351=>"000000000",
  41352=>"000000000",
  41353=>"111111001",
  41354=>"000000111",
  41355=>"111111111",
  41356=>"101101111",
  41357=>"000000010",
  41358=>"111111111",
  41359=>"000000000",
  41360=>"000010000",
  41361=>"111101100",
  41362=>"000000000",
  41363=>"011111110",
  41364=>"000000000",
  41365=>"000110000",
  41366=>"100001001",
  41367=>"000000000",
  41368=>"011011111",
  41369=>"110000011",
  41370=>"110110110",
  41371=>"111111111",
  41372=>"000100100",
  41373=>"111111111",
  41374=>"000000000",
  41375=>"000000111",
  41376=>"000010110",
  41377=>"111111000",
  41378=>"100100111",
  41379=>"110111111",
  41380=>"000000111",
  41381=>"000000000",
  41382=>"111111111",
  41383=>"000101111",
  41384=>"000000000",
  41385=>"111111110",
  41386=>"111111111",
  41387=>"111111111",
  41388=>"111111111",
  41389=>"110110000",
  41390=>"111110111",
  41391=>"110010010",
  41392=>"000000000",
  41393=>"000000100",
  41394=>"000000000",
  41395=>"000000110",
  41396=>"011001000",
  41397=>"111001111",
  41398=>"000100000",
  41399=>"100000000",
  41400=>"000000110",
  41401=>"111111111",
  41402=>"000000000",
  41403=>"000011000",
  41404=>"000000111",
  41405=>"111010111",
  41406=>"000000000",
  41407=>"000000000",
  41408=>"000111100",
  41409=>"000001111",
  41410=>"010111111",
  41411=>"000000000",
  41412=>"100100111",
  41413=>"111111011",
  41414=>"000010010",
  41415=>"111111111",
  41416=>"001111100",
  41417=>"000000000",
  41418=>"111111101",
  41419=>"000000111",
  41420=>"000101100",
  41421=>"000000000",
  41422=>"111101111",
  41423=>"000000000",
  41424=>"000000000",
  41425=>"111011011",
  41426=>"111111111",
  41427=>"111111111",
  41428=>"111111111",
  41429=>"111110000",
  41430=>"000000111",
  41431=>"110110001",
  41432=>"000001001",
  41433=>"000001001",
  41434=>"100110110",
  41435=>"111111111",
  41436=>"000001001",
  41437=>"111111111",
  41438=>"101111001",
  41439=>"111111111",
  41440=>"000100111",
  41441=>"111011100",
  41442=>"111110000",
  41443=>"111111111",
  41444=>"001011111",
  41445=>"000000000",
  41446=>"101000000",
  41447=>"110110000",
  41448=>"000000000",
  41449=>"000000000",
  41450=>"111111111",
  41451=>"100000000",
  41452=>"010010111",
  41453=>"001001011",
  41454=>"001110010",
  41455=>"111111111",
  41456=>"101000000",
  41457=>"000100111",
  41458=>"000000000",
  41459=>"000000000",
  41460=>"110111000",
  41461=>"000000110",
  41462=>"100000011",
  41463=>"000100100",
  41464=>"000111111",
  41465=>"100000000",
  41466=>"100110111",
  41467=>"001101111",
  41468=>"111111111",
  41469=>"111111111",
  41470=>"000001111",
  41471=>"111111111",
  41472=>"101101101",
  41473=>"000000000",
  41474=>"111101111",
  41475=>"000000000",
  41476=>"001001001",
  41477=>"111110000",
  41478=>"100100101",
  41479=>"111111111",
  41480=>"000000000",
  41481=>"000010000",
  41482=>"111111100",
  41483=>"111110000",
  41484=>"011011001",
  41485=>"101000000",
  41486=>"000000111",
  41487=>"001111111",
  41488=>"000000000",
  41489=>"010111111",
  41490=>"111111100",
  41491=>"000111011",
  41492=>"000000000",
  41493=>"111000000",
  41494=>"111111111",
  41495=>"000000001",
  41496=>"111111111",
  41497=>"011011000",
  41498=>"000000000",
  41499=>"001010000",
  41500=>"000000000",
  41501=>"000000111",
  41502=>"011101011",
  41503=>"000000001",
  41504=>"111111111",
  41505=>"111111000",
  41506=>"000010010",
  41507=>"000000100",
  41508=>"111111110",
  41509=>"000001000",
  41510=>"000000000",
  41511=>"111111101",
  41512=>"111111000",
  41513=>"111111110",
  41514=>"111111111",
  41515=>"100100000",
  41516=>"111111111",
  41517=>"111111111",
  41518=>"111100000",
  41519=>"011111001",
  41520=>"100111010",
  41521=>"011001001",
  41522=>"000011011",
  41523=>"000000000",
  41524=>"000110111",
  41525=>"010010011",
  41526=>"100100111",
  41527=>"111010000",
  41528=>"100000000",
  41529=>"000110110",
  41530=>"111111111",
  41531=>"011111111",
  41532=>"000010010",
  41533=>"000111110",
  41534=>"011111010",
  41535=>"011000001",
  41536=>"111000001",
  41537=>"000000000",
  41538=>"110111000",
  41539=>"001101111",
  41540=>"111001001",
  41541=>"111011011",
  41542=>"111000110",
  41543=>"111111000",
  41544=>"111110100",
  41545=>"000000000",
  41546=>"110100001",
  41547=>"000101000",
  41548=>"000101000",
  41549=>"111001000",
  41550=>"000000111",
  41551=>"000000000",
  41552=>"110100000",
  41553=>"111011011",
  41554=>"110000000",
  41555=>"001001001",
  41556=>"111111111",
  41557=>"000000110",
  41558=>"111000000",
  41559=>"010000000",
  41560=>"111111110",
  41561=>"110111111",
  41562=>"111101000",
  41563=>"110100000",
  41564=>"000111111",
  41565=>"000110110",
  41566=>"001000001",
  41567=>"111111111",
  41568=>"110110000",
  41569=>"000010010",
  41570=>"000000111",
  41571=>"000010000",
  41572=>"111111101",
  41573=>"000000000",
  41574=>"111000111",
  41575=>"111100000",
  41576=>"111111110",
  41577=>"111100000",
  41578=>"000000100",
  41579=>"000111111",
  41580=>"000011011",
  41581=>"111111111",
  41582=>"001000001",
  41583=>"000000001",
  41584=>"110110110",
  41585=>"000000011",
  41586=>"001000000",
  41587=>"000111111",
  41588=>"000000000",
  41589=>"000111111",
  41590=>"111111001",
  41591=>"000101101",
  41592=>"000000101",
  41593=>"111111111",
  41594=>"000000000",
  41595=>"110000000",
  41596=>"111111011",
  41597=>"000000000",
  41598=>"000000000",
  41599=>"000111111",
  41600=>"000000111",
  41601=>"111111111",
  41602=>"111000011",
  41603=>"111110000",
  41604=>"110000000",
  41605=>"101000001",
  41606=>"011001001",
  41607=>"111111000",
  41608=>"111001111",
  41609=>"000000000",
  41610=>"000011000",
  41611=>"111000000",
  41612=>"000000000",
  41613=>"111110110",
  41614=>"000000000",
  41615=>"100111111",
  41616=>"000000000",
  41617=>"111111111",
  41618=>"000000001",
  41619=>"100111111",
  41620=>"000000001",
  41621=>"111000001",
  41622=>"111000100",
  41623=>"000000000",
  41624=>"000000111",
  41625=>"111111111",
  41626=>"000000000",
  41627=>"000111011",
  41628=>"101101111",
  41629=>"000111111",
  41630=>"100100001",
  41631=>"000000000",
  41632=>"111001111",
  41633=>"000000110",
  41634=>"000001111",
  41635=>"100111111",
  41636=>"000000101",
  41637=>"101001111",
  41638=>"001111111",
  41639=>"111011001",
  41640=>"000000000",
  41641=>"000000111",
  41642=>"000011111",
  41643=>"110000000",
  41644=>"001111111",
  41645=>"000000000",
  41646=>"111111010",
  41647=>"001000100",
  41648=>"000000101",
  41649=>"110111111",
  41650=>"011111011",
  41651=>"111111111",
  41652=>"111111011",
  41653=>"111111000",
  41654=>"111111110",
  41655=>"111111111",
  41656=>"000000000",
  41657=>"101111111",
  41658=>"001001101",
  41659=>"001001000",
  41660=>"110110111",
  41661=>"111111100",
  41662=>"111111111",
  41663=>"000000000",
  41664=>"000000000",
  41665=>"000000000",
  41666=>"000111111",
  41667=>"000000011",
  41668=>"000011111",
  41669=>"001001000",
  41670=>"000000000",
  41671=>"100000000",
  41672=>"111111111",
  41673=>"010000000",
  41674=>"010000000",
  41675=>"111101101",
  41676=>"011000101",
  41677=>"100110110",
  41678=>"111111011",
  41679=>"111011000",
  41680=>"111111100",
  41681=>"011111111",
  41682=>"000010111",
  41683=>"000000011",
  41684=>"000000111",
  41685=>"100000000",
  41686=>"111000111",
  41687=>"000000000",
  41688=>"110111111",
  41689=>"001011011",
  41690=>"111000000",
  41691=>"000000100",
  41692=>"110011011",
  41693=>"111110100",
  41694=>"000000000",
  41695=>"101100111",
  41696=>"000000001",
  41697=>"001111111",
  41698=>"000000000",
  41699=>"111101101",
  41700=>"100101101",
  41701=>"101111110",
  41702=>"001011110",
  41703=>"111111111",
  41704=>"101101111",
  41705=>"001111111",
  41706=>"111111110",
  41707=>"100000000",
  41708=>"000000100",
  41709=>"000000000",
  41710=>"011011110",
  41711=>"011101100",
  41712=>"110000000",
  41713=>"111111000",
  41714=>"000111111",
  41715=>"001000111",
  41716=>"000000001",
  41717=>"111110111",
  41718=>"110010111",
  41719=>"011110111",
  41720=>"111111111",
  41721=>"000000000",
  41722=>"000111000",
  41723=>"000101111",
  41724=>"111000000",
  41725=>"000010010",
  41726=>"111000000",
  41727=>"111111111",
  41728=>"000111011",
  41729=>"001011011",
  41730=>"011110110",
  41731=>"000000001",
  41732=>"111110111",
  41733=>"000011111",
  41734=>"111110111",
  41735=>"111111001",
  41736=>"100000000",
  41737=>"111111010",
  41738=>"000000000",
  41739=>"000000000",
  41740=>"110110111",
  41741=>"111101111",
  41742=>"001110111",
  41743=>"111111000",
  41744=>"111000110",
  41745=>"101000100",
  41746=>"000000001",
  41747=>"000110111",
  41748=>"000000000",
  41749=>"111111111",
  41750=>"000010111",
  41751=>"100111011",
  41752=>"000001010",
  41753=>"111111111",
  41754=>"100000101",
  41755=>"111111111",
  41756=>"010011001",
  41757=>"011111111",
  41758=>"000000101",
  41759=>"111111111",
  41760=>"111110100",
  41761=>"000000000",
  41762=>"111111000",
  41763=>"101001111",
  41764=>"111111111",
  41765=>"000000011",
  41766=>"111100100",
  41767=>"100110100",
  41768=>"000000111",
  41769=>"100100111",
  41770=>"011111110",
  41771=>"000000000",
  41772=>"000000000",
  41773=>"001111111",
  41774=>"100110111",
  41775=>"000000100",
  41776=>"110111000",
  41777=>"000000111",
  41778=>"000000000",
  41779=>"000000000",
  41780=>"111110000",
  41781=>"100100110",
  41782=>"000000001",
  41783=>"111111111",
  41784=>"100000000",
  41785=>"001000111",
  41786=>"000000000",
  41787=>"000111001",
  41788=>"000001111",
  41789=>"001000110",
  41790=>"000111111",
  41791=>"001001000",
  41792=>"001011001",
  41793=>"000000000",
  41794=>"111111111",
  41795=>"000000111",
  41796=>"110000000",
  41797=>"000000010",
  41798=>"111111101",
  41799=>"111101000",
  41800=>"000000000",
  41801=>"111111110",
  41802=>"111111000",
  41803=>"000010110",
  41804=>"110110111",
  41805=>"110111111",
  41806=>"000000000",
  41807=>"000000111",
  41808=>"100100101",
  41809=>"101101111",
  41810=>"111111111",
  41811=>"100100111",
  41812=>"111010000",
  41813=>"011111001",
  41814=>"111111111",
  41815=>"000000111",
  41816=>"111011011",
  41817=>"000111000",
  41818=>"111111000",
  41819=>"110111111",
  41820=>"000101000",
  41821=>"111111111",
  41822=>"000000001",
  41823=>"011011000",
  41824=>"101101111",
  41825=>"000000111",
  41826=>"110000000",
  41827=>"001011100",
  41828=>"111111111",
  41829=>"111001111",
  41830=>"100000111",
  41831=>"000100110",
  41832=>"000000011",
  41833=>"110100100",
  41834=>"111111110",
  41835=>"011010110",
  41836=>"011111111",
  41837=>"000011101",
  41838=>"000110110",
  41839=>"000011011",
  41840=>"110000000",
  41841=>"111111110",
  41842=>"010000000",
  41843=>"001110000",
  41844=>"100100111",
  41845=>"000000000",
  41846=>"011011011",
  41847=>"000000000",
  41848=>"111111111",
  41849=>"000001000",
  41850=>"110000101",
  41851=>"101111000",
  41852=>"000001100",
  41853=>"000000000",
  41854=>"001001000",
  41855=>"000101111",
  41856=>"000100110",
  41857=>"111111100",
  41858=>"001000110",
  41859=>"000000000",
  41860=>"111111001",
  41861=>"000000100",
  41862=>"000110111",
  41863=>"111111000",
  41864=>"000000000",
  41865=>"000100111",
  41866=>"100000110",
  41867=>"111000000",
  41868=>"011110001",
  41869=>"000010010",
  41870=>"111111000",
  41871=>"000000011",
  41872=>"000000000",
  41873=>"110010000",
  41874=>"110110111",
  41875=>"000000110",
  41876=>"111111111",
  41877=>"111101000",
  41878=>"000000000",
  41879=>"111111000",
  41880=>"111111000",
  41881=>"111011110",
  41882=>"000101111",
  41883=>"000110110",
  41884=>"100000000",
  41885=>"000000000",
  41886=>"000000101",
  41887=>"000000000",
  41888=>"111101111",
  41889=>"110111111",
  41890=>"000110000",
  41891=>"111001000",
  41892=>"000000111",
  41893=>"110000000",
  41894=>"111110110",
  41895=>"111111111",
  41896=>"010000000",
  41897=>"000000110",
  41898=>"000001000",
  41899=>"011011000",
  41900=>"000000000",
  41901=>"111000111",
  41902=>"111011010",
  41903=>"111001000",
  41904=>"000001111",
  41905=>"111111101",
  41906=>"000000111",
  41907=>"000111111",
  41908=>"111111110",
  41909=>"110100111",
  41910=>"011111111",
  41911=>"000000000",
  41912=>"110010000",
  41913=>"001111111",
  41914=>"111101101",
  41915=>"111100000",
  41916=>"001001000",
  41917=>"010110000",
  41918=>"101101111",
  41919=>"010010011",
  41920=>"100100111",
  41921=>"100000000",
  41922=>"111001111",
  41923=>"000000000",
  41924=>"111000000",
  41925=>"001000110",
  41926=>"000000000",
  41927=>"000000000",
  41928=>"101100100",
  41929=>"101111000",
  41930=>"000000100",
  41931=>"000000000",
  41932=>"111111100",
  41933=>"001000111",
  41934=>"111100100",
  41935=>"111001000",
  41936=>"000000011",
  41937=>"000000100",
  41938=>"000110010",
  41939=>"010010000",
  41940=>"000000000",
  41941=>"111000111",
  41942=>"000000000",
  41943=>"110110011",
  41944=>"111000111",
  41945=>"111111111",
  41946=>"111111000",
  41947=>"111000000",
  41948=>"010111010",
  41949=>"001000000",
  41950=>"011011011",
  41951=>"001111111",
  41952=>"111111111",
  41953=>"111000000",
  41954=>"000100111",
  41955=>"101111111",
  41956=>"111010010",
  41957=>"000000000",
  41958=>"000000100",
  41959=>"111100111",
  41960=>"110110010",
  41961=>"001000100",
  41962=>"111110000",
  41963=>"000000111",
  41964=>"000000111",
  41965=>"111100000",
  41966=>"111111111",
  41967=>"000110110",
  41968=>"000101101",
  41969=>"000000000",
  41970=>"101001011",
  41971=>"011101000",
  41972=>"000110000",
  41973=>"000000111",
  41974=>"010000100",
  41975=>"011111111",
  41976=>"000000000",
  41977=>"100000000",
  41978=>"010000000",
  41979=>"111111001",
  41980=>"000000111",
  41981=>"111111111",
  41982=>"110100101",
  41983=>"000000000",
  41984=>"001001001",
  41985=>"110110111",
  41986=>"000000001",
  41987=>"000000000",
  41988=>"000100101",
  41989=>"001000000",
  41990=>"101000000",
  41991=>"111111111",
  41992=>"010000000",
  41993=>"111111000",
  41994=>"000111111",
  41995=>"000111111",
  41996=>"011000000",
  41997=>"100110111",
  41998=>"001000101",
  41999=>"100000000",
  42000=>"000111111",
  42001=>"000000001",
  42002=>"000000000",
  42003=>"000000000",
  42004=>"011001111",
  42005=>"000111111",
  42006=>"110111111",
  42007=>"110111000",
  42008=>"001001000",
  42009=>"101101011",
  42010=>"001111111",
  42011=>"110000000",
  42012=>"001011111",
  42013=>"010010111",
  42014=>"000000010",
  42015=>"110111111",
  42016=>"110111111",
  42017=>"011111000",
  42018=>"001000101",
  42019=>"111000101",
  42020=>"000000100",
  42021=>"011111111",
  42022=>"010000000",
  42023=>"000000111",
  42024=>"111100110",
  42025=>"000000000",
  42026=>"111100000",
  42027=>"111000000",
  42028=>"111111111",
  42029=>"111111111",
  42030=>"000000110",
  42031=>"001000000",
  42032=>"111111110",
  42033=>"111111011",
  42034=>"000100100",
  42035=>"101101101",
  42036=>"000110110",
  42037=>"100111110",
  42038=>"000000000",
  42039=>"111101001",
  42040=>"111111000",
  42041=>"000000000",
  42042=>"000000000",
  42043=>"111111111",
  42044=>"100000000",
  42045=>"000111111",
  42046=>"000111111",
  42047=>"000000000",
  42048=>"010011000",
  42049=>"000000000",
  42050=>"111111111",
  42051=>"011111111",
  42052=>"110110100",
  42053=>"001011011",
  42054=>"000000000",
  42055=>"111111111",
  42056=>"110110111",
  42057=>"111000000",
  42058=>"000000000",
  42059=>"111111111",
  42060=>"000000000",
  42061=>"111111010",
  42062=>"111000000",
  42063=>"000000001",
  42064=>"000000000",
  42065=>"111000011",
  42066=>"000000000",
  42067=>"001000000",
  42068=>"000000000",
  42069=>"000010110",
  42070=>"011000100",
  42071=>"110111110",
  42072=>"111100001",
  42073=>"111111101",
  42074=>"101000000",
  42075=>"100001100",
  42076=>"001000000",
  42077=>"110111111",
  42078=>"101100111",
  42079=>"010011111",
  42080=>"110111010",
  42081=>"000000111",
  42082=>"000000000",
  42083=>"000000111",
  42084=>"111100110",
  42085=>"000000111",
  42086=>"111111000",
  42087=>"111100000",
  42088=>"000111010",
  42089=>"111101111",
  42090=>"000000111",
  42091=>"111111111",
  42092=>"100100100",
  42093=>"000000000",
  42094=>"000111011",
  42095=>"000000010",
  42096=>"111111000",
  42097=>"010010111",
  42098=>"111001000",
  42099=>"100111111",
  42100=>"000001111",
  42101=>"000000001",
  42102=>"010000000",
  42103=>"001000000",
  42104=>"010111011",
  42105=>"110111111",
  42106=>"111000000",
  42107=>"011000000",
  42108=>"100110110",
  42109=>"111111111",
  42110=>"000001000",
  42111=>"011000000",
  42112=>"111111111",
  42113=>"011011111",
  42114=>"111111100",
  42115=>"000000000",
  42116=>"000000000",
  42117=>"001000000",
  42118=>"000000110",
  42119=>"000000001",
  42120=>"111100000",
  42121=>"000000000",
  42122=>"000000001",
  42123=>"000000100",
  42124=>"110000000",
  42125=>"000000000",
  42126=>"111111110",
  42127=>"000000000",
  42128=>"000000000",
  42129=>"110111000",
  42130=>"000010111",
  42131=>"111001001",
  42132=>"001111111",
  42133=>"000000001",
  42134=>"001000000",
  42135=>"111000000",
  42136=>"111000000",
  42137=>"111000000",
  42138=>"000000000",
  42139=>"000011011",
  42140=>"111100100",
  42141=>"000000000",
  42142=>"111111110",
  42143=>"111011111",
  42144=>"111111110",
  42145=>"111111111",
  42146=>"111011000",
  42147=>"000000000",
  42148=>"111011000",
  42149=>"111111111",
  42150=>"111111010",
  42151=>"000011000",
  42152=>"101111111",
  42153=>"111111111",
  42154=>"100100111",
  42155=>"000000000",
  42156=>"100000000",
  42157=>"011111100",
  42158=>"100100000",
  42159=>"111111111",
  42160=>"111111000",
  42161=>"111111111",
  42162=>"110111111",
  42163=>"111111111",
  42164=>"100111111",
  42165=>"111101000",
  42166=>"110111011",
  42167=>"000000011",
  42168=>"001001111",
  42169=>"000000000",
  42170=>"001000111",
  42171=>"110011111",
  42172=>"000000111",
  42173=>"001111110",
  42174=>"111111111",
  42175=>"010000000",
  42176=>"111111101",
  42177=>"000001101",
  42178=>"000000000",
  42179=>"011000000",
  42180=>"000000100",
  42181=>"101101000",
  42182=>"111101001",
  42183=>"111111001",
  42184=>"000110111",
  42185=>"000000011",
  42186=>"001100100",
  42187=>"000010111",
  42188=>"000000001",
  42189=>"111111111",
  42190=>"000000110",
  42191=>"101011111",
  42192=>"000111110",
  42193=>"000000000",
  42194=>"000000010",
  42195=>"111001000",
  42196=>"000010111",
  42197=>"001000000",
  42198=>"100000000",
  42199=>"111111111",
  42200=>"001000000",
  42201=>"110110100",
  42202=>"000000000",
  42203=>"111011111",
  42204=>"110111111",
  42205=>"000000000",
  42206=>"000000010",
  42207=>"100000000",
  42208=>"001101111",
  42209=>"100110111",
  42210=>"001000111",
  42211=>"000000000",
  42212=>"110111111",
  42213=>"010111111",
  42214=>"111111111",
  42215=>"000100111",
  42216=>"111111111",
  42217=>"100000000",
  42218=>"000000111",
  42219=>"111000000",
  42220=>"000110111",
  42221=>"010000000",
  42222=>"111010000",
  42223=>"111101000",
  42224=>"110000000",
  42225=>"111111000",
  42226=>"000000000",
  42227=>"010000000",
  42228=>"111110111",
  42229=>"000110110",
  42230=>"001000001",
  42231=>"000000000",
  42232=>"000000011",
  42233=>"000000000",
  42234=>"100000000",
  42235=>"011111101",
  42236=>"111100100",
  42237=>"111111111",
  42238=>"000000100",
  42239=>"000000100",
  42240=>"001000001",
  42241=>"001101111",
  42242=>"000000000",
  42243=>"000000000",
  42244=>"000000111",
  42245=>"110110100",
  42246=>"000000000",
  42247=>"011000000",
  42248=>"011010000",
  42249=>"000000001",
  42250=>"111111111",
  42251=>"001000000",
  42252=>"111111111",
  42253=>"000110000",
  42254=>"000000000",
  42255=>"100111111",
  42256=>"000000001",
  42257=>"111000000",
  42258=>"000000000",
  42259=>"111111001",
  42260=>"000000000",
  42261=>"100000000",
  42262=>"100100110",
  42263=>"000000111",
  42264=>"110110111",
  42265=>"111111111",
  42266=>"100110111",
  42267=>"111111111",
  42268=>"111111111",
  42269=>"000000000",
  42270=>"111111111",
  42271=>"000000001",
  42272=>"011000000",
  42273=>"001000000",
  42274=>"110000000",
  42275=>"111101111",
  42276=>"000000101",
  42277=>"111111111",
  42278=>"111000000",
  42279=>"010000111",
  42280=>"110100011",
  42281=>"000100111",
  42282=>"111110101",
  42283=>"000100110",
  42284=>"010010110",
  42285=>"110111110",
  42286=>"101011000",
  42287=>"111111111",
  42288=>"000000000",
  42289=>"000000000",
  42290=>"110000000",
  42291=>"000000110",
  42292=>"110110110",
  42293=>"111111100",
  42294=>"001000000",
  42295=>"000000001",
  42296=>"000010001",
  42297=>"111111111",
  42298=>"000000000",
  42299=>"111111011",
  42300=>"110111011",
  42301=>"111010110",
  42302=>"000000011",
  42303=>"111000000",
  42304=>"001000000",
  42305=>"000100000",
  42306=>"111011001",
  42307=>"001000000",
  42308=>"111111010",
  42309=>"111001010",
  42310=>"000000000",
  42311=>"000000000",
  42312=>"111110110",
  42313=>"111000000",
  42314=>"111111111",
  42315=>"000011111",
  42316=>"111111110",
  42317=>"000000000",
  42318=>"110111111",
  42319=>"100000100",
  42320=>"111001000",
  42321=>"000000000",
  42322=>"000000000",
  42323=>"000000001",
  42324=>"001000000",
  42325=>"001001001",
  42326=>"111110110",
  42327=>"111110110",
  42328=>"111001001",
  42329=>"111111111",
  42330=>"111111010",
  42331=>"000000101",
  42332=>"000110100",
  42333=>"000000000",
  42334=>"000000110",
  42335=>"110111111",
  42336=>"111000000",
  42337=>"111111111",
  42338=>"000000000",
  42339=>"111111101",
  42340=>"000100000",
  42341=>"111000000",
  42342=>"101001001",
  42343=>"000000000",
  42344=>"100110110",
  42345=>"111000000",
  42346=>"111111111",
  42347=>"000000011",
  42348=>"111111110",
  42349=>"111100110",
  42350=>"111111111",
  42351=>"111000000",
  42352=>"000000110",
  42353=>"000010000",
  42354=>"000000011",
  42355=>"001001011",
  42356=>"111111000",
  42357=>"110111101",
  42358=>"111111000",
  42359=>"000110100",
  42360=>"111111111",
  42361=>"010000111",
  42362=>"111111111",
  42363=>"100000011",
  42364=>"000101111",
  42365=>"000111010",
  42366=>"111000000",
  42367=>"011001000",
  42368=>"101101111",
  42369=>"111111111",
  42370=>"110110010",
  42371=>"000111011",
  42372=>"111111101",
  42373=>"000000000",
  42374=>"000101111",
  42375=>"111111110",
  42376=>"101000000",
  42377=>"000111111",
  42378=>"111111111",
  42379=>"000111111",
  42380=>"110010111",
  42381=>"111111111",
  42382=>"000000111",
  42383=>"011001011",
  42384=>"000010010",
  42385=>"110111110",
  42386=>"111000000",
  42387=>"011111110",
  42388=>"000110000",
  42389=>"000000000",
  42390=>"000101111",
  42391=>"000110110",
  42392=>"000000000",
  42393=>"111100110",
  42394=>"111001111",
  42395=>"000001001",
  42396=>"111111111",
  42397=>"111111111",
  42398=>"000000010",
  42399=>"000000000",
  42400=>"111111100",
  42401=>"011111111",
  42402=>"111011111",
  42403=>"001001000",
  42404=>"111001101",
  42405=>"011011000",
  42406=>"000000000",
  42407=>"010010000",
  42408=>"111111010",
  42409=>"111000000",
  42410=>"111111111",
  42411=>"110000000",
  42412=>"000000000",
  42413=>"111011111",
  42414=>"100110111",
  42415=>"000000001",
  42416=>"000000000",
  42417=>"000000000",
  42418=>"000000111",
  42419=>"111111111",
  42420=>"011010000",
  42421=>"111000001",
  42422=>"110111111",
  42423=>"000110100",
  42424=>"111111111",
  42425=>"111111111",
  42426=>"111110111",
  42427=>"101000110",
  42428=>"010011000",
  42429=>"111111111",
  42430=>"000000111",
  42431=>"000111111",
  42432=>"000000100",
  42433=>"000000000",
  42434=>"111111001",
  42435=>"000110111",
  42436=>"111111111",
  42437=>"111100100",
  42438=>"000000000",
  42439=>"000001101",
  42440=>"111100100",
  42441=>"000000000",
  42442=>"011000000",
  42443=>"011010000",
  42444=>"111000000",
  42445=>"100111111",
  42446=>"111000001",
  42447=>"000000000",
  42448=>"000000010",
  42449=>"000000110",
  42450=>"100000000",
  42451=>"111111000",
  42452=>"011111011",
  42453=>"110100100",
  42454=>"000000111",
  42455=>"111011000",
  42456=>"001000100",
  42457=>"111110000",
  42458=>"010010011",
  42459=>"110100000",
  42460=>"000000000",
  42461=>"111000000",
  42462=>"100100000",
  42463=>"111111001",
  42464=>"111001111",
  42465=>"000000000",
  42466=>"000110000",
  42467=>"001000101",
  42468=>"111100100",
  42469=>"000000000",
  42470=>"000010111",
  42471=>"000000000",
  42472=>"111111110",
  42473=>"110000000",
  42474=>"111110010",
  42475=>"001011000",
  42476=>"000000111",
  42477=>"001001001",
  42478=>"010111111",
  42479=>"000010111",
  42480=>"000000011",
  42481=>"000010000",
  42482=>"111111111",
  42483=>"000000010",
  42484=>"111111111",
  42485=>"010000111",
  42486=>"111111111",
  42487=>"000000000",
  42488=>"111111111",
  42489=>"100000011",
  42490=>"000000000",
  42491=>"111001001",
  42492=>"011111001",
  42493=>"000000111",
  42494=>"000000000",
  42495=>"111000001",
  42496=>"100111111",
  42497=>"111111111",
  42498=>"111111111",
  42499=>"011011011",
  42500=>"110111001",
  42501=>"000101111",
  42502=>"000000000",
  42503=>"000000000",
  42504=>"011000000",
  42505=>"110000000",
  42506=>"111111011",
  42507=>"110000001",
  42508=>"110000000",
  42509=>"111001000",
  42510=>"000100100",
  42511=>"111111100",
  42512=>"000000000",
  42513=>"111111111",
  42514=>"000000000",
  42515=>"100000000",
  42516=>"111000000",
  42517=>"111111111",
  42518=>"000000001",
  42519=>"111111111",
  42520=>"000000000",
  42521=>"111111101",
  42522=>"000000000",
  42523=>"100110111",
  42524=>"111111111",
  42525=>"000000100",
  42526=>"111110110",
  42527=>"100000000",
  42528=>"111011000",
  42529=>"100000000",
  42530=>"000001111",
  42531=>"111111101",
  42532=>"111000001",
  42533=>"000000000",
  42534=>"111111111",
  42535=>"000111111",
  42536=>"101111000",
  42537=>"100100110",
  42538=>"001011111",
  42539=>"011111110",
  42540=>"111111101",
  42541=>"111111111",
  42542=>"010001001",
  42543=>"111010010",
  42544=>"100110111",
  42545=>"000000000",
  42546=>"011000100",
  42547=>"000000000",
  42548=>"001001101",
  42549=>"111100000",
  42550=>"111111110",
  42551=>"000000000",
  42552=>"111111111",
  42553=>"000001000",
  42554=>"000000000",
  42555=>"000000111",
  42556=>"111000000",
  42557=>"000111011",
  42558=>"111110110",
  42559=>"100000100",
  42560=>"001001000",
  42561=>"000000010",
  42562=>"111111111",
  42563=>"010000000",
  42564=>"111111111",
  42565=>"000000000",
  42566=>"100110111",
  42567=>"011111000",
  42568=>"000000000",
  42569=>"111111111",
  42570=>"000000000",
  42571=>"101111111",
  42572=>"000000000",
  42573=>"000000000",
  42574=>"000000111",
  42575=>"000000000",
  42576=>"001011111",
  42577=>"000000000",
  42578=>"111010111",
  42579=>"111111111",
  42580=>"110110110",
  42581=>"111111111",
  42582=>"011000101",
  42583=>"000001001",
  42584=>"001101000",
  42585=>"001111111",
  42586=>"000000001",
  42587=>"110110111",
  42588=>"001001000",
  42589=>"111101001",
  42590=>"011111111",
  42591=>"111011000",
  42592=>"011011001",
  42593=>"000000000",
  42594=>"001000000",
  42595=>"000000000",
  42596=>"000000000",
  42597=>"000000000",
  42598=>"000000000",
  42599=>"000000000",
  42600=>"111111111",
  42601=>"000000111",
  42602=>"110010000",
  42603=>"111010001",
  42604=>"000111111",
  42605=>"111101000",
  42606=>"111111111",
  42607=>"000010010",
  42608=>"000000001",
  42609=>"111111111",
  42610=>"111111001",
  42611=>"000000001",
  42612=>"100101000",
  42613=>"000000100",
  42614=>"000000000",
  42615=>"000000000",
  42616=>"001000010",
  42617=>"001001111",
  42618=>"000100100",
  42619=>"111111111",
  42620=>"100100100",
  42621=>"000010000",
  42622=>"001000000",
  42623=>"110000111",
  42624=>"010111110",
  42625=>"000000111",
  42626=>"111000000",
  42627=>"000100000",
  42628=>"000011111",
  42629=>"111000000",
  42630=>"001001000",
  42631=>"101111100",
  42632=>"111111000",
  42633=>"000000000",
  42634=>"011111111",
  42635=>"111111111",
  42636=>"000000100",
  42637=>"111111111",
  42638=>"111111000",
  42639=>"000000000",
  42640=>"111111111",
  42641=>"111100100",
  42642=>"110000000",
  42643=>"100100110",
  42644=>"100000000",
  42645=>"000000100",
  42646=>"000111111",
  42647=>"100111111",
  42648=>"110010001",
  42649=>"111111111",
  42650=>"011001000",
  42651=>"000000000",
  42652=>"100111111",
  42653=>"000000001",
  42654=>"000001000",
  42655=>"111111111",
  42656=>"111111000",
  42657=>"111011001",
  42658=>"000000111",
  42659=>"000000000",
  42660=>"011111111",
  42661=>"100101111",
  42662=>"000000110",
  42663=>"111000001",
  42664=>"100000000",
  42665=>"111111111",
  42666=>"111111111",
  42667=>"111111111",
  42668=>"001111001",
  42669=>"111111110",
  42670=>"000000110",
  42671=>"001001111",
  42672=>"000000000",
  42673=>"111111010",
  42674=>"111111000",
  42675=>"111111011",
  42676=>"111111111",
  42677=>"101101111",
  42678=>"001001000",
  42679=>"000000000",
  42680=>"000000100",
  42681=>"000100111",
  42682=>"111111111",
  42683=>"000000000",
  42684=>"000101100",
  42685=>"100110000",
  42686=>"011111100",
  42687=>"111111101",
  42688=>"000011000",
  42689=>"110011110",
  42690=>"011001001",
  42691=>"010111111",
  42692=>"001000101",
  42693=>"000000111",
  42694=>"111111000",
  42695=>"001111111",
  42696=>"000011011",
  42697=>"011001000",
  42698=>"111100000",
  42699=>"000000000",
  42700=>"111101000",
  42701=>"111111111",
  42702=>"000000000",
  42703=>"111001000",
  42704=>"111111111",
  42705=>"000000000",
  42706=>"100110111",
  42707=>"111111011",
  42708=>"111111111",
  42709=>"010000100",
  42710=>"000000000",
  42711=>"110010010",
  42712=>"111110101",
  42713=>"110110000",
  42714=>"111011000",
  42715=>"110110110",
  42716=>"111111111",
  42717=>"011011000",
  42718=>"111001000",
  42719=>"111111110",
  42720=>"111111111",
  42721=>"000000000",
  42722=>"000000000",
  42723=>"000000000",
  42724=>"010011000",
  42725=>"111111000",
  42726=>"000000001",
  42727=>"111111001",
  42728=>"111111011",
  42729=>"101000000",
  42730=>"111110110",
  42731=>"001001111",
  42732=>"111111111",
  42733=>"111110110",
  42734=>"111111001",
  42735=>"000000000",
  42736=>"111111011",
  42737=>"001000001",
  42738=>"111111111",
  42739=>"000110000",
  42740=>"100110111",
  42741=>"111011000",
  42742=>"011001001",
  42743=>"111111111",
  42744=>"111011000",
  42745=>"111111000",
  42746=>"110111100",
  42747=>"000000000",
  42748=>"111111111",
  42749=>"100001011",
  42750=>"111111000",
  42751=>"111111111",
  42752=>"000000000",
  42753=>"000000000",
  42754=>"000000000",
  42755=>"111111000",
  42756=>"000001000",
  42757=>"000000000",
  42758=>"000000000",
  42759=>"100110111",
  42760=>"111111000",
  42761=>"001000000",
  42762=>"111111111",
  42763=>"110111111",
  42764=>"101000111",
  42765=>"111111111",
  42766=>"111111111",
  42767=>"000000000",
  42768=>"100100100",
  42769=>"000000011",
  42770=>"100110000",
  42771=>"100001001",
  42772=>"011000001",
  42773=>"111010011",
  42774=>"000000000",
  42775=>"001001011",
  42776=>"111111110",
  42777=>"000000000",
  42778=>"111111111",
  42779=>"000000011",
  42780=>"011001000",
  42781=>"111111111",
  42782=>"000000000",
  42783=>"000000100",
  42784=>"000111111",
  42785=>"111001000",
  42786=>"111111111",
  42787=>"100000000",
  42788=>"111000000",
  42789=>"000000000",
  42790=>"000000000",
  42791=>"111111110",
  42792=>"111101111",
  42793=>"001000100",
  42794=>"000001000",
  42795=>"000000000",
  42796=>"111111111",
  42797=>"101000000",
  42798=>"000010000",
  42799=>"000000000",
  42800=>"111110000",
  42801=>"110110000",
  42802=>"111111111",
  42803=>"000000000",
  42804=>"111111010",
  42805=>"111000000",
  42806=>"100111111",
  42807=>"111111111",
  42808=>"110000000",
  42809=>"111111111",
  42810=>"111111111",
  42811=>"100100100",
  42812=>"111111111",
  42813=>"000000000",
  42814=>"000000001",
  42815=>"111000000",
  42816=>"000000000",
  42817=>"000000000",
  42818=>"000001000",
  42819=>"111111111",
  42820=>"000000000",
  42821=>"000111111",
  42822=>"101010110",
  42823=>"110011000",
  42824=>"011111111",
  42825=>"111000000",
  42826=>"000001101",
  42827=>"111111111",
  42828=>"000000000",
  42829=>"000000000",
  42830=>"110100000",
  42831=>"000010000",
  42832=>"000000000",
  42833=>"111011001",
  42834=>"000000010",
  42835=>"000000000",
  42836=>"000100000",
  42837=>"011011011",
  42838=>"111111000",
  42839=>"000000000",
  42840=>"001111111",
  42841=>"101101111",
  42842=>"000110100",
  42843=>"111111000",
  42844=>"010000000",
  42845=>"001101111",
  42846=>"111111111",
  42847=>"110101101",
  42848=>"000000000",
  42849=>"111111111",
  42850=>"111111111",
  42851=>"111111111",
  42852=>"000000000",
  42853=>"000100111",
  42854=>"100100111",
  42855=>"111011011",
  42856=>"000000000",
  42857=>"000000000",
  42858=>"001000111",
  42859=>"000000000",
  42860=>"100100100",
  42861=>"111111110",
  42862=>"111111111",
  42863=>"000000000",
  42864=>"000000000",
  42865=>"000011000",
  42866=>"001111111",
  42867=>"100110010",
  42868=>"011001000",
  42869=>"000000000",
  42870=>"000000000",
  42871=>"111111111",
  42872=>"000000111",
  42873=>"000000000",
  42874=>"111001000",
  42875=>"100111111",
  42876=>"111000100",
  42877=>"001000000",
  42878=>"100101111",
  42879=>"111111111",
  42880=>"100111111",
  42881=>"001111111",
  42882=>"000000000",
  42883=>"111101101",
  42884=>"000000000",
  42885=>"111111111",
  42886=>"100000000",
  42887=>"111111111",
  42888=>"000000000",
  42889=>"011001000",
  42890=>"110000000",
  42891=>"000000010",
  42892=>"111111111",
  42893=>"000110000",
  42894=>"000000000",
  42895=>"111111001",
  42896=>"111000000",
  42897=>"000001001",
  42898=>"100000000",
  42899=>"001111111",
  42900=>"111111111",
  42901=>"000000000",
  42902=>"111000101",
  42903=>"000100000",
  42904=>"111111111",
  42905=>"111110000",
  42906=>"000000001",
  42907=>"000000111",
  42908=>"111111111",
  42909=>"111111111",
  42910=>"000000111",
  42911=>"101111111",
  42912=>"000111111",
  42913=>"111011000",
  42914=>"000001101",
  42915=>"000000000",
  42916=>"000000000",
  42917=>"111111111",
  42918=>"011000000",
  42919=>"010111111",
  42920=>"011011111",
  42921=>"111111111",
  42922=>"000000100",
  42923=>"111101110",
  42924=>"000000000",
  42925=>"011000111",
  42926=>"000000000",
  42927=>"001100000",
  42928=>"111000000",
  42929=>"000000111",
  42930=>"000111111",
  42931=>"000000000",
  42932=>"000001001",
  42933=>"011111111",
  42934=>"000000001",
  42935=>"000000001",
  42936=>"000000000",
  42937=>"011111101",
  42938=>"111111111",
  42939=>"111111001",
  42940=>"011000011",
  42941=>"111111111",
  42942=>"000000100",
  42943=>"110110110",
  42944=>"111110110",
  42945=>"000000001",
  42946=>"000001000",
  42947=>"000000000",
  42948=>"111111111",
  42949=>"100100110",
  42950=>"101000110",
  42951=>"100101111",
  42952=>"110110000",
  42953=>"111111111",
  42954=>"111011001",
  42955=>"111111111",
  42956=>"111111111",
  42957=>"111111111",
  42958=>"001000000",
  42959=>"000110111",
  42960=>"000000000",
  42961=>"000001011",
  42962=>"000000000",
  42963=>"001000001",
  42964=>"100100100",
  42965=>"111111001",
  42966=>"111110010",
  42967=>"100000000",
  42968=>"000000000",
  42969=>"000000000",
  42970=>"001000000",
  42971=>"000000000",
  42972=>"000000000",
  42973=>"000000000",
  42974=>"111111000",
  42975=>"001001001",
  42976=>"100000000",
  42977=>"000001001",
  42978=>"100110111",
  42979=>"000110111",
  42980=>"110000000",
  42981=>"100100110",
  42982=>"111011000",
  42983=>"000000010",
  42984=>"000000001",
  42985=>"000000110",
  42986=>"000000000",
  42987=>"001001000",
  42988=>"000000000",
  42989=>"111011001",
  42990=>"010000000",
  42991=>"000000000",
  42992=>"001111111",
  42993=>"111000000",
  42994=>"100111111",
  42995=>"000000000",
  42996=>"110100000",
  42997=>"111110110",
  42998=>"110110010",
  42999=>"111001000",
  43000=>"111111111",
  43001=>"111111111",
  43002=>"101000000",
  43003=>"111110111",
  43004=>"000000000",
  43005=>"011011000",
  43006=>"111111000",
  43007=>"111111111",
  43008=>"000000110",
  43009=>"010011000",
  43010=>"000000000",
  43011=>"000000000",
  43012=>"010111100",
  43013=>"110100000",
  43014=>"100100000",
  43015=>"000000000",
  43016=>"000000001",
  43017=>"111111111",
  43018=>"000010000",
  43019=>"000000000",
  43020=>"011010111",
  43021=>"001010000",
  43022=>"001000000",
  43023=>"000000000",
  43024=>"000000000",
  43025=>"000011111",
  43026=>"001100100",
  43027=>"111111000",
  43028=>"111111111",
  43029=>"000000111",
  43030=>"111111111",
  43031=>"010110000",
  43032=>"111111010",
  43033=>"011001110",
  43034=>"001001000",
  43035=>"000000110",
  43036=>"000000111",
  43037=>"100100000",
  43038=>"111111110",
  43039=>"000000011",
  43040=>"000000000",
  43041=>"111111111",
  43042=>"110000000",
  43043=>"100100111",
  43044=>"111111111",
  43045=>"001101101",
  43046=>"100100000",
  43047=>"001000000",
  43048=>"100101101",
  43049=>"000000000",
  43050=>"000000000",
  43051=>"011000101",
  43052=>"111111011",
  43053=>"111000000",
  43054=>"000000110",
  43055=>"000000000",
  43056=>"000101100",
  43057=>"111000000",
  43058=>"111111111",
  43059=>"111111111",
  43060=>"000000001",
  43061=>"111111011",
  43062=>"011011111",
  43063=>"000111111",
  43064=>"011110110",
  43065=>"111000000",
  43066=>"000000000",
  43067=>"000000000",
  43068=>"111101101",
  43069=>"111111111",
  43070=>"000010100",
  43071=>"000000111",
  43072=>"100100000",
  43073=>"111001000",
  43074=>"110000000",
  43075=>"000111000",
  43076=>"000000000",
  43077=>"111111000",
  43078=>"000000000",
  43079=>"100111111",
  43080=>"111111111",
  43081=>"000000101",
  43082=>"111111010",
  43083=>"000000000",
  43084=>"111000000",
  43085=>"000100011",
  43086=>"011111110",
  43087=>"000000000",
  43088=>"110000000",
  43089=>"000100111",
  43090=>"111111111",
  43091=>"101100100",
  43092=>"111000000",
  43093=>"011000000",
  43094=>"101001000",
  43095=>"111111111",
  43096=>"000000000",
  43097=>"000000000",
  43098=>"011111111",
  43099=>"111100111",
  43100=>"001001000",
  43101=>"000000000",
  43102=>"000110011",
  43103=>"000111111",
  43104=>"000000000",
  43105=>"110110110",
  43106=>"000000000",
  43107=>"111111110",
  43108=>"101101100",
  43109=>"000110010",
  43110=>"110110110",
  43111=>"111111000",
  43112=>"001011000",
  43113=>"000000011",
  43114=>"000000000",
  43115=>"000111111",
  43116=>"000000000",
  43117=>"000000000",
  43118=>"111111000",
  43119=>"111100000",
  43120=>"110111111",
  43121=>"111110100",
  43122=>"011110000",
  43123=>"000000000",
  43124=>"110101101",
  43125=>"011111111",
  43126=>"000000100",
  43127=>"000000100",
  43128=>"000111000",
  43129=>"000000000",
  43130=>"101100101",
  43131=>"000000000",
  43132=>"111111111",
  43133=>"001100100",
  43134=>"111111111",
  43135=>"010010000",
  43136=>"000000000",
  43137=>"111111111",
  43138=>"001111111",
  43139=>"111000000",
  43140=>"000010000",
  43141=>"000000000",
  43142=>"000000000",
  43143=>"000000000",
  43144=>"111111111",
  43145=>"111111111",
  43146=>"000000000",
  43147=>"011111111",
  43148=>"111110000",
  43149=>"010001000",
  43150=>"001001001",
  43151=>"000011111",
  43152=>"000000000",
  43153=>"111111110",
  43154=>"000010111",
  43155=>"111111111",
  43156=>"000000000",
  43157=>"000000001",
  43158=>"000010111",
  43159=>"111111001",
  43160=>"111111000",
  43161=>"111111111",
  43162=>"000000000",
  43163=>"110111111",
  43164=>"110111011",
  43165=>"010110100",
  43166=>"000000000",
  43167=>"111111000",
  43168=>"000000000",
  43169=>"000110110",
  43170=>"110111111",
  43171=>"000111111",
  43172=>"001111101",
  43173=>"111110010",
  43174=>"010111111",
  43175=>"010111111",
  43176=>"011011100",
  43177=>"111111111",
  43178=>"111111000",
  43179=>"110111111",
  43180=>"000000111",
  43181=>"010110110",
  43182=>"110111111",
  43183=>"011011111",
  43184=>"000010111",
  43185=>"100101101",
  43186=>"011011111",
  43187=>"000000000",
  43188=>"000000000",
  43189=>"000000000",
  43190=>"000000000",
  43191=>"111111111",
  43192=>"110111111",
  43193=>"000000000",
  43194=>"111111111",
  43195=>"000001001",
  43196=>"000000000",
  43197=>"111111111",
  43198=>"111111111",
  43199=>"000000111",
  43200=>"111111111",
  43201=>"010000111",
  43202=>"111110100",
  43203=>"111000000",
  43204=>"000000000",
  43205=>"000000011",
  43206=>"000000000",
  43207=>"111111110",
  43208=>"000100100",
  43209=>"111100110",
  43210=>"000000111",
  43211=>"000100100",
  43212=>"000000000",
  43213=>"111000000",
  43214=>"000000111",
  43215=>"011000000",
  43216=>"000000000",
  43217=>"010110110",
  43218=>"111100000",
  43219=>"011111111",
  43220=>"000010110",
  43221=>"000000000",
  43222=>"111111010",
  43223=>"000000000",
  43224=>"111111111",
  43225=>"111110111",
  43226=>"000000111",
  43227=>"111111111",
  43228=>"111111111",
  43229=>"111111111",
  43230=>"010010010",
  43231=>"000000000",
  43232=>"000011111",
  43233=>"111100000",
  43234=>"000000000",
  43235=>"000111101",
  43236=>"010001000",
  43237=>"000001011",
  43238=>"111011011",
  43239=>"110010000",
  43240=>"000000000",
  43241=>"111111111",
  43242=>"000001011",
  43243=>"111111111",
  43244=>"111011111",
  43245=>"000000000",
  43246=>"011011000",
  43247=>"001011110",
  43248=>"011001000",
  43249=>"001101001",
  43250=>"111001001",
  43251=>"000000000",
  43252=>"000000000",
  43253=>"001100101",
  43254=>"001011111",
  43255=>"100000000",
  43256=>"000000000",
  43257=>"000000001",
  43258=>"111001111",
  43259=>"000000000",
  43260=>"110110011",
  43261=>"001001100",
  43262=>"000000000",
  43263=>"111111111",
  43264=>"111111000",
  43265=>"110110011",
  43266=>"101000110",
  43267=>"000000111",
  43268=>"001001001",
  43269=>"111111000",
  43270=>"001000001",
  43271=>"111111000",
  43272=>"000000000",
  43273=>"111101101",
  43274=>"111111100",
  43275=>"000000111",
  43276=>"111001001",
  43277=>"100111111",
  43278=>"011001110",
  43279=>"000110000",
  43280=>"111111110",
  43281=>"111111111",
  43282=>"111111110",
  43283=>"111111111",
  43284=>"111111111",
  43285=>"100000000",
  43286=>"011101000",
  43287=>"000000000",
  43288=>"111111111",
  43289=>"101101111",
  43290=>"111111010",
  43291=>"000000000",
  43292=>"000001000",
  43293=>"000000101",
  43294=>"011111111",
  43295=>"011000000",
  43296=>"011011111",
  43297=>"000111110",
  43298=>"110110000",
  43299=>"000000000",
  43300=>"100100110",
  43301=>"001000000",
  43302=>"000111111",
  43303=>"111000010",
  43304=>"111111111",
  43305=>"011000000",
  43306=>"000110100",
  43307=>"000000111",
  43308=>"000000000",
  43309=>"001000000",
  43310=>"000000000",
  43311=>"001001001",
  43312=>"111111010",
  43313=>"001001000",
  43314=>"010000000",
  43315=>"111111110",
  43316=>"001111111",
  43317=>"100100000",
  43318=>"111111000",
  43319=>"001011111",
  43320=>"000010010",
  43321=>"001001001",
  43322=>"000101111",
  43323=>"100000000",
  43324=>"100000000",
  43325=>"111111011",
  43326=>"000000001",
  43327=>"000110000",
  43328=>"111011000",
  43329=>"111111111",
  43330=>"000000000",
  43331=>"111111111",
  43332=>"010100110",
  43333=>"111111111",
  43334=>"111000000",
  43335=>"000000000",
  43336=>"000100000",
  43337=>"111111100",
  43338=>"111111111",
  43339=>"110110000",
  43340=>"000111110",
  43341=>"000111111",
  43342=>"000000001",
  43343=>"111111111",
  43344=>"000011011",
  43345=>"010111111",
  43346=>"110111111",
  43347=>"111101000",
  43348=>"000000000",
  43349=>"000000011",
  43350=>"111111111",
  43351=>"011000000",
  43352=>"000000000",
  43353=>"111111111",
  43354=>"000000000",
  43355=>"111111000",
  43356=>"111000000",
  43357=>"000000000",
  43358=>"000000100",
  43359=>"000000000",
  43360=>"000000110",
  43361=>"111111111",
  43362=>"111111011",
  43363=>"100000000",
  43364=>"111110110",
  43365=>"000010010",
  43366=>"111110010",
  43367=>"011000000",
  43368=>"011000000",
  43369=>"111111111",
  43370=>"111111010",
  43371=>"000000000",
  43372=>"110100100",
  43373=>"000111011",
  43374=>"110000000",
  43375=>"000000111",
  43376=>"011111111",
  43377=>"000111111",
  43378=>"011111111",
  43379=>"100100100",
  43380=>"000000000",
  43381=>"110110000",
  43382=>"000011111",
  43383=>"110110111",
  43384=>"000000111",
  43385=>"000000000",
  43386=>"010000000",
  43387=>"010011111",
  43388=>"000000100",
  43389=>"000000000",
  43390=>"110111111",
  43391=>"100000000",
  43392=>"001011011",
  43393=>"001001011",
  43394=>"110111000",
  43395=>"010111000",
  43396=>"000000000",
  43397=>"000100101",
  43398=>"101100111",
  43399=>"000000000",
  43400=>"111110000",
  43401=>"000100111",
  43402=>"000000000",
  43403=>"000011111",
  43404=>"111111011",
  43405=>"111111111",
  43406=>"110111011",
  43407=>"000000000",
  43408=>"111111010",
  43409=>"111111111",
  43410=>"111111111",
  43411=>"111010111",
  43412=>"000111111",
  43413=>"010000000",
  43414=>"000000111",
  43415=>"111111100",
  43416=>"011000000",
  43417=>"110100110",
  43418=>"000000001",
  43419=>"101111111",
  43420=>"000100100",
  43421=>"111111110",
  43422=>"000000000",
  43423=>"111000000",
  43424=>"111111111",
  43425=>"011111111",
  43426=>"000000001",
  43427=>"111111111",
  43428=>"111111011",
  43429=>"000001000",
  43430=>"000101000",
  43431=>"000100010",
  43432=>"001001000",
  43433=>"000000000",
  43434=>"000011111",
  43435=>"000000000",
  43436=>"100111111",
  43437=>"000011001",
  43438=>"101101101",
  43439=>"000001111",
  43440=>"000110000",
  43441=>"111001000",
  43442=>"000000000",
  43443=>"111111011",
  43444=>"011111111",
  43445=>"111000101",
  43446=>"111111111",
  43447=>"001111001",
  43448=>"111111100",
  43449=>"000010111",
  43450=>"000000100",
  43451=>"000000111",
  43452=>"000000000",
  43453=>"111011101",
  43454=>"000000000",
  43455=>"011011011",
  43456=>"000011011",
  43457=>"101000000",
  43458=>"111111111",
  43459=>"111111111",
  43460=>"011001111",
  43461=>"100001011",
  43462=>"110100000",
  43463=>"101000010",
  43464=>"101000000",
  43465=>"100000111",
  43466=>"001100111",
  43467=>"101001011",
  43468=>"111000000",
  43469=>"010111111",
  43470=>"000000000",
  43471=>"000111111",
  43472=>"111111000",
  43473=>"100110111",
  43474=>"111001000",
  43475=>"000000000",
  43476=>"000000001",
  43477=>"000000001",
  43478=>"011000000",
  43479=>"111111001",
  43480=>"000000000",
  43481=>"111000000",
  43482=>"000000100",
  43483=>"000111111",
  43484=>"111111110",
  43485=>"000000100",
  43486=>"101101000",
  43487=>"110010000",
  43488=>"001101111",
  43489=>"000000000",
  43490=>"111111000",
  43491=>"101100111",
  43492=>"100111111",
  43493=>"000000000",
  43494=>"000000001",
  43495=>"100101111",
  43496=>"111111111",
  43497=>"111011000",
  43498=>"111000000",
  43499=>"000000010",
  43500=>"011011000",
  43501=>"000011011",
  43502=>"000000111",
  43503=>"000000000",
  43504=>"000000101",
  43505=>"000111111",
  43506=>"000000101",
  43507=>"000000000",
  43508=>"111111111",
  43509=>"000000000",
  43510=>"111111010",
  43511=>"100110110",
  43512=>"111101101",
  43513=>"001111111",
  43514=>"011011111",
  43515=>"111000000",
  43516=>"000001111",
  43517=>"000000000",
  43518=>"000000000",
  43519=>"000000101",
  43520=>"111110001",
  43521=>"111111010",
  43522=>"110010000",
  43523=>"000000001",
  43524=>"110110000",
  43525=>"000000000",
  43526=>"001000000",
  43527=>"000000001",
  43528=>"000100100",
  43529=>"111111110",
  43530=>"000000010",
  43531=>"101011011",
  43532=>"001001001",
  43533=>"010110110",
  43534=>"000000000",
  43535=>"101001001",
  43536=>"110110111",
  43537=>"010000010",
  43538=>"111100001",
  43539=>"000000101",
  43540=>"100111000",
  43541=>"111111101",
  43542=>"111011011",
  43543=>"100110100",
  43544=>"001001001",
  43545=>"100001001",
  43546=>"111101101",
  43547=>"011011000",
  43548=>"001001011",
  43549=>"111111101",
  43550=>"001100000",
  43551=>"110110010",
  43552=>"101001001",
  43553=>"101101100",
  43554=>"110110101",
  43555=>"111011011",
  43556=>"111111111",
  43557=>"111011000",
  43558=>"010000010",
  43559=>"001000100",
  43560=>"111110111",
  43561=>"000000000",
  43562=>"101000001",
  43563=>"000000001",
  43564=>"110111111",
  43565=>"000000000",
  43566=>"101111101",
  43567=>"110001101",
  43568=>"101001000",
  43569=>"111001111",
  43570=>"110100101",
  43571=>"000000000",
  43572=>"101100101",
  43573=>"101101101",
  43574=>"000000000",
  43575=>"110000101",
  43576=>"100111111",
  43577=>"110110010",
  43578=>"100000000",
  43579=>"000000111",
  43580=>"101101100",
  43581=>"010111000",
  43582=>"000001001",
  43583=>"101000010",
  43584=>"010010110",
  43585=>"000110010",
  43586=>"111011000",
  43587=>"010111010",
  43588=>"101001001",
  43589=>"001001100",
  43590=>"111010010",
  43591=>"010111111",
  43592=>"100100100",
  43593=>"110010000",
  43594=>"000000000",
  43595=>"001001001",
  43596=>"111111111",
  43597=>"110110000",
  43598=>"001000000",
  43599=>"000000011",
  43600=>"111101000",
  43601=>"000001001",
  43602=>"101111001",
  43603=>"100100000",
  43604=>"001001000",
  43605=>"110110110",
  43606=>"111010000",
  43607=>"101101101",
  43608=>"000100111",
  43609=>"111111111",
  43610=>"000000010",
  43611=>"110100100",
  43612=>"110110000",
  43613=>"111111111",
  43614=>"110110010",
  43615=>"111111001",
  43616=>"010000000",
  43617=>"110010010",
  43618=>"010011010",
  43619=>"000111101",
  43620=>"110110001",
  43621=>"001101101",
  43622=>"000000000",
  43623=>"110110111",
  43624=>"000011001",
  43625=>"111111111",
  43626=>"010010111",
  43627=>"011010000",
  43628=>"000000000",
  43629=>"000100101",
  43630=>"111111111",
  43631=>"111001000",
  43632=>"111010000",
  43633=>"010010111",
  43634=>"000100100",
  43635=>"100000010",
  43636=>"100100100",
  43637=>"110110110",
  43638=>"111111111",
  43639=>"011000000",
  43640=>"011001111",
  43641=>"111111111",
  43642=>"010010111",
  43643=>"000111101",
  43644=>"100100000",
  43645=>"111100100",
  43646=>"000000000",
  43647=>"000000000",
  43648=>"101101101",
  43649=>"111101101",
  43650=>"000010111",
  43651=>"001001001",
  43652=>"011110110",
  43653=>"000101111",
  43654=>"100000000",
  43655=>"000110111",
  43656=>"000110010",
  43657=>"111101001",
  43658=>"000111111",
  43659=>"101101101",
  43660=>"000001100",
  43661=>"110000000",
  43662=>"000010010",
  43663=>"111110111",
  43664=>"111101100",
  43665=>"101000000",
  43666=>"000000000",
  43667=>"000000000",
  43668=>"010110110",
  43669=>"111100000",
  43670=>"001001000",
  43671=>"000111111",
  43672=>"000101111",
  43673=>"101101111",
  43674=>"011000001",
  43675=>"000000000",
  43676=>"000000001",
  43677=>"111111000",
  43678=>"101101111",
  43679=>"101111111",
  43680=>"100111111",
  43681=>"000000110",
  43682=>"000000000",
  43683=>"011111110",
  43684=>"010110110",
  43685=>"110110110",
  43686=>"000001001",
  43687=>"100000100",
  43688=>"000000111",
  43689=>"000010110",
  43690=>"111011011",
  43691=>"001000000",
  43692=>"110111111",
  43693=>"000010110",
  43694=>"000000101",
  43695=>"000001000",
  43696=>"010111001",
  43697=>"001011100",
  43698=>"011111111",
  43699=>"011111001",
  43700=>"101111110",
  43701=>"101101101",
  43702=>"101100110",
  43703=>"000110010",
  43704=>"000101111",
  43705=>"100111111",
  43706=>"111001111",
  43707=>"000110110",
  43708=>"011000011",
  43709=>"011111111",
  43710=>"000000000",
  43711=>"111111111",
  43712=>"000000000",
  43713=>"000000011",
  43714=>"011111000",
  43715=>"010110110",
  43716=>"101101001",
  43717=>"010010010",
  43718=>"000000011",
  43719=>"000000000",
  43720=>"011111110",
  43721=>"111111111",
  43722=>"000001100",
  43723=>"000000100",
  43724=>"110111111",
  43725=>"111100100",
  43726=>"000000000",
  43727=>"111001111",
  43728=>"000000000",
  43729=>"001011000",
  43730=>"110010010",
  43731=>"101101101",
  43732=>"111101101",
  43733=>"001110110",
  43734=>"111111000",
  43735=>"001001001",
  43736=>"000000100",
  43737=>"000100110",
  43738=>"000101000",
  43739=>"000001000",
  43740=>"110111111",
  43741=>"111110010",
  43742=>"110110110",
  43743=>"110111010",
  43744=>"000000000",
  43745=>"011111111",
  43746=>"111111000",
  43747=>"110111111",
  43748=>"110110000",
  43749=>"011011011",
  43750=>"111011111",
  43751=>"000011111",
  43752=>"010110111",
  43753=>"111111011",
  43754=>"000000011",
  43755=>"111110010",
  43756=>"001001000",
  43757=>"001000000",
  43758=>"010010110",
  43759=>"011111000",
  43760=>"000111111",
  43761=>"000001001",
  43762=>"110111001",
  43763=>"000000000",
  43764=>"101101111",
  43765=>"111111110",
  43766=>"000011010",
  43767=>"010010010",
  43768=>"000011111",
  43769=>"011011000",
  43770=>"000110000",
  43771=>"000000001",
  43772=>"111111111",
  43773=>"001001000",
  43774=>"010000000",
  43775=>"111110111",
  43776=>"000101111",
  43777=>"101001100",
  43778=>"000000001",
  43779=>"110111111",
  43780=>"001000011",
  43781=>"001000000",
  43782=>"111111111",
  43783=>"011111001",
  43784=>"000000000",
  43785=>"000000000",
  43786=>"000110110",
  43787=>"111111111",
  43788=>"000101101",
  43789=>"001000000",
  43790=>"111111011",
  43791=>"101000000",
  43792=>"000000000",
  43793=>"111100000",
  43794=>"101101000",
  43795=>"100000010",
  43796=>"001000000",
  43797=>"010010010",
  43798=>"100100100",
  43799=>"101101111",
  43800=>"110110111",
  43801=>"000010110",
  43802=>"100000110",
  43803=>"111000000",
  43804=>"000011011",
  43805=>"010011111",
  43806=>"101111111",
  43807=>"010111110",
  43808=>"111100100",
  43809=>"000000000",
  43810=>"111111111",
  43811=>"110110110",
  43812=>"111111111",
  43813=>"111110110",
  43814=>"000000000",
  43815=>"111111111",
  43816=>"111111111",
  43817=>"000001100",
  43818=>"000000000",
  43819=>"101001000",
  43820=>"111011001",
  43821=>"000000000",
  43822=>"011000000",
  43823=>"000000000",
  43824=>"100111101",
  43825=>"110000000",
  43826=>"111111110",
  43827=>"110111110",
  43828=>"110110010",
  43829=>"101111101",
  43830=>"000101111",
  43831=>"111111001",
  43832=>"011111111",
  43833=>"010010111",
  43834=>"011001111",
  43835=>"000000111",
  43836=>"011000010",
  43837=>"000010000",
  43838=>"000000000",
  43839=>"000000110",
  43840=>"101101000",
  43841=>"000000110",
  43842=>"111110100",
  43843=>"001000000",
  43844=>"111011000",
  43845=>"000000000",
  43846=>"111101111",
  43847=>"111100111",
  43848=>"010011011",
  43849=>"010010000",
  43850=>"110111010",
  43851=>"001001011",
  43852=>"000011100",
  43853=>"010111111",
  43854=>"111111010",
  43855=>"011001001",
  43856=>"001001001",
  43857=>"110110010",
  43858=>"110110111",
  43859=>"110110111",
  43860=>"111111111",
  43861=>"001001001",
  43862=>"110110110",
  43863=>"000101000",
  43864=>"111111111",
  43865=>"111111011",
  43866=>"111111100",
  43867=>"101111101",
  43868=>"001111111",
  43869=>"101101111",
  43870=>"100000000",
  43871=>"110110110",
  43872=>"111011000",
  43873=>"000000101",
  43874=>"110011000",
  43875=>"111110000",
  43876=>"001001101",
  43877=>"111111111",
  43878=>"000000000",
  43879=>"001111111",
  43880=>"100110110",
  43881=>"000100000",
  43882=>"001000001",
  43883=>"001000000",
  43884=>"010010000",
  43885=>"010010011",
  43886=>"101100100",
  43887=>"000000000",
  43888=>"111111010",
  43889=>"011011011",
  43890=>"111110110",
  43891=>"100101101",
  43892=>"010110110",
  43893=>"101101111",
  43894=>"011111111",
  43895=>"100100110",
  43896=>"101101101",
  43897=>"010110111",
  43898=>"010110000",
  43899=>"100101001",
  43900=>"010111111",
  43901=>"010010110",
  43902=>"000001111",
  43903=>"000000000",
  43904=>"100100110",
  43905=>"000110110",
  43906=>"100000011",
  43907=>"001001011",
  43908=>"111111000",
  43909=>"111110000",
  43910=>"000111111",
  43911=>"111111110",
  43912=>"100000000",
  43913=>"000000010",
  43914=>"010110000",
  43915=>"110010000",
  43916=>"000010010",
  43917=>"001001000",
  43918=>"111111100",
  43919=>"010010000",
  43920=>"010000000",
  43921=>"100111111",
  43922=>"110110101",
  43923=>"110110110",
  43924=>"111111111",
  43925=>"010010000",
  43926=>"000000000",
  43927=>"100100100",
  43928=>"111111011",
  43929=>"010110111",
  43930=>"001001000",
  43931=>"001000010",
  43932=>"100101101",
  43933=>"000000000",
  43934=>"001001111",
  43935=>"111111000",
  43936=>"110000000",
  43937=>"011000000",
  43938=>"000001111",
  43939=>"110111000",
  43940=>"000000000",
  43941=>"010010000",
  43942=>"000000000",
  43943=>"011010110",
  43944=>"010010000",
  43945=>"110110111",
  43946=>"000001111",
  43947=>"101001000",
  43948=>"000000000",
  43949=>"110110010",
  43950=>"010011111",
  43951=>"001001001",
  43952=>"000110111",
  43953=>"111101111",
  43954=>"011001000",
  43955=>"001000000",
  43956=>"111111110",
  43957=>"110110111",
  43958=>"100111111",
  43959=>"111110111",
  43960=>"111111100",
  43961=>"000000000",
  43962=>"000010111",
  43963=>"100100100",
  43964=>"011011111",
  43965=>"100001101",
  43966=>"100000000",
  43967=>"110000110",
  43968=>"110110000",
  43969=>"111111111",
  43970=>"001001000",
  43971=>"111111000",
  43972=>"000000000",
  43973=>"000111101",
  43974=>"010111111",
  43975=>"001101001",
  43976=>"000100111",
  43977=>"111111111",
  43978=>"000000000",
  43979=>"110100000",
  43980=>"111111000",
  43981=>"000111111",
  43982=>"101000000",
  43983=>"111111011",
  43984=>"000000000",
  43985=>"000100011",
  43986=>"110010010",
  43987=>"001001011",
  43988=>"000000000",
  43989=>"110000000",
  43990=>"000111111",
  43991=>"110110110",
  43992=>"010111111",
  43993=>"101101001",
  43994=>"111011000",
  43995=>"000000000",
  43996=>"001011011",
  43997=>"011101000",
  43998=>"111111000",
  43999=>"110100110",
  44000=>"101101100",
  44001=>"101001111",
  44002=>"111111111",
  44003=>"100111111",
  44004=>"000000000",
  44005=>"000001111",
  44006=>"101101101",
  44007=>"000000111",
  44008=>"000000100",
  44009=>"001001001",
  44010=>"011111111",
  44011=>"000010000",
  44012=>"011011010",
  44013=>"001011011",
  44014=>"100100000",
  44015=>"010000000",
  44016=>"001001101",
  44017=>"111111001",
  44018=>"111110110",
  44019=>"000100100",
  44020=>"000000010",
  44021=>"100100111",
  44022=>"000000100",
  44023=>"100100000",
  44024=>"000000000",
  44025=>"001101111",
  44026=>"000110111",
  44027=>"101101000",
  44028=>"011001000",
  44029=>"110110010",
  44030=>"100100001",
  44031=>"101101111",
  44032=>"111010111",
  44033=>"111111000",
  44034=>"111111111",
  44035=>"100111111",
  44036=>"111000000",
  44037=>"101110111",
  44038=>"000000000",
  44039=>"000000000",
  44040=>"000000111",
  44041=>"011111101",
  44042=>"100100100",
  44043=>"011001000",
  44044=>"101000100",
  44045=>"110111001",
  44046=>"111111111",
  44047=>"000000110",
  44048=>"111111100",
  44049=>"110111111",
  44050=>"000000000",
  44051=>"000000000",
  44052=>"110110111",
  44053=>"000000000",
  44054=>"000000100",
  44055=>"011111110",
  44056=>"001001001",
  44057=>"100000001",
  44058=>"111001000",
  44059=>"000011111",
  44060=>"111101110",
  44061=>"000000000",
  44062=>"111111111",
  44063=>"111110111",
  44064=>"011111111",
  44065=>"111101000",
  44066=>"101111111",
  44067=>"000001000",
  44068=>"000001001",
  44069=>"100100111",
  44070=>"000000000",
  44071=>"011011011",
  44072=>"111111111",
  44073=>"000000000",
  44074=>"111111111",
  44075=>"000000000",
  44076=>"000000000",
  44077=>"110100100",
  44078=>"100000000",
  44079=>"111111111",
  44080=>"011111111",
  44081=>"000011000",
  44082=>"000110100",
  44083=>"011011011",
  44084=>"000000000",
  44085=>"110010010",
  44086=>"110110000",
  44087=>"000000001",
  44088=>"011000000",
  44089=>"111111000",
  44090=>"000000000",
  44091=>"111111111",
  44092=>"101101101",
  44093=>"111111111",
  44094=>"111111111",
  44095=>"000000000",
  44096=>"000000000",
  44097=>"100111111",
  44098=>"111111111",
  44099=>"000000111",
  44100=>"000000001",
  44101=>"000000000",
  44102=>"111101111",
  44103=>"111011000",
  44104=>"011011111",
  44105=>"000100000",
  44106=>"111110000",
  44107=>"001000000",
  44108=>"111111111",
  44109=>"001111011",
  44110=>"111111111",
  44111=>"011011111",
  44112=>"000000000",
  44113=>"110110111",
  44114=>"111100000",
  44115=>"011110110",
  44116=>"000000000",
  44117=>"110110111",
  44118=>"011111110",
  44119=>"010010010",
  44120=>"010010011",
  44121=>"111101101",
  44122=>"000001111",
  44123=>"011011111",
  44124=>"000000111",
  44125=>"011111111",
  44126=>"100000000",
  44127=>"100100100",
  44128=>"111111111",
  44129=>"101111011",
  44130=>"101001101",
  44131=>"111000110",
  44132=>"111111000",
  44133=>"111111011",
  44134=>"000001000",
  44135=>"000000100",
  44136=>"011000000",
  44137=>"111111011",
  44138=>"000000000",
  44139=>"000010111",
  44140=>"100111111",
  44141=>"011010000",
  44142=>"000000000",
  44143=>"000000000",
  44144=>"001111111",
  44145=>"001001011",
  44146=>"111111111",
  44147=>"111000100",
  44148=>"111111111",
  44149=>"111011011",
  44150=>"111111111",
  44151=>"000000110",
  44152=>"111101101",
  44153=>"001101111",
  44154=>"111111100",
  44155=>"000000000",
  44156=>"000000001",
  44157=>"010011000",
  44158=>"111111000",
  44159=>"010110011",
  44160=>"000110000",
  44161=>"111111111",
  44162=>"111111011",
  44163=>"111111001",
  44164=>"000000101",
  44165=>"111000000",
  44166=>"110111101",
  44167=>"100011111",
  44168=>"111011011",
  44169=>"000111111",
  44170=>"110111110",
  44171=>"111111000",
  44172=>"000111100",
  44173=>"000001001",
  44174=>"111111111",
  44175=>"000000001",
  44176=>"111111111",
  44177=>"111111111",
  44178=>"000100111",
  44179=>"111110111",
  44180=>"101001011",
  44181=>"001001111",
  44182=>"000000000",
  44183=>"000000001",
  44184=>"011001000",
  44185=>"011101110",
  44186=>"110110011",
  44187=>"111111111",
  44188=>"111111111",
  44189=>"100000000",
  44190=>"011011000",
  44191=>"000100000",
  44192=>"000000000",
  44193=>"000111111",
  44194=>"000000000",
  44195=>"111111001",
  44196=>"011111001",
  44197=>"000110111",
  44198=>"101111111",
  44199=>"100100100",
  44200=>"000000000",
  44201=>"001000001",
  44202=>"000000000",
  44203=>"000100000",
  44204=>"000000000",
  44205=>"001000000",
  44206=>"111111001",
  44207=>"001011000",
  44208=>"111111111",
  44209=>"011011000",
  44210=>"010111010",
  44211=>"111111010",
  44212=>"011111000",
  44213=>"001111001",
  44214=>"000000000",
  44215=>"100110000",
  44216=>"111111111",
  44217=>"111111010",
  44218=>"101001001",
  44219=>"000000000",
  44220=>"111111111",
  44221=>"011011110",
  44222=>"000000000",
  44223=>"000000000",
  44224=>"000000010",
  44225=>"111111111",
  44226=>"000011111",
  44227=>"111111111",
  44228=>"111111110",
  44229=>"000000001",
  44230=>"011001001",
  44231=>"001111111",
  44232=>"000000000",
  44233=>"000001001",
  44234=>"001000001",
  44235=>"111000000",
  44236=>"111111111",
  44237=>"110110000",
  44238=>"000100100",
  44239=>"000000000",
  44240=>"111010010",
  44241=>"000000000",
  44242=>"000000111",
  44243=>"111111111",
  44244=>"111111111",
  44245=>"001001001",
  44246=>"001001000",
  44247=>"000000011",
  44248=>"001001001",
  44249=>"101111011",
  44250=>"111101011",
  44251=>"111111111",
  44252=>"000000000",
  44253=>"001001001",
  44254=>"111111111",
  44255=>"001011000",
  44256=>"000000100",
  44257=>"100100110",
  44258=>"000000000",
  44259=>"000000000",
  44260=>"111111011",
  44261=>"110100100",
  44262=>"111111111",
  44263=>"111111111",
  44264=>"110110111",
  44265=>"111001111",
  44266=>"110110111",
  44267=>"100000000",
  44268=>"110110110",
  44269=>"000000000",
  44270=>"111111000",
  44271=>"000000000",
  44272=>"101110000",
  44273=>"011011000",
  44274=>"000011111",
  44275=>"000000000",
  44276=>"000000111",
  44277=>"101101110",
  44278=>"001011000",
  44279=>"000000111",
  44280=>"111111111",
  44281=>"000000000",
  44282=>"000000110",
  44283=>"000000000",
  44284=>"000111111",
  44285=>"111111110",
  44286=>"000000000",
  44287=>"110111111",
  44288=>"000000000",
  44289=>"011001000",
  44290=>"000000001",
  44291=>"111111111",
  44292=>"010011001",
  44293=>"000001000",
  44294=>"001001000",
  44295=>"111100110",
  44296=>"000000000",
  44297=>"000000000",
  44298=>"000000110",
  44299=>"111111111",
  44300=>"000000111",
  44301=>"000000010",
  44302=>"000000000",
  44303=>"111111111",
  44304=>"000100101",
  44305=>"110000000",
  44306=>"000000000",
  44307=>"000000001",
  44308=>"000011011",
  44309=>"000001001",
  44310=>"100001000",
  44311=>"111111111",
  44312=>"000001111",
  44313=>"111011000",
  44314=>"111111010",
  44315=>"000000100",
  44316=>"111001111",
  44317=>"000000000",
  44318=>"000000000",
  44319=>"100101110",
  44320=>"001000101",
  44321=>"101001001",
  44322=>"011011000",
  44323=>"110000010",
  44324=>"001001001",
  44325=>"101101111",
  44326=>"111111100",
  44327=>"001000000",
  44328=>"111111000",
  44329=>"110100100",
  44330=>"111111011",
  44331=>"000000000",
  44332=>"010111111",
  44333=>"011011010",
  44334=>"000100000",
  44335=>"000000111",
  44336=>"000000001",
  44337=>"111101000",
  44338=>"111111111",
  44339=>"110010110",
  44340=>"111100111",
  44341=>"111111001",
  44342=>"001101011",
  44343=>"000000000",
  44344=>"000001111",
  44345=>"000000000",
  44346=>"111001000",
  44347=>"110111111",
  44348=>"110100100",
  44349=>"111111000",
  44350=>"011011000",
  44351=>"111111111",
  44352=>"000000000",
  44353=>"101111111",
  44354=>"000010011",
  44355=>"000011000",
  44356=>"000000100",
  44357=>"000000000",
  44358=>"000000011",
  44359=>"111111111",
  44360=>"000000111",
  44361=>"000001000",
  44362=>"111111101",
  44363=>"110110111",
  44364=>"111011011",
  44365=>"111110110",
  44366=>"000001111",
  44367=>"110110110",
  44368=>"100000000",
  44369=>"000111000",
  44370=>"111001001",
  44371=>"000000100",
  44372=>"100000000",
  44373=>"110111111",
  44374=>"000000000",
  44375=>"000000000",
  44376=>"001001000",
  44377=>"000000000",
  44378=>"111011111",
  44379=>"111111110",
  44380=>"000000001",
  44381=>"000000001",
  44382=>"100110110",
  44383=>"000000000",
  44384=>"111111001",
  44385=>"000000000",
  44386=>"111110111",
  44387=>"011001111",
  44388=>"010111111",
  44389=>"000000001",
  44390=>"100111111",
  44391=>"000001001",
  44392=>"010010011",
  44393=>"100101000",
  44394=>"111111111",
  44395=>"000000000",
  44396=>"110111111",
  44397=>"101111011",
  44398=>"000110110",
  44399=>"000100000",
  44400=>"111111111",
  44401=>"000000000",
  44402=>"110110011",
  44403=>"100111000",
  44404=>"111111111",
  44405=>"110011001",
  44406=>"111111111",
  44407=>"100100110",
  44408=>"000000000",
  44409=>"000100111",
  44410=>"110010000",
  44411=>"001000011",
  44412=>"001001001",
  44413=>"101100000",
  44414=>"111111101",
  44415=>"111000010",
  44416=>"111111111",
  44417=>"110110111",
  44418=>"000000000",
  44419=>"100000000",
  44420=>"000000111",
  44421=>"000000000",
  44422=>"000100111",
  44423=>"000000000",
  44424=>"100111000",
  44425=>"000000001",
  44426=>"111111111",
  44427=>"000000000",
  44428=>"111111111",
  44429=>"001001000",
  44430=>"011011001",
  44431=>"111111111",
  44432=>"000100111",
  44433=>"001000000",
  44434=>"000000000",
  44435=>"011011011",
  44436=>"000000000",
  44437=>"000000000",
  44438=>"000000001",
  44439=>"011011011",
  44440=>"111110110",
  44441=>"000001000",
  44442=>"111101000",
  44443=>"011001000",
  44444=>"000100111",
  44445=>"111111111",
  44446=>"100100100",
  44447=>"000010000",
  44448=>"000000000",
  44449=>"110100100",
  44450=>"000000110",
  44451=>"111111111",
  44452=>"000110111",
  44453=>"000000000",
  44454=>"000000000",
  44455=>"000000000",
  44456=>"000000011",
  44457=>"111110110",
  44458=>"111011111",
  44459=>"000000000",
  44460=>"000011111",
  44461=>"001000000",
  44462=>"000000000",
  44463=>"001001000",
  44464=>"111111111",
  44465=>"100100000",
  44466=>"111111011",
  44467=>"111111111",
  44468=>"000011111",
  44469=>"001101100",
  44470=>"111111101",
  44471=>"011111000",
  44472=>"000000011",
  44473=>"011111111",
  44474=>"111001000",
  44475=>"000011011",
  44476=>"000000000",
  44477=>"001000101",
  44478=>"111000001",
  44479=>"001011111",
  44480=>"111111111",
  44481=>"100100000",
  44482=>"000000000",
  44483=>"011110110",
  44484=>"001000000",
  44485=>"000000011",
  44486=>"001001000",
  44487=>"100000001",
  44488=>"110000000",
  44489=>"011011111",
  44490=>"011000000",
  44491=>"011011000",
  44492=>"111000000",
  44493=>"111001000",
  44494=>"001001001",
  44495=>"001101111",
  44496=>"100000001",
  44497=>"000011011",
  44498=>"111111111",
  44499=>"100111111",
  44500=>"100100110",
  44501=>"111111101",
  44502=>"000111111",
  44503=>"111111011",
  44504=>"001001111",
  44505=>"011111011",
  44506=>"000000000",
  44507=>"101001001",
  44508=>"000111100",
  44509=>"000000111",
  44510=>"000110100",
  44511=>"111111111",
  44512=>"000101111",
  44513=>"000000001",
  44514=>"000000000",
  44515=>"000111111",
  44516=>"000001000",
  44517=>"111111111",
  44518=>"111111000",
  44519=>"000000000",
  44520=>"011001001",
  44521=>"001011111",
  44522=>"011011011",
  44523=>"000000000",
  44524=>"111111000",
  44525=>"100000100",
  44526=>"110000000",
  44527=>"101001000",
  44528=>"111110110",
  44529=>"000000000",
  44530=>"000000000",
  44531=>"110110111",
  44532=>"000000000",
  44533=>"110111111",
  44534=>"111111111",
  44535=>"000010000",
  44536=>"000000000",
  44537=>"000100100",
  44538=>"000111111",
  44539=>"111111111",
  44540=>"001000000",
  44541=>"000111011",
  44542=>"000011111",
  44543=>"000000000",
  44544=>"111111011",
  44545=>"100001000",
  44546=>"000000000",
  44547=>"001011011",
  44548=>"110101000",
  44549=>"101101101",
  44550=>"011001001",
  44551=>"101111111",
  44552=>"001011001",
  44553=>"000001101",
  44554=>"111100000",
  44555=>"111111111",
  44556=>"100000000",
  44557=>"111000000",
  44558=>"000000000",
  44559=>"111100111",
  44560=>"000000111",
  44561=>"111000111",
  44562=>"111100001",
  44563=>"000001111",
  44564=>"000000000",
  44565=>"111111101",
  44566=>"110010010",
  44567=>"000000100",
  44568=>"011011011",
  44569=>"111111111",
  44570=>"000100101",
  44571=>"011000111",
  44572=>"111111111",
  44573=>"011000000",
  44574=>"011001001",
  44575=>"010000000",
  44576=>"110000011",
  44577=>"111111010",
  44578=>"000011000",
  44579=>"100100110",
  44580=>"010010110",
  44581=>"000000000",
  44582=>"100000000",
  44583=>"001111001",
  44584=>"001101111",
  44585=>"101101001",
  44586=>"100000000",
  44587=>"110110110",
  44588=>"111101001",
  44589=>"111111101",
  44590=>"001000000",
  44591=>"101111111",
  44592=>"100100000",
  44593=>"000001011",
  44594=>"000110110",
  44595=>"111011000",
  44596=>"101101101",
  44597=>"110110100",
  44598=>"111001000",
  44599=>"000000000",
  44600=>"100000000",
  44601=>"110111000",
  44602=>"000000101",
  44603=>"011000000",
  44604=>"101101110",
  44605=>"110000000",
  44606=>"110110001",
  44607=>"011011001",
  44608=>"001001000",
  44609=>"001100100",
  44610=>"010110011",
  44611=>"100000000",
  44612=>"011001001",
  44613=>"011111111",
  44614=>"000000000",
  44615=>"111100111",
  44616=>"111111001",
  44617=>"000000000",
  44618=>"111111101",
  44619=>"000000111",
  44620=>"001001001",
  44621=>"110100111",
  44622=>"101101101",
  44623=>"000100111",
  44624=>"000001001",
  44625=>"001101101",
  44626=>"111000000",
  44627=>"011110100",
  44628=>"111101001",
  44629=>"001010000",
  44630=>"110010011",
  44631=>"110110010",
  44632=>"000000110",
  44633=>"100000110",
  44634=>"100010111",
  44635=>"100000001",
  44636=>"110010010",
  44637=>"100111111",
  44638=>"000000000",
  44639=>"100100111",
  44640=>"000010010",
  44641=>"101101101",
  44642=>"111011001",
  44643=>"011101001",
  44644=>"001011010",
  44645=>"001001001",
  44646=>"100110110",
  44647=>"110000000",
  44648=>"111110110",
  44649=>"001000111",
  44650=>"001001010",
  44651=>"010000001",
  44652=>"010000000",
  44653=>"011111111",
  44654=>"000000010",
  44655=>"000000100",
  44656=>"101001101",
  44657=>"100000000",
  44658=>"101101101",
  44659=>"001011111",
  44660=>"011111101",
  44661=>"000000010",
  44662=>"101101101",
  44663=>"110111100",
  44664=>"100101111",
  44665=>"110111111",
  44666=>"110000010",
  44667=>"000111111",
  44668=>"100100101",
  44669=>"110100000",
  44670=>"110110010",
  44671=>"111111100",
  44672=>"001001000",
  44673=>"001000100",
  44674=>"101000110",
  44675=>"000101101",
  44676=>"100110010",
  44677=>"000000000",
  44678=>"100000000",
  44679=>"111110110",
  44680=>"000000111",
  44681=>"000100000",
  44682=>"000001011",
  44683=>"111111111",
  44684=>"111111111",
  44685=>"100110011",
  44686=>"101001101",
  44687=>"110100111",
  44688=>"001001100",
  44689=>"001101101",
  44690=>"111001111",
  44691=>"011010010",
  44692=>"100110110",
  44693=>"111111010",
  44694=>"000101000",
  44695=>"101101101",
  44696=>"101000000",
  44697=>"000001001",
  44698=>"010010110",
  44699=>"001101100",
  44700=>"110110110",
  44701=>"011011110",
  44702=>"111111111",
  44703=>"000000000",
  44704=>"110000001",
  44705=>"101111111",
  44706=>"011011111",
  44707=>"110000101",
  44708=>"110010000",
  44709=>"111111110",
  44710=>"001111001",
  44711=>"001000000",
  44712=>"001111100",
  44713=>"000000001",
  44714=>"001000000",
  44715=>"000110000",
  44716=>"000110111",
  44717=>"100100100",
  44718=>"111010000",
  44719=>"000000000",
  44720=>"001011111",
  44721=>"100100111",
  44722=>"111111111",
  44723=>"111101000",
  44724=>"000010000",
  44725=>"111110010",
  44726=>"000000000",
  44727=>"100001011",
  44728=>"100010110",
  44729=>"110111110",
  44730=>"110110100",
  44731=>"110110110",
  44732=>"111111111",
  44733=>"010110110",
  44734=>"000010111",
  44735=>"000010110",
  44736=>"000001011",
  44737=>"111000000",
  44738=>"000000010",
  44739=>"110110110",
  44740=>"001001000",
  44741=>"000011000",
  44742=>"110110111",
  44743=>"110100100",
  44744=>"000111111",
  44745=>"000100100",
  44746=>"101100100",
  44747=>"011111111",
  44748=>"000000100",
  44749=>"011100100",
  44750=>"111111101",
  44751=>"010010000",
  44752=>"111111111",
  44753=>"001001101",
  44754=>"010010010",
  44755=>"000000100",
  44756=>"111011000",
  44757=>"110011011",
  44758=>"000000000",
  44759=>"000110110",
  44760=>"000011000",
  44761=>"000100100",
  44762=>"100110100",
  44763=>"111111111",
  44764=>"000000010",
  44765=>"000000010",
  44766=>"111111101",
  44767=>"110110000",
  44768=>"000000010",
  44769=>"101111100",
  44770=>"110010000",
  44771=>"000000001",
  44772=>"011011111",
  44773=>"011001001",
  44774=>"110110110",
  44775=>"111111111",
  44776=>"101101110",
  44777=>"000110001",
  44778=>"100000000",
  44779=>"111111001",
  44780=>"010000000",
  44781=>"000000000",
  44782=>"111011111",
  44783=>"110111111",
  44784=>"010011011",
  44785=>"011000000",
  44786=>"110111111",
  44787=>"110110011",
  44788=>"000111111",
  44789=>"000011010",
  44790=>"001010111",
  44791=>"001000000",
  44792=>"000000000",
  44793=>"000000001",
  44794=>"001101111",
  44795=>"000001101",
  44796=>"000010100",
  44797=>"001000100",
  44798=>"111111110",
  44799=>"111100110",
  44800=>"100000001",
  44801=>"111111001",
  44802=>"111111111",
  44803=>"110100100",
  44804=>"000000000",
  44805=>"001110111",
  44806=>"110110010",
  44807=>"110111111",
  44808=>"110010010",
  44809=>"000000000",
  44810=>"000000100",
  44811=>"100000000",
  44812=>"011001011",
  44813=>"000000010",
  44814=>"111011110",
  44815=>"011111111",
  44816=>"110110010",
  44817=>"111111111",
  44818=>"000111111",
  44819=>"000000111",
  44820=>"110110010",
  44821=>"101000001",
  44822=>"100101101",
  44823=>"111110110",
  44824=>"111111111",
  44825=>"011000000",
  44826=>"000001011",
  44827=>"011001001",
  44828=>"110100110",
  44829=>"011001011",
  44830=>"001101001",
  44831=>"111001111",
  44832=>"000011000",
  44833=>"101101101",
  44834=>"000001001",
  44835=>"111111111",
  44836=>"110110000",
  44837=>"100111100",
  44838=>"111011000",
  44839=>"010110100",
  44840=>"110110110",
  44841=>"111011011",
  44842=>"101111111",
  44843=>"000000100",
  44844=>"111001011",
  44845=>"011100100",
  44846=>"000110000",
  44847=>"000000000",
  44848=>"001001111",
  44849=>"110111101",
  44850=>"010000000",
  44851=>"011011011",
  44852=>"000000000",
  44853=>"000000111",
  44854=>"100100100",
  44855=>"000001111",
  44856=>"111111100",
  44857=>"101100100",
  44858=>"110010011",
  44859=>"000000000",
  44860=>"111110111",
  44861=>"111011001",
  44862=>"110110010",
  44863=>"000000011",
  44864=>"101100100",
  44865=>"000000110",
  44866=>"000010111",
  44867=>"000000000",
  44868=>"001001110",
  44869=>"000000000",
  44870=>"000000000",
  44871=>"111000001",
  44872=>"000000000",
  44873=>"100000010",
  44874=>"110110110",
  44875=>"011010000",
  44876=>"110110110",
  44877=>"111111001",
  44878=>"111011000",
  44879=>"000000000",
  44880=>"011011111",
  44881=>"011011001",
  44882=>"000001111",
  44883=>"000001011",
  44884=>"100101111",
  44885=>"011010000",
  44886=>"110110110",
  44887=>"000000011",
  44888=>"000111011",
  44889=>"000101111",
  44890=>"111010111",
  44891=>"111111111",
  44892=>"000100000",
  44893=>"000000000",
  44894=>"001000000",
  44895=>"100100100",
  44896=>"011111111",
  44897=>"001001001",
  44898=>"100101100",
  44899=>"100111111",
  44900=>"110100100",
  44901=>"110110100",
  44902=>"101101111",
  44903=>"101111001",
  44904=>"100001001",
  44905=>"000110110",
  44906=>"111111111",
  44907=>"001001001",
  44908=>"010011001",
  44909=>"110100100",
  44910=>"000001000",
  44911=>"100100100",
  44912=>"110000000",
  44913=>"000100111",
  44914=>"111100101",
  44915=>"011011001",
  44916=>"011010010",
  44917=>"010011000",
  44918=>"000000001",
  44919=>"001000001",
  44920=>"001111111",
  44921=>"000000000",
  44922=>"000100101",
  44923=>"100100010",
  44924=>"010010111",
  44925=>"110010010",
  44926=>"100000000",
  44927=>"111111111",
  44928=>"110110110",
  44929=>"010010010",
  44930=>"000000000",
  44931=>"000001111",
  44932=>"010011001",
  44933=>"000000000",
  44934=>"001000000",
  44935=>"110011001",
  44936=>"001000000",
  44937=>"010000000",
  44938=>"001101111",
  44939=>"000000000",
  44940=>"111111111",
  44941=>"000000000",
  44942=>"110110000",
  44943=>"011111111",
  44944=>"000001001",
  44945=>"110101111",
  44946=>"000000000",
  44947=>"000000000",
  44948=>"101110101",
  44949=>"010010000",
  44950=>"111000000",
  44951=>"110100100",
  44952=>"101001101",
  44953=>"111011011",
  44954=>"010000110",
  44955=>"101001111",
  44956=>"001101101",
  44957=>"111000000",
  44958=>"110110100",
  44959=>"011010010",
  44960=>"000000000",
  44961=>"000000000",
  44962=>"111111111",
  44963=>"000000000",
  44964=>"100100110",
  44965=>"001101111",
  44966=>"001111010",
  44967=>"101101101",
  44968=>"110100000",
  44969=>"010011000",
  44970=>"111001001",
  44971=>"111101101",
  44972=>"000011000",
  44973=>"111000111",
  44974=>"000100111",
  44975=>"011011011",
  44976=>"111111010",
  44977=>"100000000",
  44978=>"000000000",
  44979=>"101101101",
  44980=>"100100111",
  44981=>"011011011",
  44982=>"100111111",
  44983=>"000100000",
  44984=>"000100110",
  44985=>"110111111",
  44986=>"111111011",
  44987=>"000000111",
  44988=>"001001000",
  44989=>"000000000",
  44990=>"101101101",
  44991=>"110100100",
  44992=>"001111111",
  44993=>"001101001",
  44994=>"001101111",
  44995=>"010011110",
  44996=>"101111110",
  44997=>"001001101",
  44998=>"100000111",
  44999=>"100000100",
  45000=>"110000100",
  45001=>"011000000",
  45002=>"000000000",
  45003=>"000000000",
  45004=>"101111000",
  45005=>"100000100",
  45006=>"111111111",
  45007=>"111001001",
  45008=>"000000000",
  45009=>"011011001",
  45010=>"111111111",
  45011=>"000111111",
  45012=>"000100111",
  45013=>"000000011",
  45014=>"101101101",
  45015=>"111101101",
  45016=>"101101001",
  45017=>"001101111",
  45018=>"111110010",
  45019=>"110000001",
  45020=>"011001000",
  45021=>"000011111",
  45022=>"000110110",
  45023=>"010010010",
  45024=>"111111101",
  45025=>"010000100",
  45026=>"011111111",
  45027=>"111001111",
  45028=>"110000100",
  45029=>"100100110",
  45030=>"101111111",
  45031=>"000000100",
  45032=>"110110110",
  45033=>"110111100",
  45034=>"001111111",
  45035=>"000011000",
  45036=>"111011111",
  45037=>"011010011",
  45038=>"101101101",
  45039=>"111100001",
  45040=>"000010011",
  45041=>"101011101",
  45042=>"011110111",
  45043=>"001000101",
  45044=>"110011011",
  45045=>"111111011",
  45046=>"100000001",
  45047=>"111000000",
  45048=>"001111100",
  45049=>"011011000",
  45050=>"110111111",
  45051=>"101001001",
  45052=>"100111100",
  45053=>"110000000",
  45054=>"100000111",
  45055=>"000000000",
  45056=>"000000000",
  45057=>"001111111",
  45058=>"000000111",
  45059=>"000000000",
  45060=>"000001001",
  45061=>"000100100",
  45062=>"000000000",
  45063=>"101000000",
  45064=>"111111001",
  45065=>"001000000",
  45066=>"000000000",
  45067=>"111111111",
  45068=>"000000111",
  45069=>"000000000",
  45070=>"000000000",
  45071=>"000000000",
  45072=>"000100101",
  45073=>"100000101",
  45074=>"000010001",
  45075=>"111111111",
  45076=>"000000110",
  45077=>"000000000",
  45078=>"110110111",
  45079=>"111111001",
  45080=>"100110110",
  45081=>"001010011",
  45082=>"111000000",
  45083=>"000000000",
  45084=>"100000000",
  45085=>"100111001",
  45086=>"111011111",
  45087=>"000011000",
  45088=>"000000001",
  45089=>"111111111",
  45090=>"000000000",
  45091=>"000000000",
  45092=>"110110001",
  45093=>"011000000",
  45094=>"000000000",
  45095=>"000000011",
  45096=>"111111111",
  45097=>"000000000",
  45098=>"000000000",
  45099=>"111111110",
  45100=>"111111111",
  45101=>"011111100",
  45102=>"001100110",
  45103=>"000000000",
  45104=>"000000000",
  45105=>"000000000",
  45106=>"111111111",
  45107=>"111110010",
  45108=>"111111111",
  45109=>"011011000",
  45110=>"000100000",
  45111=>"010000000",
  45112=>"110110000",
  45113=>"111111111",
  45114=>"000000000",
  45115=>"101111110",
  45116=>"000000001",
  45117=>"000000111",
  45118=>"110111111",
  45119=>"001000000",
  45120=>"000011001",
  45121=>"100000111",
  45122=>"111111111",
  45123=>"111111101",
  45124=>"110110000",
  45125=>"000000000",
  45126=>"001000000",
  45127=>"100000000",
  45128=>"000000001",
  45129=>"000000000",
  45130=>"111111111",
  45131=>"111111111",
  45132=>"110111111",
  45133=>"111111111",
  45134=>"111001101",
  45135=>"001011111",
  45136=>"111111111",
  45137=>"111111011",
  45138=>"111110010",
  45139=>"010100000",
  45140=>"000000000",
  45141=>"001000000",
  45142=>"111110001",
  45143=>"011001000",
  45144=>"000000000",
  45145=>"000000001",
  45146=>"111100111",
  45147=>"000010011",
  45148=>"111111111",
  45149=>"111111111",
  45150=>"000011010",
  45151=>"100100100",
  45152=>"000000000",
  45153=>"000000000",
  45154=>"000010000",
  45155=>"001000101",
  45156=>"111000000",
  45157=>"000000000",
  45158=>"111110000",
  45159=>"111111110",
  45160=>"111111111",
  45161=>"111111111",
  45162=>"111111000",
  45163=>"110110000",
  45164=>"111111110",
  45165=>"000000000",
  45166=>"111111111",
  45167=>"000000000",
  45168=>"111000000",
  45169=>"111111111",
  45170=>"111101101",
  45171=>"001000101",
  45172=>"111111111",
  45173=>"111100000",
  45174=>"110100011",
  45175=>"110111100",
  45176=>"000000000",
  45177=>"000000000",
  45178=>"000000000",
  45179=>"111111111",
  45180=>"110100100",
  45181=>"000000000",
  45182=>"010000000",
  45183=>"111111000",
  45184=>"000000000",
  45185=>"111111111",
  45186=>"000000000",
  45187=>"100111001",
  45188=>"111110111",
  45189=>"000000000",
  45190=>"000000000",
  45191=>"000000111",
  45192=>"101111111",
  45193=>"011011101",
  45194=>"000000111",
  45195=>"000000000",
  45196=>"000000110",
  45197=>"000000000",
  45198=>"111111111",
  45199=>"111111111",
  45200=>"110111111",
  45201=>"000000000",
  45202=>"000011111",
  45203=>"000000000",
  45204=>"011000000",
  45205=>"111111110",
  45206=>"001111111",
  45207=>"000110110",
  45208=>"000111111",
  45209=>"000000100",
  45210=>"001001001",
  45211=>"100000000",
  45212=>"011000000",
  45213=>"000110111",
  45214=>"111110111",
  45215=>"111111111",
  45216=>"000011000",
  45217=>"001001111",
  45218=>"111111111",
  45219=>"000000010",
  45220=>"000000000",
  45221=>"111111111",
  45222=>"111100101",
  45223=>"010111110",
  45224=>"111011111",
  45225=>"000000000",
  45226=>"000111011",
  45227=>"111111111",
  45228=>"110111000",
  45229=>"100000000",
  45230=>"101111111",
  45231=>"000000000",
  45232=>"111100101",
  45233=>"000001000",
  45234=>"110111111",
  45235=>"111000011",
  45236=>"010000000",
  45237=>"111111111",
  45238=>"000000000",
  45239=>"011011111",
  45240=>"111110100",
  45241=>"011001001",
  45242=>"000000000",
  45243=>"010110111",
  45244=>"100110000",
  45245=>"111111111",
  45246=>"000000000",
  45247=>"111111111",
  45248=>"000000000",
  45249=>"111111111",
  45250=>"000000010",
  45251=>"110111000",
  45252=>"000000000",
  45253=>"000000000",
  45254=>"110000100",
  45255=>"000100111",
  45256=>"111110000",
  45257=>"011001000",
  45258=>"100111111",
  45259=>"000100000",
  45260=>"111111111",
  45261=>"000000000",
  45262=>"000000110",
  45263=>"000011000",
  45264=>"000000000",
  45265=>"000000000",
  45266=>"011000000",
  45267=>"010010000",
  45268=>"000000000",
  45269=>"000000001",
  45270=>"111000000",
  45271=>"111000000",
  45272=>"110110111",
  45273=>"111011011",
  45274=>"000000110",
  45275=>"111111100",
  45276=>"001110111",
  45277=>"000000001",
  45278=>"111111111",
  45279=>"110100000",
  45280=>"000000000",
  45281=>"111111000",
  45282=>"000000000",
  45283=>"111111111",
  45284=>"000111111",
  45285=>"011011000",
  45286=>"100000110",
  45287=>"000110000",
  45288=>"111111111",
  45289=>"110111001",
  45290=>"111110010",
  45291=>"110100100",
  45292=>"000000101",
  45293=>"000000000",
  45294=>"000001011",
  45295=>"000110100",
  45296=>"000000111",
  45297=>"000000011",
  45298=>"111111001",
  45299=>"000000000",
  45300=>"111111111",
  45301=>"011011011",
  45302=>"000000000",
  45303=>"000000100",
  45304=>"000000000",
  45305=>"000000001",
  45306=>"011001010",
  45307=>"101000000",
  45308=>"111001101",
  45309=>"000001001",
  45310=>"010000111",
  45311=>"000000000",
  45312=>"001000000",
  45313=>"111111111",
  45314=>"111111111",
  45315=>"000000000",
  45316=>"000000000",
  45317=>"111110000",
  45318=>"111000001",
  45319=>"001101111",
  45320=>"111110111",
  45321=>"000000000",
  45322=>"000000000",
  45323=>"111111001",
  45324=>"111111111",
  45325=>"000000000",
  45326=>"100000000",
  45327=>"000100100",
  45328=>"111111111",
  45329=>"000000001",
  45330=>"000000001",
  45331=>"000000010",
  45332=>"000000000",
  45333=>"000000000",
  45334=>"011000000",
  45335=>"000001001",
  45336=>"111110000",
  45337=>"001000000",
  45338=>"000000001",
  45339=>"111111010",
  45340=>"001001000",
  45341=>"011011000",
  45342=>"000000000",
  45343=>"001111000",
  45344=>"000000000",
  45345=>"001111111",
  45346=>"111110111",
  45347=>"011001000",
  45348=>"111111111",
  45349=>"111111111",
  45350=>"111111111",
  45351=>"111111111",
  45352=>"100100001",
  45353=>"000000001",
  45354=>"000000000",
  45355=>"000111111",
  45356=>"000000000",
  45357=>"000000000",
  45358=>"110111111",
  45359=>"000000000",
  45360=>"111111111",
  45361=>"111111111",
  45362=>"010111111",
  45363=>"111100111",
  45364=>"000111111",
  45365=>"111101111",
  45366=>"111011000",
  45367=>"111100111",
  45368=>"000000100",
  45369=>"000000000",
  45370=>"111111000",
  45371=>"011111000",
  45372=>"111111111",
  45373=>"111101100",
  45374=>"101000101",
  45375=>"011010000",
  45376=>"000010000",
  45377=>"010111111",
  45378=>"000000001",
  45379=>"110110111",
  45380=>"111000000",
  45381=>"111011000",
  45382=>"010010011",
  45383=>"000000000",
  45384=>"000000111",
  45385=>"011011111",
  45386=>"111111100",
  45387=>"110110110",
  45388=>"000000110",
  45389=>"000000000",
  45390=>"111111111",
  45391=>"111110100",
  45392=>"111111111",
  45393=>"110111101",
  45394=>"000000000",
  45395=>"000000000",
  45396=>"000000000",
  45397=>"011011011",
  45398=>"111111111",
  45399=>"001001000",
  45400=>"000000011",
  45401=>"111111111",
  45402=>"000100100",
  45403=>"001111111",
  45404=>"011011000",
  45405=>"111111111",
  45406=>"000010000",
  45407=>"111111111",
  45408=>"001000000",
  45409=>"110111111",
  45410=>"111110111",
  45411=>"111111111",
  45412=>"100000000",
  45413=>"000000000",
  45414=>"000111111",
  45415=>"000000001",
  45416=>"001001011",
  45417=>"111111111",
  45418=>"110000101",
  45419=>"000000000",
  45420=>"011011111",
  45421=>"000011010",
  45422=>"000000000",
  45423=>"000000110",
  45424=>"001110011",
  45425=>"000000100",
  45426=>"000001111",
  45427=>"111110000",
  45428=>"011011111",
  45429=>"000000000",
  45430=>"011111000",
  45431=>"000000000",
  45432=>"010010000",
  45433=>"001111111",
  45434=>"000000000",
  45435=>"110111111",
  45436=>"000000001",
  45437=>"100100000",
  45438=>"000000101",
  45439=>"000000111",
  45440=>"110000000",
  45441=>"000100101",
  45442=>"000000000",
  45443=>"000000000",
  45444=>"110000000",
  45445=>"000010010",
  45446=>"111100000",
  45447=>"000001111",
  45448=>"000010011",
  45449=>"111111111",
  45450=>"000000000",
  45451=>"111110000",
  45452=>"101111111",
  45453=>"100110011",
  45454=>"111111111",
  45455=>"000000000",
  45456=>"000000000",
  45457=>"111111010",
  45458=>"001000100",
  45459=>"000111111",
  45460=>"110111111",
  45461=>"000000000",
  45462=>"000011001",
  45463=>"000000110",
  45464=>"101101111",
  45465=>"110000000",
  45466=>"000000000",
  45467=>"111111111",
  45468=>"111111000",
  45469=>"000000000",
  45470=>"111000000",
  45471=>"000000000",
  45472=>"000100001",
  45473=>"001011000",
  45474=>"111111000",
  45475=>"111011111",
  45476=>"111111101",
  45477=>"111111111",
  45478=>"110111110",
  45479=>"111111111",
  45480=>"111100000",
  45481=>"011011010",
  45482=>"111111111",
  45483=>"111000000",
  45484=>"000011000",
  45485=>"000100100",
  45486=>"001000000",
  45487=>"111111011",
  45488=>"010000000",
  45489=>"111111000",
  45490=>"111111111",
  45491=>"000000010",
  45492=>"011000110",
  45493=>"100101101",
  45494=>"111111111",
  45495=>"111111011",
  45496=>"000000010",
  45497=>"110111111",
  45498=>"000000100",
  45499=>"000001111",
  45500=>"100000000",
  45501=>"100000111",
  45502=>"000000000",
  45503=>"001011010",
  45504=>"111100111",
  45505=>"011000011",
  45506=>"000000000",
  45507=>"000000000",
  45508=>"111100000",
  45509=>"000000011",
  45510=>"111000000",
  45511=>"000000000",
  45512=>"000001011",
  45513=>"100100000",
  45514=>"000000111",
  45515=>"000000000",
  45516=>"011000011",
  45517=>"111111000",
  45518=>"011001000",
  45519=>"111111100",
  45520=>"001110100",
  45521=>"000000000",
  45522=>"000000001",
  45523=>"000000000",
  45524=>"111110111",
  45525=>"000111111",
  45526=>"000000000",
  45527=>"000111001",
  45528=>"001010010",
  45529=>"000001000",
  45530=>"100111110",
  45531=>"111111111",
  45532=>"111111011",
  45533=>"111100100",
  45534=>"111111011",
  45535=>"011111011",
  45536=>"001000000",
  45537=>"111111111",
  45538=>"011011001",
  45539=>"111001001",
  45540=>"001011110",
  45541=>"111000111",
  45542=>"001000001",
  45543=>"000000000",
  45544=>"001100000",
  45545=>"111111111",
  45546=>"111000000",
  45547=>"111111000",
  45548=>"111111000",
  45549=>"111111111",
  45550=>"100111111",
  45551=>"111110100",
  45552=>"000111111",
  45553=>"000000000",
  45554=>"001001111",
  45555=>"000000000",
  45556=>"111111111",
  45557=>"010000000",
  45558=>"000000000",
  45559=>"001000110",
  45560=>"110110001",
  45561=>"000010011",
  45562=>"001011000",
  45563=>"100111111",
  45564=>"111111010",
  45565=>"111110111",
  45566=>"000010110",
  45567=>"110110110",
  45568=>"001001111",
  45569=>"111111111",
  45570=>"111000000",
  45571=>"000000111",
  45572=>"000000100",
  45573=>"101000101",
  45574=>"011111111",
  45575=>"101000001",
  45576=>"010011000",
  45577=>"101000000",
  45578=>"000000000",
  45579=>"110001011",
  45580=>"100001101",
  45581=>"000000001",
  45582=>"000000111",
  45583=>"000000000",
  45584=>"111000000",
  45585=>"000011011",
  45586=>"000111111",
  45587=>"111000001",
  45588=>"111111111",
  45589=>"000001000",
  45590=>"000000101",
  45591=>"000000001",
  45592=>"111110110",
  45593=>"011000000",
  45594=>"111110110",
  45595=>"001000000",
  45596=>"000110110",
  45597=>"110110111",
  45598=>"000010010",
  45599=>"000101111",
  45600=>"111010000",
  45601=>"111101000",
  45602=>"100010100",
  45603=>"000100111",
  45604=>"000001111",
  45605=>"000000000",
  45606=>"111000100",
  45607=>"111000000",
  45608=>"111111111",
  45609=>"111111011",
  45610=>"000000000",
  45611=>"100111111",
  45612=>"111011000",
  45613=>"101101110",
  45614=>"110111110",
  45615=>"001000010",
  45616=>"000000100",
  45617=>"000000011",
  45618=>"011111010",
  45619=>"100100100",
  45620=>"000100111",
  45621=>"111111111",
  45622=>"100000000",
  45623=>"000000000",
  45624=>"000001101",
  45625=>"111001001",
  45626=>"111111111",
  45627=>"000000000",
  45628=>"111100100",
  45629=>"111000100",
  45630=>"000000000",
  45631=>"110111010",
  45632=>"001000000",
  45633=>"000110110",
  45634=>"010111111",
  45635=>"111000000",
  45636=>"100100110",
  45637=>"000111111",
  45638=>"000000000",
  45639=>"111111111",
  45640=>"111111110",
  45641=>"001000001",
  45642=>"011001011",
  45643=>"111111111",
  45644=>"111111000",
  45645=>"111001111",
  45646=>"111111010",
  45647=>"100100110",
  45648=>"100000000",
  45649=>"000000000",
  45650=>"111010000",
  45651=>"001001111",
  45652=>"000000011",
  45653=>"000000100",
  45654=>"100000111",
  45655=>"110111111",
  45656=>"110111111",
  45657=>"000000000",
  45658=>"000000000",
  45659=>"111111100",
  45660=>"000000001",
  45661=>"000000010",
  45662=>"000000110",
  45663=>"100100000",
  45664=>"100000000",
  45665=>"100000000",
  45666=>"011111110",
  45667=>"010010000",
  45668=>"000011111",
  45669=>"100000011",
  45670=>"101101110",
  45671=>"000000111",
  45672=>"000010000",
  45673=>"111000000",
  45674=>"011000000",
  45675=>"000111011",
  45676=>"000001101",
  45677=>"111111111",
  45678=>"001001001",
  45679=>"011010000",
  45680=>"111111001",
  45681=>"101100111",
  45682=>"100110000",
  45683=>"111111001",
  45684=>"110100000",
  45685=>"010110111",
  45686=>"000000000",
  45687=>"000000000",
  45688=>"010000000",
  45689=>"100000111",
  45690=>"001000000",
  45691=>"000000001",
  45692=>"111110110",
  45693=>"111111010",
  45694=>"111111011",
  45695=>"000000000",
  45696=>"110111010",
  45697=>"111011000",
  45698=>"111011000",
  45699=>"100000100",
  45700=>"111111111",
  45701=>"011111000",
  45702=>"111111111",
  45703=>"010010000",
  45704=>"100011011",
  45705=>"110110111",
  45706=>"000100111",
  45707=>"111111110",
  45708=>"010000111",
  45709=>"000110000",
  45710=>"111111000",
  45711=>"010011111",
  45712=>"111111110",
  45713=>"101011111",
  45714=>"011000000",
  45715=>"001001111",
  45716=>"001111111",
  45717=>"000000110",
  45718=>"000000000",
  45719=>"100100000",
  45720=>"000000100",
  45721=>"000100110",
  45722=>"111111010",
  45723=>"000000000",
  45724=>"111110100",
  45725=>"111000011",
  45726=>"110110000",
  45727=>"001011011",
  45728=>"110000000",
  45729=>"111111011",
  45730=>"010000010",
  45731=>"111111011",
  45732=>"000000000",
  45733=>"111000000",
  45734=>"001000111",
  45735=>"100100101",
  45736=>"000000001",
  45737=>"001000000",
  45738=>"000001011",
  45739=>"111011111",
  45740=>"101000000",
  45741=>"100111100",
  45742=>"110110111",
  45743=>"000000000",
  45744=>"111000000",
  45745=>"000000001",
  45746=>"111111111",
  45747=>"000000000",
  45748=>"111101101",
  45749=>"111111101",
  45750=>"110111111",
  45751=>"111111001",
  45752=>"010110110",
  45753=>"000000001",
  45754=>"000011000",
  45755=>"100010111",
  45756=>"110110100",
  45757=>"111111011",
  45758=>"111111110",
  45759=>"111000100",
  45760=>"111110100",
  45761=>"000000000",
  45762=>"111011011",
  45763=>"001001111",
  45764=>"111111110",
  45765=>"100111111",
  45766=>"000000000",
  45767=>"011001101",
  45768=>"000000000",
  45769=>"110111100",
  45770=>"101000000",
  45771=>"001001001",
  45772=>"100000101",
  45773=>"111100000",
  45774=>"000000100",
  45775=>"101001000",
  45776=>"111111111",
  45777=>"011000000",
  45778=>"000111010",
  45779=>"000000001",
  45780=>"000000000",
  45781=>"111110110",
  45782=>"000000100",
  45783=>"001000000",
  45784=>"011111111",
  45785=>"110110110",
  45786=>"001001111",
  45787=>"000111111",
  45788=>"111011111",
  45789=>"110100110",
  45790=>"000010000",
  45791=>"111011000",
  45792=>"000000111",
  45793=>"001111111",
  45794=>"111001111",
  45795=>"110110111",
  45796=>"011111000",
  45797=>"000111000",
  45798=>"000000001",
  45799=>"111111111",
  45800=>"001000000",
  45801=>"111111111",
  45802=>"111111111",
  45803=>"111111011",
  45804=>"110111010",
  45805=>"111001000",
  45806=>"111111011",
  45807=>"000110000",
  45808=>"000000000",
  45809=>"111000010",
  45810=>"000000000",
  45811=>"100000000",
  45812=>"010011011",
  45813=>"011010001",
  45814=>"111100111",
  45815=>"000111111",
  45816=>"001000001",
  45817=>"000000000",
  45818=>"100000000",
  45819=>"101101111",
  45820=>"001111111",
  45821=>"110110100",
  45822=>"111111011",
  45823=>"011111111",
  45824=>"000000001",
  45825=>"100101101",
  45826=>"001001000",
  45827=>"111110100",
  45828=>"000111111",
  45829=>"110111110",
  45830=>"000000000",
  45831=>"000000111",
  45832=>"110000000",
  45833=>"111111111",
  45834=>"000000100",
  45835=>"011111111",
  45836=>"001000000",
  45837=>"100111100",
  45838=>"100111111",
  45839=>"111111001",
  45840=>"000000001",
  45841=>"100100000",
  45842=>"001000010",
  45843=>"000000000",
  45844=>"000000000",
  45845=>"000000000",
  45846=>"111111111",
  45847=>"100111111",
  45848=>"011000110",
  45849=>"111111111",
  45850=>"000000111",
  45851=>"011000000",
  45852=>"100110100",
  45853=>"000000100",
  45854=>"000000000",
  45855=>"111001010",
  45856=>"100001000",
  45857=>"111001000",
  45858=>"111011001",
  45859=>"001000111",
  45860=>"000000000",
  45861=>"111111111",
  45862=>"000000101",
  45863=>"000001000",
  45864=>"011011010",
  45865=>"000000000",
  45866=>"000000000",
  45867=>"000000110",
  45868=>"000101111",
  45869=>"001110000",
  45870=>"011010010",
  45871=>"100000001",
  45872=>"001011111",
  45873=>"111111110",
  45874=>"100010000",
  45875=>"011011011",
  45876=>"000000000",
  45877=>"000000000",
  45878=>"001000000",
  45879=>"010010011",
  45880=>"100001100",
  45881=>"101000001",
  45882=>"111001000",
  45883=>"111111011",
  45884=>"110100110",
  45885=>"100100111",
  45886=>"000101111",
  45887=>"000110110",
  45888=>"111000111",
  45889=>"000001111",
  45890=>"100010111",
  45891=>"100111111",
  45892=>"000111111",
  45893=>"111111100",
  45894=>"011111111",
  45895=>"000000001",
  45896=>"000001011",
  45897=>"000110010",
  45898=>"001011010",
  45899=>"000000110",
  45900=>"111111111",
  45901=>"011011001",
  45902=>"100000110",
  45903=>"110111100",
  45904=>"111111111",
  45905=>"111000110",
  45906=>"001000000",
  45907=>"101001000",
  45908=>"000000000",
  45909=>"001011011",
  45910=>"000010111",
  45911=>"111111111",
  45912=>"000000001",
  45913=>"111010000",
  45914=>"011000000",
  45915=>"000000111",
  45916=>"000000100",
  45917=>"000111011",
  45918=>"111010010",
  45919=>"110111111",
  45920=>"111101111",
  45921=>"000000101",
  45922=>"111111111",
  45923=>"110100101",
  45924=>"111111111",
  45925=>"111000111",
  45926=>"000000000",
  45927=>"110100100",
  45928=>"100100111",
  45929=>"001011000",
  45930=>"000000000",
  45931=>"110100100",
  45932=>"100000000",
  45933=>"110100100",
  45934=>"000000111",
  45935=>"111110000",
  45936=>"011111111",
  45937=>"111111111",
  45938=>"011000010",
  45939=>"110110110",
  45940=>"000011001",
  45941=>"000000111",
  45942=>"010000100",
  45943=>"000001111",
  45944=>"000000001",
  45945=>"000000000",
  45946=>"000000000",
  45947=>"111111111",
  45948=>"111111111",
  45949=>"010111111",
  45950=>"101111000",
  45951=>"000000000",
  45952=>"000000101",
  45953=>"111111111",
  45954=>"000011011",
  45955=>"101000000",
  45956=>"000001111",
  45957=>"000000000",
  45958=>"000000000",
  45959=>"000001001",
  45960=>"000000001",
  45961=>"111111000",
  45962=>"000000100",
  45963=>"000101111",
  45964=>"111111111",
  45965=>"111111101",
  45966=>"100100111",
  45967=>"000000000",
  45968=>"000001111",
  45969=>"110110000",
  45970=>"001000000",
  45971=>"111011011",
  45972=>"000000000",
  45973=>"000000000",
  45974=>"111111110",
  45975=>"101011000",
  45976=>"001111111",
  45977=>"000000000",
  45978=>"000000100",
  45979=>"000111111",
  45980=>"100000000",
  45981=>"110010000",
  45982=>"110000000",
  45983=>"101100100",
  45984=>"111111111",
  45985=>"110111000",
  45986=>"111110111",
  45987=>"111111011",
  45988=>"100000100",
  45989=>"111111010",
  45990=>"000000011",
  45991=>"111101101",
  45992=>"000000000",
  45993=>"111110111",
  45994=>"000000100",
  45995=>"100000111",
  45996=>"001001001",
  45997=>"000001000",
  45998=>"000000001",
  45999=>"111111111",
  46000=>"001001000",
  46001=>"001000010",
  46002=>"111011011",
  46003=>"111000000",
  46004=>"000010000",
  46005=>"111111001",
  46006=>"111111110",
  46007=>"111111111",
  46008=>"111000000",
  46009=>"111111111",
  46010=>"000000000",
  46011=>"000110110",
  46012=>"000100111",
  46013=>"101101111",
  46014=>"000000111",
  46015=>"100101001",
  46016=>"111111000",
  46017=>"000000111",
  46018=>"111111101",
  46019=>"011010000",
  46020=>"100101111",
  46021=>"000000100",
  46022=>"101101111",
  46023=>"111101101",
  46024=>"111100111",
  46025=>"011111011",
  46026=>"100000000",
  46027=>"000000110",
  46028=>"111111111",
  46029=>"111001111",
  46030=>"000000001",
  46031=>"011000000",
  46032=>"000000000",
  46033=>"010011111",
  46034=>"111011011",
  46035=>"111111011",
  46036=>"110101101",
  46037=>"000111111",
  46038=>"111000011",
  46039=>"001011011",
  46040=>"100100110",
  46041=>"011000000",
  46042=>"000000000",
  46043=>"000001011",
  46044=>"000000000",
  46045=>"111111111",
  46046=>"111111111",
  46047=>"000100000",
  46048=>"010010000",
  46049=>"001001001",
  46050=>"000000111",
  46051=>"111111000",
  46052=>"111111111",
  46053=>"010111111",
  46054=>"110111000",
  46055=>"111111111",
  46056=>"111000110",
  46057=>"111000000",
  46058=>"000000000",
  46059=>"111111100",
  46060=>"000000000",
  46061=>"111100100",
  46062=>"000000000",
  46063=>"110000000",
  46064=>"000001101",
  46065=>"011011011",
  46066=>"000000010",
  46067=>"111100100",
  46068=>"000000000",
  46069=>"010110010",
  46070=>"000000000",
  46071=>"111110110",
  46072=>"010111000",
  46073=>"000010010",
  46074=>"011111111",
  46075=>"011000000",
  46076=>"111111101",
  46077=>"111111000",
  46078=>"111010010",
  46079=>"000000111",
  46080=>"000000000",
  46081=>"000000011",
  46082=>"111111010",
  46083=>"000000000",
  46084=>"000000000",
  46085=>"010110011",
  46086=>"101111111",
  46087=>"111111111",
  46088=>"100110111",
  46089=>"111000101",
  46090=>"111111111",
  46091=>"000110111",
  46092=>"111000000",
  46093=>"000000100",
  46094=>"000000000",
  46095=>"111011111",
  46096=>"000000000",
  46097=>"011001111",
  46098=>"111000000",
  46099=>"111111111",
  46100=>"111111111",
  46101=>"000000000",
  46102=>"111111101",
  46103=>"001001001",
  46104=>"111111110",
  46105=>"111000011",
  46106=>"000111111",
  46107=>"000111101",
  46108=>"111111111",
  46109=>"000000000",
  46110=>"000000100",
  46111=>"000000000",
  46112=>"111111111",
  46113=>"110111111",
  46114=>"111111111",
  46115=>"001000000",
  46116=>"100101111",
  46117=>"000000000",
  46118=>"000000000",
  46119=>"000001111",
  46120=>"110100010",
  46121=>"000000000",
  46122=>"000000000",
  46123=>"111111111",
  46124=>"111111111",
  46125=>"000011111",
  46126=>"001001111",
  46127=>"100000111",
  46128=>"001111011",
  46129=>"000000101",
  46130=>"000000001",
  46131=>"100110110",
  46132=>"000000000",
  46133=>"000011010",
  46134=>"111111111",
  46135=>"111111111",
  46136=>"000000111",
  46137=>"111111111",
  46138=>"000000000",
  46139=>"111001111",
  46140=>"111111011",
  46141=>"111000000",
  46142=>"000000011",
  46143=>"111100000",
  46144=>"101000000",
  46145=>"111111111",
  46146=>"111111111",
  46147=>"100000000",
  46148=>"111111100",
  46149=>"001001111",
  46150=>"000000110",
  46151=>"000001111",
  46152=>"001000001",
  46153=>"011111111",
  46154=>"100101111",
  46155=>"111001001",
  46156=>"000000111",
  46157=>"101001111",
  46158=>"110100100",
  46159=>"000000000",
  46160=>"111111111",
  46161=>"000000000",
  46162=>"110110110",
  46163=>"111111111",
  46164=>"111111111",
  46165=>"111000000",
  46166=>"100110000",
  46167=>"111111111",
  46168=>"001000101",
  46169=>"010000000",
  46170=>"000000100",
  46171=>"100000000",
  46172=>"111111111",
  46173=>"111100000",
  46174=>"000000000",
  46175=>"111100101",
  46176=>"111000000",
  46177=>"111111111",
  46178=>"111001011",
  46179=>"000000000",
  46180=>"001000100",
  46181=>"000000001",
  46182=>"100000000",
  46183=>"000000000",
  46184=>"000000000",
  46185=>"111111000",
  46186=>"100101001",
  46187=>"001001101",
  46188=>"000010110",
  46189=>"110111100",
  46190=>"111111111",
  46191=>"010000000",
  46192=>"111111111",
  46193=>"000111101",
  46194=>"111111111",
  46195=>"000000000",
  46196=>"111111111",
  46197=>"000001011",
  46198=>"101111111",
  46199=>"111111111",
  46200=>"011011111",
  46201=>"111111111",
  46202=>"000000001",
  46203=>"111111111",
  46204=>"100000100",
  46205=>"001001001",
  46206=>"110110100",
  46207=>"000000000",
  46208=>"111111111",
  46209=>"111111010",
  46210=>"000000000",
  46211=>"000101101",
  46212=>"111111111",
  46213=>"011011111",
  46214=>"000000001",
  46215=>"000000000",
  46216=>"000001000",
  46217=>"111111111",
  46218=>"000000000",
  46219=>"111111111",
  46220=>"111001011",
  46221=>"000000000",
  46222=>"110100000",
  46223=>"000000000",
  46224=>"000000001",
  46225=>"001011111",
  46226=>"000000000",
  46227=>"111000000",
  46228=>"111110111",
  46229=>"001000111",
  46230=>"000000000",
  46231=>"000000000",
  46232=>"111111000",
  46233=>"101111111",
  46234=>"011111111",
  46235=>"111100110",
  46236=>"111111111",
  46237=>"111000111",
  46238=>"000000100",
  46239=>"111000111",
  46240=>"111111111",
  46241=>"000000000",
  46242=>"111111110",
  46243=>"100001111",
  46244=>"111110110",
  46245=>"111111111",
  46246=>"000111111",
  46247=>"001001001",
  46248=>"111011000",
  46249=>"111111111",
  46250=>"111011011",
  46251=>"110111111",
  46252=>"111111001",
  46253=>"000000110",
  46254=>"011000000",
  46255=>"001000000",
  46256=>"111111000",
  46257=>"111101111",
  46258=>"010010000",
  46259=>"000000111",
  46260=>"111111101",
  46261=>"000000000",
  46262=>"000000010",
  46263=>"101000000",
  46264=>"111010011",
  46265=>"000011010",
  46266=>"000000010",
  46267=>"110000000",
  46268=>"000000000",
  46269=>"001001101",
  46270=>"100100100",
  46271=>"111111111",
  46272=>"000000000",
  46273=>"111101111",
  46274=>"111111111",
  46275=>"111111111",
  46276=>"000011000",
  46277=>"111111111",
  46278=>"111011000",
  46279=>"000000111",
  46280=>"001111010",
  46281=>"111001111",
  46282=>"100000100",
  46283=>"111111111",
  46284=>"111101101",
  46285=>"000000101",
  46286=>"000000111",
  46287=>"000000001",
  46288=>"000000000",
  46289=>"010111011",
  46290=>"101001111",
  46291=>"111001001",
  46292=>"000000000",
  46293=>"111111111",
  46294=>"000000100",
  46295=>"000000000",
  46296=>"000000000",
  46297=>"111100110",
  46298=>"110101000",
  46299=>"010100111",
  46300=>"010110110",
  46301=>"000100111",
  46302=>"111111111",
  46303=>"111111111",
  46304=>"000000000",
  46305=>"000011111",
  46306=>"000111110",
  46307=>"111100110",
  46308=>"000000100",
  46309=>"001001001",
  46310=>"000000110",
  46311=>"111111100",
  46312=>"101101111",
  46313=>"111111111",
  46314=>"110111111",
  46315=>"100100111",
  46316=>"111000000",
  46317=>"111111111",
  46318=>"000000000",
  46319=>"000000000",
  46320=>"111111111",
  46321=>"111100110",
  46322=>"011011111",
  46323=>"000000000",
  46324=>"111000100",
  46325=>"100000000",
  46326=>"111111000",
  46327=>"000000000",
  46328=>"111111111",
  46329=>"000000000",
  46330=>"110000000",
  46331=>"000000000",
  46332=>"000000000",
  46333=>"000010010",
  46334=>"111111000",
  46335=>"100100000",
  46336=>"111001000",
  46337=>"000000000",
  46338=>"000111111",
  46339=>"000000111",
  46340=>"111111111",
  46341=>"111000000",
  46342=>"101100000",
  46343=>"000000011",
  46344=>"100100111",
  46345=>"000000001",
  46346=>"000000000",
  46347=>"110111111",
  46348=>"111101010",
  46349=>"111111111",
  46350=>"111000000",
  46351=>"000000000",
  46352=>"110000111",
  46353=>"100111111",
  46354=>"000000001",
  46355=>"011110100",
  46356=>"001001000",
  46357=>"111111011",
  46358=>"000000000",
  46359=>"000000000",
  46360=>"111110100",
  46361=>"000000000",
  46362=>"000000000",
  46363=>"101111110",
  46364=>"011001011",
  46365=>"111000110",
  46366=>"000000000",
  46367=>"010000011",
  46368=>"000000011",
  46369=>"000001001",
  46370=>"111101111",
  46371=>"000000000",
  46372=>"000000000",
  46373=>"011011111",
  46374=>"000000000",
  46375=>"111000000",
  46376=>"000000111",
  46377=>"100000000",
  46378=>"000000000",
  46379=>"111111111",
  46380=>"001000000",
  46381=>"100000000",
  46382=>"111111111",
  46383=>"111110111",
  46384=>"111111011",
  46385=>"111101001",
  46386=>"111111111",
  46387=>"000000000",
  46388=>"111111111",
  46389=>"000000101",
  46390=>"111111111",
  46391=>"000000000",
  46392=>"000000000",
  46393=>"000000000",
  46394=>"000100111",
  46395=>"010110111",
  46396=>"111111111",
  46397=>"000000000",
  46398=>"000000000",
  46399=>"111111111",
  46400=>"010000000",
  46401=>"001000111",
  46402=>"000000101",
  46403=>"111000000",
  46404=>"111111111",
  46405=>"000000000",
  46406=>"111100111",
  46407=>"000000010",
  46408=>"100110111",
  46409=>"010110111",
  46410=>"000000001",
  46411=>"000000000",
  46412=>"101111000",
  46413=>"111111111",
  46414=>"110010000",
  46415=>"110101000",
  46416=>"111101100",
  46417=>"000000000",
  46418=>"011111111",
  46419=>"000000000",
  46420=>"000000000",
  46421=>"011111011",
  46422=>"110000000",
  46423=>"000000000",
  46424=>"000000000",
  46425=>"111111111",
  46426=>"000011111",
  46427=>"111001000",
  46428=>"110110000",
  46429=>"110110000",
  46430=>"000000001",
  46431=>"001011110",
  46432=>"111111111",
  46433=>"111000111",
  46434=>"000001011",
  46435=>"000010111",
  46436=>"000000000",
  46437=>"000100100",
  46438=>"111111111",
  46439=>"000000000",
  46440=>"000000000",
  46441=>"000000010",
  46442=>"000111111",
  46443=>"000000000",
  46444=>"000000000",
  46445=>"101101111",
  46446=>"000001001",
  46447=>"000000011",
  46448=>"100111111",
  46449=>"111111111",
  46450=>"111111111",
  46451=>"000000000",
  46452=>"000000000",
  46453=>"111111111",
  46454=>"000000000",
  46455=>"000000000",
  46456=>"111111111",
  46457=>"000111110",
  46458=>"000001000",
  46459=>"100100100",
  46460=>"111111110",
  46461=>"100000000",
  46462=>"010110110",
  46463=>"000000000",
  46464=>"001001001",
  46465=>"000000000",
  46466=>"000110110",
  46467=>"111111111",
  46468=>"111111111",
  46469=>"000000000",
  46470=>"111101101",
  46471=>"111110110",
  46472=>"111111111",
  46473=>"111111111",
  46474=>"100110011",
  46475=>"010010010",
  46476=>"111011011",
  46477=>"111001001",
  46478=>"101000000",
  46479=>"000000000",
  46480=>"111111111",
  46481=>"100000000",
  46482=>"111111111",
  46483=>"111111111",
  46484=>"000000000",
  46485=>"000001001",
  46486=>"001000000",
  46487=>"000011010",
  46488=>"001001000",
  46489=>"001111111",
  46490=>"101101111",
  46491=>"000000001",
  46492=>"111000000",
  46493=>"000000000",
  46494=>"000000000",
  46495=>"000011000",
  46496=>"110100000",
  46497=>"001011001",
  46498=>"111100000",
  46499=>"111111111",
  46500=>"111110000",
  46501=>"000010000",
  46502=>"110110000",
  46503=>"111111101",
  46504=>"111111111",
  46505=>"111001000",
  46506=>"111110110",
  46507=>"011011011",
  46508=>"000000000",
  46509=>"111110110",
  46510=>"000000001",
  46511=>"100100111",
  46512=>"000000001",
  46513=>"011000000",
  46514=>"000111110",
  46515=>"110110100",
  46516=>"111000100",
  46517=>"000000000",
  46518=>"101111000",
  46519=>"000100111",
  46520=>"000000000",
  46521=>"001000010",
  46522=>"111011000",
  46523=>"111100100",
  46524=>"001010000",
  46525=>"111111111",
  46526=>"000100100",
  46527=>"000000001",
  46528=>"110110111",
  46529=>"011111111",
  46530=>"111111111",
  46531=>"111111111",
  46532=>"000101001",
  46533=>"100100111",
  46534=>"111111011",
  46535=>"000000000",
  46536=>"111111110",
  46537=>"110111000",
  46538=>"000000000",
  46539=>"000000111",
  46540=>"000000000",
  46541=>"000000000",
  46542=>"000001001",
  46543=>"001101001",
  46544=>"000110110",
  46545=>"000100100",
  46546=>"000001011",
  46547=>"111111011",
  46548=>"110100000",
  46549=>"000000000",
  46550=>"110100110",
  46551=>"001000000",
  46552=>"000000001",
  46553=>"111000000",
  46554=>"111111111",
  46555=>"001011111",
  46556=>"001000001",
  46557=>"000000000",
  46558=>"001001011",
  46559=>"011001011",
  46560=>"010111110",
  46561=>"101111111",
  46562=>"010010000",
  46563=>"111100100",
  46564=>"000000001",
  46565=>"111111111",
  46566=>"110010000",
  46567=>"111111110",
  46568=>"000000000",
  46569=>"111011111",
  46570=>"000000000",
  46571=>"100111111",
  46572=>"111000011",
  46573=>"000000000",
  46574=>"111111111",
  46575=>"000100111",
  46576=>"000000001",
  46577=>"111000111",
  46578=>"000000001",
  46579=>"000110111",
  46580=>"000000000",
  46581=>"000000000",
  46582=>"011011011",
  46583=>"111001111",
  46584=>"000011111",
  46585=>"000100110",
  46586=>"001111111",
  46587=>"000000000",
  46588=>"000111000",
  46589=>"111110000",
  46590=>"110111111",
  46591=>"011011000",
  46592=>"001001101",
  46593=>"001110000",
  46594=>"000100111",
  46595=>"111111110",
  46596=>"111011011",
  46597=>"110000001",
  46598=>"000000000",
  46599=>"000000111",
  46600=>"111001001",
  46601=>"101101100",
  46602=>"111111111",
  46603=>"111010010",
  46604=>"110110110",
  46605=>"001000011",
  46606=>"110111111",
  46607=>"000000000",
  46608=>"000000000",
  46609=>"111111000",
  46610=>"111111100",
  46611=>"001001011",
  46612=>"000000000",
  46613=>"110111111",
  46614=>"111001110",
  46615=>"011001001",
  46616=>"001100010",
  46617=>"011111100",
  46618=>"000010000",
  46619=>"110110010",
  46620=>"111011010",
  46621=>"101000000",
  46622=>"011000000",
  46623=>"011011100",
  46624=>"100100100",
  46625=>"000000000",
  46626=>"111111111",
  46627=>"011111011",
  46628=>"111110000",
  46629=>"000001111",
  46630=>"111111111",
  46631=>"000011111",
  46632=>"101111110",
  46633=>"111111111",
  46634=>"111101001",
  46635=>"010000101",
  46636=>"000011011",
  46637=>"000011111",
  46638=>"100100000",
  46639=>"011011000",
  46640=>"011111111",
  46641=>"100100100",
  46642=>"011011011",
  46643=>"111101101",
  46644=>"000000111",
  46645=>"001001001",
  46646=>"111111111",
  46647=>"001001111",
  46648=>"000000000",
  46649=>"111010000",
  46650=>"000000000",
  46651=>"000000000",
  46652=>"100000111",
  46653=>"111111010",
  46654=>"010001110",
  46655=>"111111011",
  46656=>"110110010",
  46657=>"111111111",
  46658=>"000010111",
  46659=>"110011110",
  46660=>"110110110",
  46661=>"000100110",
  46662=>"111110010",
  46663=>"000111011",
  46664=>"000000001",
  46665=>"000000000",
  46666=>"111111111",
  46667=>"000000110",
  46668=>"010000000",
  46669=>"001110001",
  46670=>"000000001",
  46671=>"111111111",
  46672=>"111000000",
  46673=>"111111101",
  46674=>"000000011",
  46675=>"001001101",
  46676=>"111111111",
  46677=>"011111010",
  46678=>"001000011",
  46679=>"111111111",
  46680=>"001110100",
  46681=>"000000000",
  46682=>"000000111",
  46683=>"000001001",
  46684=>"000000000",
  46685=>"000000100",
  46686=>"111100110",
  46687=>"110100110",
  46688=>"111111101",
  46689=>"011011001",
  46690=>"111000010",
  46691=>"111111111",
  46692=>"111111100",
  46693=>"000000000",
  46694=>"111111011",
  46695=>"110110000",
  46696=>"000000000",
  46697=>"111111111",
  46698=>"110100111",
  46699=>"111111111",
  46700=>"000111111",
  46701=>"000000000",
  46702=>"000000100",
  46703=>"101111111",
  46704=>"111111111",
  46705=>"010010110",
  46706=>"000000000",
  46707=>"110111111",
  46708=>"000000000",
  46709=>"111111110",
  46710=>"000000000",
  46711=>"110111010",
  46712=>"111000100",
  46713=>"000000000",
  46714=>"100100000",
  46715=>"111000000",
  46716=>"111111000",
  46717=>"000010111",
  46718=>"111000011",
  46719=>"111111111",
  46720=>"000100000",
  46721=>"001000000",
  46722=>"000100111",
  46723=>"100100110",
  46724=>"111111110",
  46725=>"111000000",
  46726=>"011000111",
  46727=>"000000000",
  46728=>"111101000",
  46729=>"110110110",
  46730=>"111100000",
  46731=>"111111000",
  46732=>"100100111",
  46733=>"011011000",
  46734=>"000000000",
  46735=>"000000000",
  46736=>"111011111",
  46737=>"111111111",
  46738=>"010010111",
  46739=>"000000011",
  46740=>"111111011",
  46741=>"111111111",
  46742=>"111110111",
  46743=>"000000000",
  46744=>"111101111",
  46745=>"101000000",
  46746=>"111111110",
  46747=>"000000011",
  46748=>"111111111",
  46749=>"110000000",
  46750=>"011000110",
  46751=>"000000000",
  46752=>"000000110",
  46753=>"000001011",
  46754=>"011111111",
  46755=>"111000000",
  46756=>"001001000",
  46757=>"101000010",
  46758=>"111111111",
  46759=>"000000111",
  46760=>"111001011",
  46761=>"111001000",
  46762=>"001000000",
  46763=>"111111111",
  46764=>"100110111",
  46765=>"010010011",
  46766=>"000000000",
  46767=>"111001000",
  46768=>"011000000",
  46769=>"000000000",
  46770=>"111111011",
  46771=>"111000111",
  46772=>"100000000",
  46773=>"101000000",
  46774=>"111111111",
  46775=>"111111001",
  46776=>"110100111",
  46777=>"000000000",
  46778=>"001000000",
  46779=>"001001111",
  46780=>"010000000",
  46781=>"111111111",
  46782=>"011000000",
  46783=>"100000000",
  46784=>"000000000",
  46785=>"011001000",
  46786=>"111000000",
  46787=>"111000000",
  46788=>"000000000",
  46789=>"111111111",
  46790=>"000000100",
  46791=>"100110111",
  46792=>"111000000",
  46793=>"111000000",
  46794=>"001000110",
  46795=>"111111111",
  46796=>"000010111",
  46797=>"001100100",
  46798=>"100110111",
  46799=>"101111000",
  46800=>"000100111",
  46801=>"100000100",
  46802=>"111111111",
  46803=>"000000000",
  46804=>"000111111",
  46805=>"000101001",
  46806=>"000000000",
  46807=>"011111111",
  46808=>"110111110",
  46809=>"111111110",
  46810=>"111111111",
  46811=>"011010010",
  46812=>"000000000",
  46813=>"001001001",
  46814=>"110010010",
  46815=>"000000110",
  46816=>"111111011",
  46817=>"101000000",
  46818=>"000000000",
  46819=>"001000110",
  46820=>"111111111",
  46821=>"000100111",
  46822=>"111000000",
  46823=>"000000000",
  46824=>"000000000",
  46825=>"111111011",
  46826=>"111111111",
  46827=>"110010111",
  46828=>"110110000",
  46829=>"110111100",
  46830=>"111100100",
  46831=>"111110110",
  46832=>"111111000",
  46833=>"000000111",
  46834=>"111101111",
  46835=>"111111010",
  46836=>"100111111",
  46837=>"000001001",
  46838=>"111111100",
  46839=>"111010000",
  46840=>"000111111",
  46841=>"000000000",
  46842=>"110100111",
  46843=>"010000000",
  46844=>"001000000",
  46845=>"100010111",
  46846=>"001001000",
  46847=>"111111111",
  46848=>"100100100",
  46849=>"111000000",
  46850=>"000000000",
  46851=>"000011111",
  46852=>"111111111",
  46853=>"111111111",
  46854=>"000000000",
  46855=>"110110111",
  46856=>"111111111",
  46857=>"111000000",
  46858=>"111000000",
  46859=>"000000110",
  46860=>"111111011",
  46861=>"111111111",
  46862=>"110111110",
  46863=>"000000011",
  46864=>"000000000",
  46865=>"110111111",
  46866=>"000001110",
  46867=>"000000000",
  46868=>"001101111",
  46869=>"000000111",
  46870=>"001011001",
  46871=>"101101000",
  46872=>"001001000",
  46873=>"100000000",
  46874=>"000000111",
  46875=>"111111111",
  46876=>"100110110",
  46877=>"000010011",
  46878=>"111111111",
  46879=>"110000111",
  46880=>"000000111",
  46881=>"111111111",
  46882=>"110110110",
  46883=>"101101011",
  46884=>"000100000",
  46885=>"001001001",
  46886=>"111110100",
  46887=>"111111000",
  46888=>"000000000",
  46889=>"000000000",
  46890=>"000000000",
  46891=>"111111111",
  46892=>"111111111",
  46893=>"010110000",
  46894=>"000000000",
  46895=>"000000000",
  46896=>"011011000",
  46897=>"111111111",
  46898=>"000001011",
  46899=>"011000111",
  46900=>"101001000",
  46901=>"110110110",
  46902=>"111111111",
  46903=>"101111111",
  46904=>"000000100",
  46905=>"000000000",
  46906=>"000000000",
  46907=>"000110110",
  46908=>"110111111",
  46909=>"111111111",
  46910=>"111000001",
  46911=>"000000000",
  46912=>"111000101",
  46913=>"011001111",
  46914=>"101101111",
  46915=>"000000000",
  46916=>"100000000",
  46917=>"000000110",
  46918=>"101111111",
  46919=>"001000111",
  46920=>"111111111",
  46921=>"000100100",
  46922=>"111111111",
  46923=>"111110110",
  46924=>"111111111",
  46925=>"110110111",
  46926=>"101110110",
  46927=>"000001001",
  46928=>"000000110",
  46929=>"000000110",
  46930=>"111111111",
  46931=>"101111111",
  46932=>"000000100",
  46933=>"000000100",
  46934=>"111111111",
  46935=>"000000000",
  46936=>"111111111",
  46937=>"111011011",
  46938=>"000000001",
  46939=>"100100100",
  46940=>"000000010",
  46941=>"000000000",
  46942=>"000000000",
  46943=>"111110111",
  46944=>"111011111",
  46945=>"111111111",
  46946=>"111000000",
  46947=>"111111111",
  46948=>"000000110",
  46949=>"111111111",
  46950=>"000001001",
  46951=>"000100000",
  46952=>"001000000",
  46953=>"111111011",
  46954=>"111100000",
  46955=>"111111110",
  46956=>"011001001",
  46957=>"000000100",
  46958=>"000000000",
  46959=>"111111111",
  46960=>"000000000",
  46961=>"111111111",
  46962=>"001000000",
  46963=>"101110110",
  46964=>"111100100",
  46965=>"111111111",
  46966=>"000000111",
  46967=>"011001001",
  46968=>"111111111",
  46969=>"110110110",
  46970=>"000000000",
  46971=>"101011011",
  46972=>"111111111",
  46973=>"011011000",
  46974=>"000100110",
  46975=>"111111111",
  46976=>"001011011",
  46977=>"001111111",
  46978=>"001011011",
  46979=>"000000000",
  46980=>"111111000",
  46981=>"000000101",
  46982=>"100000111",
  46983=>"100000000",
  46984=>"000000000",
  46985=>"111111100",
  46986=>"111110000",
  46987=>"111111111",
  46988=>"000000000",
  46989=>"000000000",
  46990=>"011111111",
  46991=>"111101101",
  46992=>"101110110",
  46993=>"111111110",
  46994=>"011010000",
  46995=>"001011011",
  46996=>"000000000",
  46997=>"000000000",
  46998=>"101111111",
  46999=>"011001111",
  47000=>"010000100",
  47001=>"101110111",
  47002=>"111111110",
  47003=>"111111110",
  47004=>"111111111",
  47005=>"111111110",
  47006=>"101111111",
  47007=>"110001011",
  47008=>"111110110",
  47009=>"010010000",
  47010=>"000000110",
  47011=>"111111111",
  47012=>"001001111",
  47013=>"000000000",
  47014=>"000000000",
  47015=>"000000110",
  47016=>"111110000",
  47017=>"000100111",
  47018=>"000110111",
  47019=>"000000011",
  47020=>"100100100",
  47021=>"000000000",
  47022=>"100000000",
  47023=>"110000110",
  47024=>"111111010",
  47025=>"010000000",
  47026=>"111001001",
  47027=>"111111111",
  47028=>"111111111",
  47029=>"101101111",
  47030=>"111000000",
  47031=>"001000000",
  47032=>"011011110",
  47033=>"000010010",
  47034=>"100111111",
  47035=>"111000000",
  47036=>"000111110",
  47037=>"111111111",
  47038=>"111111111",
  47039=>"011111111",
  47040=>"111111111",
  47041=>"000000101",
  47042=>"000000101",
  47043=>"111100000",
  47044=>"111001111",
  47045=>"111111111",
  47046=>"111110110",
  47047=>"111111110",
  47048=>"100100111",
  47049=>"001011111",
  47050=>"100100110",
  47051=>"000000110",
  47052=>"000010111",
  47053=>"000000000",
  47054=>"110110110",
  47055=>"000000000",
  47056=>"111001001",
  47057=>"111111111",
  47058=>"000001000",
  47059=>"000111111",
  47060=>"000000000",
  47061=>"111111111",
  47062=>"000000000",
  47063=>"111111111",
  47064=>"000000000",
  47065=>"111001111",
  47066=>"111111001",
  47067=>"111111010",
  47068=>"000001011",
  47069=>"111111011",
  47070=>"000100111",
  47071=>"001000000",
  47072=>"110110110",
  47073=>"111111111",
  47074=>"111111100",
  47075=>"001110110",
  47076=>"111001000",
  47077=>"110110111",
  47078=>"110110000",
  47079=>"100100111",
  47080=>"111111111",
  47081=>"111111001",
  47082=>"111111000",
  47083=>"110000011",
  47084=>"110101111",
  47085=>"000000100",
  47086=>"000000000",
  47087=>"101000000",
  47088=>"100111111",
  47089=>"000000000",
  47090=>"000000000",
  47091=>"111110110",
  47092=>"011110000",
  47093=>"111111111",
  47094=>"110100000",
  47095=>"000100100",
  47096=>"111001000",
  47097=>"100110011",
  47098=>"111111111",
  47099=>"110110111",
  47100=>"110111111",
  47101=>"001001000",
  47102=>"000000000",
  47103=>"001000000",
  47104=>"111111111",
  47105=>"111010111",
  47106=>"001000001",
  47107=>"101001001",
  47108=>"011011001",
  47109=>"011011011",
  47110=>"001000001",
  47111=>"110100111",
  47112=>"110111111",
  47113=>"111010000",
  47114=>"111111111",
  47115=>"101001101",
  47116=>"001000000",
  47117=>"010011000",
  47118=>"100000000",
  47119=>"111111111",
  47120=>"000111110",
  47121=>"111010011",
  47122=>"001000000",
  47123=>"000111111",
  47124=>"000000000",
  47125=>"110111111",
  47126=>"111101111",
  47127=>"001000000",
  47128=>"111111011",
  47129=>"101001001",
  47130=>"000000111",
  47131=>"101000000",
  47132=>"111111111",
  47133=>"111111111",
  47134=>"100010000",
  47135=>"111111110",
  47136=>"101100100",
  47137=>"111111001",
  47138=>"100111000",
  47139=>"111001001",
  47140=>"010000010",
  47141=>"111010001",
  47142=>"001001001",
  47143=>"001111111",
  47144=>"100000010",
  47145=>"000000111",
  47146=>"001001101",
  47147=>"000011010",
  47148=>"000000111",
  47149=>"101100000",
  47150=>"001010011",
  47151=>"011000000",
  47152=>"111111110",
  47153=>"101101101",
  47154=>"100100000",
  47155=>"000100000",
  47156=>"100100101",
  47157=>"111101001",
  47158=>"000111111",
  47159=>"111111001",
  47160=>"110111000",
  47161=>"000010010",
  47162=>"000000000",
  47163=>"110000100",
  47164=>"000000101",
  47165=>"001111111",
  47166=>"100100111",
  47167=>"111111111",
  47168=>"011111010",
  47169=>"000010010",
  47170=>"010000110",
  47171=>"001011110",
  47172=>"001111001",
  47173=>"001100100",
  47174=>"001000000",
  47175=>"111100111",
  47176=>"011011111",
  47177=>"110000101",
  47178=>"110111111",
  47179=>"011011001",
  47180=>"001000110",
  47181=>"100000000",
  47182=>"011001000",
  47183=>"000000111",
  47184=>"000000000",
  47185=>"111111000",
  47186=>"000001111",
  47187=>"001001000",
  47188=>"101101101",
  47189=>"000110111",
  47190=>"000100100",
  47191=>"001001000",
  47192=>"000000000",
  47193=>"000000111",
  47194=>"010111101",
  47195=>"000100100",
  47196=>"000000000",
  47197=>"110111111",
  47198=>"000000000",
  47199=>"010111111",
  47200=>"001000000",
  47201=>"000010011",
  47202=>"001001101",
  47203=>"111000000",
  47204=>"101000000",
  47205=>"000111111",
  47206=>"111111001",
  47207=>"000000111",
  47208=>"000000100",
  47209=>"111110110",
  47210=>"010111111",
  47211=>"000000000",
  47212=>"011001001",
  47213=>"000001001",
  47214=>"000000000",
  47215=>"111110000",
  47216=>"000000011",
  47217=>"110110001",
  47218=>"000000110",
  47219=>"111111111",
  47220=>"101101111",
  47221=>"010110100",
  47222=>"111111111",
  47223=>"000000000",
  47224=>"000000001",
  47225=>"111111111",
  47226=>"001000100",
  47227=>"000000000",
  47228=>"011011001",
  47229=>"101001001",
  47230=>"000000000",
  47231=>"000000001",
  47232=>"110000000",
  47233=>"001000000",
  47234=>"000000000",
  47235=>"000000100",
  47236=>"000111100",
  47237=>"111111111",
  47238=>"111111110",
  47239=>"111001000",
  47240=>"000010010",
  47241=>"000110110",
  47242=>"100000000",
  47243=>"000000000",
  47244=>"010110111",
  47245=>"011111111",
  47246=>"101101101",
  47247=>"000101101",
  47248=>"111000111",
  47249=>"111001111",
  47250=>"110011010",
  47251=>"000001001",
  47252=>"111011000",
  47253=>"101100100",
  47254=>"000000100",
  47255=>"000000000",
  47256=>"100100000",
  47257=>"010000110",
  47258=>"000111100",
  47259=>"010111110",
  47260=>"100100100",
  47261=>"100110111",
  47262=>"100100000",
  47263=>"000111101",
  47264=>"000000000",
  47265=>"111111010",
  47266=>"000111110",
  47267=>"000111111",
  47268=>"011001101",
  47269=>"000000000",
  47270=>"001111111",
  47271=>"100100100",
  47272=>"000011110",
  47273=>"000010111",
  47274=>"000010111",
  47275=>"101111111",
  47276=>"010000000",
  47277=>"110110110",
  47278=>"110100110",
  47279=>"000000000",
  47280=>"000000000",
  47281=>"000000100",
  47282=>"111111111",
  47283=>"100100000",
  47284=>"010000000",
  47285=>"111111000",
  47286=>"111001000",
  47287=>"110110111",
  47288=>"110000000",
  47289=>"111011011",
  47290=>"111000101",
  47291=>"111000111",
  47292=>"000000000",
  47293=>"001110111",
  47294=>"000111111",
  47295=>"000111111",
  47296=>"111100100",
  47297=>"000001000",
  47298=>"111111011",
  47299=>"000111111",
  47300=>"110111111",
  47301=>"000000000",
  47302=>"001111001",
  47303=>"111111111",
  47304=>"000111111",
  47305=>"000111111",
  47306=>"000000000",
  47307=>"111111001",
  47308=>"100111000",
  47309=>"000001000",
  47310=>"000000111",
  47311=>"111000000",
  47312=>"111011000",
  47313=>"101001001",
  47314=>"010000010",
  47315=>"000000000",
  47316=>"111111101",
  47317=>"000000000",
  47318=>"111010010",
  47319=>"000000111",
  47320=>"001000010",
  47321=>"111111000",
  47322=>"000000000",
  47323=>"000010111",
  47324=>"111101000",
  47325=>"001111111",
  47326=>"000111000",
  47327=>"111111000",
  47328=>"100101111",
  47329=>"110000000",
  47330=>"000000000",
  47331=>"110111111",
  47332=>"000000001",
  47333=>"001001011",
  47334=>"000010010",
  47335=>"000101000",
  47336=>"000000011",
  47337=>"001101111",
  47338=>"001100100",
  47339=>"111000110",
  47340=>"110010000",
  47341=>"000000000",
  47342=>"111001000",
  47343=>"111000000",
  47344=>"001000000",
  47345=>"000000000",
  47346=>"000010110",
  47347=>"000100111",
  47348=>"001000010",
  47349=>"100111110",
  47350=>"101111111",
  47351=>"110110111",
  47352=>"111000001",
  47353=>"000100000",
  47354=>"100111111",
  47355=>"111111000",
  47356=>"100101101",
  47357=>"000000001",
  47358=>"110011001",
  47359=>"000000001",
  47360=>"110110110",
  47361=>"000000100",
  47362=>"001101000",
  47363=>"111111111",
  47364=>"000111111",
  47365=>"111111001",
  47366=>"110111110",
  47367=>"111001010",
  47368=>"000000000",
  47369=>"101111111",
  47370=>"000000000",
  47371=>"000101000",
  47372=>"101001001",
  47373=>"111010010",
  47374=>"111111011",
  47375=>"101001001",
  47376=>"000000011",
  47377=>"101101111",
  47378=>"000000000",
  47379=>"000000000",
  47380=>"000110110",
  47381=>"000110111",
  47382=>"111111111",
  47383=>"000000110",
  47384=>"000011001",
  47385=>"111111000",
  47386=>"011001000",
  47387=>"011111111",
  47388=>"100110110",
  47389=>"110111111",
  47390=>"000111010",
  47391=>"111000000",
  47392=>"111011011",
  47393=>"110111111",
  47394=>"010010011",
  47395=>"010000111",
  47396=>"000000000",
  47397=>"101100100",
  47398=>"111101100",
  47399=>"111000011",
  47400=>"000000000",
  47401=>"111111111",
  47402=>"111111110",
  47403=>"111010111",
  47404=>"111111000",
  47405=>"000011011",
  47406=>"011000111",
  47407=>"000000110",
  47408=>"001111111",
  47409=>"101101101",
  47410=>"111001000",
  47411=>"111010000",
  47412=>"010010000",
  47413=>"111111000",
  47414=>"000000000",
  47415=>"011000111",
  47416=>"000100101",
  47417=>"000001111",
  47418=>"001000011",
  47419=>"111111000",
  47420=>"100001001",
  47421=>"000000111",
  47422=>"011001000",
  47423=>"111100111",
  47424=>"000010000",
  47425=>"111001001",
  47426=>"101111111",
  47427=>"101000000",
  47428=>"111111111",
  47429=>"000000111",
  47430=>"001000111",
  47431=>"001000111",
  47432=>"000000001",
  47433=>"011010010",
  47434=>"000000010",
  47435=>"000001001",
  47436=>"011111000",
  47437=>"010000000",
  47438=>"000000000",
  47439=>"000000001",
  47440=>"001111111",
  47441=>"000000011",
  47442=>"000110111",
  47443=>"111101000",
  47444=>"010111111",
  47445=>"011011011",
  47446=>"111111010",
  47447=>"011111111",
  47448=>"100000101",
  47449=>"000000111",
  47450=>"111111111",
  47451=>"000110011",
  47452=>"000111111",
  47453=>"111111101",
  47454=>"000000011",
  47455=>"000101111",
  47456=>"000000000",
  47457=>"000011111",
  47458=>"111101111",
  47459=>"001000000",
  47460=>"000100000",
  47461=>"011000000",
  47462=>"110000000",
  47463=>"001000011",
  47464=>"000000000",
  47465=>"000101111",
  47466=>"000000000",
  47467=>"000001011",
  47468=>"001001001",
  47469=>"000000110",
  47470=>"111100000",
  47471=>"000000000",
  47472=>"111011000",
  47473=>"011001001",
  47474=>"111000000",
  47475=>"110111101",
  47476=>"000001001",
  47477=>"001000100",
  47478=>"100100111",
  47479=>"010000100",
  47480=>"010110110",
  47481=>"011111111",
  47482=>"000000000",
  47483=>"001000000",
  47484=>"000010111",
  47485=>"000001111",
  47486=>"111010111",
  47487=>"000100100",
  47488=>"111000000",
  47489=>"011111111",
  47490=>"000001001",
  47491=>"011111111",
  47492=>"000011000",
  47493=>"110000110",
  47494=>"000000010",
  47495=>"000000110",
  47496=>"111001111",
  47497=>"101101111",
  47498=>"011110110",
  47499=>"000010110",
  47500=>"110011111",
  47501=>"100100000",
  47502=>"110000000",
  47503=>"000000000",
  47504=>"000111111",
  47505=>"001111011",
  47506=>"010000000",
  47507=>"001000000",
  47508=>"111000111",
  47509=>"111010000",
  47510=>"100001001",
  47511=>"100001011",
  47512=>"000000111",
  47513=>"000010010",
  47514=>"000000001",
  47515=>"100100100",
  47516=>"000111111",
  47517=>"010111110",
  47518=>"111011011",
  47519=>"000111111",
  47520=>"001101111",
  47521=>"011111111",
  47522=>"111101001",
  47523=>"000000000",
  47524=>"000001111",
  47525=>"111111111",
  47526=>"001000011",
  47527=>"111111011",
  47528=>"000000000",
  47529=>"000111101",
  47530=>"110101000",
  47531=>"111010000",
  47532=>"010111011",
  47533=>"111011111",
  47534=>"110110110",
  47535=>"100110000",
  47536=>"011000000",
  47537=>"111001111",
  47538=>"111111100",
  47539=>"011101101",
  47540=>"111000100",
  47541=>"101110111",
  47542=>"000000111",
  47543=>"001000000",
  47544=>"111011011",
  47545=>"111111111",
  47546=>"101101001",
  47547=>"100000001",
  47548=>"000000000",
  47549=>"001011111",
  47550=>"111101000",
  47551=>"110110100",
  47552=>"111111111",
  47553=>"000000001",
  47554=>"111111111",
  47555=>"000000010",
  47556=>"110100100",
  47557=>"111011111",
  47558=>"000000000",
  47559=>"010000000",
  47560=>"100111010",
  47561=>"000000111",
  47562=>"000000100",
  47563=>"000010111",
  47564=>"000010100",
  47565=>"000111100",
  47566=>"110010010",
  47567=>"000000000",
  47568=>"000110010",
  47569=>"000111001",
  47570=>"000000000",
  47571=>"011011001",
  47572=>"011111111",
  47573=>"000000100",
  47574=>"000000000",
  47575=>"110000000",
  47576=>"000000101",
  47577=>"000111111",
  47578=>"111111111",
  47579=>"111111111",
  47580=>"100000000",
  47581=>"000001111",
  47582=>"111111000",
  47583=>"110000010",
  47584=>"100000010",
  47585=>"011000111",
  47586=>"111101111",
  47587=>"111100000",
  47588=>"010010010",
  47589=>"010111111",
  47590=>"011011110",
  47591=>"000000000",
  47592=>"111100110",
  47593=>"111111110",
  47594=>"000110111",
  47595=>"111111111",
  47596=>"000110110",
  47597=>"000110010",
  47598=>"100100101",
  47599=>"111001001",
  47600=>"111000101",
  47601=>"111000100",
  47602=>"001011011",
  47603=>"000000001",
  47604=>"000000000",
  47605=>"011001000",
  47606=>"101000001",
  47607=>"110110100",
  47608=>"110110110",
  47609=>"001000000",
  47610=>"001001001",
  47611=>"000000111",
  47612=>"111111111",
  47613=>"011111110",
  47614=>"010011111",
  47615=>"111000000",
  47616=>"011011001",
  47617=>"101000000",
  47618=>"000100111",
  47619=>"000000000",
  47620=>"000000000",
  47621=>"111011111",
  47622=>"000000000",
  47623=>"111111111",
  47624=>"111101000",
  47625=>"000000111",
  47626=>"111111111",
  47627=>"000000000",
  47628=>"111111010",
  47629=>"100110111",
  47630=>"110000001",
  47631=>"000000000",
  47632=>"111010000",
  47633=>"000000000",
  47634=>"000010111",
  47635=>"011000111",
  47636=>"111000101",
  47637=>"000000111",
  47638=>"110111011",
  47639=>"000000011",
  47640=>"000000001",
  47641=>"100100000",
  47642=>"000000010",
  47643=>"010000101",
  47644=>"111100000",
  47645=>"000000111",
  47646=>"000100101",
  47647=>"110111111",
  47648=>"010011001",
  47649=>"111011111",
  47650=>"110110111",
  47651=>"111111111",
  47652=>"001000000",
  47653=>"001010010",
  47654=>"110000101",
  47655=>"111111000",
  47656=>"111000000",
  47657=>"111111010",
  47658=>"000000000",
  47659=>"101000000",
  47660=>"111111111",
  47661=>"011111000",
  47662=>"001111110",
  47663=>"001000000",
  47664=>"000100111",
  47665=>"000111111",
  47666=>"111100100",
  47667=>"111111011",
  47668=>"000111110",
  47669=>"100111110",
  47670=>"011001000",
  47671=>"000110110",
  47672=>"110000001",
  47673=>"110000001",
  47674=>"000000000",
  47675=>"000101100",
  47676=>"111111000",
  47677=>"011011000",
  47678=>"010100110",
  47679=>"100100111",
  47680=>"010111111",
  47681=>"011001000",
  47682=>"111110000",
  47683=>"111111000",
  47684=>"000101111",
  47685=>"100110100",
  47686=>"111111000",
  47687=>"000011000",
  47688=>"000000001",
  47689=>"000000000",
  47690=>"111111111",
  47691=>"110000110",
  47692=>"000111111",
  47693=>"000000001",
  47694=>"111111111",
  47695=>"110000000",
  47696=>"000000110",
  47697=>"000011111",
  47698=>"111110111",
  47699=>"111001111",
  47700=>"100100000",
  47701=>"000000000",
  47702=>"000000001",
  47703=>"110111000",
  47704=>"000000000",
  47705=>"111111111",
  47706=>"001001000",
  47707=>"010000000",
  47708=>"000000000",
  47709=>"000001111",
  47710=>"111100000",
  47711=>"100000000",
  47712=>"110111111",
  47713=>"010010110",
  47714=>"000000000",
  47715=>"000000000",
  47716=>"000000001",
  47717=>"000000000",
  47718=>"110111111",
  47719=>"000000111",
  47720=>"111000000",
  47721=>"111101100",
  47722=>"111010000",
  47723=>"000001001",
  47724=>"011011111",
  47725=>"000000100",
  47726=>"011000001",
  47727=>"100101000",
  47728=>"100000110",
  47729=>"110110000",
  47730=>"101111000",
  47731=>"000111111",
  47732=>"110111001",
  47733=>"010110110",
  47734=>"000000000",
  47735=>"100110110",
  47736=>"000000111",
  47737=>"010111111",
  47738=>"100110101",
  47739=>"110111111",
  47740=>"010110111",
  47741=>"000000111",
  47742=>"010111110",
  47743=>"100111111",
  47744=>"111111111",
  47745=>"110110000",
  47746=>"111000000",
  47747=>"111000010",
  47748=>"111011011",
  47749=>"111111000",
  47750=>"111110010",
  47751=>"000000000",
  47752=>"001111111",
  47753=>"111011011",
  47754=>"100011111",
  47755=>"111111000",
  47756=>"000000000",
  47757=>"110000010",
  47758=>"110100100",
  47759=>"000110000",
  47760=>"000111111",
  47761=>"000000000",
  47762=>"110000110",
  47763=>"000000000",
  47764=>"000000000",
  47765=>"000000111",
  47766=>"111101111",
  47767=>"111001111",
  47768=>"111001110",
  47769=>"111000111",
  47770=>"000000000",
  47771=>"000101101",
  47772=>"111000000",
  47773=>"100110110",
  47774=>"111111000",
  47775=>"000110000",
  47776=>"111111000",
  47777=>"111111000",
  47778=>"000000000",
  47779=>"001000111",
  47780=>"100001001",
  47781=>"100000111",
  47782=>"000111000",
  47783=>"000011111",
  47784=>"110111000",
  47785=>"000111111",
  47786=>"111101111",
  47787=>"000110111",
  47788=>"110000000",
  47789=>"100001001",
  47790=>"111111111",
  47791=>"000000010",
  47792=>"101000000",
  47793=>"000010110",
  47794=>"111111011",
  47795=>"011000000",
  47796=>"111000000",
  47797=>"110111111",
  47798=>"110111000",
  47799=>"111111000",
  47800=>"111111111",
  47801=>"000111000",
  47802=>"110110110",
  47803=>"110000001",
  47804=>"100000001",
  47805=>"110111000",
  47806=>"111111111",
  47807=>"011010000",
  47808=>"111000001",
  47809=>"000000100",
  47810=>"000000100",
  47811=>"111001000",
  47812=>"111111111",
  47813=>"111110000",
  47814=>"010111111",
  47815=>"110111000",
  47816=>"001110000",
  47817=>"111000000",
  47818=>"111110000",
  47819=>"111111001",
  47820=>"100000111",
  47821=>"000100000",
  47822=>"000000000",
  47823=>"110010000",
  47824=>"111001000",
  47825=>"000000000",
  47826=>"100110000",
  47827=>"111110000",
  47828=>"110100010",
  47829=>"111001000",
  47830=>"000001000",
  47831=>"000100111",
  47832=>"001000010",
  47833=>"111111111",
  47834=>"000000000",
  47835=>"110000000",
  47836=>"110011000",
  47837=>"111000000",
  47838=>"011111111",
  47839=>"110000001",
  47840=>"011000000",
  47841=>"111111000",
  47842=>"000000101",
  47843=>"110000101",
  47844=>"000000110",
  47845=>"111001001",
  47846=>"000000000",
  47847=>"110110111",
  47848=>"111000000",
  47849=>"000001101",
  47850=>"111110111",
  47851=>"100000000",
  47852=>"100111111",
  47853=>"011001111",
  47854=>"110000000",
  47855=>"000000000",
  47856=>"000010100",
  47857=>"000000111",
  47858=>"001001001",
  47859=>"110010000",
  47860=>"111000000",
  47861=>"011001001",
  47862=>"100100101",
  47863=>"111101100",
  47864=>"011000000",
  47865=>"111111000",
  47866=>"000000100",
  47867=>"111101000",
  47868=>"000000100",
  47869=>"111000101",
  47870=>"111011110",
  47871=>"000000000",
  47872=>"000000100",
  47873=>"110110000",
  47874=>"111100000",
  47875=>"110001001",
  47876=>"000000111",
  47877=>"101110111",
  47878=>"110111111",
  47879=>"111010000",
  47880=>"000000000",
  47881=>"000100000",
  47882=>"000000000",
  47883=>"110000000",
  47884=>"111011111",
  47885=>"111110110",
  47886=>"100100000",
  47887=>"000100100",
  47888=>"000010110",
  47889=>"110000000",
  47890=>"000000111",
  47891=>"111000000",
  47892=>"011111111",
  47893=>"111001000",
  47894=>"101111111",
  47895=>"000001000",
  47896=>"000110110",
  47897=>"011000101",
  47898=>"111110111",
  47899=>"010010000",
  47900=>"100000110",
  47901=>"111111011",
  47902=>"000011111",
  47903=>"000000000",
  47904=>"000001001",
  47905=>"000000111",
  47906=>"010011111",
  47907=>"100110111",
  47908=>"111011000",
  47909=>"011010000",
  47910=>"111011010",
  47911=>"010001000",
  47912=>"001001000",
  47913=>"010111000",
  47914=>"000000000",
  47915=>"011011101",
  47916=>"111000000",
  47917=>"000110111",
  47918=>"000000010",
  47919=>"110000000",
  47920=>"000111111",
  47921=>"010000000",
  47922=>"000010010",
  47923=>"001100111",
  47924=>"111101110",
  47925=>"111101000",
  47926=>"101111111",
  47927=>"111111011",
  47928=>"111000000",
  47929=>"111000000",
  47930=>"111000000",
  47931=>"000101111",
  47932=>"100000001",
  47933=>"110010011",
  47934=>"111110111",
  47935=>"111110000",
  47936=>"110000000",
  47937=>"000110100",
  47938=>"110010111",
  47939=>"101111110",
  47940=>"111111111",
  47941=>"000000000",
  47942=>"100110000",
  47943=>"111111000",
  47944=>"111010001",
  47945=>"110000000",
  47946=>"001111010",
  47947=>"010011011",
  47948=>"000000001",
  47949=>"000101111",
  47950=>"110000000",
  47951=>"011011101",
  47952=>"000100100",
  47953=>"000000001",
  47954=>"110110110",
  47955=>"111011000",
  47956=>"100000000",
  47957=>"010100001",
  47958=>"111010000",
  47959=>"111110111",
  47960=>"111100000",
  47961=>"101000010",
  47962=>"100100111",
  47963=>"111000001",
  47964=>"000000000",
  47965=>"000000111",
  47966=>"010010110",
  47967=>"000000111",
  47968=>"001001111",
  47969=>"010111111",
  47970=>"011111111",
  47971=>"111111000",
  47972=>"110110100",
  47973=>"111110110",
  47974=>"111111000",
  47975=>"111111111",
  47976=>"100110111",
  47977=>"000000101",
  47978=>"111111011",
  47979=>"111100010",
  47980=>"000001111",
  47981=>"110111111",
  47982=>"111111111",
  47983=>"111000001",
  47984=>"000000111",
  47985=>"001000001",
  47986=>"000000100",
  47987=>"011000100",
  47988=>"111100111",
  47989=>"111111110",
  47990=>"110000001",
  47991=>"111000000",
  47992=>"111110000",
  47993=>"000001111",
  47994=>"001111000",
  47995=>"110110111",
  47996=>"111001000",
  47997=>"110011011",
  47998=>"000011010",
  47999=>"111111101",
  48000=>"000000110",
  48001=>"111111111",
  48002=>"000111111",
  48003=>"111111000",
  48004=>"111010000",
  48005=>"111100000",
  48006=>"000000110",
  48007=>"001000000",
  48008=>"000110111",
  48009=>"111111100",
  48010=>"000001101",
  48011=>"111000000",
  48012=>"001101111",
  48013=>"011001001",
  48014=>"111001111",
  48015=>"111000000",
  48016=>"000001111",
  48017=>"111111000",
  48018=>"011001110",
  48019=>"111111101",
  48020=>"100100111",
  48021=>"000110100",
  48022=>"111100000",
  48023=>"111101000",
  48024=>"101001001",
  48025=>"110110110",
  48026=>"111111111",
  48027=>"110110000",
  48028=>"100000000",
  48029=>"010000111",
  48030=>"010110110",
  48031=>"000010000",
  48032=>"000000101",
  48033=>"000000011",
  48034=>"111000000",
  48035=>"011000101",
  48036=>"111010110",
  48037=>"101111000",
  48038=>"011111110",
  48039=>"000000111",
  48040=>"111111001",
  48041=>"000101111",
  48042=>"000000111",
  48043=>"110110110",
  48044=>"000000000",
  48045=>"100000110",
  48046=>"110010000",
  48047=>"000000011",
  48048=>"110000000",
  48049=>"000000110",
  48050=>"000111111",
  48051=>"111111000",
  48052=>"111111111",
  48053=>"111111000",
  48054=>"011001011",
  48055=>"000110110",
  48056=>"101000000",
  48057=>"111101000",
  48058=>"011001011",
  48059=>"111000111",
  48060=>"110100111",
  48061=>"111000000",
  48062=>"101001001",
  48063=>"110100111",
  48064=>"111101001",
  48065=>"000101111",
  48066=>"110000111",
  48067=>"011011011",
  48068=>"111110101",
  48069=>"111000000",
  48070=>"111111000",
  48071=>"001001000",
  48072=>"000000000",
  48073=>"111010000",
  48074=>"111000000",
  48075=>"110001111",
  48076=>"100100000",
  48077=>"000111111",
  48078=>"101000000",
  48079=>"100110110",
  48080=>"111011111",
  48081=>"011011000",
  48082=>"111111111",
  48083=>"111111111",
  48084=>"000000110",
  48085=>"110110101",
  48086=>"000011001",
  48087=>"011001000",
  48088=>"110000000",
  48089=>"111010110",
  48090=>"000100111",
  48091=>"111111100",
  48092=>"001000000",
  48093=>"110000110",
  48094=>"000000100",
  48095=>"110111011",
  48096=>"111111000",
  48097=>"111000000",
  48098=>"111110111",
  48099=>"000000110",
  48100=>"111110111",
  48101=>"000000000",
  48102=>"001011111",
  48103=>"001001111",
  48104=>"111100110",
  48105=>"000001001",
  48106=>"011000000",
  48107=>"111000000",
  48108=>"000000011",
  48109=>"010010011",
  48110=>"000111111",
  48111=>"111111000",
  48112=>"010010000",
  48113=>"000000111",
  48114=>"100000100",
  48115=>"100000000",
  48116=>"110000000",
  48117=>"000000000",
  48118=>"111110000",
  48119=>"111001110",
  48120=>"111000111",
  48121=>"010110100",
  48122=>"100000001",
  48123=>"111000011",
  48124=>"110100001",
  48125=>"000110111",
  48126=>"101110010",
  48127=>"000000111",
  48128=>"011001000",
  48129=>"000000110",
  48130=>"101000001",
  48131=>"000000000",
  48132=>"000000111",
  48133=>"000000001",
  48134=>"000000000",
  48135=>"000111111",
  48136=>"101101100",
  48137=>"101111111",
  48138=>"111111101",
  48139=>"111001000",
  48140=>"000000010",
  48141=>"111011011",
  48142=>"111111011",
  48143=>"110111111",
  48144=>"000100111",
  48145=>"000000011",
  48146=>"001000011",
  48147=>"100100111",
  48148=>"000110110",
  48149=>"100001010",
  48150=>"011111111",
  48151=>"111111110",
  48152=>"111111011",
  48153=>"111111111",
  48154=>"101000000",
  48155=>"000000100",
  48156=>"111111011",
  48157=>"000000000",
  48158=>"010111110",
  48159=>"010000111",
  48160=>"000000000",
  48161=>"111111000",
  48162=>"011110000",
  48163=>"111111111",
  48164=>"111111101",
  48165=>"100111111",
  48166=>"100000000",
  48167=>"111111111",
  48168=>"000000000",
  48169=>"000000000",
  48170=>"001001000",
  48171=>"111000000",
  48172=>"111111111",
  48173=>"000110110",
  48174=>"000001111",
  48175=>"001000111",
  48176=>"011111000",
  48177=>"000000000",
  48178=>"100000100",
  48179=>"111011111",
  48180=>"000100000",
  48181=>"010101000",
  48182=>"000110111",
  48183=>"111111000",
  48184=>"111111111",
  48185=>"111111111",
  48186=>"001001000",
  48187=>"100100111",
  48188=>"111111000",
  48189=>"011111111",
  48190=>"011011001",
  48191=>"111111111",
  48192=>"001011111",
  48193=>"000000000",
  48194=>"010111010",
  48195=>"111111011",
  48196=>"111111011",
  48197=>"000000110",
  48198=>"000111111",
  48199=>"000000111",
  48200=>"111111111",
  48201=>"111101101",
  48202=>"010000000",
  48203=>"101101000",
  48204=>"111011000",
  48205=>"000000000",
  48206=>"111111111",
  48207=>"000000000",
  48208=>"001010000",
  48209=>"110000000",
  48210=>"111111111",
  48211=>"000000010",
  48212=>"010000000",
  48213=>"111000000",
  48214=>"111111000",
  48215=>"000000000",
  48216=>"010010001",
  48217=>"111100101",
  48218=>"100101111",
  48219=>"000000000",
  48220=>"111011011",
  48221=>"111111111",
  48222=>"000110100",
  48223=>"011001111",
  48224=>"111111101",
  48225=>"111111111",
  48226=>"000000111",
  48227=>"001101111",
  48228=>"111001000",
  48229=>"101000111",
  48230=>"001111000",
  48231=>"000000000",
  48232=>"000000110",
  48233=>"000101111",
  48234=>"110000000",
  48235=>"000000000",
  48236=>"100101001",
  48237=>"111111001",
  48238=>"000000111",
  48239=>"000100110",
  48240=>"000000000",
  48241=>"111111111",
  48242=>"000000011",
  48243=>"000111111",
  48244=>"001000000",
  48245=>"111000010",
  48246=>"111001010",
  48247=>"000000000",
  48248=>"100000000",
  48249=>"011011000",
  48250=>"011001000",
  48251=>"100000111",
  48252=>"110110100",
  48253=>"111011011",
  48254=>"111111110",
  48255=>"000011111",
  48256=>"111110110",
  48257=>"111111111",
  48258=>"000110111",
  48259=>"000100101",
  48260=>"001001001",
  48261=>"111111111",
  48262=>"111111000",
  48263=>"000111111",
  48264=>"111100000",
  48265=>"000111111",
  48266=>"001001111",
  48267=>"100100100",
  48268=>"010010000",
  48269=>"111111011",
  48270=>"111111000",
  48271=>"000010011",
  48272=>"111111000",
  48273=>"000000110",
  48274=>"111100111",
  48275=>"001011111",
  48276=>"011110000",
  48277=>"010111111",
  48278=>"111100100",
  48279=>"111111000",
  48280=>"000000100",
  48281=>"000001000",
  48282=>"000000000",
  48283=>"110111111",
  48284=>"100000111",
  48285=>"001111110",
  48286=>"111111000",
  48287=>"000111111",
  48288=>"000000000",
  48289=>"111111100",
  48290=>"001000000",
  48291=>"111110000",
  48292=>"000000000",
  48293=>"000000111",
  48294=>"001000011",
  48295=>"000000000",
  48296=>"000000101",
  48297=>"111111111",
  48298=>"000100111",
  48299=>"111111110",
  48300=>"111111111",
  48301=>"110110000",
  48302=>"000000000",
  48303=>"001111111",
  48304=>"000011000",
  48305=>"100011011",
  48306=>"000110010",
  48307=>"111111000",
  48308=>"010010000",
  48309=>"000001001",
  48310=>"110011001",
  48311=>"111000011",
  48312=>"000000000",
  48313=>"000000111",
  48314=>"000000000",
  48315=>"111111000",
  48316=>"000000011",
  48317=>"111110000",
  48318=>"000110111",
  48319=>"110111111",
  48320=>"001000000",
  48321=>"101111111",
  48322=>"000001011",
  48323=>"000001111",
  48324=>"100100000",
  48325=>"000000000",
  48326=>"101100000",
  48327=>"011000000",
  48328=>"111111011",
  48329=>"000000111",
  48330=>"000000001",
  48331=>"000000000",
  48332=>"000001101",
  48333=>"011011000",
  48334=>"000000011",
  48335=>"001111111",
  48336=>"111100110",
  48337=>"100000100",
  48338=>"001011011",
  48339=>"011111111",
  48340=>"000000001",
  48341=>"110110001",
  48342=>"000000111",
  48343=>"000000000",
  48344=>"011000000",
  48345=>"110000100",
  48346=>"100100000",
  48347=>"111111011",
  48348=>"111111001",
  48349=>"111101001",
  48350=>"111111000",
  48351=>"000000000",
  48352=>"000000000",
  48353=>"000111110",
  48354=>"000011111",
  48355=>"000000000",
  48356=>"000000110",
  48357=>"000000000",
  48358=>"110100000",
  48359=>"111011000",
  48360=>"111111111",
  48361=>"111011000",
  48362=>"001001101",
  48363=>"000000000",
  48364=>"111111111",
  48365=>"110111111",
  48366=>"011011111",
  48367=>"000000011",
  48368=>"110111000",
  48369=>"110000100",
  48370=>"111111001",
  48371=>"000000000",
  48372=>"111111000",
  48373=>"100100110",
  48374=>"111101101",
  48375=>"000000011",
  48376=>"111111110",
  48377=>"011111111",
  48378=>"111111111",
  48379=>"100100111",
  48380=>"000100000",
  48381=>"101111111",
  48382=>"010010000",
  48383=>"111111111",
  48384=>"001001111",
  48385=>"000000000",
  48386=>"000000000",
  48387=>"111111111",
  48388=>"000000000",
  48389=>"110100100",
  48390=>"111111000",
  48391=>"111111000",
  48392=>"000011111",
  48393=>"000000001",
  48394=>"000000000",
  48395=>"000000000",
  48396=>"110110000",
  48397=>"011000000",
  48398=>"111011111",
  48399=>"001000001",
  48400=>"111111011",
  48401=>"001001100",
  48402=>"100100000",
  48403=>"111110000",
  48404=>"111011111",
  48405=>"111100000",
  48406=>"001000000",
  48407=>"000000000",
  48408=>"111101000",
  48409=>"000101111",
  48410=>"000110000",
  48411=>"110000111",
  48412=>"111001011",
  48413=>"000000111",
  48414=>"111010000",
  48415=>"111111111",
  48416=>"110111011",
  48417=>"101101100",
  48418=>"000000000",
  48419=>"000001001",
  48420=>"100111111",
  48421=>"000011000",
  48422=>"000000111",
  48423=>"000100111",
  48424=>"101111111",
  48425=>"011011000",
  48426=>"110110100",
  48427=>"100000000",
  48428=>"000001000",
  48429=>"001101111",
  48430=>"000111111",
  48431=>"111000000",
  48432=>"000001000",
  48433=>"000001111",
  48434=>"001100110",
  48435=>"000110111",
  48436=>"111111110",
  48437=>"011001000",
  48438=>"111111110",
  48439=>"000000000",
  48440=>"000011000",
  48441=>"110000000",
  48442=>"111111100",
  48443=>"000100111",
  48444=>"011110110",
  48445=>"000000000",
  48446=>"001111111",
  48447=>"111111000",
  48448=>"111111111",
  48449=>"111111001",
  48450=>"000011011",
  48451=>"001000000",
  48452=>"011001000",
  48453=>"000000000",
  48454=>"000111110",
  48455=>"000000000",
  48456=>"000100110",
  48457=>"111111111",
  48458=>"011100000",
  48459=>"011111011",
  48460=>"011011011",
  48461=>"111111000",
  48462=>"011000000",
  48463=>"111111000",
  48464=>"000000000",
  48465=>"111000011",
  48466=>"111110001",
  48467=>"111111000",
  48468=>"000000100",
  48469=>"001001001",
  48470=>"001011001",
  48471=>"001111111",
  48472=>"000011111",
  48473=>"001000111",
  48474=>"111111010",
  48475=>"000000101",
  48476=>"101101111",
  48477=>"000000000",
  48478=>"000000000",
  48479=>"111001000",
  48480=>"111111111",
  48481=>"001001011",
  48482=>"001011111",
  48483=>"000000111",
  48484=>"111101000",
  48485=>"001001011",
  48486=>"010000000",
  48487=>"000000000",
  48488=>"111110010",
  48489=>"111111101",
  48490=>"000000110",
  48491=>"100110110",
  48492=>"010010010",
  48493=>"101111011",
  48494=>"111111111",
  48495=>"000111111",
  48496=>"111111110",
  48497=>"110111000",
  48498=>"001111111",
  48499=>"001011000",
  48500=>"000000000",
  48501=>"000000100",
  48502=>"000000111",
  48503=>"000000100",
  48504=>"000000111",
  48505=>"100000111",
  48506=>"000010000",
  48507=>"111111000",
  48508=>"111111010",
  48509=>"011010000",
  48510=>"001111110",
  48511=>"001111111",
  48512=>"000000000",
  48513=>"000010110",
  48514=>"000000111",
  48515=>"000000001",
  48516=>"001011111",
  48517=>"111001010",
  48518=>"100000001",
  48519=>"000100111",
  48520=>"000100110",
  48521=>"011001001",
  48522=>"000000000",
  48523=>"001001111",
  48524=>"111111111",
  48525=>"100110110",
  48526=>"100000000",
  48527=>"111101111",
  48528=>"000000001",
  48529=>"111011101",
  48530=>"000000101",
  48531=>"001011111",
  48532=>"111100111",
  48533=>"000000000",
  48534=>"111000000",
  48535=>"000000000",
  48536=>"111001001",
  48537=>"100110011",
  48538=>"111011001",
  48539=>"001001001",
  48540=>"100000000",
  48541=>"111111111",
  48542=>"100000000",
  48543=>"000111111",
  48544=>"000000000",
  48545=>"110110010",
  48546=>"001111111",
  48547=>"000100101",
  48548=>"111111111",
  48549=>"000000111",
  48550=>"001110111",
  48551=>"100111111",
  48552=>"000001001",
  48553=>"111111100",
  48554=>"111000000",
  48555=>"001011110",
  48556=>"100100100",
  48557=>"001001000",
  48558=>"100100111",
  48559=>"111000000",
  48560=>"000000000",
  48561=>"000000000",
  48562=>"110110100",
  48563=>"111111000",
  48564=>"101110110",
  48565=>"111111111",
  48566=>"111111111",
  48567=>"100000111",
  48568=>"000000111",
  48569=>"101100000",
  48570=>"000100110",
  48571=>"011111000",
  48572=>"100000011",
  48573=>"001000000",
  48574=>"101001111",
  48575=>"000000001",
  48576=>"111110000",
  48577=>"001000000",
  48578=>"011111111",
  48579=>"111111111",
  48580=>"000000101",
  48581=>"001011001",
  48582=>"111110010",
  48583=>"111000000",
  48584=>"000000111",
  48585=>"000000000",
  48586=>"010111101",
  48587=>"110111111",
  48588=>"010100111",
  48589=>"111111000",
  48590=>"111111010",
  48591=>"000000100",
  48592=>"001001111",
  48593=>"000111111",
  48594=>"011110010",
  48595=>"111100010",
  48596=>"001011000",
  48597=>"100111101",
  48598=>"111110000",
  48599=>"000000000",
  48600=>"000011000",
  48601=>"101000000",
  48602=>"000000111",
  48603=>"000000000",
  48604=>"000000000",
  48605=>"111111000",
  48606=>"111111111",
  48607=>"000000000",
  48608=>"000100000",
  48609=>"111111111",
  48610=>"000000000",
  48611=>"111111000",
  48612=>"111111100",
  48613=>"001010000",
  48614=>"011111111",
  48615=>"100110111",
  48616=>"011001000",
  48617=>"100000111",
  48618=>"001000000",
  48619=>"111111000",
  48620=>"111111111",
  48621=>"001001001",
  48622=>"011000000",
  48623=>"111111111",
  48624=>"000000000",
  48625=>"111111111",
  48626=>"111111111",
  48627=>"001111111",
  48628=>"000000000",
  48629=>"000000100",
  48630=>"010010110",
  48631=>"011011000",
  48632=>"111111001",
  48633=>"001001011",
  48634=>"111110000",
  48635=>"000000100",
  48636=>"111111111",
  48637=>"000000111",
  48638=>"000000000",
  48639=>"000000000",
  48640=>"000001001",
  48641=>"111010010",
  48642=>"111110000",
  48643=>"000111111",
  48644=>"010111111",
  48645=>"000000000",
  48646=>"000000000",
  48647=>"111011011",
  48648=>"111111111",
  48649=>"000000000",
  48650=>"111111111",
  48651=>"001111110",
  48652=>"100000011",
  48653=>"101000011",
  48654=>"000100110",
  48655=>"111001011",
  48656=>"111001001",
  48657=>"111111000",
  48658=>"110111111",
  48659=>"111111111",
  48660=>"110000111",
  48661=>"001001000",
  48662=>"110110001",
  48663=>"011001001",
  48664=>"111111000",
  48665=>"111111110",
  48666=>"011111001",
  48667=>"111011000",
  48668=>"000100110",
  48669=>"010000000",
  48670=>"111110001",
  48671=>"110100100",
  48672=>"000000000",
  48673=>"110110110",
  48674=>"111110000",
  48675=>"101000000",
  48676=>"000000000",
  48677=>"001001001",
  48678=>"110110110",
  48679=>"000101001",
  48680=>"001111101",
  48681=>"010010010",
  48682=>"111111111",
  48683=>"111110000",
  48684=>"111111111",
  48685=>"101111111",
  48686=>"101000111",
  48687=>"011010111",
  48688=>"000110000",
  48689=>"101001011",
  48690=>"001101011",
  48691=>"011111011",
  48692=>"111011001",
  48693=>"000000111",
  48694=>"100101000",
  48695=>"001111111",
  48696=>"000000111",
  48697=>"000001101",
  48698=>"001000000",
  48699=>"011111111",
  48700=>"101000000",
  48701=>"000000001",
  48702=>"000110111",
  48703=>"000000111",
  48704=>"000000101",
  48705=>"000001001",
  48706=>"000000111",
  48707=>"111111111",
  48708=>"001011000",
  48709=>"011001111",
  48710=>"000111011",
  48711=>"000000000",
  48712=>"111111001",
  48713=>"001001000",
  48714=>"111111111",
  48715=>"000000000",
  48716=>"000100110",
  48717=>"111011101",
  48718=>"001000101",
  48719=>"111001000",
  48720=>"011001000",
  48721=>"100111111",
  48722=>"001000000",
  48723=>"001001001",
  48724=>"000000111",
  48725=>"110000000",
  48726=>"011010111",
  48727=>"000000000",
  48728=>"110110111",
  48729=>"000000000",
  48730=>"111111111",
  48731=>"111010111",
  48732=>"110111110",
  48733=>"000000101",
  48734=>"111111110",
  48735=>"000000111",
  48736=>"110111110",
  48737=>"110111111",
  48738=>"111111111",
  48739=>"000010011",
  48740=>"000111111",
  48741=>"011001101",
  48742=>"000000110",
  48743=>"000000111",
  48744=>"000000100",
  48745=>"001001001",
  48746=>"000000000",
  48747=>"001001100",
  48748=>"111111111",
  48749=>"000000001",
  48750=>"111011000",
  48751=>"111101000",
  48752=>"100110110",
  48753=>"100101001",
  48754=>"001001001",
  48755=>"010000001",
  48756=>"010010010",
  48757=>"111000001",
  48758=>"000000011",
  48759=>"111111111",
  48760=>"111111111",
  48761=>"111110000",
  48762=>"000000000",
  48763=>"111111111",
  48764=>"111111111",
  48765=>"000000000",
  48766=>"100000001",
  48767=>"000000001",
  48768=>"101000000",
  48769=>"111111000",
  48770=>"010010110",
  48771=>"001000011",
  48772=>"000001001",
  48773=>"000000000",
  48774=>"000001111",
  48775=>"000001000",
  48776=>"001001001",
  48777=>"000001001",
  48778=>"001000100",
  48779=>"000111111",
  48780=>"011101101",
  48781=>"111111111",
  48782=>"110000111",
  48783=>"101101101",
  48784=>"111101111",
  48785=>"001000000",
  48786=>"011000111",
  48787=>"110110110",
  48788=>"010110001",
  48789=>"101001011",
  48790=>"111001111",
  48791=>"000001000",
  48792=>"001001000",
  48793=>"000000000",
  48794=>"010000111",
  48795=>"001000000",
  48796=>"000010000",
  48797=>"000000111",
  48798=>"110110110",
  48799=>"000000000",
  48800=>"010110001",
  48801=>"001111101",
  48802=>"000000001",
  48803=>"010111110",
  48804=>"000000000",
  48805=>"110111111",
  48806=>"010010000",
  48807=>"010010111",
  48808=>"111101011",
  48809=>"000000000",
  48810=>"111111100",
  48811=>"000000011",
  48812=>"001001101",
  48813=>"110100110",
  48814=>"110110000",
  48815=>"111111111",
  48816=>"100000111",
  48817=>"000000100",
  48818=>"010111111",
  48819=>"111000000",
  48820=>"111110110",
  48821=>"111101111",
  48822=>"000000000",
  48823=>"111111000",
  48824=>"000000000",
  48825=>"000000000",
  48826=>"001101100",
  48827=>"010010111",
  48828=>"000000000",
  48829=>"001001000",
  48830=>"000100111",
  48831=>"000000000",
  48832=>"000000000",
  48833=>"000100110",
  48834=>"001001111",
  48835=>"110111010",
  48836=>"111000000",
  48837=>"010000001",
  48838=>"000111010",
  48839=>"111111000",
  48840=>"111111001",
  48841=>"001000001",
  48842=>"000100000",
  48843=>"111100000",
  48844=>"110001010",
  48845=>"111110111",
  48846=>"111011011",
  48847=>"111110111",
  48848=>"111000011",
  48849=>"000000000",
  48850=>"111011111",
  48851=>"110110111",
  48852=>"100000001",
  48853=>"111111001",
  48854=>"100000000",
  48855=>"011111110",
  48856=>"110110001",
  48857=>"001111101",
  48858=>"000000111",
  48859=>"111111111",
  48860=>"111111111",
  48861=>"100100111",
  48862=>"111111111",
  48863=>"000000001",
  48864=>"000000000",
  48865=>"111111010",
  48866=>"111111101",
  48867=>"010001000",
  48868=>"000000100",
  48869=>"111111111",
  48870=>"001000000",
  48871=>"000000101",
  48872=>"100000000",
  48873=>"000100001",
  48874=>"000000001",
  48875=>"010000000",
  48876=>"111101101",
  48877=>"000000000",
  48878=>"111111111",
  48879=>"001001001",
  48880=>"100100111",
  48881=>"000000111",
  48882=>"001000000",
  48883=>"000000100",
  48884=>"111111001",
  48885=>"000000010",
  48886=>"111111010",
  48887=>"000000001",
  48888=>"001000000",
  48889=>"111011000",
  48890=>"010010110",
  48891=>"000000100",
  48892=>"111101100",
  48893=>"010000010",
  48894=>"010110001",
  48895=>"111111111",
  48896=>"100101111",
  48897=>"111111101",
  48898=>"100100000",
  48899=>"001000000",
  48900=>"011111111",
  48901=>"100000110",
  48902=>"000100100",
  48903=>"111111111",
  48904=>"000000111",
  48905=>"001000001",
  48906=>"111000000",
  48907=>"000000000",
  48908=>"001001011",
  48909=>"001111100",
  48910=>"100111010",
  48911=>"000000111",
  48912=>"000000110",
  48913=>"100101000",
  48914=>"011001111",
  48915=>"000000001",
  48916=>"101001000",
  48917=>"111000000",
  48918=>"101001110",
  48919=>"111111111",
  48920=>"000010000",
  48921=>"111111000",
  48922=>"110000000",
  48923=>"100100000",
  48924=>"000000110",
  48925=>"000000000",
  48926=>"111111111",
  48927=>"000001001",
  48928=>"000110011",
  48929=>"100110111",
  48930=>"000000111",
  48931=>"000000010",
  48932=>"011110111",
  48933=>"101000001",
  48934=>"111111101",
  48935=>"010101111",
  48936=>"000111111",
  48937=>"000100100",
  48938=>"000000001",
  48939=>"000000110",
  48940=>"001000000",
  48941=>"000000111",
  48942=>"011011111",
  48943=>"111101111",
  48944=>"111111000",
  48945=>"111111111",
  48946=>"111001111",
  48947=>"111110111",
  48948=>"111111001",
  48949=>"110100111",
  48950=>"111011000",
  48951=>"001000001",
  48952=>"111111111",
  48953=>"111011111",
  48954=>"110111101",
  48955=>"101111111",
  48956=>"010000000",
  48957=>"101001000",
  48958=>"111110110",
  48959=>"000110001",
  48960=>"111000000",
  48961=>"000100100",
  48962=>"111111111",
  48963=>"000111111",
  48964=>"101111011",
  48965=>"001010011",
  48966=>"000000000",
  48967=>"000100100",
  48968=>"111111011",
  48969=>"000011000",
  48970=>"110000000",
  48971=>"010011011",
  48972=>"011000001",
  48973=>"111011001",
  48974=>"000100001",
  48975=>"111101101",
  48976=>"000000101",
  48977=>"010100111",
  48978=>"001000111",
  48979=>"000000000",
  48980=>"000000000",
  48981=>"110110010",
  48982=>"010001111",
  48983=>"000000000",
  48984=>"000000000",
  48985=>"111110011",
  48986=>"010000111",
  48987=>"001001001",
  48988=>"111111111",
  48989=>"001000000",
  48990=>"111001001",
  48991=>"001101100",
  48992=>"000101001",
  48993=>"010010011",
  48994=>"111011000",
  48995=>"100000000",
  48996=>"111011000",
  48997=>"011111001",
  48998=>"001111000",
  48999=>"111111110",
  49000=>"101110111",
  49001=>"000000010",
  49002=>"000110111",
  49003=>"001000000",
  49004=>"111111110",
  49005=>"000000000",
  49006=>"000000000",
  49007=>"111100101",
  49008=>"000000000",
  49009=>"111111111",
  49010=>"000011010",
  49011=>"111111000",
  49012=>"100000110",
  49013=>"001111111",
  49014=>"011111110",
  49015=>"111111111",
  49016=>"111100111",
  49017=>"000010011",
  49018=>"111110110",
  49019=>"110000100",
  49020=>"001000000",
  49021=>"110110000",
  49022=>"111010000",
  49023=>"111111111",
  49024=>"111111111",
  49025=>"110010001",
  49026=>"101000000",
  49027=>"011011011",
  49028=>"010111001",
  49029=>"100000000",
  49030=>"000011111",
  49031=>"001001000",
  49032=>"011000000",
  49033=>"111110101",
  49034=>"111011011",
  49035=>"000001000",
  49036=>"111111100",
  49037=>"111111111",
  49038=>"111111101",
  49039=>"111101101",
  49040=>"010111011",
  49041=>"110100100",
  49042=>"000011010",
  49043=>"111000000",
  49044=>"111111111",
  49045=>"000000000",
  49046=>"001001001",
  49047=>"001100111",
  49048=>"100111110",
  49049=>"011111110",
  49050=>"000000000",
  49051=>"000000000",
  49052=>"000000100",
  49053=>"001111111",
  49054=>"001101111",
  49055=>"000000001",
  49056=>"111110000",
  49057=>"110110000",
  49058=>"000000110",
  49059=>"011111111",
  49060=>"111111111",
  49061=>"000000011",
  49062=>"010111111",
  49063=>"000000000",
  49064=>"111110000",
  49065=>"110110010",
  49066=>"111111111",
  49067=>"000000000",
  49068=>"111111000",
  49069=>"110111001",
  49070=>"100000111",
  49071=>"010110000",
  49072=>"000000111",
  49073=>"111111111",
  49074=>"001001011",
  49075=>"110111111",
  49076=>"111110111",
  49077=>"000000000",
  49078=>"000100101",
  49079=>"000000111",
  49080=>"111111111",
  49081=>"111111111",
  49082=>"111001000",
  49083=>"000000001",
  49084=>"101111111",
  49085=>"111111110",
  49086=>"001001111",
  49087=>"100111110",
  49088=>"100000000",
  49089=>"011011111",
  49090=>"111111111",
  49091=>"001011111",
  49092=>"111110011",
  49093=>"100110111",
  49094=>"110110000",
  49095=>"000000110",
  49096=>"111111111",
  49097=>"010000001",
  49098=>"001000000",
  49099=>"011111111",
  49100=>"111010011",
  49101=>"111101000",
  49102=>"000110110",
  49103=>"010100111",
  49104=>"001000111",
  49105=>"001100100",
  49106=>"000110110",
  49107=>"111111001",
  49108=>"000000000",
  49109=>"111111111",
  49110=>"000000111",
  49111=>"000000000",
  49112=>"101110110",
  49113=>"000000000",
  49114=>"000000111",
  49115=>"111101111",
  49116=>"100111111",
  49117=>"100101001",
  49118=>"111110000",
  49119=>"000000101",
  49120=>"010100000",
  49121=>"001111000",
  49122=>"100000001",
  49123=>"100111001",
  49124=>"111010010",
  49125=>"011011011",
  49126=>"001000000",
  49127=>"000000000",
  49128=>"000111111",
  49129=>"000000000",
  49130=>"111111111",
  49131=>"000000000",
  49132=>"111101111",
  49133=>"001001000",
  49134=>"111110011",
  49135=>"111111111",
  49136=>"000000001",
  49137=>"000000000",
  49138=>"111111111",
  49139=>"000000001",
  49140=>"000000001",
  49141=>"000100100",
  49142=>"110001111",
  49143=>"100000000",
  49144=>"111001001",
  49145=>"100100111",
  49146=>"000001111",
  49147=>"110111111",
  49148=>"000000111",
  49149=>"111110001",
  49150=>"000001000",
  49151=>"101000001",
  49152=>"000100000",
  49153=>"001000000",
  49154=>"000000101",
  49155=>"111001101",
  49156=>"000001111",
  49157=>"000000000",
  49158=>"111111111",
  49159=>"011111111",
  49160=>"111000000",
  49161=>"111111111",
  49162=>"100100000",
  49163=>"000000111",
  49164=>"000011001",
  49165=>"111111001",
  49166=>"001111111",
  49167=>"111000000",
  49168=>"111011000",
  49169=>"111111111",
  49170=>"111111111",
  49171=>"000000101",
  49172=>"000000110",
  49173=>"110100110",
  49174=>"111111011",
  49175=>"100011001",
  49176=>"001000010",
  49177=>"011001000",
  49178=>"000000000",
  49179=>"000000000",
  49180=>"000110100",
  49181=>"111111111",
  49182=>"111110110",
  49183=>"111100100",
  49184=>"010000000",
  49185=>"000100000",
  49186=>"111111111",
  49187=>"111111111",
  49188=>"001001001",
  49189=>"000000011",
  49190=>"111100000",
  49191=>"111111111",
  49192=>"100101111",
  49193=>"111111111",
  49194=>"000111111",
  49195=>"111111111",
  49196=>"111010011",
  49197=>"001001111",
  49198=>"010110000",
  49199=>"000000110",
  49200=>"101000011",
  49201=>"000000000",
  49202=>"110111011",
  49203=>"000000000",
  49204=>"000101111",
  49205=>"010000011",
  49206=>"101000100",
  49207=>"110110110",
  49208=>"000111111",
  49209=>"111111111",
  49210=>"111111111",
  49211=>"111111000",
  49212=>"111000100",
  49213=>"100100000",
  49214=>"000001011",
  49215=>"000000111",
  49216=>"000011000",
  49217=>"010111110",
  49218=>"001111101",
  49219=>"111101111",
  49220=>"001000000",
  49221=>"000100110",
  49222=>"000110111",
  49223=>"111111111",
  49224=>"100100000",
  49225=>"111111111",
  49226=>"111111000",
  49227=>"110100000",
  49228=>"011111111",
  49229=>"111100001",
  49230=>"111100100",
  49231=>"111111111",
  49232=>"111111000",
  49233=>"000111111",
  49234=>"000000010",
  49235=>"000000100",
  49236=>"001001000",
  49237=>"000000111",
  49238=>"111111100",
  49239=>"000010010",
  49240=>"101111101",
  49241=>"100000100",
  49242=>"111111110",
  49243=>"111111111",
  49244=>"001111111",
  49245=>"100101000",
  49246=>"000000000",
  49247=>"111001000",
  49248=>"000100111",
  49249=>"000000000",
  49250=>"000000001",
  49251=>"011000000",
  49252=>"111111011",
  49253=>"000000000",
  49254=>"100100111",
  49255=>"111111111",
  49256=>"111111111",
  49257=>"000000100",
  49258=>"000111111",
  49259=>"111111111",
  49260=>"000110011",
  49261=>"111111111",
  49262=>"111111111",
  49263=>"010000000",
  49264=>"000111111",
  49265=>"000000000",
  49266=>"111111100",
  49267=>"111111111",
  49268=>"000000000",
  49269=>"111111001",
  49270=>"000000000",
  49271=>"000000000",
  49272=>"010010000",
  49273=>"000000001",
  49274=>"000000000",
  49275=>"000001001",
  49276=>"000110010",
  49277=>"000000000",
  49278=>"000000000",
  49279=>"111111000",
  49280=>"111111111",
  49281=>"110100110",
  49282=>"100111111",
  49283=>"000100000",
  49284=>"000011011",
  49285=>"000000111",
  49286=>"000000001",
  49287=>"111111111",
  49288=>"111111111",
  49289=>"111010000",
  49290=>"111111111",
  49291=>"000000000",
  49292=>"101111000",
  49293=>"001000100",
  49294=>"110110110",
  49295=>"111111101",
  49296=>"000000111",
  49297=>"111100000",
  49298=>"000000000",
  49299=>"000111111",
  49300=>"000000011",
  49301=>"111111000",
  49302=>"111111111",
  49303=>"111111111",
  49304=>"000000101",
  49305=>"101000000",
  49306=>"100100111",
  49307=>"000001000",
  49308=>"000000110",
  49309=>"000111000",
  49310=>"100000000",
  49311=>"111000000",
  49312=>"000000000",
  49313=>"111100100",
  49314=>"111111111",
  49315=>"000111111",
  49316=>"001111111",
  49317=>"000000000",
  49318=>"111110000",
  49319=>"010000110",
  49320=>"000111111",
  49321=>"000000000",
  49322=>"111100000",
  49323=>"000000000",
  49324=>"111111111",
  49325=>"111111111",
  49326=>"000100111",
  49327=>"000111111",
  49328=>"001111111",
  49329=>"011011001",
  49330=>"010110010",
  49331=>"111111111",
  49332=>"111000000",
  49333=>"000111111",
  49334=>"101111111",
  49335=>"111111000",
  49336=>"111111001",
  49337=>"111111011",
  49338=>"000000000",
  49339=>"100111111",
  49340=>"000000000",
  49341=>"111111110",
  49342=>"000111111",
  49343=>"000001000",
  49344=>"111111111",
  49345=>"001011011",
  49346=>"111111001",
  49347=>"110010000",
  49348=>"000000000",
  49349=>"000111111",
  49350=>"110110111",
  49351=>"111111111",
  49352=>"111111111",
  49353=>"111011000",
  49354=>"000000000",
  49355=>"111111111",
  49356=>"100100000",
  49357=>"111111111",
  49358=>"001011111",
  49359=>"111111111",
  49360=>"111111111",
  49361=>"111000100",
  49362=>"000111111",
  49363=>"111111111",
  49364=>"000000011",
  49365=>"111000000",
  49366=>"100100000",
  49367=>"111111111",
  49368=>"101111111",
  49369=>"000000001",
  49370=>"111111100",
  49371=>"001000000",
  49372=>"111111111",
  49373=>"000000000",
  49374=>"000101111",
  49375=>"000000000",
  49376=>"100100000",
  49377=>"000100111",
  49378=>"111111111",
  49379=>"111111110",
  49380=>"000000000",
  49381=>"111111111",
  49382=>"001000000",
  49383=>"000001111",
  49384=>"111101000",
  49385=>"000000000",
  49386=>"000000000",
  49387=>"001000111",
  49388=>"011111111",
  49389=>"111111000",
  49390=>"000000111",
  49391=>"111000000",
  49392=>"110010000",
  49393=>"010111111",
  49394=>"000111111",
  49395=>"100100000",
  49396=>"000000011",
  49397=>"100000110",
  49398=>"000111100",
  49399=>"111000111",
  49400=>"110111111",
  49401=>"000011000",
  49402=>"000000000",
  49403=>"000001111",
  49404=>"111111100",
  49405=>"000001001",
  49406=>"111100100",
  49407=>"111000000",
  49408=>"111111111",
  49409=>"001000100",
  49410=>"000010000",
  49411=>"000100000",
  49412=>"100110110",
  49413=>"000101111",
  49414=>"111111111",
  49415=>"010111111",
  49416=>"000000011",
  49417=>"000000000",
  49418=>"111010000",
  49419=>"110110111",
  49420=>"000000000",
  49421=>"000000111",
  49422=>"000000000",
  49423=>"111111000",
  49424=>"000000000",
  49425=>"000111101",
  49426=>"111111101",
  49427=>"001011011",
  49428=>"111111111",
  49429=>"000011111",
  49430=>"001001001",
  49431=>"000000111",
  49432=>"111100100",
  49433=>"111111111",
  49434=>"000000000",
  49435=>"100111111",
  49436=>"011111001",
  49437=>"000000000",
  49438=>"100000000",
  49439=>"100100100",
  49440=>"111111000",
  49441=>"101111111",
  49442=>"111000000",
  49443=>"111111111",
  49444=>"000000011",
  49445=>"111001000",
  49446=>"100110110",
  49447=>"000000000",
  49448=>"000000100",
  49449=>"000000000",
  49450=>"000111000",
  49451=>"110110000",
  49452=>"111010110",
  49453=>"000011000",
  49454=>"111111011",
  49455=>"000010011",
  49456=>"110110000",
  49457=>"000100000",
  49458=>"111110111",
  49459=>"000011111",
  49460=>"010011011",
  49461=>"000000000",
  49462=>"000111111",
  49463=>"000111111",
  49464=>"000000000",
  49465=>"011011111",
  49466=>"000000000",
  49467=>"011000000",
  49468=>"000111111",
  49469=>"000000100",
  49470=>"100000000",
  49471=>"111000000",
  49472=>"000000000",
  49473=>"111000000",
  49474=>"000111111",
  49475=>"111111111",
  49476=>"111001011",
  49477=>"000110110",
  49478=>"011111000",
  49479=>"000111011",
  49480=>"000000000",
  49481=>"111111011",
  49482=>"000111101",
  49483=>"111011000",
  49484=>"111110000",
  49485=>"111111110",
  49486=>"111101101",
  49487=>"111111111",
  49488=>"000000000",
  49489=>"101100111",
  49490=>"111111000",
  49491=>"111001010",
  49492=>"000111111",
  49493=>"011011011",
  49494=>"110101110",
  49495=>"000000001",
  49496=>"111111111",
  49497=>"000000000",
  49498=>"110000000",
  49499=>"110000111",
  49500=>"000000000",
  49501=>"110000000",
  49502=>"111000000",
  49503=>"001001000",
  49504=>"000100111",
  49505=>"000000000",
  49506=>"111111111",
  49507=>"000011000",
  49508=>"000000111",
  49509=>"000000000",
  49510=>"111111100",
  49511=>"000111111",
  49512=>"000100100",
  49513=>"111111100",
  49514=>"000011010",
  49515=>"000010000",
  49516=>"111111111",
  49517=>"000000000",
  49518=>"111111000",
  49519=>"000000000",
  49520=>"000000000",
  49521=>"111011000",
  49522=>"111101111",
  49523=>"000000111",
  49524=>"111111111",
  49525=>"000000000",
  49526=>"000110000",
  49527=>"000000000",
  49528=>"111111001",
  49529=>"111000000",
  49530=>"111110000",
  49531=>"000000010",
  49532=>"111111100",
  49533=>"111111111",
  49534=>"001011011",
  49535=>"111111000",
  49536=>"001001001",
  49537=>"111001000",
  49538=>"000001001",
  49539=>"000000111",
  49540=>"000111001",
  49541=>"000000000",
  49542=>"100000000",
  49543=>"111001000",
  49544=>"111000000",
  49545=>"000000111",
  49546=>"110010000",
  49547=>"111111111",
  49548=>"111111001",
  49549=>"000000000",
  49550=>"100001101",
  49551=>"000111111",
  49552=>"000001001",
  49553=>"111000000",
  49554=>"111111111",
  49555=>"000110110",
  49556=>"011011111",
  49557=>"001001000",
  49558=>"111111111",
  49559=>"000010010",
  49560=>"000111111",
  49561=>"111010010",
  49562=>"000000000",
  49563=>"101111111",
  49564=>"101000111",
  49565=>"000111111",
  49566=>"000110111",
  49567=>"000110111",
  49568=>"111101000",
  49569=>"101100000",
  49570=>"111110010",
  49571=>"111111000",
  49572=>"000000101",
  49573=>"100111111",
  49574=>"111000000",
  49575=>"111111001",
  49576=>"111111111",
  49577=>"000000111",
  49578=>"000001111",
  49579=>"110100000",
  49580=>"111110010",
  49581=>"001000101",
  49582=>"111000000",
  49583=>"111111100",
  49584=>"001000000",
  49585=>"000111000",
  49586=>"111111111",
  49587=>"000111111",
  49588=>"000111111",
  49589=>"000000000",
  49590=>"101001101",
  49591=>"000011111",
  49592=>"100000000",
  49593=>"010111111",
  49594=>"000000000",
  49595=>"000000000",
  49596=>"000000000",
  49597=>"000001000",
  49598=>"101101000",
  49599=>"111010110",
  49600=>"000111111",
  49601=>"000000000",
  49602=>"000000000",
  49603=>"000111000",
  49604=>"000000000",
  49605=>"011111000",
  49606=>"111111111",
  49607=>"110000100",
  49608=>"000000100",
  49609=>"000000000",
  49610=>"000000000",
  49611=>"111111111",
  49612=>"000000000",
  49613=>"110000000",
  49614=>"111101101",
  49615=>"100100100",
  49616=>"000000000",
  49617=>"000110110",
  49618=>"111110100",
  49619=>"000000110",
  49620=>"000000000",
  49621=>"000000000",
  49622=>"001011111",
  49623=>"100110111",
  49624=>"111011000",
  49625=>"111011000",
  49626=>"000000000",
  49627=>"000010000",
  49628=>"000111111",
  49629=>"000000100",
  49630=>"111011000",
  49631=>"101101001",
  49632=>"000001011",
  49633=>"000000000",
  49634=>"001000000",
  49635=>"000000001",
  49636=>"010000000",
  49637=>"000000000",
  49638=>"111111111",
  49639=>"110000000",
  49640=>"000111111",
  49641=>"111111111",
  49642=>"000111100",
  49643=>"001111000",
  49644=>"000110111",
  49645=>"000111001",
  49646=>"111001000",
  49647=>"000000111",
  49648=>"000000000",
  49649=>"110100110",
  49650=>"001000000",
  49651=>"000000000",
  49652=>"101111111",
  49653=>"101111100",
  49654=>"000011000",
  49655=>"000001111",
  49656=>"000110100",
  49657=>"010011011",
  49658=>"000111111",
  49659=>"111101111",
  49660=>"000100101",
  49661=>"111111110",
  49662=>"011111111",
  49663=>"110000000",
  49664=>"011011011",
  49665=>"000000000",
  49666=>"000000000",
  49667=>"010000010",
  49668=>"110111111",
  49669=>"011001001",
  49670=>"111111100",
  49671=>"000000000",
  49672=>"111111110",
  49673=>"001111111",
  49674=>"110011011",
  49675=>"100110100",
  49676=>"000011111",
  49677=>"000000110",
  49678=>"000000000",
  49679=>"101111111",
  49680=>"000010000",
  49681=>"100100100",
  49682=>"110000000",
  49683=>"001111111",
  49684=>"110000000",
  49685=>"001001001",
  49686=>"110101000",
  49687=>"111111111",
  49688=>"111111000",
  49689=>"110110100",
  49690=>"000000000",
  49691=>"001001001",
  49692=>"000000000",
  49693=>"111111111",
  49694=>"000000000",
  49695=>"000000000",
  49696=>"000001111",
  49697=>"111110100",
  49698=>"111111110",
  49699=>"111000000",
  49700=>"100000111",
  49701=>"111111000",
  49702=>"001001000",
  49703=>"001111111",
  49704=>"111111111",
  49705=>"000111111",
  49706=>"000000000",
  49707=>"000010000",
  49708=>"011111011",
  49709=>"000000000",
  49710=>"011011101",
  49711=>"111111111",
  49712=>"000000000",
  49713=>"100100101",
  49714=>"110000000",
  49715=>"001000000",
  49716=>"011011011",
  49717=>"000001101",
  49718=>"111111110",
  49719=>"110110110",
  49720=>"000000000",
  49721=>"001111001",
  49722=>"000111111",
  49723=>"111011000",
  49724=>"000000000",
  49725=>"001000000",
  49726=>"111001000",
  49727=>"001010000",
  49728=>"001001001",
  49729=>"010010010",
  49730=>"100110110",
  49731=>"111111001",
  49732=>"111100111",
  49733=>"001001100",
  49734=>"111111111",
  49735=>"000001111",
  49736=>"001000001",
  49737=>"001001011",
  49738=>"111111111",
  49739=>"000000001",
  49740=>"000001000",
  49741=>"110110000",
  49742=>"000000100",
  49743=>"111111111",
  49744=>"111001011",
  49745=>"001111111",
  49746=>"000000000",
  49747=>"001001000",
  49748=>"111111001",
  49749=>"011000111",
  49750=>"111101111",
  49751=>"111111111",
  49752=>"001101101",
  49753=>"000000010",
  49754=>"000000000",
  49755=>"111111010",
  49756=>"000000000",
  49757=>"011011000",
  49758=>"011011000",
  49759=>"001011000",
  49760=>"011000001",
  49761=>"000100100",
  49762=>"000000011",
  49763=>"110110000",
  49764=>"111100100",
  49765=>"000000000",
  49766=>"111000010",
  49767=>"111111111",
  49768=>"110110000",
  49769=>"100001111",
  49770=>"000000000",
  49771=>"010011010",
  49772=>"111001000",
  49773=>"000000011",
  49774=>"000000000",
  49775=>"111111111",
  49776=>"011011000",
  49777=>"000000000",
  49778=>"111111111",
  49779=>"000000000",
  49780=>"100111011",
  49781=>"101111111",
  49782=>"000000000",
  49783=>"111111111",
  49784=>"000111111",
  49785=>"111001000",
  49786=>"000000011",
  49787=>"000100000",
  49788=>"110010110",
  49789=>"000000000",
  49790=>"111111111",
  49791=>"000111111",
  49792=>"111111111",
  49793=>"111111011",
  49794=>"111001000",
  49795=>"000000000",
  49796=>"000000000",
  49797=>"001000011",
  49798=>"011111000",
  49799=>"111011000",
  49800=>"000000011",
  49801=>"000110111",
  49802=>"101110100",
  49803=>"011001000",
  49804=>"011000000",
  49805=>"110110100",
  49806=>"111111111",
  49807=>"110111000",
  49808=>"111111001",
  49809=>"011001000",
  49810=>"000000000",
  49811=>"001000000",
  49812=>"000000000",
  49813=>"111111111",
  49814=>"111111111",
  49815=>"011111011",
  49816=>"011000000",
  49817=>"001000000",
  49818=>"000000000",
  49819=>"110111111",
  49820=>"000000000",
  49821=>"100001001",
  49822=>"000000000",
  49823=>"000000000",
  49824=>"011000000",
  49825=>"000000101",
  49826=>"000000000",
  49827=>"000111111",
  49828=>"110111101",
  49829=>"111011111",
  49830=>"101000000",
  49831=>"001101001",
  49832=>"001000000",
  49833=>"000000000",
  49834=>"000001010",
  49835=>"111111111",
  49836=>"111111111",
  49837=>"010110110",
  49838=>"011011000",
  49839=>"111000101",
  49840=>"111111111",
  49841=>"101101111",
  49842=>"001101001",
  49843=>"000000111",
  49844=>"000010011",
  49845=>"111110101",
  49846=>"111111011",
  49847=>"111111100",
  49848=>"000101110",
  49849=>"001000000",
  49850=>"011000000",
  49851=>"001010100",
  49852=>"010000000",
  49853=>"111001101",
  49854=>"110000000",
  49855=>"000001000",
  49856=>"111011111",
  49857=>"000000000",
  49858=>"000111111",
  49859=>"000000000",
  49860=>"011111111",
  49861=>"000000000",
  49862=>"111111111",
  49863=>"001101111",
  49864=>"000110111",
  49865=>"111111111",
  49866=>"000111111",
  49867=>"111011001",
  49868=>"000000000",
  49869=>"111001001",
  49870=>"000000000",
  49871=>"000000000",
  49872=>"111110100",
  49873=>"111111111",
  49874=>"100000101",
  49875=>"000000000",
  49876=>"111111111",
  49877=>"100101111",
  49878=>"011000000",
  49879=>"000000000",
  49880=>"011000010",
  49881=>"111111110",
  49882=>"011111111",
  49883=>"111111111",
  49884=>"110111001",
  49885=>"111111111",
  49886=>"000000000",
  49887=>"001101010",
  49888=>"000000000",
  49889=>"000010000",
  49890=>"111111011",
  49891=>"111000000",
  49892=>"000111111",
  49893=>"001000011",
  49894=>"111111111",
  49895=>"011001001",
  49896=>"111111111",
  49897=>"111111111",
  49898=>"110110110",
  49899=>"000011111",
  49900=>"100000000",
  49901=>"000000001",
  49902=>"111111000",
  49903=>"000000000",
  49904=>"111000000",
  49905=>"111100111",
  49906=>"110110001",
  49907=>"001001001",
  49908=>"111111111",
  49909=>"110110110",
  49910=>"001000000",
  49911=>"111111001",
  49912=>"000000110",
  49913=>"000000000",
  49914=>"000011111",
  49915=>"101110000",
  49916=>"000001111",
  49917=>"000000000",
  49918=>"000101011",
  49919=>"000100000",
  49920=>"111001000",
  49921=>"001111001",
  49922=>"110111111",
  49923=>"111111111",
  49924=>"111111111",
  49925=>"110110111",
  49926=>"111111100",
  49927=>"000001000",
  49928=>"001001000",
  49929=>"000000000",
  49930=>"000000000",
  49931=>"001000000",
  49932=>"110000010",
  49933=>"011011001",
  49934=>"111100000",
  49935=>"110000000",
  49936=>"000000000",
  49937=>"100000111",
  49938=>"111111111",
  49939=>"000000000",
  49940=>"000000100",
  49941=>"000000000",
  49942=>"000000000",
  49943=>"000000001",
  49944=>"000000000",
  49945=>"000000000",
  49946=>"000000000",
  49947=>"111110000",
  49948=>"000000000",
  49949=>"000000000",
  49950=>"000000000",
  49951=>"111000000",
  49952=>"001000000",
  49953=>"011011111",
  49954=>"000000000",
  49955=>"000000000",
  49956=>"111111111",
  49957=>"000000111",
  49958=>"111000000",
  49959=>"000000110",
  49960=>"111101000",
  49961=>"100111111",
  49962=>"000000000",
  49963=>"000000000",
  49964=>"000000000",
  49965=>"110110100",
  49966=>"000111000",
  49967=>"000000000",
  49968=>"000000000",
  49969=>"000000000",
  49970=>"000000001",
  49971=>"110000000",
  49972=>"000000000",
  49973=>"011011001",
  49974=>"000000000",
  49975=>"000000000",
  49976=>"001000000",
  49977=>"111111111",
  49978=>"111111111",
  49979=>"000000000",
  49980=>"000111000",
  49981=>"001001111",
  49982=>"111111101",
  49983=>"110110000",
  49984=>"010010000",
  49985=>"000000000",
  49986=>"001111111",
  49987=>"011111111",
  49988=>"011000000",
  49989=>"111111111",
  49990=>"111101111",
  49991=>"111101111",
  49992=>"100000001",
  49993=>"111111111",
  49994=>"000000000",
  49995=>"000000001",
  49996=>"111110110",
  49997=>"000000000",
  49998=>"111000000",
  49999=>"111111111",
  50000=>"111001101",
  50001=>"111111111",
  50002=>"111111001",
  50003=>"111110111",
  50004=>"111111110",
  50005=>"001000001",
  50006=>"011011000",
  50007=>"000001111",
  50008=>"111111110",
  50009=>"000010000",
  50010=>"011111100",
  50011=>"011111001",
  50012=>"111110000",
  50013=>"111111111",
  50014=>"110111111",
  50015=>"110000011",
  50016=>"000000100",
  50017=>"000000101",
  50018=>"000000000",
  50019=>"000000111",
  50020=>"000001101",
  50021=>"001000000",
  50022=>"000000111",
  50023=>"001000000",
  50024=>"111110100",
  50025=>"011000111",
  50026=>"111101100",
  50027=>"000000000",
  50028=>"000000000",
  50029=>"001001000",
  50030=>"000000000",
  50031=>"000011001",
  50032=>"000000000",
  50033=>"100110111",
  50034=>"111111111",
  50035=>"100100111",
  50036=>"100100001",
  50037=>"000001000",
  50038=>"111110000",
  50039=>"000000011",
  50040=>"111111111",
  50041=>"000000000",
  50042=>"000011111",
  50043=>"111111111",
  50044=>"100000100",
  50045=>"011011111",
  50046=>"110111111",
  50047=>"000000110",
  50048=>"111111000",
  50049=>"011010010",
  50050=>"100111101",
  50051=>"000000000",
  50052=>"000000000",
  50053=>"000000000",
  50054=>"110111111",
  50055=>"000000000",
  50056=>"111111111",
  50057=>"111111110",
  50058=>"111011111",
  50059=>"000011111",
  50060=>"111111111",
  50061=>"111111111",
  50062=>"011001000",
  50063=>"000000000",
  50064=>"010000000",
  50065=>"001001001",
  50066=>"011111111",
  50067=>"111111111",
  50068=>"111111111",
  50069=>"000011011",
  50070=>"000000101",
  50071=>"101101000",
  50072=>"000001001",
  50073=>"111111000",
  50074=>"111111111",
  50075=>"000100100",
  50076=>"111111111",
  50077=>"000000000",
  50078=>"111000011",
  50079=>"000000000",
  50080=>"000000000",
  50081=>"011111011",
  50082=>"000000000",
  50083=>"111111111",
  50084=>"011111111",
  50085=>"011111001",
  50086=>"111111111",
  50087=>"111111111",
  50088=>"000000000",
  50089=>"001110111",
  50090=>"001001000",
  50091=>"100000100",
  50092=>"010111001",
  50093=>"000000000",
  50094=>"000111111",
  50095=>"111111111",
  50096=>"111111011",
  50097=>"111110111",
  50098=>"000001011",
  50099=>"111111110",
  50100=>"111111100",
  50101=>"111111111",
  50102=>"000000000",
  50103=>"000000000",
  50104=>"111010000",
  50105=>"000010100",
  50106=>"000000000",
  50107=>"011111111",
  50108=>"111010000",
  50109=>"001001000",
  50110=>"000000000",
  50111=>"101101000",
  50112=>"111101110",
  50113=>"111111111",
  50114=>"000111111",
  50115=>"111111111",
  50116=>"111101111",
  50117=>"001001000",
  50118=>"011111111",
  50119=>"001011001",
  50120=>"001001011",
  50121=>"110101011",
  50122=>"111001111",
  50123=>"000000001",
  50124=>"110111000",
  50125=>"000001001",
  50126=>"000000000",
  50127=>"100000000",
  50128=>"110110111",
  50129=>"000000000",
  50130=>"110010110",
  50131=>"111111111",
  50132=>"011000000",
  50133=>"111111000",
  50134=>"010000101",
  50135=>"001001001",
  50136=>"000000000",
  50137=>"010111111",
  50138=>"111111111",
  50139=>"111001000",
  50140=>"010010011",
  50141=>"011011111",
  50142=>"000000000",
  50143=>"101101111",
  50144=>"011111111",
  50145=>"000001111",
  50146=>"000000000",
  50147=>"111111111",
  50148=>"000001111",
  50149=>"110110110",
  50150=>"011100110",
  50151=>"000111111",
  50152=>"001000100",
  50153=>"111001000",
  50154=>"011011000",
  50155=>"111111111",
  50156=>"100000110",
  50157=>"001001001",
  50158=>"000000110",
  50159=>"100110111",
  50160=>"100000000",
  50161=>"000110111",
  50162=>"111001111",
  50163=>"010000000",
  50164=>"000000111",
  50165=>"001011111",
  50166=>"011000000",
  50167=>"000100100",
  50168=>"000000000",
  50169=>"010000000",
  50170=>"100000000",
  50171=>"111111111",
  50172=>"000000000",
  50173=>"000001001",
  50174=>"001001001",
  50175=>"001000001",
  50176=>"111111111",
  50177=>"111000000",
  50178=>"001111111",
  50179=>"000000100",
  50180=>"111111000",
  50181=>"111110111",
  50182=>"000000000",
  50183=>"111011111",
  50184=>"111000111",
  50185=>"001111111",
  50186=>"111000000",
  50187=>"111111111",
  50188=>"000010001",
  50189=>"111111111",
  50190=>"110100111",
  50191=>"111111000",
  50192=>"001011111",
  50193=>"000010111",
  50194=>"000100111",
  50195=>"000101111",
  50196=>"111000000",
  50197=>"111000111",
  50198=>"111111111",
  50199=>"110110111",
  50200=>"000000001",
  50201=>"000010010",
  50202=>"010000000",
  50203=>"111100111",
  50204=>"000000000",
  50205=>"111111111",
  50206=>"111111111",
  50207=>"001111110",
  50208=>"000111000",
  50209=>"110110110",
  50210=>"101000101",
  50211=>"111111111",
  50212=>"000111000",
  50213=>"000001111",
  50214=>"010000000",
  50215=>"111011111",
  50216=>"111111110",
  50217=>"000101111",
  50218=>"011111111",
  50219=>"111111111",
  50220=>"101000000",
  50221=>"000001011",
  50222=>"110110000",
  50223=>"111111111",
  50224=>"110000000",
  50225=>"000000001",
  50226=>"000000000",
  50227=>"000000111",
  50228=>"010011010",
  50229=>"010010111",
  50230=>"000000111",
  50231=>"000100111",
  50232=>"111110000",
  50233=>"000101100",
  50234=>"111000000",
  50235=>"000110000",
  50236=>"000000001",
  50237=>"111111001",
  50238=>"000000111",
  50239=>"110000000",
  50240=>"000100110",
  50241=>"001001000",
  50242=>"111111011",
  50243=>"110111111",
  50244=>"000101111",
  50245=>"111110111",
  50246=>"000000111",
  50247=>"100110110",
  50248=>"000110111",
  50249=>"000001111",
  50250=>"010011011",
  50251=>"000000111",
  50252=>"110110011",
  50253=>"001111001",
  50254=>"111111111",
  50255=>"111000101",
  50256=>"111111111",
  50257=>"111111111",
  50258=>"000010011",
  50259=>"110111111",
  50260=>"000000110",
  50261=>"111000000",
  50262=>"000000000",
  50263=>"100000000",
  50264=>"111111111",
  50265=>"000000000",
  50266=>"000000111",
  50267=>"100100100",
  50268=>"000000000",
  50269=>"110100100",
  50270=>"000000000",
  50271=>"100100100",
  50272=>"000110000",
  50273=>"111000000",
  50274=>"001000111",
  50275=>"111000000",
  50276=>"000100110",
  50277=>"000000000",
  50278=>"000000111",
  50279=>"000000010",
  50280=>"100111111",
  50281=>"000011111",
  50282=>"000110000",
  50283=>"000101111",
  50284=>"100000110",
  50285=>"100100000",
  50286=>"111000111",
  50287=>"111111010",
  50288=>"111111000",
  50289=>"111011111",
  50290=>"110110110",
  50291=>"000000000",
  50292=>"011001001",
  50293=>"110110111",
  50294=>"000000111",
  50295=>"111110110",
  50296=>"111000000",
  50297=>"000000010",
  50298=>"000000000",
  50299=>"000000011",
  50300=>"000011111",
  50301=>"000000000",
  50302=>"000000000",
  50303=>"000000000",
  50304=>"000000000",
  50305=>"111111111",
  50306=>"111000000",
  50307=>"011111000",
  50308=>"100100100",
  50309=>"000000000",
  50310=>"000110001",
  50311=>"000000000",
  50312=>"000111111",
  50313=>"001000000",
  50314=>"111000000",
  50315=>"000011111",
  50316=>"000111111",
  50317=>"111111111",
  50318=>"000000000",
  50319=>"111111101",
  50320=>"000000111",
  50321=>"010010010",
  50322=>"000000000",
  50323=>"000000000",
  50324=>"000110111",
  50325=>"001111110",
  50326=>"111101001",
  50327=>"100100100",
  50328=>"000000100",
  50329=>"000000000",
  50330=>"001101111",
  50331=>"000000000",
  50332=>"100100111",
  50333=>"100010111",
  50334=>"011111111",
  50335=>"100000000",
  50336=>"111111010",
  50337=>"111100111",
  50338=>"000000001",
  50339=>"000011111",
  50340=>"100100100",
  50341=>"010110101",
  50342=>"111111111",
  50343=>"111001001",
  50344=>"000111001",
  50345=>"110010010",
  50346=>"000000000",
  50347=>"000000111",
  50348=>"000000000",
  50349=>"001001000",
  50350=>"000000000",
  50351=>"000000000",
  50352=>"000000000",
  50353=>"000010110",
  50354=>"111111111",
  50355=>"111000000",
  50356=>"100100000",
  50357=>"111101001",
  50358=>"000000001",
  50359=>"000011000",
  50360=>"101111111",
  50361=>"111001111",
  50362=>"100110101",
  50363=>"000000101",
  50364=>"111010000",
  50365=>"111111001",
  50366=>"111111111",
  50367=>"000000000",
  50368=>"000001111",
  50369=>"000000000",
  50370=>"011111000",
  50371=>"000000000",
  50372=>"001001111",
  50373=>"111000110",
  50374=>"000000000",
  50375=>"000000000",
  50376=>"100000000",
  50377=>"111111000",
  50378=>"000100100",
  50379=>"110000000",
  50380=>"000000000",
  50381=>"111111110",
  50382=>"001111011",
  50383=>"000000110",
  50384=>"100100000",
  50385=>"111000000",
  50386=>"011000000",
  50387=>"100000000",
  50388=>"011011010",
  50389=>"111111100",
  50390=>"111111111",
  50391=>"100000011",
  50392=>"011110111",
  50393=>"111111001",
  50394=>"000000000",
  50395=>"111001000",
  50396=>"000000000",
  50397=>"000000000",
  50398=>"000000111",
  50399=>"111101001",
  50400=>"011000000",
  50401=>"111101111",
  50402=>"111111111",
  50403=>"000000000",
  50404=>"001111111",
  50405=>"000000000",
  50406=>"000000000",
  50407=>"101000001",
  50408=>"001001000",
  50409=>"100100111",
  50410=>"111100100",
  50411=>"111000011",
  50412=>"000000000",
  50413=>"111101000",
  50414=>"000100100",
  50415=>"111000000",
  50416=>"110111000",
  50417=>"111100000",
  50418=>"111111111",
  50419=>"111111111",
  50420=>"000000000",
  50421=>"000011001",
  50422=>"000111000",
  50423=>"111111111",
  50424=>"001111111",
  50425=>"111111010",
  50426=>"000000000",
  50427=>"000000010",
  50428=>"101100100",
  50429=>"000010111",
  50430=>"001111111",
  50431=>"100001000",
  50432=>"101101101",
  50433=>"001100111",
  50434=>"010010111",
  50435=>"000000000",
  50436=>"111011000",
  50437=>"000000111",
  50438=>"100000000",
  50439=>"011011110",
  50440=>"000000111",
  50441=>"000000111",
  50442=>"110110111",
  50443=>"000111111",
  50444=>"111101101",
  50445=>"000000000",
  50446=>"000001111",
  50447=>"000100000",
  50448=>"000000111",
  50449=>"000000111",
  50450=>"111001000",
  50451=>"000111111",
  50452=>"000101000",
  50453=>"010111111",
  50454=>"110110000",
  50455=>"000010111",
  50456=>"111011110",
  50457=>"000011001",
  50458=>"001000010",
  50459=>"110000000",
  50460=>"111111111",
  50461=>"111100000",
  50462=>"001111011",
  50463=>"000111111",
  50464=>"011100110",
  50465=>"001011111",
  50466=>"111111111",
  50467=>"110100000",
  50468=>"110111111",
  50469=>"000000000",
  50470=>"000110100",
  50471=>"111111010",
  50472=>"001001000",
  50473=>"011011001",
  50474=>"111000001",
  50475=>"111111000",
  50476=>"100100000",
  50477=>"111101111",
  50478=>"000000000",
  50479=>"000111111",
  50480=>"010111111",
  50481=>"000000000",
  50482=>"111111111",
  50483=>"000110110",
  50484=>"000000000",
  50485=>"111000000",
  50486=>"000000110",
  50487=>"111111101",
  50488=>"111000000",
  50489=>"110000101",
  50490=>"111101111",
  50491=>"111111111",
  50492=>"000000111",
  50493=>"001101000",
  50494=>"100000000",
  50495=>"010110000",
  50496=>"000000111",
  50497=>"100111111",
  50498=>"000000000",
  50499=>"001000011",
  50500=>"111001111",
  50501=>"111111111",
  50502=>"111111111",
  50503=>"110100000",
  50504=>"111100111",
  50505=>"000000000",
  50506=>"110110011",
  50507=>"100000100",
  50508=>"000101111",
  50509=>"000000011",
  50510=>"000111011",
  50511=>"111111110",
  50512=>"110110100",
  50513=>"001111000",
  50514=>"000000000",
  50515=>"111111000",
  50516=>"111111111",
  50517=>"111110111",
  50518=>"110111111",
  50519=>"000000000",
  50520=>"000111111",
  50521=>"101101111",
  50522=>"000000000",
  50523=>"111111111",
  50524=>"111111011",
  50525=>"001000000",
  50526=>"111000000",
  50527=>"000001111",
  50528=>"000000011",
  50529=>"000000000",
  50530=>"111111111",
  50531=>"111001001",
  50532=>"111111100",
  50533=>"000000000",
  50534=>"111111111",
  50535=>"100000111",
  50536=>"011000110",
  50537=>"000000000",
  50538=>"011000000",
  50539=>"000000010",
  50540=>"000001011",
  50541=>"100100110",
  50542=>"111111011",
  50543=>"000000000",
  50544=>"111111111",
  50545=>"101111100",
  50546=>"111100000",
  50547=>"001000000",
  50548=>"111111100",
  50549=>"111110011",
  50550=>"000000000",
  50551=>"000001111",
  50552=>"000000000",
  50553=>"111111000",
  50554=>"000000000",
  50555=>"000000000",
  50556=>"100000000",
  50557=>"000000000",
  50558=>"011000011",
  50559=>"000000000",
  50560=>"111111011",
  50561=>"111001001",
  50562=>"111111111",
  50563=>"111000000",
  50564=>"111111110",
  50565=>"111100111",
  50566=>"000000000",
  50567=>"111111000",
  50568=>"000000110",
  50569=>"111000000",
  50570=>"000000100",
  50571=>"000001101",
  50572=>"000000111",
  50573=>"000000111",
  50574=>"000000001",
  50575=>"010000000",
  50576=>"111111111",
  50577=>"101001001",
  50578=>"001111111",
  50579=>"000100000",
  50580=>"111111111",
  50581=>"000110000",
  50582=>"111111111",
  50583=>"110100111",
  50584=>"111111111",
  50585=>"000100100",
  50586=>"000000001",
  50587=>"110100000",
  50588=>"100000011",
  50589=>"111111011",
  50590=>"000100111",
  50591=>"000000101",
  50592=>"111100000",
  50593=>"110110110",
  50594=>"111001000",
  50595=>"000000101",
  50596=>"110000000",
  50597=>"111000000",
  50598=>"000111111",
  50599=>"111111000",
  50600=>"000000000",
  50601=>"000100101",
  50602=>"111000000",
  50603=>"010111111",
  50604=>"000000000",
  50605=>"001011011",
  50606=>"011011000",
  50607=>"111111000",
  50608=>"000000111",
  50609=>"000000000",
  50610=>"011111111",
  50611=>"000001000",
  50612=>"000111111",
  50613=>"101011001",
  50614=>"111111111",
  50615=>"000000000",
  50616=>"000000000",
  50617=>"000000001",
  50618=>"000000000",
  50619=>"000000000",
  50620=>"111111111",
  50621=>"001001001",
  50622=>"111111110",
  50623=>"011000111",
  50624=>"111101101",
  50625=>"111011000",
  50626=>"010010000",
  50627=>"000001000",
  50628=>"000000000",
  50629=>"000000000",
  50630=>"010111111",
  50631=>"000000111",
  50632=>"000000100",
  50633=>"000111111",
  50634=>"000000000",
  50635=>"000110111",
  50636=>"000000010",
  50637=>"011111111",
  50638=>"000111111",
  50639=>"111011000",
  50640=>"100111111",
  50641=>"000111111",
  50642=>"000001110",
  50643=>"110000000",
  50644=>"111111111",
  50645=>"000000000",
  50646=>"000000111",
  50647=>"001000001",
  50648=>"000000000",
  50649=>"111111111",
  50650=>"000111111",
  50651=>"000000001",
  50652=>"000011011",
  50653=>"111011000",
  50654=>"111110111",
  50655=>"111011001",
  50656=>"010111111",
  50657=>"100000000",
  50658=>"000000001",
  50659=>"001000011",
  50660=>"000000000",
  50661=>"000001101",
  50662=>"111111000",
  50663=>"101000111",
  50664=>"000000011",
  50665=>"111111110",
  50666=>"111000000",
  50667=>"000000111",
  50668=>"100000111",
  50669=>"010000000",
  50670=>"011011011",
  50671=>"010000000",
  50672=>"110110100",
  50673=>"111111000",
  50674=>"000110101",
  50675=>"000000010",
  50676=>"111000000",
  50677=>"011000000",
  50678=>"001000000",
  50679=>"000001111",
  50680=>"000111111",
  50681=>"111100000",
  50682=>"111111100",
  50683=>"111111101",
  50684=>"010110111",
  50685=>"111111111",
  50686=>"000000011",
  50687=>"000000000",
  50688=>"111111110",
  50689=>"100100000",
  50690=>"111000000",
  50691=>"100000110",
  50692=>"001010110",
  50693=>"100110100",
  50694=>"000000000",
  50695=>"100111111",
  50696=>"111110010",
  50697=>"111111111",
  50698=>"000000111",
  50699=>"011111111",
  50700=>"000000000",
  50701=>"111111000",
  50702=>"000111111",
  50703=>"111111111",
  50704=>"110100101",
  50705=>"010100010",
  50706=>"000000000",
  50707=>"111111110",
  50708=>"000100100",
  50709=>"011000000",
  50710=>"000100111",
  50711=>"011011011",
  50712=>"101000101",
  50713=>"100101001",
  50714=>"111100000",
  50715=>"000101110",
  50716=>"111111011",
  50717=>"111000000",
  50718=>"001111111",
  50719=>"000111111",
  50720=>"000000010",
  50721=>"110010110",
  50722=>"011001001",
  50723=>"011001110",
  50724=>"000000000",
  50725=>"111111111",
  50726=>"000011111",
  50727=>"000000000",
  50728=>"111110111",
  50729=>"001000000",
  50730=>"001001001",
  50731=>"111111111",
  50732=>"111111111",
  50733=>"111011000",
  50734=>"000000000",
  50735=>"000000000",
  50736=>"000101111",
  50737=>"011001000",
  50738=>"111001001",
  50739=>"000000000",
  50740=>"000000011",
  50741=>"100101011",
  50742=>"111111111",
  50743=>"111111011",
  50744=>"000111111",
  50745=>"110111001",
  50746=>"111000000",
  50747=>"111111110",
  50748=>"111111000",
  50749=>"111001000",
  50750=>"011001000",
  50751=>"111111011",
  50752=>"111111111",
  50753=>"010011111",
  50754=>"001111111",
  50755=>"000000100",
  50756=>"001011111",
  50757=>"010000000",
  50758=>"000011111",
  50759=>"110000111",
  50760=>"111011011",
  50761=>"111111001",
  50762=>"000110111",
  50763=>"100101011",
  50764=>"100100100",
  50765=>"101000000",
  50766=>"000100111",
  50767=>"111110011",
  50768=>"111111111",
  50769=>"110101001",
  50770=>"001000111",
  50771=>"000000000",
  50772=>"111111111",
  50773=>"111111000",
  50774=>"000000000",
  50775=>"100110110",
  50776=>"010110110",
  50777=>"111101000",
  50778=>"000000110",
  50779=>"100111110",
  50780=>"000111110",
  50781=>"001111111",
  50782=>"100000101",
  50783=>"000000000",
  50784=>"011010010",
  50785=>"110111111",
  50786=>"111011000",
  50787=>"001111111",
  50788=>"001000011",
  50789=>"100000100",
  50790=>"111011111",
  50791=>"000000000",
  50792=>"000000011",
  50793=>"000000000",
  50794=>"000001111",
  50795=>"010010000",
  50796=>"111011110",
  50797=>"000010000",
  50798=>"111001000",
  50799=>"000010110",
  50800=>"111011111",
  50801=>"111111011",
  50802=>"000000001",
  50803=>"000001011",
  50804=>"111111111",
  50805=>"000000111",
  50806=>"111011011",
  50807=>"000000000",
  50808=>"101100001",
  50809=>"111111111",
  50810=>"000000011",
  50811=>"111111000",
  50812=>"101101101",
  50813=>"001011001",
  50814=>"000000100",
  50815=>"011000000",
  50816=>"111100000",
  50817=>"111000000",
  50818=>"000000111",
  50819=>"100000111",
  50820=>"011100111",
  50821=>"111010111",
  50822=>"000000110",
  50823=>"000000000",
  50824=>"111000000",
  50825=>"101100100",
  50826=>"000000001",
  50827=>"111011111",
  50828=>"111000000",
  50829=>"100111101",
  50830=>"111101000",
  50831=>"011000101",
  50832=>"000000000",
  50833=>"111111111",
  50834=>"111101000",
  50835=>"000001011",
  50836=>"110001001",
  50837=>"000000111",
  50838=>"111000000",
  50839=>"111101111",
  50840=>"001000000",
  50841=>"111111111",
  50842=>"000000110",
  50843=>"111111111",
  50844=>"000000111",
  50845=>"001001001",
  50846=>"111111111",
  50847=>"001000000",
  50848=>"010000000",
  50849=>"111101101",
  50850=>"111100000",
  50851=>"111111111",
  50852=>"000000000",
  50853=>"111111111",
  50854=>"111001111",
  50855=>"011110100",
  50856=>"000001111",
  50857=>"000101101",
  50858=>"001000111",
  50859=>"110110111",
  50860=>"111111111",
  50861=>"100111111",
  50862=>"000000111",
  50863=>"101111111",
  50864=>"000000111",
  50865=>"001111111",
  50866=>"010111111",
  50867=>"000000000",
  50868=>"101000000",
  50869=>"000000011",
  50870=>"000000011",
  50871=>"000000000",
  50872=>"111111111",
  50873=>"111111111",
  50874=>"101000001",
  50875=>"001001001",
  50876=>"111100111",
  50877=>"001001000",
  50878=>"000010111",
  50879=>"000000000",
  50880=>"000000000",
  50881=>"111111111",
  50882=>"001001010",
  50883=>"000111111",
  50884=>"000000001",
  50885=>"111111111",
  50886=>"000111111",
  50887=>"101101100",
  50888=>"000001111",
  50889=>"111000011",
  50890=>"001000111",
  50891=>"000000000",
  50892=>"100111111",
  50893=>"000000000",
  50894=>"001001000",
  50895=>"000000000",
  50896=>"100000111",
  50897=>"001000000",
  50898=>"000100110",
  50899=>"000000000",
  50900=>"111000000",
  50901=>"110000101",
  50902=>"111001000",
  50903=>"101111011",
  50904=>"000011000",
  50905=>"111111111",
  50906=>"000000000",
  50907=>"001111111",
  50908=>"000010000",
  50909=>"111110111",
  50910=>"000000011",
  50911=>"100100001",
  50912=>"111000000",
  50913=>"000000000",
  50914=>"000000000",
  50915=>"111001000",
  50916=>"111100100",
  50917=>"000000100",
  50918=>"000000000",
  50919=>"111111111",
  50920=>"001000010",
  50921=>"000100000",
  50922=>"111110000",
  50923=>"011000000",
  50924=>"000000000",
  50925=>"111001000",
  50926=>"111001001",
  50927=>"111000000",
  50928=>"000000011",
  50929=>"111111100",
  50930=>"110000000",
  50931=>"000000000",
  50932=>"000000110",
  50933=>"000001000",
  50934=>"000111100",
  50935=>"000000000",
  50936=>"111110110",
  50937=>"000011011",
  50938=>"111001001",
  50939=>"101111111",
  50940=>"111111111",
  50941=>"111111111",
  50942=>"000001111",
  50943=>"001000000",
  50944=>"101111111",
  50945=>"111100110",
  50946=>"011111111",
  50947=>"101000000",
  50948=>"000001111",
  50949=>"001001011",
  50950=>"000000010",
  50951=>"000000001",
  50952=>"000000011",
  50953=>"111111111",
  50954=>"111100000",
  50955=>"011000111",
  50956=>"110111111",
  50957=>"111011001",
  50958=>"001000111",
  50959=>"111111111",
  50960=>"000000111",
  50961=>"000000001",
  50962=>"111110011",
  50963=>"111000000",
  50964=>"010111000",
  50965=>"000000111",
  50966=>"100000111",
  50967=>"000000000",
  50968=>"111111111",
  50969=>"000000001",
  50970=>"000001111",
  50971=>"000111111",
  50972=>"001101110",
  50973=>"011111111",
  50974=>"111111111",
  50975=>"010011111",
  50976=>"100111000",
  50977=>"001111111",
  50978=>"000111110",
  50979=>"111111000",
  50980=>"111000000",
  50981=>"100000000",
  50982=>"111111100",
  50983=>"000001000",
  50984=>"001110100",
  50985=>"011011011",
  50986=>"001100100",
  50987=>"000000000",
  50988=>"000000111",
  50989=>"101111111",
  50990=>"000000000",
  50991=>"000000000",
  50992=>"111101101",
  50993=>"111111111",
  50994=>"000111111",
  50995=>"111000000",
  50996=>"110000000",
  50997=>"000100001",
  50998=>"000000000",
  50999=>"000000000",
  51000=>"000000000",
  51001=>"000111111",
  51002=>"111001000",
  51003=>"111111000",
  51004=>"110000101",
  51005=>"100000100",
  51006=>"000000001",
  51007=>"011111111",
  51008=>"111101011",
  51009=>"000000011",
  51010=>"111111111",
  51011=>"111001000",
  51012=>"111101101",
  51013=>"111001001",
  51014=>"000111001",
  51015=>"000000100",
  51016=>"000000111",
  51017=>"000000111",
  51018=>"101001000",
  51019=>"111011000",
  51020=>"000001111",
  51021=>"111100000",
  51022=>"000000000",
  51023=>"001011001",
  51024=>"000111111",
  51025=>"100000000",
  51026=>"111111111",
  51027=>"010110100",
  51028=>"000000000",
  51029=>"011000100",
  51030=>"111000000",
  51031=>"111011111",
  51032=>"101000110",
  51033=>"000000111",
  51034=>"111111111",
  51035=>"111000111",
  51036=>"111000000",
  51037=>"000000011",
  51038=>"000001000",
  51039=>"101111111",
  51040=>"111111000",
  51041=>"000000000",
  51042=>"101111001",
  51043=>"100000000",
  51044=>"000011111",
  51045=>"001000000",
  51046=>"110100000",
  51047=>"111111111",
  51048=>"111111001",
  51049=>"100111111",
  51050=>"111111111",
  51051=>"111111110",
  51052=>"000110110",
  51053=>"000100111",
  51054=>"011011011",
  51055=>"011000000",
  51056=>"111111111",
  51057=>"111001111",
  51058=>"000000000",
  51059=>"000100111",
  51060=>"000011110",
  51061=>"001111111",
  51062=>"111101100",
  51063=>"000000101",
  51064=>"111111011",
  51065=>"111000000",
  51066=>"000110111",
  51067=>"110110111",
  51068=>"011111011",
  51069=>"110110111",
  51070=>"000100000",
  51071=>"100100000",
  51072=>"111011011",
  51073=>"000000111",
  51074=>"111110010",
  51075=>"001000101",
  51076=>"000000111",
  51077=>"110000010",
  51078=>"111111111",
  51079=>"111001000",
  51080=>"001000011",
  51081=>"100100100",
  51082=>"111111111",
  51083=>"000111100",
  51084=>"100111111",
  51085=>"111111111",
  51086=>"000110111",
  51087=>"000000111",
  51088=>"000111111",
  51089=>"000000111",
  51090=>"111111000",
  51091=>"111100100",
  51092=>"000000000",
  51093=>"000000101",
  51094=>"111011011",
  51095=>"100000000",
  51096=>"111001011",
  51097=>"101101111",
  51098=>"111111110",
  51099=>"001111011",
  51100=>"001111111",
  51101=>"000011010",
  51102=>"001000000",
  51103=>"000011111",
  51104=>"000000000",
  51105=>"110111001",
  51106=>"011000111",
  51107=>"000000000",
  51108=>"000000000",
  51109=>"011000010",
  51110=>"111110111",
  51111=>"111110111",
  51112=>"001000000",
  51113=>"110100000",
  51114=>"101000000",
  51115=>"110000000",
  51116=>"000000000",
  51117=>"001111101",
  51118=>"101111111",
  51119=>"000000001",
  51120=>"100000000",
  51121=>"111111000",
  51122=>"011011000",
  51123=>"000000000",
  51124=>"000011111",
  51125=>"000111000",
  51126=>"000000111",
  51127=>"000011111",
  51128=>"011000000",
  51129=>"000000010",
  51130=>"000000111",
  51131=>"000111111",
  51132=>"010010111",
  51133=>"000111111",
  51134=>"000000001",
  51135=>"111011111",
  51136=>"000000000",
  51137=>"111111110",
  51138=>"111111111",
  51139=>"101001001",
  51140=>"000000000",
  51141=>"000001001",
  51142=>"100100101",
  51143=>"100000000",
  51144=>"000001011",
  51145=>"000000011",
  51146=>"000000000",
  51147=>"000000111",
  51148=>"000010010",
  51149=>"001111111",
  51150=>"111000000",
  51151=>"011011111",
  51152=>"001111111",
  51153=>"111010000",
  51154=>"000000000",
  51155=>"010010111",
  51156=>"011000001",
  51157=>"111001001",
  51158=>"111111110",
  51159=>"000000011",
  51160=>"100101111",
  51161=>"111111111",
  51162=>"111011011",
  51163=>"001001000",
  51164=>"001001001",
  51165=>"000111111",
  51166=>"111110110",
  51167=>"000000111",
  51168=>"111000110",
  51169=>"001001011",
  51170=>"000000000",
  51171=>"111000001",
  51172=>"111111111",
  51173=>"111111000",
  51174=>"010111111",
  51175=>"011000000",
  51176=>"111111111",
  51177=>"110111100",
  51178=>"101100100",
  51179=>"111110110",
  51180=>"001000000",
  51181=>"001001001",
  51182=>"111001011",
  51183=>"000000011",
  51184=>"111001000",
  51185=>"111110111",
  51186=>"110000000",
  51187=>"111111111",
  51188=>"000000000",
  51189=>"000001001",
  51190=>"000000000",
  51191=>"001001000",
  51192=>"110000010",
  51193=>"000111111",
  51194=>"000000111",
  51195=>"000000000",
  51196=>"111111011",
  51197=>"000000100",
  51198=>"110110100",
  51199=>"000000000",
  51200=>"000001001",
  51201=>"111111111",
  51202=>"110000000",
  51203=>"111111111",
  51204=>"000001000",
  51205=>"100110111",
  51206=>"001000000",
  51207=>"000000000",
  51208=>"111001000",
  51209=>"111010000",
  51210=>"111111110",
  51211=>"001000111",
  51212=>"111101111",
  51213=>"111111111",
  51214=>"010100111",
  51215=>"111000000",
  51216=>"000000000",
  51217=>"000110011",
  51218=>"001000000",
  51219=>"011011111",
  51220=>"000000100",
  51221=>"011000110",
  51222=>"111111011",
  51223=>"111111101",
  51224=>"111100000",
  51225=>"111111111",
  51226=>"011001000",
  51227=>"011111111",
  51228=>"101111111",
  51229=>"010110111",
  51230=>"000111111",
  51231=>"000111001",
  51232=>"000001001",
  51233=>"011111110",
  51234=>"110110111",
  51235=>"011011111",
  51236=>"111110111",
  51237=>"111000000",
  51238=>"111010010",
  51239=>"100001000",
  51240=>"101100000",
  51241=>"010000000",
  51242=>"000000011",
  51243=>"000111111",
  51244=>"111111000",
  51245=>"110111110",
  51246=>"000000000",
  51247=>"111110111",
  51248=>"111111000",
  51249=>"000000000",
  51250=>"100100110",
  51251=>"100100111",
  51252=>"110110000",
  51253=>"111010000",
  51254=>"000000000",
  51255=>"111111000",
  51256=>"000101111",
  51257=>"111111111",
  51258=>"000000000",
  51259=>"111001001",
  51260=>"111000000",
  51261=>"111110100",
  51262=>"111111111",
  51263=>"111111100",
  51264=>"110000010",
  51265=>"111111111",
  51266=>"000000000",
  51267=>"111111110",
  51268=>"000001001",
  51269=>"100000000",
  51270=>"000000000",
  51271=>"000000110",
  51272=>"111111111",
  51273=>"101101111",
  51274=>"111111111",
  51275=>"111111000",
  51276=>"111111111",
  51277=>"101111111",
  51278=>"000000100",
  51279=>"000000111",
  51280=>"111110110",
  51281=>"111010000",
  51282=>"111110010",
  51283=>"100111110",
  51284=>"111111111",
  51285=>"000000000",
  51286=>"011111111",
  51287=>"111111111",
  51288=>"111111111",
  51289=>"111100111",
  51290=>"111010010",
  51291=>"110110111",
  51292=>"000110110",
  51293=>"111111111",
  51294=>"000100111",
  51295=>"000000001",
  51296=>"000111010",
  51297=>"111010000",
  51298=>"011001011",
  51299=>"000000000",
  51300=>"000100100",
  51301=>"000000000",
  51302=>"111111111",
  51303=>"000111111",
  51304=>"111111100",
  51305=>"000000000",
  51306=>"111111111",
  51307=>"000001011",
  51308=>"111111111",
  51309=>"000000110",
  51310=>"000000111",
  51311=>"000000000",
  51312=>"111111001",
  51313=>"000000000",
  51314=>"111110110",
  51315=>"000000000",
  51316=>"011011000",
  51317=>"111111110",
  51318=>"000000111",
  51319=>"001000000",
  51320=>"010010010",
  51321=>"000000000",
  51322=>"000000000",
  51323=>"000010000",
  51324=>"110110110",
  51325=>"111110100",
  51326=>"000000000",
  51327=>"111111111",
  51328=>"111000000",
  51329=>"111101001",
  51330=>"111111111",
  51331=>"000000110",
  51332=>"111111000",
  51333=>"000000001",
  51334=>"111111110",
  51335=>"000000000",
  51336=>"000000000",
  51337=>"110000100",
  51338=>"000000000",
  51339=>"000000101",
  51340=>"111101000",
  51341=>"000000001",
  51342=>"111111000",
  51343=>"000000001",
  51344=>"000000000",
  51345=>"100000000",
  51346=>"000010000",
  51347=>"000111111",
  51348=>"111111111",
  51349=>"011011000",
  51350=>"000001111",
  51351=>"101100100",
  51352=>"110000111",
  51353=>"111111000",
  51354=>"101001111",
  51355=>"111111111",
  51356=>"111110111",
  51357=>"000000111",
  51358=>"011111111",
  51359=>"111111111",
  51360=>"111111111",
  51361=>"000100100",
  51362=>"000000000",
  51363=>"111111111",
  51364=>"110110001",
  51365=>"111111110",
  51366=>"001111111",
  51367=>"111111001",
  51368=>"100000100",
  51369=>"000010011",
  51370=>"111000101",
  51371=>"000111111",
  51372=>"011010111",
  51373=>"111111111",
  51374=>"000000100",
  51375=>"111001001",
  51376=>"111110000",
  51377=>"111111111",
  51378=>"011111111",
  51379=>"000000001",
  51380=>"111111111",
  51381=>"000000011",
  51382=>"000000111",
  51383=>"011011111",
  51384=>"000000111",
  51385=>"100100111",
  51386=>"000110000",
  51387=>"111011011",
  51388=>"111100111",
  51389=>"111101111",
  51390=>"111111111",
  51391=>"111101011",
  51392=>"001000110",
  51393=>"011001001",
  51394=>"111111111",
  51395=>"111101101",
  51396=>"111111111",
  51397=>"111111111",
  51398=>"000000000",
  51399=>"000000000",
  51400=>"111111111",
  51401=>"001001000",
  51402=>"111011110",
  51403=>"000000000",
  51404=>"000000110",
  51405=>"010010110",
  51406=>"111111110",
  51407=>"000000000",
  51408=>"000010000",
  51409=>"110111111",
  51410=>"110111111",
  51411=>"000000011",
  51412=>"001000111",
  51413=>"110110000",
  51414=>"000000000",
  51415=>"000000000",
  51416=>"000000000",
  51417=>"000000000",
  51418=>"000000000",
  51419=>"011000111",
  51420=>"111111111",
  51421=>"111110111",
  51422=>"111011101",
  51423=>"111110000",
  51424=>"000000000",
  51425=>"000000000",
  51426=>"110000000",
  51427=>"000111111",
  51428=>"001000000",
  51429=>"111011101",
  51430=>"000000000",
  51431=>"011111101",
  51432=>"000000000",
  51433=>"011011111",
  51434=>"100101111",
  51435=>"000101100",
  51436=>"111011111",
  51437=>"111111111",
  51438=>"111111100",
  51439=>"000000000",
  51440=>"111111111",
  51441=>"011000000",
  51442=>"111111111",
  51443=>"110111101",
  51444=>"110111111",
  51445=>"000000000",
  51446=>"001000000",
  51447=>"000000000",
  51448=>"111111000",
  51449=>"111111011",
  51450=>"000000111",
  51451=>"110110000",
  51452=>"111111111",
  51453=>"001000000",
  51454=>"011111111",
  51455=>"000001001",
  51456=>"011000001",
  51457=>"011111111",
  51458=>"000011011",
  51459=>"011000000",
  51460=>"111001001",
  51461=>"111100000",
  51462=>"000000000",
  51463=>"000000100",
  51464=>"000000101",
  51465=>"111000000",
  51466=>"111000000",
  51467=>"100000100",
  51468=>"011111001",
  51469=>"111111111",
  51470=>"000000000",
  51471=>"000000000",
  51472=>"000000000",
  51473=>"000000000",
  51474=>"001001000",
  51475=>"100011111",
  51476=>"011011011",
  51477=>"001000000",
  51478=>"011011001",
  51479=>"001001001",
  51480=>"111101000",
  51481=>"000001110",
  51482=>"000000110",
  51483=>"111110110",
  51484=>"111111111",
  51485=>"111111100",
  51486=>"111111111",
  51487=>"100000000",
  51488=>"011011011",
  51489=>"000001001",
  51490=>"000110000",
  51491=>"000000001",
  51492=>"111111111",
  51493=>"111100001",
  51494=>"000100000",
  51495=>"000001000",
  51496=>"111111000",
  51497=>"100010000",
  51498=>"110110101",
  51499=>"111111111",
  51500=>"000000000",
  51501=>"110110000",
  51502=>"111111011",
  51503=>"111100000",
  51504=>"111111110",
  51505=>"100000000",
  51506=>"010110111",
  51507=>"000000000",
  51508=>"111111111",
  51509=>"111011111",
  51510=>"111111011",
  51511=>"110111111",
  51512=>"100100111",
  51513=>"111001000",
  51514=>"111111111",
  51515=>"111111111",
  51516=>"111111111",
  51517=>"000000101",
  51518=>"101111101",
  51519=>"111111111",
  51520=>"000000000",
  51521=>"000110110",
  51522=>"000000100",
  51523=>"000000100",
  51524=>"111001111",
  51525=>"000000000",
  51526=>"100100011",
  51527=>"111000000",
  51528=>"010011010",
  51529=>"111111111",
  51530=>"110000000",
  51531=>"011011000",
  51532=>"111111111",
  51533=>"111111000",
  51534=>"000000011",
  51535=>"111111001",
  51536=>"111101111",
  51537=>"000000000",
  51538=>"001011001",
  51539=>"111111111",
  51540=>"000000000",
  51541=>"001000001",
  51542=>"110111001",
  51543=>"000000000",
  51544=>"000000000",
  51545=>"111111111",
  51546=>"000000000",
  51547=>"000000111",
  51548=>"111001000",
  51549=>"010000111",
  51550=>"111111111",
  51551=>"000000000",
  51552=>"110111011",
  51553=>"000000000",
  51554=>"001111101",
  51555=>"111111111",
  51556=>"001001101",
  51557=>"111111011",
  51558=>"000000111",
  51559=>"000000000",
  51560=>"110100000",
  51561=>"000100000",
  51562=>"111111111",
  51563=>"100110111",
  51564=>"111111110",
  51565=>"000000110",
  51566=>"001111011",
  51567=>"011000000",
  51568=>"000100100",
  51569=>"100000000",
  51570=>"111011000",
  51571=>"000000011",
  51572=>"000000000",
  51573=>"100000100",
  51574=>"111111110",
  51575=>"000000111",
  51576=>"111101111",
  51577=>"000010111",
  51578=>"000110100",
  51579=>"111111011",
  51580=>"000000010",
  51581=>"010010111",
  51582=>"011111111",
  51583=>"101111111",
  51584=>"111001001",
  51585=>"110000000",
  51586=>"011001001",
  51587=>"111111011",
  51588=>"111111100",
  51589=>"000100111",
  51590=>"111111110",
  51591=>"000100000",
  51592=>"011100100",
  51593=>"111111001",
  51594=>"111011001",
  51595=>"111111100",
  51596=>"000000100",
  51597=>"010110111",
  51598=>"100000000",
  51599=>"000000001",
  51600=>"111000000",
  51601=>"111111111",
  51602=>"000000000",
  51603=>"111111111",
  51604=>"000000000",
  51605=>"111111000",
  51606=>"111011111",
  51607=>"100000000",
  51608=>"001000000",
  51609=>"101000111",
  51610=>"001000000",
  51611=>"100110101",
  51612=>"101000100",
  51613=>"111111000",
  51614=>"101000000",
  51615=>"000010110",
  51616=>"000000000",
  51617=>"000000100",
  51618=>"111111111",
  51619=>"000011000",
  51620=>"111100100",
  51621=>"110111111",
  51622=>"001111001",
  51623=>"000000110",
  51624=>"111111111",
  51625=>"111111111",
  51626=>"111111111",
  51627=>"000000001",
  51628=>"000000000",
  51629=>"111111011",
  51630=>"111111111",
  51631=>"000000000",
  51632=>"000100111",
  51633=>"010110111",
  51634=>"000000000",
  51635=>"000000110",
  51636=>"011000001",
  51637=>"111010110",
  51638=>"111111111",
  51639=>"111111101",
  51640=>"100000110",
  51641=>"011000000",
  51642=>"111000000",
  51643=>"111111111",
  51644=>"000011111",
  51645=>"111110000",
  51646=>"111011111",
  51647=>"111001111",
  51648=>"001011111",
  51649=>"000000000",
  51650=>"000000000",
  51651=>"000110010",
  51652=>"001000110",
  51653=>"111111011",
  51654=>"111111111",
  51655=>"110100110",
  51656=>"110111111",
  51657=>"000000000",
  51658=>"111111111",
  51659=>"000000011",
  51660=>"100111000",
  51661=>"111111011",
  51662=>"011011111",
  51663=>"000000000",
  51664=>"000000000",
  51665=>"111111111",
  51666=>"111111100",
  51667=>"000000000",
  51668=>"101000101",
  51669=>"001101110",
  51670=>"011111111",
  51671=>"111011011",
  51672=>"011000000",
  51673=>"111111111",
  51674=>"001111010",
  51675=>"000101111",
  51676=>"001011001",
  51677=>"111111111",
  51678=>"111111111",
  51679=>"111111111",
  51680=>"111011001",
  51681=>"100111111",
  51682=>"000000110",
  51683=>"110000110",
  51684=>"000000000",
  51685=>"000000000",
  51686=>"000000000",
  51687=>"111111111",
  51688=>"111011000",
  51689=>"111000111",
  51690=>"110111111",
  51691=>"100110000",
  51692=>"111011011",
  51693=>"001100110",
  51694=>"000000000",
  51695=>"000010111",
  51696=>"000000000",
  51697=>"000000000",
  51698=>"110110110",
  51699=>"111110000",
  51700=>"000000100",
  51701=>"011100100",
  51702=>"000000100",
  51703=>"110000000",
  51704=>"011111111",
  51705=>"111111111",
  51706=>"000111110",
  51707=>"101001111",
  51708=>"011011111",
  51709=>"111111111",
  51710=>"111010110",
  51711=>"000010110",
  51712=>"111100110",
  51713=>"011000000",
  51714=>"111000001",
  51715=>"111000110",
  51716=>"000000001",
  51717=>"100000000",
  51718=>"000000111",
  51719=>"000000000",
  51720=>"000010000",
  51721=>"010111111",
  51722=>"000000000",
  51723=>"000011111",
  51724=>"000000010",
  51725=>"001111111",
  51726=>"111111000",
  51727=>"111110110",
  51728=>"111111111",
  51729=>"011000000",
  51730=>"000000101",
  51731=>"111111111",
  51732=>"111000000",
  51733=>"111101111",
  51734=>"000000001",
  51735=>"110000110",
  51736=>"000000110",
  51737=>"011010000",
  51738=>"000101111",
  51739=>"011001001",
  51740=>"000000000",
  51741=>"000100000",
  51742=>"001001001",
  51743=>"000110000",
  51744=>"000110111",
  51745=>"111111110",
  51746=>"011111110",
  51747=>"111111111",
  51748=>"001000111",
  51749=>"000101111",
  51750=>"111111101",
  51751=>"000111111",
  51752=>"111111111",
  51753=>"000000000",
  51754=>"111111110",
  51755=>"100100100",
  51756=>"111111000",
  51757=>"111101000",
  51758=>"001111000",
  51759=>"000001000",
  51760=>"001000000",
  51761=>"000011111",
  51762=>"000000000",
  51763=>"001000000",
  51764=>"000000100",
  51765=>"000111110",
  51766=>"000000000",
  51767=>"101000100",
  51768=>"111111110",
  51769=>"111111101",
  51770=>"000000000",
  51771=>"111000000",
  51772=>"000000000",
  51773=>"001000000",
  51774=>"000001101",
  51775=>"111011000",
  51776=>"000000000",
  51777=>"111101100",
  51778=>"000000000",
  51779=>"100000000",
  51780=>"100110110",
  51781=>"110111111",
  51782=>"000110111",
  51783=>"000000000",
  51784=>"000000100",
  51785=>"001001111",
  51786=>"000000000",
  51787=>"111111111",
  51788=>"000000110",
  51789=>"100100100",
  51790=>"110010000",
  51791=>"000111111",
  51792=>"111111111",
  51793=>"111111000",
  51794=>"000100111",
  51795=>"011110000",
  51796=>"111111000",
  51797=>"111111111",
  51798=>"000111111",
  51799=>"111111000",
  51800=>"101000111",
  51801=>"110111111",
  51802=>"101111001",
  51803=>"101000100",
  51804=>"000000000",
  51805=>"000000000",
  51806=>"011110100",
  51807=>"111111110",
  51808=>"000000000",
  51809=>"000000000",
  51810=>"000000000",
  51811=>"111111000",
  51812=>"110111000",
  51813=>"111011000",
  51814=>"111000000",
  51815=>"000001001",
  51816=>"000111000",
  51817=>"111111111",
  51818=>"000011111",
  51819=>"111111011",
  51820=>"001111101",
  51821=>"111111110",
  51822=>"000000000",
  51823=>"110111000",
  51824=>"111011001",
  51825=>"000001000",
  51826=>"010110111",
  51827=>"000000111",
  51828=>"111100111",
  51829=>"000001111",
  51830=>"111111111",
  51831=>"111111111",
  51832=>"111000110",
  51833=>"111011000",
  51834=>"100111111",
  51835=>"000000000",
  51836=>"110111100",
  51837=>"000000111",
  51838=>"101111111",
  51839=>"000000010",
  51840=>"100000111",
  51841=>"000001111",
  51842=>"111011000",
  51843=>"110100110",
  51844=>"111111110",
  51845=>"000000111",
  51846=>"000000111",
  51847=>"000000111",
  51848=>"000000011",
  51849=>"111111000",
  51850=>"001111010",
  51851=>"000000111",
  51852=>"000000110",
  51853=>"000101111",
  51854=>"100100111",
  51855=>"000110000",
  51856=>"000100100",
  51857=>"000110111",
  51858=>"011000000",
  51859=>"000000110",
  51860=>"111111000",
  51861=>"111111111",
  51862=>"001001111",
  51863=>"000000000",
  51864=>"000000000",
  51865=>"000000111",
  51866=>"000000000",
  51867=>"011011000",
  51868=>"000000000",
  51869=>"111010000",
  51870=>"111111011",
  51871=>"000000100",
  51872=>"000000000",
  51873=>"111111111",
  51874=>"000111111",
  51875=>"000000000",
  51876=>"000001111",
  51877=>"001101111",
  51878=>"101111111",
  51879=>"000111110",
  51880=>"000001111",
  51881=>"000000000",
  51882=>"000000000",
  51883=>"110110000",
  51884=>"111111000",
  51885=>"000000001",
  51886=>"000000001",
  51887=>"111111000",
  51888=>"000000000",
  51889=>"000100000",
  51890=>"111111111",
  51891=>"111111110",
  51892=>"010000000",
  51893=>"000000111",
  51894=>"110000000",
  51895=>"111111010",
  51896=>"000100111",
  51897=>"111101111",
  51898=>"100101111",
  51899=>"111111001",
  51900=>"101100000",
  51901=>"010000011",
  51902=>"111101111",
  51903=>"000000010",
  51904=>"000011111",
  51905=>"111111111",
  51906=>"010000000",
  51907=>"111111011",
  51908=>"000000000",
  51909=>"111111111",
  51910=>"000110101",
  51911=>"000000001",
  51912=>"000100111",
  51913=>"000001001",
  51914=>"000000111",
  51915=>"111111111",
  51916=>"000000000",
  51917=>"110111111",
  51918=>"000111010",
  51919=>"000111111",
  51920=>"001000000",
  51921=>"111110000",
  51922=>"000000100",
  51923=>"110111110",
  51924=>"111111110",
  51925=>"000000111",
  51926=>"111110110",
  51927=>"111111111",
  51928=>"111111111",
  51929=>"011001101",
  51930=>"000000111",
  51931=>"110111000",
  51932=>"000000100",
  51933=>"111101100",
  51934=>"000011000",
  51935=>"101011000",
  51936=>"000000000",
  51937=>"000000000",
  51938=>"001110000",
  51939=>"001000000",
  51940=>"000000000",
  51941=>"111111001",
  51942=>"111001000",
  51943=>"000000011",
  51944=>"000000000",
  51945=>"111111110",
  51946=>"000000111",
  51947=>"111111000",
  51948=>"110111110",
  51949=>"000000100",
  51950=>"000000111",
  51951=>"111001111",
  51952=>"111111111",
  51953=>"101101001",
  51954=>"001011111",
  51955=>"000001000",
  51956=>"111111000",
  51957=>"111111111",
  51958=>"000100100",
  51959=>"000000000",
  51960=>"111111000",
  51961=>"111001000",
  51962=>"111111110",
  51963=>"011011101",
  51964=>"100110000",
  51965=>"100000000",
  51966=>"110111111",
  51967=>"110000000",
  51968=>"000000000",
  51969=>"100000111",
  51970=>"111111010",
  51971=>"111110000",
  51972=>"000111111",
  51973=>"000000001",
  51974=>"000000101",
  51975=>"000110111",
  51976=>"111111111",
  51977=>"000000000",
  51978=>"111111111",
  51979=>"111111000",
  51980=>"001001001",
  51981=>"111110000",
  51982=>"001011011",
  51983=>"111111111",
  51984=>"111101001",
  51985=>"000000000",
  51986=>"111100110",
  51987=>"111000001",
  51988=>"111111111",
  51989=>"000111100",
  51990=>"011111000",
  51991=>"000001111",
  51992=>"101111100",
  51993=>"111111000",
  51994=>"100111000",
  51995=>"110110111",
  51996=>"111111000",
  51997=>"000000010",
  51998=>"111011111",
  51999=>"011000011",
  52000=>"000000000",
  52001=>"000010011",
  52002=>"011000000",
  52003=>"011000000",
  52004=>"011000000",
  52005=>"000000000",
  52006=>"101111100",
  52007=>"000000000",
  52008=>"111111111",
  52009=>"111110000",
  52010=>"011000000",
  52011=>"000000111",
  52012=>"001111111",
  52013=>"100101000",
  52014=>"111000111",
  52015=>"111111000",
  52016=>"000001001",
  52017=>"110110110",
  52018=>"000000000",
  52019=>"111111000",
  52020=>"000000000",
  52021=>"111000010",
  52022=>"110000111",
  52023=>"000000000",
  52024=>"000000000",
  52025=>"101000101",
  52026=>"111110101",
  52027=>"111111111",
  52028=>"000000000",
  52029=>"000000000",
  52030=>"110100000",
  52031=>"000000010",
  52032=>"111000000",
  52033=>"011111000",
  52034=>"011000101",
  52035=>"000000011",
  52036=>"000100110",
  52037=>"100000000",
  52038=>"111101100",
  52039=>"111111111",
  52040=>"111111111",
  52041=>"001000000",
  52042=>"111011000",
  52043=>"100000000",
  52044=>"000000111",
  52045=>"111110000",
  52046=>"111111111",
  52047=>"000000000",
  52048=>"000000000",
  52049=>"001000111",
  52050=>"010010100",
  52051=>"100101001",
  52052=>"000101111",
  52053=>"001000000",
  52054=>"100000000",
  52055=>"010000000",
  52056=>"111111111",
  52057=>"001000111",
  52058=>"110110111",
  52059=>"011111011",
  52060=>"000000001",
  52061=>"000100110",
  52062=>"000000100",
  52063=>"001111100",
  52064=>"000000001",
  52065=>"111000000",
  52066=>"000000110",
  52067=>"111111111",
  52068=>"111111111",
  52069=>"011111010",
  52070=>"000000010",
  52071=>"000000000",
  52072=>"000000001",
  52073=>"000000000",
  52074=>"000001111",
  52075=>"111111111",
  52076=>"000000000",
  52077=>"000001111",
  52078=>"111100000",
  52079=>"010001111",
  52080=>"100100111",
  52081=>"000000000",
  52082=>"000111111",
  52083=>"111111111",
  52084=>"010100000",
  52085=>"000000101",
  52086=>"111111111",
  52087=>"001101000",
  52088=>"000000100",
  52089=>"010111110",
  52090=>"000110110",
  52091=>"100000000",
  52092=>"000000111",
  52093=>"111111111",
  52094=>"100110000",
  52095=>"111111110",
  52096=>"111000000",
  52097=>"111111111",
  52098=>"100111111",
  52099=>"110100000",
  52100=>"010010000",
  52101=>"000001000",
  52102=>"110010000",
  52103=>"111000000",
  52104=>"100100111",
  52105=>"001000111",
  52106=>"000000100",
  52107=>"000001001",
  52108=>"000110111",
  52109=>"111111111",
  52110=>"111101001",
  52111=>"000000000",
  52112=>"111111110",
  52113=>"001000011",
  52114=>"000000110",
  52115=>"110000011",
  52116=>"000000000",
  52117=>"011111000",
  52118=>"100110111",
  52119=>"001000110",
  52120=>"000000001",
  52121=>"111111011",
  52122=>"000000001",
  52123=>"001000000",
  52124=>"000000111",
  52125=>"000001001",
  52126=>"000000011",
  52127=>"000000110",
  52128=>"000000100",
  52129=>"000100001",
  52130=>"101101111",
  52131=>"111000000",
  52132=>"111010001",
  52133=>"111111111",
  52134=>"000000111",
  52135=>"000000000",
  52136=>"000000000",
  52137=>"111100000",
  52138=>"001000000",
  52139=>"111111110",
  52140=>"000000110",
  52141=>"000000111",
  52142=>"000000100",
  52143=>"000111111",
  52144=>"000000000",
  52145=>"000000000",
  52146=>"000011111",
  52147=>"110000000",
  52148=>"111111011",
  52149=>"001101111",
  52150=>"101000001",
  52151=>"000000110",
  52152=>"100100100",
  52153=>"111111111",
  52154=>"000000000",
  52155=>"111111111",
  52156=>"000001111",
  52157=>"000000001",
  52158=>"111111000",
  52159=>"111001001",
  52160=>"000000000",
  52161=>"000000000",
  52162=>"000000111",
  52163=>"111111111",
  52164=>"000111111",
  52165=>"001000110",
  52166=>"000000000",
  52167=>"111111111",
  52168=>"101000111",
  52169=>"110110000",
  52170=>"000000111",
  52171=>"101001111",
  52172=>"000000000",
  52173=>"111110000",
  52174=>"000000111",
  52175=>"111000111",
  52176=>"000000101",
  52177=>"111111100",
  52178=>"111111011",
  52179=>"000000000",
  52180=>"000111111",
  52181=>"111111000",
  52182=>"100000000",
  52183=>"000100000",
  52184=>"111111110",
  52185=>"111111110",
  52186=>"110110111",
  52187=>"111111111",
  52188=>"110110111",
  52189=>"001000000",
  52190=>"111111111",
  52191=>"100000011",
  52192=>"001001111",
  52193=>"110111111",
  52194=>"000000011",
  52195=>"111111001",
  52196=>"000000001",
  52197=>"111111000",
  52198=>"111100000",
  52199=>"000010110",
  52200=>"011000011",
  52201=>"011000000",
  52202=>"110000000",
  52203=>"001001000",
  52204=>"111111110",
  52205=>"000000000",
  52206=>"000000111",
  52207=>"001000000",
  52208=>"000000111",
  52209=>"000000000",
  52210=>"000111100",
  52211=>"001011111",
  52212=>"101111111",
  52213=>"101111111",
  52214=>"000000000",
  52215=>"000000110",
  52216=>"000110110",
  52217=>"100000001",
  52218=>"110111000",
  52219=>"111111111",
  52220=>"001000100",
  52221=>"111111000",
  52222=>"000011000",
  52223=>"000000111",
  52224=>"111111111",
  52225=>"000010000",
  52226=>"000000000",
  52227=>"100111111",
  52228=>"111000110",
  52229=>"111000000",
  52230=>"110111001",
  52231=>"111111111",
  52232=>"000000101",
  52233=>"000000100",
  52234=>"000000110",
  52235=>"000100111",
  52236=>"000110110",
  52237=>"000000000",
  52238=>"101000000",
  52239=>"001001001",
  52240=>"110010110",
  52241=>"111111111",
  52242=>"000000000",
  52243=>"000000000",
  52244=>"000000000",
  52245=>"000000000",
  52246=>"000000000",
  52247=>"111101111",
  52248=>"111111111",
  52249=>"111111011",
  52250=>"010000000",
  52251=>"001011001",
  52252=>"000000000",
  52253=>"010000000",
  52254=>"100000100",
  52255=>"011000101",
  52256=>"101111000",
  52257=>"000000000",
  52258=>"000110000",
  52259=>"110100001",
  52260=>"010000111",
  52261=>"000000100",
  52262=>"001111111",
  52263=>"101111111",
  52264=>"000011111",
  52265=>"000000000",
  52266=>"110111011",
  52267=>"100110110",
  52268=>"000010011",
  52269=>"010011000",
  52270=>"111111111",
  52271=>"000001111",
  52272=>"111111111",
  52273=>"101101111",
  52274=>"000000001",
  52275=>"000110010",
  52276=>"101001001",
  52277=>"110110000",
  52278=>"000000000",
  52279=>"111111111",
  52280=>"000000111",
  52281=>"000010111",
  52282=>"000000000",
  52283=>"111111111",
  52284=>"111111110",
  52285=>"111111000",
  52286=>"100110110",
  52287=>"100000000",
  52288=>"101111000",
  52289=>"111101101",
  52290=>"110000000",
  52291=>"001001000",
  52292=>"110110100",
  52293=>"101111111",
  52294=>"111111000",
  52295=>"111111111",
  52296=>"000000000",
  52297=>"011011001",
  52298=>"011111111",
  52299=>"001011001",
  52300=>"111111111",
  52301=>"111101111",
  52302=>"011000000",
  52303=>"110111111",
  52304=>"000000000",
  52305=>"000000011",
  52306=>"000000000",
  52307=>"110000000",
  52308=>"000000000",
  52309=>"001011111",
  52310=>"000000111",
  52311=>"101101100",
  52312=>"111111101",
  52313=>"000000000",
  52314=>"011111000",
  52315=>"100000100",
  52316=>"000000000",
  52317=>"111111101",
  52318=>"111111101",
  52319=>"011011001",
  52320=>"000000000",
  52321=>"011000000",
  52322=>"000000110",
  52323=>"000000000",
  52324=>"111111001",
  52325=>"000000101",
  52326=>"001000000",
  52327=>"000110000",
  52328=>"111111011",
  52329=>"000000000",
  52330=>"000011000",
  52331=>"000001000",
  52332=>"111111000",
  52333=>"111111111",
  52334=>"000000001",
  52335=>"000111001",
  52336=>"000011000",
  52337=>"000110111",
  52338=>"001001101",
  52339=>"111111111",
  52340=>"000000000",
  52341=>"010000000",
  52342=>"000000000",
  52343=>"111111001",
  52344=>"100100100",
  52345=>"001111111",
  52346=>"111111111",
  52347=>"000000100",
  52348=>"111111010",
  52349=>"101100101",
  52350=>"110010111",
  52351=>"111110000",
  52352=>"000001111",
  52353=>"100100000",
  52354=>"000000001",
  52355=>"011011011",
  52356=>"000000000",
  52357=>"000000011",
  52358=>"001000000",
  52359=>"000100110",
  52360=>"000000000",
  52361=>"111100000",
  52362=>"001101111",
  52363=>"111000011",
  52364=>"000010010",
  52365=>"110111110",
  52366=>"111111001",
  52367=>"000000000",
  52368=>"000000000",
  52369=>"111110100",
  52370=>"110000111",
  52371=>"100100001",
  52372=>"001000000",
  52373=>"111111101",
  52374=>"000000000",
  52375=>"011011011",
  52376=>"010110010",
  52377=>"000000000",
  52378=>"111110010",
  52379=>"111111000",
  52380=>"111111010",
  52381=>"000010110",
  52382=>"111111111",
  52383=>"000001011",
  52384=>"111111001",
  52385=>"110110010",
  52386=>"001000000",
  52387=>"000000000",
  52388=>"110100111",
  52389=>"111110111",
  52390=>"010110010",
  52391=>"111100100",
  52392=>"110110000",
  52393=>"000111111",
  52394=>"000000000",
  52395=>"111111111",
  52396=>"111111010",
  52397=>"001011111",
  52398=>"111111000",
  52399=>"000000011",
  52400=>"000111111",
  52401=>"111111111",
  52402=>"111111000",
  52403=>"000000000",
  52404=>"111101001",
  52405=>"111111111",
  52406=>"000000000",
  52407=>"101111011",
  52408=>"111111111",
  52409=>"000000000",
  52410=>"111101101",
  52411=>"101111101",
  52412=>"111111111",
  52413=>"001001001",
  52414=>"000000000",
  52415=>"000000000",
  52416=>"011000000",
  52417=>"000000111",
  52418=>"111111111",
  52419=>"000000000",
  52420=>"000000000",
  52421=>"111111111",
  52422=>"111111111",
  52423=>"111111111",
  52424=>"000111111",
  52425=>"100100100",
  52426=>"000000001",
  52427=>"101011000",
  52428=>"011000000",
  52429=>"001000011",
  52430=>"010111011",
  52431=>"111111001",
  52432=>"000001011",
  52433=>"000010010",
  52434=>"000010000",
  52435=>"000000000",
  52436=>"000000000",
  52437=>"100111111",
  52438=>"000000000",
  52439=>"111011000",
  52440=>"111111111",
  52441=>"111000000",
  52442=>"000000000",
  52443=>"011001111",
  52444=>"111111111",
  52445=>"111111111",
  52446=>"111001011",
  52447=>"111111011",
  52448=>"000000000",
  52449=>"000000001",
  52450=>"111111111",
  52451=>"110111011",
  52452=>"000000111",
  52453=>"000010010",
  52454=>"111100101",
  52455=>"111111111",
  52456=>"000000000",
  52457=>"001001000",
  52458=>"010010111",
  52459=>"000000000",
  52460=>"000010111",
  52461=>"011000000",
  52462=>"110110111",
  52463=>"111111111",
  52464=>"011111111",
  52465=>"011011111",
  52466=>"001011111",
  52467=>"000011000",
  52468=>"000000000",
  52469=>"110110100",
  52470=>"011011111",
  52471=>"010001000",
  52472=>"110000000",
  52473=>"000000000",
  52474=>"000101001",
  52475=>"000010111",
  52476=>"110111111",
  52477=>"000000000",
  52478=>"000000101",
  52479=>"000111111",
  52480=>"000001011",
  52481=>"111011101",
  52482=>"000000100",
  52483=>"000000000",
  52484=>"011001001",
  52485=>"000011011",
  52486=>"000000110",
  52487=>"000001111",
  52488=>"000110110",
  52489=>"010010000",
  52490=>"000000011",
  52491=>"011011001",
  52492=>"000000000",
  52493=>"000011000",
  52494=>"111111010",
  52495=>"111111110",
  52496=>"000111111",
  52497=>"000100010",
  52498=>"000000000",
  52499=>"001011011",
  52500=>"011010000",
  52501=>"111111111",
  52502=>"100110000",
  52503=>"001000111",
  52504=>"111111001",
  52505=>"111111111",
  52506=>"111111001",
  52507=>"010010000",
  52508=>"111101000",
  52509=>"000000000",
  52510=>"000000010",
  52511=>"000010000",
  52512=>"111011011",
  52513=>"000111111",
  52514=>"000010010",
  52515=>"011001000",
  52516=>"000000000",
  52517=>"111111111",
  52518=>"111011001",
  52519=>"001000001",
  52520=>"111110100",
  52521=>"111111011",
  52522=>"000111111",
  52523=>"000010010",
  52524=>"100000000",
  52525=>"110001000",
  52526=>"111010000",
  52527=>"000000000",
  52528=>"000011011",
  52529=>"000000100",
  52530=>"110111111",
  52531=>"111011001",
  52532=>"110010010",
  52533=>"001000000",
  52534=>"100100000",
  52535=>"011110010",
  52536=>"000000000",
  52537=>"000000111",
  52538=>"111111111",
  52539=>"010000001",
  52540=>"111111011",
  52541=>"111111111",
  52542=>"111111111",
  52543=>"000000000",
  52544=>"000000000",
  52545=>"100101111",
  52546=>"000110000",
  52547=>"000000000",
  52548=>"101100000",
  52549=>"010111011",
  52550=>"000000000",
  52551=>"111111111",
  52552=>"000000000",
  52553=>"000111011",
  52554=>"110111111",
  52555=>"111011000",
  52556=>"110100000",
  52557=>"000000000",
  52558=>"111011000",
  52559=>"000000000",
  52560=>"011111011",
  52561=>"111111101",
  52562=>"000000000",
  52563=>"101001111",
  52564=>"111010110",
  52565=>"011011111",
  52566=>"100000000",
  52567=>"111100000",
  52568=>"000011111",
  52569=>"111111010",
  52570=>"111111111",
  52571=>"000111111",
  52572=>"000001111",
  52573=>"110000000",
  52574=>"001000000",
  52575=>"000000100",
  52576=>"101001111",
  52577=>"000000000",
  52578=>"000000001",
  52579=>"111111111",
  52580=>"000000000",
  52581=>"111010000",
  52582=>"100111111",
  52583=>"000000111",
  52584=>"111111101",
  52585=>"111110000",
  52586=>"110100111",
  52587=>"000001000",
  52588=>"000110110",
  52589=>"000000000",
  52590=>"000000000",
  52591=>"000111111",
  52592=>"000000000",
  52593=>"111010111",
  52594=>"000101111",
  52595=>"111111110",
  52596=>"111111001",
  52597=>"011010000",
  52598=>"000100111",
  52599=>"000000000",
  52600=>"111111111",
  52601=>"000010100",
  52602=>"100100100",
  52603=>"000000000",
  52604=>"110010111",
  52605=>"000000000",
  52606=>"000001000",
  52607=>"000000000",
  52608=>"110110111",
  52609=>"000000111",
  52610=>"110110110",
  52611=>"000000000",
  52612=>"111111111",
  52613=>"000000000",
  52614=>"111011011",
  52615=>"000000011",
  52616=>"000000000",
  52617=>"000000001",
  52618=>"000000110",
  52619=>"000111010",
  52620=>"111111111",
  52621=>"110000100",
  52622=>"000010111",
  52623=>"000000001",
  52624=>"000000000",
  52625=>"111111111",
  52626=>"000000000",
  52627=>"100100100",
  52628=>"111111011",
  52629=>"000000000",
  52630=>"110000000",
  52631=>"101001001",
  52632=>"110000111",
  52633=>"001000110",
  52634=>"000000000",
  52635=>"111111111",
  52636=>"000000111",
  52637=>"110100000",
  52638=>"100000000",
  52639=>"111111111",
  52640=>"111111111",
  52641=>"100000011",
  52642=>"101100101",
  52643=>"000000000",
  52644=>"111111111",
  52645=>"111111111",
  52646=>"100000000",
  52647=>"111111000",
  52648=>"000111110",
  52649=>"100110000",
  52650=>"000000000",
  52651=>"100000000",
  52652=>"000000000",
  52653=>"111011111",
  52654=>"000000011",
  52655=>"111111111",
  52656=>"011111111",
  52657=>"000000111",
  52658=>"000111101",
  52659=>"000000000",
  52660=>"111111111",
  52661=>"101101101",
  52662=>"000100111",
  52663=>"000100111",
  52664=>"000000011",
  52665=>"110110111",
  52666=>"111100000",
  52667=>"011000101",
  52668=>"111111111",
  52669=>"001001101",
  52670=>"001001000",
  52671=>"110000000",
  52672=>"000000100",
  52673=>"111111111",
  52674=>"111111000",
  52675=>"111111110",
  52676=>"111110101",
  52677=>"001101111",
  52678=>"011111111",
  52679=>"111111111",
  52680=>"000000001",
  52681=>"101111111",
  52682=>"000001000",
  52683=>"000000111",
  52684=>"111011000",
  52685=>"111111111",
  52686=>"011000010",
  52687=>"011000000",
  52688=>"011011000",
  52689=>"000000000",
  52690=>"100001001",
  52691=>"111110111",
  52692=>"000010011",
  52693=>"000000000",
  52694=>"000000000",
  52695=>"000001011",
  52696=>"000111111",
  52697=>"011011001",
  52698=>"000000110",
  52699=>"111011111",
  52700=>"000000000",
  52701=>"000111111",
  52702=>"111111010",
  52703=>"110100100",
  52704=>"111111000",
  52705=>"111101110",
  52706=>"000000000",
  52707=>"000000000",
  52708=>"000111000",
  52709=>"000000111",
  52710=>"011111011",
  52711=>"011111111",
  52712=>"001000000",
  52713=>"100000001",
  52714=>"111110110",
  52715=>"111111111",
  52716=>"111111111",
  52717=>"101000000",
  52718=>"100100000",
  52719=>"011010010",
  52720=>"111111111",
  52721=>"000000000",
  52722=>"011001011",
  52723=>"110010000",
  52724=>"000000000",
  52725=>"000000001",
  52726=>"010000000",
  52727=>"000101101",
  52728=>"001000000",
  52729=>"011110110",
  52730=>"001000000",
  52731=>"000000000",
  52732=>"110111011",
  52733=>"000000111",
  52734=>"000000000",
  52735=>"111000000",
  52736=>"001011001",
  52737=>"111001000",
  52738=>"001000000",
  52739=>"000110111",
  52740=>"000001001",
  52741=>"110001111",
  52742=>"111111111",
  52743=>"111111000",
  52744=>"111111001",
  52745=>"000000100",
  52746=>"000100101",
  52747=>"111100111",
  52748=>"101000000",
  52749=>"000000000",
  52750=>"000000000",
  52751=>"101000001",
  52752=>"111111111",
  52753=>"010000000",
  52754=>"000000010",
  52755=>"111111111",
  52756=>"110111000",
  52757=>"101000000",
  52758=>"000000000",
  52759=>"000000001",
  52760=>"100000111",
  52761=>"100110000",
  52762=>"000000111",
  52763=>"000000010",
  52764=>"100101111",
  52765=>"000111111",
  52766=>"111111111",
  52767=>"000000101",
  52768=>"111110110",
  52769=>"110110000",
  52770=>"100000100",
  52771=>"111100100",
  52772=>"111111011",
  52773=>"000000000",
  52774=>"111110000",
  52775=>"000000000",
  52776=>"000111111",
  52777=>"111010000",
  52778=>"000001001",
  52779=>"000000000",
  52780=>"111000011",
  52781=>"000000000",
  52782=>"111001000",
  52783=>"011000000",
  52784=>"100111111",
  52785=>"111111111",
  52786=>"001100100",
  52787=>"111111100",
  52788=>"000111111",
  52789=>"111110000",
  52790=>"111111100",
  52791=>"000001111",
  52792=>"001001000",
  52793=>"100000000",
  52794=>"101000101",
  52795=>"111111000",
  52796=>"000000111",
  52797=>"000000000",
  52798=>"000110111",
  52799=>"001111111",
  52800=>"111101111",
  52801=>"000011100",
  52802=>"000100010",
  52803=>"001011110",
  52804=>"001011101",
  52805=>"011111010",
  52806=>"000011111",
  52807=>"111111111",
  52808=>"100110111",
  52809=>"111111111",
  52810=>"000011111",
  52811=>"011011111",
  52812=>"111111111",
  52813=>"011000000",
  52814=>"000000000",
  52815=>"101001101",
  52816=>"000001000",
  52817=>"011011000",
  52818=>"111111000",
  52819=>"011011011",
  52820=>"000000000",
  52821=>"010111111",
  52822=>"111000111",
  52823=>"000000001",
  52824=>"100111100",
  52825=>"000000001",
  52826=>"000110010",
  52827=>"110101000",
  52828=>"110111000",
  52829=>"001001000",
  52830=>"000000001",
  52831=>"111100000",
  52832=>"111111111",
  52833=>"110000000",
  52834=>"111100111",
  52835=>"001000011",
  52836=>"000001000",
  52837=>"111111000",
  52838=>"000011111",
  52839=>"111111111",
  52840=>"110000000",
  52841=>"001010000",
  52842=>"001000001",
  52843=>"000111111",
  52844=>"000111111",
  52845=>"111111111",
  52846=>"000000111",
  52847=>"011111111",
  52848=>"000111111",
  52849=>"000000111",
  52850=>"100111111",
  52851=>"000000111",
  52852=>"111100100",
  52853=>"000000000",
  52854=>"000000100",
  52855=>"111100111",
  52856=>"000000000",
  52857=>"000000001",
  52858=>"000000000",
  52859=>"000000000",
  52860=>"110110010",
  52861=>"000010110",
  52862=>"000000111",
  52863=>"100110111",
  52864=>"001000000",
  52865=>"100110110",
  52866=>"111000110",
  52867=>"100000100",
  52868=>"001101001",
  52869=>"100000111",
  52870=>"101111000",
  52871=>"000000000",
  52872=>"111111111",
  52873=>"000000001",
  52874=>"101001010",
  52875=>"101000011",
  52876=>"000101000",
  52877=>"000000110",
  52878=>"111111111",
  52879=>"111011000",
  52880=>"000111111",
  52881=>"010000011",
  52882=>"011001001",
  52883=>"001001000",
  52884=>"000011000",
  52885=>"111111000",
  52886=>"000001111",
  52887=>"001000000",
  52888=>"000110100",
  52889=>"111111000",
  52890=>"000110111",
  52891=>"001000000",
  52892=>"000000100",
  52893=>"101000000",
  52894=>"111111111",
  52895=>"000000111",
  52896=>"111000000",
  52897=>"111010000",
  52898=>"000001000",
  52899=>"111111111",
  52900=>"111000000",
  52901=>"011010000",
  52902=>"000000000",
  52903=>"111110100",
  52904=>"000000111",
  52905=>"011000000",
  52906=>"000000111",
  52907=>"100100111",
  52908=>"000001111",
  52909=>"101001000",
  52910=>"111111000",
  52911=>"111111000",
  52912=>"000000000",
  52913=>"001001001",
  52914=>"111111111",
  52915=>"011000000",
  52916=>"111000000",
  52917=>"000111000",
  52918=>"111111111",
  52919=>"111111111",
  52920=>"000111101",
  52921=>"111111111",
  52922=>"100000000",
  52923=>"111000000",
  52924=>"000000000",
  52925=>"111111100",
  52926=>"000111010",
  52927=>"111111100",
  52928=>"111100100",
  52929=>"000001111",
  52930=>"111111111",
  52931=>"010111000",
  52932=>"111111010",
  52933=>"000000011",
  52934=>"000111111",
  52935=>"111101100",
  52936=>"000000000",
  52937=>"101001111",
  52938=>"101111111",
  52939=>"000000000",
  52940=>"000110101",
  52941=>"000100111",
  52942=>"011010000",
  52943=>"110000000",
  52944=>"011000000",
  52945=>"001000101",
  52946=>"011000000",
  52947=>"000010111",
  52948=>"000111111",
  52949=>"111111111",
  52950=>"101000000",
  52951=>"000111111",
  52952=>"000000000",
  52953=>"111111000",
  52954=>"000000000",
  52955=>"110000001",
  52956=>"111011011",
  52957=>"110110010",
  52958=>"011111000",
  52959=>"000000000",
  52960=>"001000100",
  52961=>"000111111",
  52962=>"111000000",
  52963=>"101000101",
  52964=>"000110110",
  52965=>"010000000",
  52966=>"111010000",
  52967=>"111101111",
  52968=>"111100000",
  52969=>"111111111",
  52970=>"100100100",
  52971=>"111000000",
  52972=>"111111111",
  52973=>"000000000",
  52974=>"111000111",
  52975=>"000000000",
  52976=>"000000001",
  52977=>"111000101",
  52978=>"111100000",
  52979=>"110110000",
  52980=>"011001001",
  52981=>"011111000",
  52982=>"111110100",
  52983=>"110111111",
  52984=>"111000000",
  52985=>"111001000",
  52986=>"000000111",
  52987=>"000000000",
  52988=>"001111111",
  52989=>"111011011",
  52990=>"111001111",
  52991=>"011011110",
  52992=>"110100111",
  52993=>"000000100",
  52994=>"000110000",
  52995=>"000001111",
  52996=>"110000000",
  52997=>"000000100",
  52998=>"111110000",
  52999=>"000101111",
  53000=>"110100101",
  53001=>"011000000",
  53002=>"000000000",
  53003=>"000000000",
  53004=>"111111111",
  53005=>"000000111",
  53006=>"100000000",
  53007=>"110000000",
  53008=>"111011000",
  53009=>"111000000",
  53010=>"000000111",
  53011=>"110011111",
  53012=>"111111100",
  53013=>"000000000",
  53014=>"001111101",
  53015=>"000000110",
  53016=>"000010110",
  53017=>"011011001",
  53018=>"010010011",
  53019=>"000000000",
  53020=>"101101000",
  53021=>"000000000",
  53022=>"110111111",
  53023=>"111110000",
  53024=>"000100100",
  53025=>"111111000",
  53026=>"110111111",
  53027=>"000100101",
  53028=>"111111111",
  53029=>"111000100",
  53030=>"111110000",
  53031=>"100011111",
  53032=>"100010111",
  53033=>"100110110",
  53034=>"000101100",
  53035=>"000100111",
  53036=>"000000011",
  53037=>"010000000",
  53038=>"000000110",
  53039=>"100000000",
  53040=>"111111111",
  53041=>"111010111",
  53042=>"000000000",
  53043=>"111111111",
  53044=>"000000000",
  53045=>"110100111",
  53046=>"111111111",
  53047=>"111100000",
  53048=>"000000000",
  53049=>"111000000",
  53050=>"110111111",
  53051=>"111000000",
  53052=>"111100100",
  53053=>"111011011",
  53054=>"111101000",
  53055=>"010000000",
  53056=>"111000000",
  53057=>"001001000",
  53058=>"100000100",
  53059=>"000000001",
  53060=>"000110111",
  53061=>"111111000",
  53062=>"010001000",
  53063=>"100100001",
  53064=>"111111011",
  53065=>"001000000",
  53066=>"000001000",
  53067=>"000111111",
  53068=>"011000000",
  53069=>"101111111",
  53070=>"111001000",
  53071=>"000000111",
  53072=>"011001000",
  53073=>"000000000",
  53074=>"001111110",
  53075=>"111111111",
  53076=>"000000000",
  53077=>"011011011",
  53078=>"000000001",
  53079=>"101000000",
  53080=>"000111111",
  53081=>"000000000",
  53082=>"001111101",
  53083=>"110100110",
  53084=>"000000111",
  53085=>"000110110",
  53086=>"111111010",
  53087=>"000110110",
  53088=>"000000000",
  53089=>"000111000",
  53090=>"100111011",
  53091=>"000100000",
  53092=>"100111111",
  53093=>"000111111",
  53094=>"110110111",
  53095=>"000000000",
  53096=>"000110111",
  53097=>"011111000",
  53098=>"000000111",
  53099=>"111100101",
  53100=>"000011000",
  53101=>"110000000",
  53102=>"111111111",
  53103=>"101001111",
  53104=>"111000111",
  53105=>"111011111",
  53106=>"000110100",
  53107=>"100001101",
  53108=>"111010011",
  53109=>"000100100",
  53110=>"111111111",
  53111=>"110110010",
  53112=>"001001000",
  53113=>"000000001",
  53114=>"001001000",
  53115=>"100000100",
  53116=>"010000111",
  53117=>"010000000",
  53118=>"111011000",
  53119=>"100001000",
  53120=>"000000111",
  53121=>"010110111",
  53122=>"110111000",
  53123=>"000000000",
  53124=>"000000000",
  53125=>"000010111",
  53126=>"111111111",
  53127=>"111011011",
  53128=>"000000111",
  53129=>"010000000",
  53130=>"001010110",
  53131=>"111111000",
  53132=>"111111101",
  53133=>"111100110",
  53134=>"111111111",
  53135=>"111111111",
  53136=>"111111000",
  53137=>"110110100",
  53138=>"001011000",
  53139=>"111001000",
  53140=>"000000001",
  53141=>"011000000",
  53142=>"111101111",
  53143=>"111000000",
  53144=>"001111000",
  53145=>"110111101",
  53146=>"000000000",
  53147=>"111111111",
  53148=>"111110110",
  53149=>"111111100",
  53150=>"000110100",
  53151=>"111011010",
  53152=>"000000000",
  53153=>"110000110",
  53154=>"110000101",
  53155=>"000000111",
  53156=>"101101111",
  53157=>"001001000",
  53158=>"000000001",
  53159=>"000111101",
  53160=>"000000000",
  53161=>"000010011",
  53162=>"111001101",
  53163=>"110000000",
  53164=>"000000011",
  53165=>"111001000",
  53166=>"111111111",
  53167=>"111000111",
  53168=>"000001101",
  53169=>"000111111",
  53170=>"111011111",
  53171=>"011001000",
  53172=>"110111111",
  53173=>"111111000",
  53174=>"000000010",
  53175=>"111111111",
  53176=>"101111000",
  53177=>"001000101",
  53178=>"111111011",
  53179=>"111111011",
  53180=>"011111111",
  53181=>"000001000",
  53182=>"101111000",
  53183=>"100111100",
  53184=>"000000011",
  53185=>"110110000",
  53186=>"111000000",
  53187=>"101101110",
  53188=>"001101111",
  53189=>"011000111",
  53190=>"111111110",
  53191=>"000101000",
  53192=>"110000100",
  53193=>"111100100",
  53194=>"001000000",
  53195=>"000000110",
  53196=>"101000000",
  53197=>"111011110",
  53198=>"100000000",
  53199=>"111000100",
  53200=>"001000111",
  53201=>"111000010",
  53202=>"010011001",
  53203=>"101111111",
  53204=>"000010111",
  53205=>"111000111",
  53206=>"111111000",
  53207=>"001000000",
  53208=>"111101111",
  53209=>"000000000",
  53210=>"000000111",
  53211=>"101000100",
  53212=>"100100111",
  53213=>"111111111",
  53214=>"111111111",
  53215=>"110000001",
  53216=>"000001111",
  53217=>"110111000",
  53218=>"000000000",
  53219=>"111110000",
  53220=>"111111111",
  53221=>"001111111",
  53222=>"110000000",
  53223=>"111000000",
  53224=>"110000011",
  53225=>"111000000",
  53226=>"000000000",
  53227=>"100101100",
  53228=>"000100110",
  53229=>"110100000",
  53230=>"101000111",
  53231=>"100111111",
  53232=>"000000000",
  53233=>"010000110",
  53234=>"111100000",
  53235=>"000100000",
  53236=>"110000100",
  53237=>"000001011",
  53238=>"111000100",
  53239=>"010111000",
  53240=>"000000111",
  53241=>"111100000",
  53242=>"111111111",
  53243=>"000000000",
  53244=>"000000101",
  53245=>"111011000",
  53246=>"111110000",
  53247=>"000000001",
  53248=>"000000000",
  53249=>"000110111",
  53250=>"111111111",
  53251=>"000000000",
  53252=>"111111111",
  53253=>"100100110",
  53254=>"111100100",
  53255=>"111111111",
  53256=>"111110111",
  53257=>"000100111",
  53258=>"111111111",
  53259=>"000111111",
  53260=>"110110111",
  53261=>"000001000",
  53262=>"111111101",
  53263=>"000000000",
  53264=>"111111111",
  53265=>"111111111",
  53266=>"111111111",
  53267=>"111111110",
  53268=>"000000001",
  53269=>"000000110",
  53270=>"011000000",
  53271=>"000000000",
  53272=>"111111111",
  53273=>"100000100",
  53274=>"000000111",
  53275=>"100100100",
  53276=>"111111111",
  53277=>"000000010",
  53278=>"111110100",
  53279=>"011000000",
  53280=>"111111111",
  53281=>"000011011",
  53282=>"000000000",
  53283=>"111110111",
  53284=>"111100000",
  53285=>"111111101",
  53286=>"111101001",
  53287=>"011111111",
  53288=>"111110110",
  53289=>"000000000",
  53290=>"011110000",
  53291=>"111111111",
  53292=>"110111111",
  53293=>"111111111",
  53294=>"011111001",
  53295=>"000011111",
  53296=>"111111111",
  53297=>"001001000",
  53298=>"100001100",
  53299=>"111111111",
  53300=>"000000000",
  53301=>"100110110",
  53302=>"000000000",
  53303=>"000111111",
  53304=>"111111111",
  53305=>"000000000",
  53306=>"000110011",
  53307=>"111111100",
  53308=>"110100000",
  53309=>"111000000",
  53310=>"111110110",
  53311=>"000001011",
  53312=>"000000000",
  53313=>"111111111",
  53314=>"111000000",
  53315=>"011000000",
  53316=>"100100100",
  53317=>"100100110",
  53318=>"000000000",
  53319=>"000111111",
  53320=>"000000100",
  53321=>"111111111",
  53322=>"111111111",
  53323=>"000000000",
  53324=>"111111100",
  53325=>"001000011",
  53326=>"111100111",
  53327=>"111111110",
  53328=>"111111011",
  53329=>"011011011",
  53330=>"111111111",
  53331=>"100100100",
  53332=>"001001000",
  53333=>"111111001",
  53334=>"111011111",
  53335=>"010000000",
  53336=>"111111111",
  53337=>"000100000",
  53338=>"111111011",
  53339=>"110010110",
  53340=>"000000000",
  53341=>"111111110",
  53342=>"000011000",
  53343=>"001111111",
  53344=>"100000000",
  53345=>"000000000",
  53346=>"100100000",
  53347=>"000000000",
  53348=>"110000000",
  53349=>"001011111",
  53350=>"111111111",
  53351=>"111111111",
  53352=>"111111111",
  53353=>"111111111",
  53354=>"001011000",
  53355=>"000000001",
  53356=>"111111011",
  53357=>"000000001",
  53358=>"111111111",
  53359=>"111111100",
  53360=>"110111111",
  53361=>"001011111",
  53362=>"111111111",
  53363=>"111111001",
  53364=>"000001000",
  53365=>"111111111",
  53366=>"000000000",
  53367=>"111111111",
  53368=>"101111111",
  53369=>"000000000",
  53370=>"000000000",
  53371=>"000000000",
  53372=>"111111111",
  53373=>"001001000",
  53374=>"100000001",
  53375=>"011000000",
  53376=>"111111111",
  53377=>"111110110",
  53378=>"111010100",
  53379=>"110111000",
  53380=>"000000000",
  53381=>"001111111",
  53382=>"110110110",
  53383=>"001001000",
  53384=>"111000000",
  53385=>"111101111",
  53386=>"000000000",
  53387=>"010111111",
  53388=>"111111111",
  53389=>"111111111",
  53390=>"111111111",
  53391=>"000000000",
  53392=>"000000000",
  53393=>"000000000",
  53394=>"111011010",
  53395=>"111111111",
  53396=>"110000000",
  53397=>"111111111",
  53398=>"111000000",
  53399=>"011111111",
  53400=>"111000000",
  53401=>"111011011",
  53402=>"111000000",
  53403=>"110010000",
  53404=>"001001111",
  53405=>"000000000",
  53406=>"110001011",
  53407=>"111111111",
  53408=>"111111000",
  53409=>"111110111",
  53410=>"000011000",
  53411=>"110110111",
  53412=>"101101111",
  53413=>"110000001",
  53414=>"000000000",
  53415=>"110100111",
  53416=>"000110110",
  53417=>"110110110",
  53418=>"111111101",
  53419=>"110111110",
  53420=>"100000000",
  53421=>"111111111",
  53422=>"110000001",
  53423=>"111111000",
  53424=>"000000000",
  53425=>"111111111",
  53426=>"110110000",
  53427=>"000110110",
  53428=>"001000100",
  53429=>"111111111",
  53430=>"111111111",
  53431=>"110000000",
  53432=>"000000001",
  53433=>"001111000",
  53434=>"011111011",
  53435=>"110000000",
  53436=>"111111111",
  53437=>"111111111",
  53438=>"000000100",
  53439=>"000000000",
  53440=>"111111100",
  53441=>"110100001",
  53442=>"111111010",
  53443=>"000000000",
  53444=>"000001011",
  53445=>"111011001",
  53446=>"111111111",
  53447=>"000111111",
  53448=>"001000000",
  53449=>"111111111",
  53450=>"000000000",
  53451=>"100000000",
  53452=>"111111111",
  53453=>"000100001",
  53454=>"110000000",
  53455=>"000000000",
  53456=>"000100100",
  53457=>"111111111",
  53458=>"000000001",
  53459=>"111111111",
  53460=>"010000000",
  53461=>"111111110",
  53462=>"011111111",
  53463=>"100000000",
  53464=>"000000000",
  53465=>"011111000",
  53466=>"000000000",
  53467=>"110111011",
  53468=>"000001000",
  53469=>"111000000",
  53470=>"000000000",
  53471=>"010000111",
  53472=>"000000001",
  53473=>"011001011",
  53474=>"111111111",
  53475=>"011011001",
  53476=>"000000000",
  53477=>"000110101",
  53478=>"111011011",
  53479=>"111001000",
  53480=>"000000111",
  53481=>"000000000",
  53482=>"000100111",
  53483=>"111111111",
  53484=>"111111111",
  53485=>"111111111",
  53486=>"110111111",
  53487=>"000000000",
  53488=>"000111000",
  53489=>"111100111",
  53490=>"111100111",
  53491=>"111111011",
  53492=>"000000000",
  53493=>"110111110",
  53494=>"101111111",
  53495=>"111011011",
  53496=>"000111000",
  53497=>"111111010",
  53498=>"000001001",
  53499=>"000000000",
  53500=>"100101101",
  53501=>"101111111",
  53502=>"111000000",
  53503=>"111000000",
  53504=>"000001011",
  53505=>"111110110",
  53506=>"000000101",
  53507=>"000000000",
  53508=>"110010111",
  53509=>"000110111",
  53510=>"000000000",
  53511=>"001001000",
  53512=>"111000000",
  53513=>"111111111",
  53514=>"111110111",
  53515=>"111110011",
  53516=>"000000000",
  53517=>"000111001",
  53518=>"111111111",
  53519=>"010111111",
  53520=>"010110111",
  53521=>"111111111",
  53522=>"000100100",
  53523=>"111110010",
  53524=>"111110000",
  53525=>"000000110",
  53526=>"001011001",
  53527=>"110010000",
  53528=>"100000000",
  53529=>"011000000",
  53530=>"100000000",
  53531=>"011111111",
  53532=>"001000001",
  53533=>"011011000",
  53534=>"111111111",
  53535=>"100100111",
  53536=>"000001000",
  53537=>"000000001",
  53538=>"000001001",
  53539=>"100000001",
  53540=>"000000000",
  53541=>"110111111",
  53542=>"010000000",
  53543=>"001001011",
  53544=>"111111111",
  53545=>"000000010",
  53546=>"000000110",
  53547=>"010111001",
  53548=>"000000000",
  53549=>"100111111",
  53550=>"111111111",
  53551=>"000000000",
  53552=>"111001111",
  53553=>"111011000",
  53554=>"010111111",
  53555=>"000010111",
  53556=>"111111111",
  53557=>"111111011",
  53558=>"000000000",
  53559=>"000100111",
  53560=>"000000110",
  53561=>"000000000",
  53562=>"111000010",
  53563=>"011000100",
  53564=>"111111111",
  53565=>"111110110",
  53566=>"111000011",
  53567=>"000000000",
  53568=>"111011000",
  53569=>"110000000",
  53570=>"100100100",
  53571=>"000000000",
  53572=>"000100110",
  53573=>"000000000",
  53574=>"000000000",
  53575=>"100100100",
  53576=>"111000100",
  53577=>"111101111",
  53578=>"000010111",
  53579=>"100000000",
  53580=>"001001000",
  53581=>"001100000",
  53582=>"011000000",
  53583=>"111110111",
  53584=>"100100000",
  53585=>"011000000",
  53586=>"100010000",
  53587=>"010000000",
  53588=>"110011000",
  53589=>"001111011",
  53590=>"000000011",
  53591=>"111101101",
  53592=>"000000000",
  53593=>"001011000",
  53594=>"000000000",
  53595=>"000000000",
  53596=>"111111000",
  53597=>"111111111",
  53598=>"101111111",
  53599=>"000000000",
  53600=>"000000000",
  53601=>"000000000",
  53602=>"110011011",
  53603=>"111111111",
  53604=>"110111100",
  53605=>"000000010",
  53606=>"000111111",
  53607=>"000000110",
  53608=>"111111110",
  53609=>"000000111",
  53610=>"111111111",
  53611=>"000000000",
  53612=>"100000000",
  53613=>"011000000",
  53614=>"000000000",
  53615=>"000000000",
  53616=>"111111111",
  53617=>"111100110",
  53618=>"111111111",
  53619=>"011000000",
  53620=>"001000000",
  53621=>"111010000",
  53622=>"111111111",
  53623=>"001000001",
  53624=>"100110111",
  53625=>"000000000",
  53626=>"100110010",
  53627=>"111100010",
  53628=>"000100111",
  53629=>"111111111",
  53630=>"110110110",
  53631=>"111111111",
  53632=>"111111111",
  53633=>"010000000",
  53634=>"000000001",
  53635=>"000000000",
  53636=>"111111111",
  53637=>"000000000",
  53638=>"111111111",
  53639=>"100100101",
  53640=>"111111100",
  53641=>"000000000",
  53642=>"111111000",
  53643=>"011111001",
  53644=>"111111111",
  53645=>"000000000",
  53646=>"111011111",
  53647=>"110101111",
  53648=>"111111111",
  53649=>"011011110",
  53650=>"000000000",
  53651=>"111110100",
  53652=>"011011000",
  53653=>"000000000",
  53654=>"110100000",
  53655=>"111111111",
  53656=>"111000000",
  53657=>"001000111",
  53658=>"000000000",
  53659=>"111111111",
  53660=>"001001000",
  53661=>"000000000",
  53662=>"010011000",
  53663=>"000000000",
  53664=>"111001101",
  53665=>"100100111",
  53666=>"001000001",
  53667=>"111111111",
  53668=>"111111111",
  53669=>"111111111",
  53670=>"110111011",
  53671=>"111000011",
  53672=>"111100100",
  53673=>"000000001",
  53674=>"011111001",
  53675=>"000000000",
  53676=>"001000000",
  53677=>"111111111",
  53678=>"111000000",
  53679=>"000000111",
  53680=>"000000110",
  53681=>"011001000",
  53682=>"111111111",
  53683=>"110110010",
  53684=>"110100111",
  53685=>"111111111",
  53686=>"110111111",
  53687=>"100100000",
  53688=>"011010110",
  53689=>"110110110",
  53690=>"101000111",
  53691=>"011011111",
  53692=>"000000000",
  53693=>"111111111",
  53694=>"000010111",
  53695=>"011001011",
  53696=>"000000000",
  53697=>"111111110",
  53698=>"011111011",
  53699=>"111111111",
  53700=>"111111111",
  53701=>"111111111",
  53702=>"011011011",
  53703=>"000000111",
  53704=>"110000000",
  53705=>"010011111",
  53706=>"111111111",
  53707=>"000011001",
  53708=>"000000000",
  53709=>"000111010",
  53710=>"111111100",
  53711=>"111111111",
  53712=>"110000000",
  53713=>"000000000",
  53714=>"111111011",
  53715=>"000000000",
  53716=>"000001001",
  53717=>"000000000",
  53718=>"000000000",
  53719=>"011111111",
  53720=>"110010010",
  53721=>"000000010",
  53722=>"111010111",
  53723=>"111111111",
  53724=>"101100000",
  53725=>"000001001",
  53726=>"111111110",
  53727=>"011111111",
  53728=>"000000000",
  53729=>"111111011",
  53730=>"110010000",
  53731=>"000111111",
  53732=>"111111001",
  53733=>"010000000",
  53734=>"110111111",
  53735=>"111111000",
  53736=>"110110100",
  53737=>"100101000",
  53738=>"000111100",
  53739=>"111111000",
  53740=>"000100101",
  53741=>"011011111",
  53742=>"010011011",
  53743=>"011110000",
  53744=>"000000000",
  53745=>"011011001",
  53746=>"110111111",
  53747=>"000101100",
  53748=>"111111111",
  53749=>"000001000",
  53750=>"000001000",
  53751=>"100110111",
  53752=>"000001111",
  53753=>"110110000",
  53754=>"111110000",
  53755=>"000000000",
  53756=>"000000000",
  53757=>"111001101",
  53758=>"000000000",
  53759=>"011011111",
  53760=>"000000000",
  53761=>"011000000",
  53762=>"000111111",
  53763=>"000000000",
  53764=>"000001111",
  53765=>"111001001",
  53766=>"000000111",
  53767=>"111111111",
  53768=>"000000110",
  53769=>"111111111",
  53770=>"111111111",
  53771=>"111111000",
  53772=>"110110111",
  53773=>"101111111",
  53774=>"000000000",
  53775=>"111111111",
  53776=>"010000100",
  53777=>"101111111",
  53778=>"111111110",
  53779=>"000000000",
  53780=>"100000000",
  53781=>"110010001",
  53782=>"111111111",
  53783=>"111001111",
  53784=>"000000000",
  53785=>"000000001",
  53786=>"000000010",
  53787=>"100110100",
  53788=>"000000000",
  53789=>"111000000",
  53790=>"000000111",
  53791=>"101111111",
  53792=>"001101111",
  53793=>"100101111",
  53794=>"011011111",
  53795=>"000000111",
  53796=>"111111011",
  53797=>"001111110",
  53798=>"100100000",
  53799=>"111001011",
  53800=>"100001111",
  53801=>"100000000",
  53802=>"010111110",
  53803=>"000000011",
  53804=>"111111111",
  53805=>"100001000",
  53806=>"111111100",
  53807=>"000000000",
  53808=>"111111110",
  53809=>"111111001",
  53810=>"011001111",
  53811=>"111111000",
  53812=>"101101111",
  53813=>"111111111",
  53814=>"111101000",
  53815=>"100111011",
  53816=>"000000000",
  53817=>"100100000",
  53818=>"001111111",
  53819=>"111001111",
  53820=>"111111111",
  53821=>"111110110",
  53822=>"000000000",
  53823=>"100000000",
  53824=>"000000100",
  53825=>"110010011",
  53826=>"111001011",
  53827=>"100000111",
  53828=>"000000001",
  53829=>"111111110",
  53830=>"000000111",
  53831=>"111111111",
  53832=>"000001001",
  53833=>"001011111",
  53834=>"100100100",
  53835=>"111111111",
  53836=>"001000110",
  53837=>"111000000",
  53838=>"001111111",
  53839=>"110111111",
  53840=>"110111111",
  53841=>"011000000",
  53842=>"000100001",
  53843=>"010110111",
  53844=>"000001111",
  53845=>"111100000",
  53846=>"000000000",
  53847=>"101111111",
  53848=>"111101101",
  53849=>"101101111",
  53850=>"010111011",
  53851=>"001001001",
  53852=>"110111111",
  53853=>"111000000",
  53854=>"001001001",
  53855=>"011000000",
  53856=>"000000000",
  53857=>"000000000",
  53858=>"000011000",
  53859=>"110111111",
  53860=>"111000000",
  53861=>"101111111",
  53862=>"000000000",
  53863=>"000000000",
  53864=>"011001000",
  53865=>"000100100",
  53866=>"111011000",
  53867=>"011111111",
  53868=>"000000000",
  53869=>"111000000",
  53870=>"000111111",
  53871=>"000000000",
  53872=>"000111011",
  53873=>"000000000",
  53874=>"011011101",
  53875=>"011111111",
  53876=>"000000000",
  53877=>"000000000",
  53878=>"000000000",
  53879=>"000000000",
  53880=>"000000000",
  53881=>"110100110",
  53882=>"111000000",
  53883=>"011000000",
  53884=>"111110000",
  53885=>"000000000",
  53886=>"000000000",
  53887=>"100000000",
  53888=>"010111111",
  53889=>"000000000",
  53890=>"000000000",
  53891=>"111001000",
  53892=>"101001000",
  53893=>"000000000",
  53894=>"000000000",
  53895=>"000111111",
  53896=>"111111111",
  53897=>"000000000",
  53898=>"000000000",
  53899=>"011111111",
  53900=>"111111111",
  53901=>"111101111",
  53902=>"000000000",
  53903=>"000111000",
  53904=>"001001111",
  53905=>"111011011",
  53906=>"000000000",
  53907=>"111111111",
  53908=>"000000000",
  53909=>"011111111",
  53910=>"000000000",
  53911=>"000000000",
  53912=>"100101000",
  53913=>"111111111",
  53914=>"111111001",
  53915=>"110000000",
  53916=>"000101111",
  53917=>"001000000",
  53918=>"111111111",
  53919=>"000000000",
  53920=>"000000000",
  53921=>"000000000",
  53922=>"111111111",
  53923=>"110111111",
  53924=>"000000000",
  53925=>"111111111",
  53926=>"000000011",
  53927=>"110111111",
  53928=>"100110000",
  53929=>"110000111",
  53930=>"000100000",
  53931=>"101000000",
  53932=>"111011001",
  53933=>"110011110",
  53934=>"000000000",
  53935=>"000000111",
  53936=>"000000000",
  53937=>"111111101",
  53938=>"111111111",
  53939=>"110110101",
  53940=>"101100000",
  53941=>"000110100",
  53942=>"001000000",
  53943=>"000111111",
  53944=>"111111000",
  53945=>"000011011",
  53946=>"001001000",
  53947=>"111111111",
  53948=>"111111111",
  53949=>"000000000",
  53950=>"111101111",
  53951=>"111101000",
  53952=>"100111111",
  53953=>"001001001",
  53954=>"110110000",
  53955=>"000000100",
  53956=>"000011010",
  53957=>"000000000",
  53958=>"111111111",
  53959=>"101101101",
  53960=>"111111000",
  53961=>"111000000",
  53962=>"100100100",
  53963=>"011000000",
  53964=>"000000000",
  53965=>"111111111",
  53966=>"000011111",
  53967=>"111111011",
  53968=>"010011000",
  53969=>"110111001",
  53970=>"000100111",
  53971=>"001101111",
  53972=>"100100101",
  53973=>"011001011",
  53974=>"001000000",
  53975=>"001001000",
  53976=>"111111000",
  53977=>"110000001",
  53978=>"000000000",
  53979=>"111101101",
  53980=>"111001000",
  53981=>"111000000",
  53982=>"111001000",
  53983=>"000000000",
  53984=>"000000000",
  53985=>"000000000",
  53986=>"011111000",
  53987=>"110111111",
  53988=>"000000000",
  53989=>"000000000",
  53990=>"111111110",
  53991=>"000000111",
  53992=>"000000000",
  53993=>"001111111",
  53994=>"000000111",
  53995=>"111101000",
  53996=>"000000000",
  53997=>"111111111",
  53998=>"000000000",
  53999=>"000000001",
  54000=>"111111011",
  54001=>"000000001",
  54002=>"000011000",
  54003=>"000000000",
  54004=>"000011111",
  54005=>"111100000",
  54006=>"111111111",
  54007=>"001001000",
  54008=>"111111111",
  54009=>"001000100",
  54010=>"111111111",
  54011=>"000000000",
  54012=>"111111001",
  54013=>"000110010",
  54014=>"111110000",
  54015=>"111001000",
  54016=>"000000000",
  54017=>"011111000",
  54018=>"000000000",
  54019=>"100000111",
  54020=>"000000000",
  54021=>"111111111",
  54022=>"000000000",
  54023=>"000000000",
  54024=>"011000000",
  54025=>"111111111",
  54026=>"000001100",
  54027=>"000000111",
  54028=>"001001101",
  54029=>"100100111",
  54030=>"111111111",
  54031=>"001111111",
  54032=>"011000000",
  54033=>"100111101",
  54034=>"001001111",
  54035=>"000111111",
  54036=>"000000011",
  54037=>"000011111",
  54038=>"011011111",
  54039=>"000000000",
  54040=>"000000000",
  54041=>"000111111",
  54042=>"111111111",
  54043=>"111111000",
  54044=>"000000000",
  54045=>"000100000",
  54046=>"000000000",
  54047=>"111111111",
  54048=>"000000000",
  54049=>"111111111",
  54050=>"011000000",
  54051=>"111111111",
  54052=>"111110000",
  54053=>"101000000",
  54054=>"000111000",
  54055=>"111010000",
  54056=>"000000000",
  54057=>"000000100",
  54058=>"010000000",
  54059=>"011111111",
  54060=>"011011011",
  54061=>"100100000",
  54062=>"110101111",
  54063=>"111111000",
  54064=>"111111011",
  54065=>"101000101",
  54066=>"000000000",
  54067=>"100111011",
  54068=>"010000001",
  54069=>"000111111",
  54070=>"000000000",
  54071=>"110111111",
  54072=>"000000000",
  54073=>"000000000",
  54074=>"111111101",
  54075=>"111001001",
  54076=>"000000000",
  54077=>"111111111",
  54078=>"000100100",
  54079=>"111111111",
  54080=>"000110011",
  54081=>"000001111",
  54082=>"111111011",
  54083=>"000000000",
  54084=>"000000000",
  54085=>"000100000",
  54086=>"001000001",
  54087=>"001001001",
  54088=>"111100100",
  54089=>"000111111",
  54090=>"110111001",
  54091=>"010000000",
  54092=>"000000000",
  54093=>"111111111",
  54094=>"111000001",
  54095=>"111111010",
  54096=>"001111110",
  54097=>"100100111",
  54098=>"000000000",
  54099=>"111101101",
  54100=>"111000000",
  54101=>"011011011",
  54102=>"111001000",
  54103=>"100111111",
  54104=>"110100000",
  54105=>"000000001",
  54106=>"000111111",
  54107=>"000000000",
  54108=>"000000000",
  54109=>"000000000",
  54110=>"111111001",
  54111=>"110111000",
  54112=>"000000000",
  54113=>"000000001",
  54114=>"100101001",
  54115=>"000000000",
  54116=>"111111111",
  54117=>"101111001",
  54118=>"000000000",
  54119=>"011000001",
  54120=>"001011111",
  54121=>"111011111",
  54122=>"000000111",
  54123=>"000100001",
  54124=>"111111111",
  54125=>"100111111",
  54126=>"111111111",
  54127=>"010111111",
  54128=>"000111000",
  54129=>"111111101",
  54130=>"111011111",
  54131=>"111111111",
  54132=>"111111000",
  54133=>"000011001",
  54134=>"000100111",
  54135=>"000000011",
  54136=>"011011111",
  54137=>"000000000",
  54138=>"111001001",
  54139=>"000000000",
  54140=>"100111111",
  54141=>"000000011",
  54142=>"000000100",
  54143=>"111111111",
  54144=>"100000000",
  54145=>"111111111",
  54146=>"111111011",
  54147=>"000000000",
  54148=>"111111110",
  54149=>"111111110",
  54150=>"101000000",
  54151=>"000000000",
  54152=>"000000111",
  54153=>"110111100",
  54154=>"111111000",
  54155=>"001011111",
  54156=>"000000000",
  54157=>"000000000",
  54158=>"111011001",
  54159=>"010111010",
  54160=>"011111111",
  54161=>"000000100",
  54162=>"111111111",
  54163=>"000000000",
  54164=>"000000000",
  54165=>"000011000",
  54166=>"000011111",
  54167=>"000000000",
  54168=>"000100000",
  54169=>"101000000",
  54170=>"000100111",
  54171=>"111001111",
  54172=>"000111011",
  54173=>"000000100",
  54174=>"000001000",
  54175=>"111111111",
  54176=>"000000100",
  54177=>"011111000",
  54178=>"110001000",
  54179=>"111011011",
  54180=>"100000000",
  54181=>"111111110",
  54182=>"111111011",
  54183=>"111111111",
  54184=>"000000111",
  54185=>"001000000",
  54186=>"000000000",
  54187=>"010011000",
  54188=>"011001000",
  54189=>"110000000",
  54190=>"100100000",
  54191=>"111100000",
  54192=>"000000101",
  54193=>"111111111",
  54194=>"111111111",
  54195=>"111111111",
  54196=>"111011001",
  54197=>"111100001",
  54198=>"000000001",
  54199=>"111100000",
  54200=>"111000000",
  54201=>"111111111",
  54202=>"111111111",
  54203=>"111111111",
  54204=>"000000101",
  54205=>"110010111",
  54206=>"011011000",
  54207=>"011000000",
  54208=>"000000001",
  54209=>"111111111",
  54210=>"110010000",
  54211=>"111111111",
  54212=>"111100000",
  54213=>"111111011",
  54214=>"000000000",
  54215=>"111111111",
  54216=>"000111001",
  54217=>"000100000",
  54218=>"111111111",
  54219=>"110100110",
  54220=>"100001000",
  54221=>"001001000",
  54222=>"001000000",
  54223=>"110100000",
  54224=>"111111011",
  54225=>"111111111",
  54226=>"111111111",
  54227=>"001000111",
  54228=>"000000000",
  54229=>"111111000",
  54230=>"111000000",
  54231=>"011000100",
  54232=>"000000000",
  54233=>"111001101",
  54234=>"011000000",
  54235=>"100100100",
  54236=>"000000000",
  54237=>"010000101",
  54238=>"000000000",
  54239=>"111111010",
  54240=>"111011011",
  54241=>"101111000",
  54242=>"001001111",
  54243=>"000000001",
  54244=>"000001000",
  54245=>"111110111",
  54246=>"111111000",
  54247=>"111110000",
  54248=>"000000000",
  54249=>"111111111",
  54250=>"000000000",
  54251=>"100110110",
  54252=>"110000000",
  54253=>"000000000",
  54254=>"111111111",
  54255=>"110110000",
  54256=>"000001000",
  54257=>"111111111",
  54258=>"000000001",
  54259=>"000000000",
  54260=>"011000000",
  54261=>"111111100",
  54262=>"000111111",
  54263=>"010000000",
  54264=>"000111111",
  54265=>"010000000",
  54266=>"000000000",
  54267=>"000000000",
  54268=>"111111001",
  54269=>"010111000",
  54270=>"100000000",
  54271=>"000000110",
  54272=>"111111001",
  54273=>"101001111",
  54274=>"111111000",
  54275=>"111110111",
  54276=>"000000000",
  54277=>"000010000",
  54278=>"101101111",
  54279=>"111111101",
  54280=>"111100111",
  54281=>"011111000",
  54282=>"000000010",
  54283=>"001000000",
  54284=>"111101111",
  54285=>"101110111",
  54286=>"000000111",
  54287=>"101101111",
  54288=>"000000000",
  54289=>"111111110",
  54290=>"111111000",
  54291=>"110101000",
  54292=>"011011011",
  54293=>"000100100",
  54294=>"111111111",
  54295=>"011011011",
  54296=>"111111111",
  54297=>"111010000",
  54298=>"000000101",
  54299=>"000010010",
  54300=>"111000000",
  54301=>"010011000",
  54302=>"111011111",
  54303=>"110110100",
  54304=>"100101111",
  54305=>"111111111",
  54306=>"000011011",
  54307=>"111111111",
  54308=>"101001000",
  54309=>"111111100",
  54310=>"000000000",
  54311=>"000100100",
  54312=>"000000000",
  54313=>"000000000",
  54314=>"000000000",
  54315=>"000010010",
  54316=>"110111111",
  54317=>"000000000",
  54318=>"111011010",
  54319=>"100101101",
  54320=>"110111111",
  54321=>"111111111",
  54322=>"000001011",
  54323=>"001011011",
  54324=>"111110110",
  54325=>"111111111",
  54326=>"010110111",
  54327=>"111111111",
  54328=>"000011111",
  54329=>"000000000",
  54330=>"000000000",
  54331=>"000000000",
  54332=>"111111111",
  54333=>"111100100",
  54334=>"111111110",
  54335=>"011010000",
  54336=>"000010110",
  54337=>"111101100",
  54338=>"011111111",
  54339=>"000000100",
  54340=>"010011110",
  54341=>"001111111",
  54342=>"011111010",
  54343=>"111111111",
  54344=>"111111011",
  54345=>"000000101",
  54346=>"001000001",
  54347=>"111111111",
  54348=>"000000000",
  54349=>"110000000",
  54350=>"111110100",
  54351=>"101111011",
  54352=>"000000100",
  54353=>"000000111",
  54354=>"000000111",
  54355=>"000010000",
  54356=>"000000000",
  54357=>"111111111",
  54358=>"101001000",
  54359=>"111111111",
  54360=>"000100110",
  54361=>"111111100",
  54362=>"111111111",
  54363=>"001001111",
  54364=>"111100111",
  54365=>"000011110",
  54366=>"111111000",
  54367=>"000110110",
  54368=>"100100111",
  54369=>"111111011",
  54370=>"100110111",
  54371=>"111111111",
  54372=>"000000000",
  54373=>"111111111",
  54374=>"111111111",
  54375=>"111111011",
  54376=>"000000111",
  54377=>"000000001",
  54378=>"011110111",
  54379=>"000110110",
  54380=>"110110110",
  54381=>"000111111",
  54382=>"000000000",
  54383=>"111111011",
  54384=>"111111111",
  54385=>"110111111",
  54386=>"000000000",
  54387=>"000001111",
  54388=>"000111111",
  54389=>"111101001",
  54390=>"111001111",
  54391=>"111111000",
  54392=>"000000000",
  54393=>"111000000",
  54394=>"000000111",
  54395=>"111101000",
  54396=>"001001001",
  54397=>"000011001",
  54398=>"110111111",
  54399=>"100111111",
  54400=>"111111000",
  54401=>"111011110",
  54402=>"111011111",
  54403=>"111111100",
  54404=>"001000111",
  54405=>"000000000",
  54406=>"111111111",
  54407=>"001100111",
  54408=>"111111111",
  54409=>"000011111",
  54410=>"100101111",
  54411=>"011111111",
  54412=>"000000000",
  54413=>"001001011",
  54414=>"001001110",
  54415=>"101101111",
  54416=>"111101111",
  54417=>"001001010",
  54418=>"010011010",
  54419=>"111011111",
  54420=>"111111110",
  54421=>"010110000",
  54422=>"000000000",
  54423=>"000111000",
  54424=>"110000011",
  54425=>"111111111",
  54426=>"000110111",
  54427=>"111111111",
  54428=>"111111010",
  54429=>"000000000",
  54430=>"110100100",
  54431=>"111111000",
  54432=>"111110000",
  54433=>"111100100",
  54434=>"000000000",
  54435=>"111111111",
  54436=>"111100100",
  54437=>"101000110",
  54438=>"000100000",
  54439=>"011111111",
  54440=>"011011011",
  54441=>"111111111",
  54442=>"111111010",
  54443=>"101111111",
  54444=>"101111111",
  54445=>"111100100",
  54446=>"000001000",
  54447=>"001000100",
  54448=>"000000101",
  54449=>"110100000",
  54450=>"101101111",
  54451=>"111111110",
  54452=>"100001011",
  54453=>"101001000",
  54454=>"100000000",
  54455=>"111100110",
  54456=>"000000000",
  54457=>"000000000",
  54458=>"010110110",
  54459=>"101001000",
  54460=>"010111011",
  54461=>"000000100",
  54462=>"011011010",
  54463=>"011011001",
  54464=>"010111111",
  54465=>"000000010",
  54466=>"000110111",
  54467=>"110111010",
  54468=>"111111111",
  54469=>"000000000",
  54470=>"110000000",
  54471=>"000110000",
  54472=>"000000010",
  54473=>"100111111",
  54474=>"111111101",
  54475=>"000000000",
  54476=>"000101100",
  54477=>"110100000",
  54478=>"111001000",
  54479=>"111111111",
  54480=>"111111000",
  54481=>"011010011",
  54482=>"011000100",
  54483=>"111111011",
  54484=>"111111111",
  54485=>"111111111",
  54486=>"000000000",
  54487=>"000110111",
  54488=>"111111110",
  54489=>"110111010",
  54490=>"000000110",
  54491=>"110111101",
  54492=>"110111111",
  54493=>"001001001",
  54494=>"110111111",
  54495=>"000000000",
  54496=>"000000000",
  54497=>"000000000",
  54498=>"111111100",
  54499=>"111111111",
  54500=>"011111000",
  54501=>"000011100",
  54502=>"000000100",
  54503=>"110100000",
  54504=>"000000100",
  54505=>"110110100",
  54506=>"000000000",
  54507=>"100000001",
  54508=>"000000100",
  54509=>"000100000",
  54510=>"011010000",
  54511=>"000000111",
  54512=>"000000000",
  54513=>"111101101",
  54514=>"110100110",
  54515=>"000000101",
  54516=>"001001001",
  54517=>"001001011",
  54518=>"110111111",
  54519=>"000000000",
  54520=>"000000000",
  54521=>"001000000",
  54522=>"000000111",
  54523=>"111100000",
  54524=>"000001111",
  54525=>"110110000",
  54526=>"111111111",
  54527=>"000000000",
  54528=>"100000101",
  54529=>"100100000",
  54530=>"111111111",
  54531=>"111010000",
  54532=>"111111111",
  54533=>"010110110",
  54534=>"000000000",
  54535=>"111111111",
  54536=>"110110011",
  54537=>"000100110",
  54538=>"000111000",
  54539=>"001000110",
  54540=>"000000110",
  54541=>"000000000",
  54542=>"111111111",
  54543=>"001001100",
  54544=>"001000100",
  54545=>"000000000",
  54546=>"111001000",
  54547=>"100001111",
  54548=>"111100000",
  54549=>"111111110",
  54550=>"111011000",
  54551=>"000110100",
  54552=>"011011111",
  54553=>"111111001",
  54554=>"011011010",
  54555=>"111110000",
  54556=>"000000111",
  54557=>"110111111",
  54558=>"111111111",
  54559=>"111000000",
  54560=>"000001001",
  54561=>"110111010",
  54562=>"000000110",
  54563=>"000000000",
  54564=>"110110110",
  54565=>"110100000",
  54566=>"111001000",
  54567=>"111111111",
  54568=>"000000010",
  54569=>"001111111",
  54570=>"001011110",
  54571=>"010011000",
  54572=>"110000000",
  54573=>"100000000",
  54574=>"000100000",
  54575=>"000000000",
  54576=>"000111111",
  54577=>"010010000",
  54578=>"000000000",
  54579=>"111000000",
  54580=>"101000100",
  54581=>"001011011",
  54582=>"000000010",
  54583=>"111111111",
  54584=>"000000000",
  54585=>"111111111",
  54586=>"001000011",
  54587=>"100101111",
  54588=>"101111101",
  54589=>"101111110",
  54590=>"001001111",
  54591=>"100111111",
  54592=>"111111111",
  54593=>"111111111",
  54594=>"111111111",
  54595=>"000000000",
  54596=>"000110110",
  54597=>"000110111",
  54598=>"111111000",
  54599=>"001101111",
  54600=>"000111111",
  54601=>"000000000",
  54602=>"100110110",
  54603=>"001001011",
  54604=>"111010000",
  54605=>"111001000",
  54606=>"111111111",
  54607=>"000000000",
  54608=>"011111101",
  54609=>"100100100",
  54610=>"111111111",
  54611=>"000000000",
  54612=>"010111111",
  54613=>"111111101",
  54614=>"111111111",
  54615=>"000100000",
  54616=>"011011010",
  54617=>"000000000",
  54618=>"100100100",
  54619=>"100101101",
  54620=>"100110100",
  54621=>"000000000",
  54622=>"111110000",
  54623=>"100101001",
  54624=>"011011101",
  54625=>"000000000",
  54626=>"111101111",
  54627=>"111111111",
  54628=>"001001001",
  54629=>"000001001",
  54630=>"000000010",
  54631=>"111111111",
  54632=>"111111111",
  54633=>"000000000",
  54634=>"000000000",
  54635=>"110110111",
  54636=>"000000100",
  54637=>"110111111",
  54638=>"000010010",
  54639=>"000000101",
  54640=>"111111111",
  54641=>"111111111",
  54642=>"111111111",
  54643=>"101100100",
  54644=>"011111111",
  54645=>"101111111",
  54646=>"000000000",
  54647=>"111101100",
  54648=>"111111111",
  54649=>"100000000",
  54650=>"000001001",
  54651=>"111111111",
  54652=>"111110111",
  54653=>"110001000",
  54654=>"000000000",
  54655=>"111111111",
  54656=>"111011001",
  54657=>"000011100",
  54658=>"110010000",
  54659=>"000000000",
  54660=>"010110111",
  54661=>"000000000",
  54662=>"110000000",
  54663=>"001000000",
  54664=>"000000011",
  54665=>"100100110",
  54666=>"001111111",
  54667=>"111000000",
  54668=>"111111111",
  54669=>"111101100",
  54670=>"100111111",
  54671=>"000010000",
  54672=>"111111110",
  54673=>"001011011",
  54674=>"111111110",
  54675=>"101001011",
  54676=>"111111111",
  54677=>"101101101",
  54678=>"111111111",
  54679=>"000011001",
  54680=>"111101111",
  54681=>"100000111",
  54682=>"111111111",
  54683=>"011000011",
  54684=>"111111001",
  54685=>"011000000",
  54686=>"111000000",
  54687=>"111110110",
  54688=>"000000000",
  54689=>"111111110",
  54690=>"000000101",
  54691=>"000000111",
  54692=>"000000111",
  54693=>"111110110",
  54694=>"101111111",
  54695=>"010111100",
  54696=>"001000110",
  54697=>"110000000",
  54698=>"000000111",
  54699=>"111111111",
  54700=>"010010000",
  54701=>"111111011",
  54702=>"000110111",
  54703=>"000111000",
  54704=>"111000000",
  54705=>"111111111",
  54706=>"101000000",
  54707=>"010111110",
  54708=>"110110110",
  54709=>"000011111",
  54710=>"111111110",
  54711=>"011010000",
  54712=>"111001111",
  54713=>"000010111",
  54714=>"111000000",
  54715=>"000001001",
  54716=>"111011011",
  54717=>"011111110",
  54718=>"000000000",
  54719=>"111011111",
  54720=>"000000000",
  54721=>"111111111",
  54722=>"000000000",
  54723=>"111111111",
  54724=>"111011000",
  54725=>"111111111",
  54726=>"111111111",
  54727=>"010010111",
  54728=>"110000100",
  54729=>"001111111",
  54730=>"000100100",
  54731=>"000000000",
  54732=>"000100111",
  54733=>"000000000",
  54734=>"101000100",
  54735=>"000111111",
  54736=>"111111111",
  54737=>"100110110",
  54738=>"000100111",
  54739=>"001000000",
  54740=>"000000001",
  54741=>"110010011",
  54742=>"000000000",
  54743=>"111100110",
  54744=>"100100100",
  54745=>"110111111",
  54746=>"000000000",
  54747=>"001000000",
  54748=>"000100111",
  54749=>"000110111",
  54750=>"010111110",
  54751=>"001001101",
  54752=>"111111111",
  54753=>"011111111",
  54754=>"000111111",
  54755=>"000000000",
  54756=>"011001111",
  54757=>"000000000",
  54758=>"000110110",
  54759=>"010010010",
  54760=>"111110100",
  54761=>"111111110",
  54762=>"100000001",
  54763=>"111111011",
  54764=>"111111110",
  54765=>"011001000",
  54766=>"101000001",
  54767=>"110000000",
  54768=>"000000000",
  54769=>"110000110",
  54770=>"111100100",
  54771=>"100111111",
  54772=>"111110111",
  54773=>"011111000",
  54774=>"000000100",
  54775=>"000110111",
  54776=>"111111010",
  54777=>"110100000",
  54778=>"000000000",
  54779=>"000000101",
  54780=>"111000000",
  54781=>"000010000",
  54782=>"000000000",
  54783=>"001001001",
  54784=>"111111100",
  54785=>"000000110",
  54786=>"111111000",
  54787=>"000000000",
  54788=>"111110111",
  54789=>"000000001",
  54790=>"111001101",
  54791=>"101101101",
  54792=>"111111111",
  54793=>"100110000",
  54794=>"110110111",
  54795=>"100110111",
  54796=>"100111110",
  54797=>"111111111",
  54798=>"000000000",
  54799=>"000000000",
  54800=>"111111111",
  54801=>"000000000",
  54802=>"010110110",
  54803=>"111111111",
  54804=>"110000111",
  54805=>"000000001",
  54806=>"000000000",
  54807=>"011001111",
  54808=>"110111110",
  54809=>"000000111",
  54810=>"000000111",
  54811=>"000000000",
  54812=>"111111011",
  54813=>"000000000",
  54814=>"100110110",
  54815=>"111011111",
  54816=>"011111111",
  54817=>"111000000",
  54818=>"111110110",
  54819=>"010110111",
  54820=>"000011011",
  54821=>"100000001",
  54822=>"111100000",
  54823=>"000000000",
  54824=>"001101011",
  54825=>"000000110",
  54826=>"000000000",
  54827=>"000000110",
  54828=>"101111111",
  54829=>"000000000",
  54830=>"110110000",
  54831=>"000100110",
  54832=>"001000000",
  54833=>"111111101",
  54834=>"011001111",
  54835=>"111111110",
  54836=>"111111111",
  54837=>"101111011",
  54838=>"000000001",
  54839=>"000000000",
  54840=>"001000110",
  54841=>"000000100",
  54842=>"000000000",
  54843=>"000000000",
  54844=>"111111011",
  54845=>"111000000",
  54846=>"000100110",
  54847=>"001000000",
  54848=>"100100111",
  54849=>"000000010",
  54850=>"000000111",
  54851=>"111110111",
  54852=>"100100000",
  54853=>"000000000",
  54854=>"111100100",
  54855=>"000000000",
  54856=>"001001101",
  54857=>"000000000",
  54858=>"000000000",
  54859=>"100000000",
  54860=>"001111111",
  54861=>"111111000",
  54862=>"000000000",
  54863=>"000000110",
  54864=>"011000000",
  54865=>"011111111",
  54866=>"000000110",
  54867=>"111000000",
  54868=>"111111111",
  54869=>"000001011",
  54870=>"111101100",
  54871=>"000000000",
  54872=>"000000111",
  54873=>"101001000",
  54874=>"010000000",
  54875=>"110110010",
  54876=>"000000000",
  54877=>"000000001",
  54878=>"111000001",
  54879=>"001101111",
  54880=>"000000000",
  54881=>"000000001",
  54882=>"111011111",
  54883=>"000000000",
  54884=>"110110111",
  54885=>"000010000",
  54886=>"011111011",
  54887=>"000000000",
  54888=>"000001001",
  54889=>"111111111",
  54890=>"000000000",
  54891=>"111011011",
  54892=>"100110110",
  54893=>"110110111",
  54894=>"100100110",
  54895=>"000110100",
  54896=>"000000000",
  54897=>"000000101",
  54898=>"011011001",
  54899=>"011001001",
  54900=>"111101101",
  54901=>"000000000",
  54902=>"000011111",
  54903=>"111111011",
  54904=>"000000011",
  54905=>"000000000",
  54906=>"111110110",
  54907=>"000100000",
  54908=>"110111110",
  54909=>"000000011",
  54910=>"111111111",
  54911=>"011110111",
  54912=>"111111110",
  54913=>"000110110",
  54914=>"111111101",
  54915=>"111101101",
  54916=>"100000000",
  54917=>"000100111",
  54918=>"000000000",
  54919=>"000000000",
  54920=>"001000000",
  54921=>"000111111",
  54922=>"000000000",
  54923=>"111011000",
  54924=>"111111111",
  54925=>"110000000",
  54926=>"111000000",
  54927=>"011011011",
  54928=>"000000000",
  54929=>"000000001",
  54930=>"000111111",
  54931=>"100100000",
  54932=>"111111001",
  54933=>"111100000",
  54934=>"111111111",
  54935=>"000000000",
  54936=>"011000101",
  54937=>"101001111",
  54938=>"001000000",
  54939=>"000011011",
  54940=>"111000000",
  54941=>"101100110",
  54942=>"111111111",
  54943=>"010011010",
  54944=>"111111000",
  54945=>"101110110",
  54946=>"011011111",
  54947=>"011010010",
  54948=>"111111111",
  54949=>"000001111",
  54950=>"110010111",
  54951=>"011011010",
  54952=>"000000110",
  54953=>"111111111",
  54954=>"111111111",
  54955=>"000000000",
  54956=>"001001111",
  54957=>"111111111",
  54958=>"111111111",
  54959=>"011111111",
  54960=>"000011001",
  54961=>"111111111",
  54962=>"011010000",
  54963=>"111111111",
  54964=>"110111111",
  54965=>"101111111",
  54966=>"111001001",
  54967=>"011111110",
  54968=>"001011111",
  54969=>"000000000",
  54970=>"001001000",
  54971=>"110010000",
  54972=>"000100100",
  54973=>"001000000",
  54974=>"111111111",
  54975=>"110110111",
  54976=>"111110000",
  54977=>"111111111",
  54978=>"000111110",
  54979=>"111111111",
  54980=>"011011000",
  54981=>"000000000",
  54982=>"111111000",
  54983=>"000000000",
  54984=>"000001000",
  54985=>"111100100",
  54986=>"001101001",
  54987=>"011111111",
  54988=>"000000000",
  54989=>"111000000",
  54990=>"011000001",
  54991=>"111111110",
  54992=>"000000111",
  54993=>"000110000",
  54994=>"111110111",
  54995=>"000000000",
  54996=>"000001000",
  54997=>"000110111",
  54998=>"000010111",
  54999=>"111111000",
  55000=>"000110110",
  55001=>"111000000",
  55002=>"100110000",
  55003=>"000011011",
  55004=>"110001011",
  55005=>"001000100",
  55006=>"011111111",
  55007=>"111100000",
  55008=>"000000000",
  55009=>"000000000",
  55010=>"011000000",
  55011=>"011000000",
  55012=>"110010110",
  55013=>"001000011",
  55014=>"111000001",
  55015=>"111111011",
  55016=>"000000110",
  55017=>"000000000",
  55018=>"000000000",
  55019=>"111111111",
  55020=>"111111111",
  55021=>"111010000",
  55022=>"000000010",
  55023=>"111011000",
  55024=>"101001001",
  55025=>"100000111",
  55026=>"000000000",
  55027=>"000000000",
  55028=>"111111110",
  55029=>"000000000",
  55030=>"000000000",
  55031=>"000000000",
  55032=>"000000111",
  55033=>"111101001",
  55034=>"111001000",
  55035=>"011111010",
  55036=>"110101011",
  55037=>"011001011",
  55038=>"011000000",
  55039=>"000000001",
  55040=>"000000000",
  55041=>"001001001",
  55042=>"111101111",
  55043=>"111110110",
  55044=>"100100111",
  55045=>"110000000",
  55046=>"111101111",
  55047=>"000000011",
  55048=>"000000000",
  55049=>"000000000",
  55050=>"011000000",
  55051=>"000000000",
  55052=>"000000000",
  55053=>"010011001",
  55054=>"111100100",
  55055=>"000000000",
  55056=>"000000110",
  55057=>"000000001",
  55058=>"000000001",
  55059=>"000101100",
  55060=>"111111000",
  55061=>"111111111",
  55062=>"011010000",
  55063=>"111111011",
  55064=>"101001001",
  55065=>"000100101",
  55066=>"000000111",
  55067=>"111111011",
  55068=>"000000000",
  55069=>"000000000",
  55070=>"000110110",
  55071=>"111000111",
  55072=>"100101111",
  55073=>"001000000",
  55074=>"110100100",
  55075=>"000000000",
  55076=>"000000111",
  55077=>"111011011",
  55078=>"110111111",
  55079=>"111100101",
  55080=>"011000000",
  55081=>"000000011",
  55082=>"000000111",
  55083=>"111110111",
  55084=>"111110000",
  55085=>"100001101",
  55086=>"111111011",
  55087=>"000000000",
  55088=>"000000000",
  55089=>"011000000",
  55090=>"001111111",
  55091=>"011111100",
  55092=>"111111110",
  55093=>"000000000",
  55094=>"000000000",
  55095=>"000000000",
  55096=>"110000000",
  55097=>"111110111",
  55098=>"011001001",
  55099=>"001001001",
  55100=>"000000000",
  55101=>"011000000",
  55102=>"011111000",
  55103=>"000000000",
  55104=>"001111000",
  55105=>"000000001",
  55106=>"111000010",
  55107=>"111111111",
  55108=>"011011111",
  55109=>"011010111",
  55110=>"111101100",
  55111=>"111111111",
  55112=>"111111111",
  55113=>"100000000",
  55114=>"001000000",
  55115=>"110110111",
  55116=>"011111110",
  55117=>"000111000",
  55118=>"101000000",
  55119=>"100110110",
  55120=>"111011001",
  55121=>"000001001",
  55122=>"000000000",
  55123=>"111101111",
  55124=>"000000001",
  55125=>"001000001",
  55126=>"111111100",
  55127=>"111101001",
  55128=>"100001000",
  55129=>"000011011",
  55130=>"000011011",
  55131=>"111111111",
  55132=>"000100000",
  55133=>"101101111",
  55134=>"000000000",
  55135=>"000000110",
  55136=>"101000111",
  55137=>"001001001",
  55138=>"001011011",
  55139=>"111111111",
  55140=>"111010000",
  55141=>"001000000",
  55142=>"000000000",
  55143=>"111111110",
  55144=>"001011011",
  55145=>"000000000",
  55146=>"000100000",
  55147=>"000000001",
  55148=>"111111000",
  55149=>"000000000",
  55150=>"000110110",
  55151=>"111011011",
  55152=>"010000000",
  55153=>"111111011",
  55154=>"111111111",
  55155=>"100110110",
  55156=>"101100100",
  55157=>"100000010",
  55158=>"111111000",
  55159=>"010010000",
  55160=>"111111111",
  55161=>"000000011",
  55162=>"010111011",
  55163=>"001000000",
  55164=>"111111111",
  55165=>"110110010",
  55166=>"000000000",
  55167=>"000000000",
  55168=>"111111000",
  55169=>"111111111",
  55170=>"111100000",
  55171=>"000000111",
  55172=>"111111111",
  55173=>"010010000",
  55174=>"000100000",
  55175=>"110110110",
  55176=>"000000000",
  55177=>"000110000",
  55178=>"110100111",
  55179=>"000110110",
  55180=>"111011111",
  55181=>"000000000",
  55182=>"011000011",
  55183=>"000111111",
  55184=>"110111010",
  55185=>"000000000",
  55186=>"000000000",
  55187=>"010000001",
  55188=>"111111111",
  55189=>"000111011",
  55190=>"111101100",
  55191=>"101011001",
  55192=>"000000110",
  55193=>"011001001",
  55194=>"111111111",
  55195=>"000010010",
  55196=>"111011011",
  55197=>"000000000",
  55198=>"000001000",
  55199=>"100000000",
  55200=>"111111111",
  55201=>"011001001",
  55202=>"111011011",
  55203=>"101111000",
  55204=>"000000000",
  55205=>"100000000",
  55206=>"000000000",
  55207=>"000111111",
  55208=>"000000001",
  55209=>"110110100",
  55210=>"000111111",
  55211=>"000010000",
  55212=>"000000000",
  55213=>"011101100",
  55214=>"011001011",
  55215=>"111111111",
  55216=>"000000000",
  55217=>"111110110",
  55218=>"001000000",
  55219=>"001000000",
  55220=>"111000000",
  55221=>"111101111",
  55222=>"000000000",
  55223=>"111011111",
  55224=>"111100111",
  55225=>"110110111",
  55226=>"001000001",
  55227=>"110110111",
  55228=>"111110111",
  55229=>"000000000",
  55230=>"111111111",
  55231=>"010010000",
  55232=>"111010000",
  55233=>"111111111",
  55234=>"111111111",
  55235=>"111111111",
  55236=>"000000000",
  55237=>"001000100",
  55238=>"000000000",
  55239=>"011111011",
  55240=>"101000111",
  55241=>"000001111",
  55242=>"100000000",
  55243=>"010011111",
  55244=>"000000000",
  55245=>"111111111",
  55246=>"011001001",
  55247=>"111010010",
  55248=>"000000000",
  55249=>"000000000",
  55250=>"111111111",
  55251=>"111111111",
  55252=>"000000001",
  55253=>"011111111",
  55254=>"000000000",
  55255=>"110011011",
  55256=>"111111111",
  55257=>"111111111",
  55258=>"000000000",
  55259=>"111011000",
  55260=>"000000000",
  55261=>"111111111",
  55262=>"011010011",
  55263=>"000010000",
  55264=>"111001000",
  55265=>"111111111",
  55266=>"000000000",
  55267=>"111011000",
  55268=>"101101111",
  55269=>"111111101",
  55270=>"000000001",
  55271=>"111100100",
  55272=>"000000000",
  55273=>"011001111",
  55274=>"111111110",
  55275=>"111111111",
  55276=>"111111111",
  55277=>"100100100",
  55278=>"000010000",
  55279=>"100000000",
  55280=>"111111001",
  55281=>"000000000",
  55282=>"111111111",
  55283=>"011000000",
  55284=>"110010010",
  55285=>"111111111",
  55286=>"010000011",
  55287=>"110000110",
  55288=>"000001111",
  55289=>"001000001",
  55290=>"111111111",
  55291=>"001111111",
  55292=>"111111111",
  55293=>"111111111",
  55294=>"111011011",
  55295=>"010111111",
  55296=>"110111111",
  55297=>"111110110",
  55298=>"111111111",
  55299=>"111011000",
  55300=>"000000011",
  55301=>"001000000",
  55302=>"001001001",
  55303=>"000000000",
  55304=>"101001001",
  55305=>"010010111",
  55306=>"000000000",
  55307=>"011000000",
  55308=>"111111111",
  55309=>"000110011",
  55310=>"111100000",
  55311=>"000000111",
  55312=>"001000000",
  55313=>"111111111",
  55314=>"111101000",
  55315=>"111111111",
  55316=>"111111111",
  55317=>"000000110",
  55318=>"110111111",
  55319=>"110000011",
  55320=>"000111000",
  55321=>"001001001",
  55322=>"111111111",
  55323=>"001001000",
  55324=>"000000000",
  55325=>"000000000",
  55326=>"100100010",
  55327=>"110110000",
  55328=>"110110111",
  55329=>"111111111",
  55330=>"100110110",
  55331=>"111111111",
  55332=>"111111100",
  55333=>"000111001",
  55334=>"000000000",
  55335=>"000000000",
  55336=>"111110000",
  55337=>"000000000",
  55338=>"100100000",
  55339=>"111110000",
  55340=>"100000010",
  55341=>"111111111",
  55342=>"101001001",
  55343=>"001110000",
  55344=>"110110010",
  55345=>"101100000",
  55346=>"011111001",
  55347=>"011111111",
  55348=>"000100100",
  55349=>"000000100",
  55350=>"000000000",
  55351=>"011011001",
  55352=>"011001000",
  55353=>"010110000",
  55354=>"000000000",
  55355=>"011111110",
  55356=>"100100100",
  55357=>"111111001",
  55358=>"111111100",
  55359=>"000000000",
  55360=>"000110110",
  55361=>"100111111",
  55362=>"000000000",
  55363=>"010111000",
  55364=>"111111111",
  55365=>"000000000",
  55366=>"001100111",
  55367=>"111111111",
  55368=>"010000000",
  55369=>"001000000",
  55370=>"111111111",
  55371=>"111111111",
  55372=>"000000000",
  55373=>"110111000",
  55374=>"101111111",
  55375=>"111111111",
  55376=>"000000000",
  55377=>"101111111",
  55378=>"111110100",
  55379=>"111011111",
  55380=>"111111111",
  55381=>"000010010",
  55382=>"110111001",
  55383=>"111111111",
  55384=>"011011111",
  55385=>"001000111",
  55386=>"111111111",
  55387=>"111000000",
  55388=>"000000001",
  55389=>"111111000",
  55390=>"111111111",
  55391=>"100111111",
  55392=>"000100000",
  55393=>"100110111",
  55394=>"111111111",
  55395=>"000000000",
  55396=>"110111000",
  55397=>"000000000",
  55398=>"000000000",
  55399=>"000000001",
  55400=>"111110000",
  55401=>"111111111",
  55402=>"000000000",
  55403=>"110100100",
  55404=>"010001001",
  55405=>"110000111",
  55406=>"111000000",
  55407=>"111110111",
  55408=>"110111110",
  55409=>"001001000",
  55410=>"101100111",
  55411=>"000000000",
  55412=>"100110000",
  55413=>"010001011",
  55414=>"110110110",
  55415=>"000000000",
  55416=>"110111110",
  55417=>"010000000",
  55418=>"000000000",
  55419=>"111000000",
  55420=>"000000000",
  55421=>"000000000",
  55422=>"000000000",
  55423=>"111111111",
  55424=>"000000000",
  55425=>"000010111",
  55426=>"000000010",
  55427=>"011011001",
  55428=>"111111111",
  55429=>"111111010",
  55430=>"000000111",
  55431=>"110100111",
  55432=>"111111100",
  55433=>"000110111",
  55434=>"111000001",
  55435=>"000000000",
  55436=>"101001001",
  55437=>"111111011",
  55438=>"000110111",
  55439=>"000000000",
  55440=>"111111100",
  55441=>"111111111",
  55442=>"000000000",
  55443=>"010010001",
  55444=>"100100000",
  55445=>"100000000",
  55446=>"000111000",
  55447=>"111111111",
  55448=>"111111111",
  55449=>"000000000",
  55450=>"101111111",
  55451=>"100100000",
  55452=>"111111111",
  55453=>"110010110",
  55454=>"111110110",
  55455=>"111010010",
  55456=>"110000111",
  55457=>"000000000",
  55458=>"010010000",
  55459=>"011110111",
  55460=>"100000011",
  55461=>"111010010",
  55462=>"111111111",
  55463=>"010000000",
  55464=>"000100000",
  55465=>"111111111",
  55466=>"000000000",
  55467=>"011011010",
  55468=>"000110010",
  55469=>"110110110",
  55470=>"010001000",
  55471=>"111111000",
  55472=>"111111111",
  55473=>"110010001",
  55474=>"110000110",
  55475=>"001000000",
  55476=>"110111110",
  55477=>"110110000",
  55478=>"000000000",
  55479=>"111111111",
  55480=>"010011000",
  55481=>"000000000",
  55482=>"011001001",
  55483=>"110100000",
  55484=>"101101101",
  55485=>"110111110",
  55486=>"111000000",
  55487=>"111110110",
  55488=>"000000000",
  55489=>"100000000",
  55490=>"000100000",
  55491=>"000000000",
  55492=>"000000000",
  55493=>"111010111",
  55494=>"010111111",
  55495=>"010010001",
  55496=>"111000000",
  55497=>"000000000",
  55498=>"101101111",
  55499=>"001101101",
  55500=>"000110010",
  55501=>"000100110",
  55502=>"100100000",
  55503=>"111111111",
  55504=>"000000000",
  55505=>"000000100",
  55506=>"111001111",
  55507=>"000000000",
  55508=>"110111111",
  55509=>"011000000",
  55510=>"111111111",
  55511=>"000000000",
  55512=>"010111011",
  55513=>"000000010",
  55514=>"111111111",
  55515=>"000010000",
  55516=>"111111000",
  55517=>"000000000",
  55518=>"000000000",
  55519=>"110110010",
  55520=>"001000110",
  55521=>"111001111",
  55522=>"111101100",
  55523=>"100111111",
  55524=>"111101101",
  55525=>"101111111",
  55526=>"111110100",
  55527=>"100100111",
  55528=>"000000000",
  55529=>"111111111",
  55530=>"100000000",
  55531=>"100000010",
  55532=>"000000000",
  55533=>"000000110",
  55534=>"001001000",
  55535=>"011111111",
  55536=>"000011011",
  55537=>"000110110",
  55538=>"111111111",
  55539=>"101101011",
  55540=>"001111011",
  55541=>"111111011",
  55542=>"000000110",
  55543=>"000001011",
  55544=>"111110010",
  55545=>"101001101",
  55546=>"000000000",
  55547=>"100100100",
  55548=>"011001001",
  55549=>"010011011",
  55550=>"000000110",
  55551=>"001100100",
  55552=>"010110000",
  55553=>"010010010",
  55554=>"111111111",
  55555=>"110110110",
  55556=>"101000000",
  55557=>"010110110",
  55558=>"111111110",
  55559=>"111100000",
  55560=>"000000000",
  55561=>"111000000",
  55562=>"100000000",
  55563=>"101101111",
  55564=>"111111111",
  55565=>"011011011",
  55566=>"111111111",
  55567=>"100000110",
  55568=>"111110111",
  55569=>"000000000",
  55570=>"111111111",
  55571=>"111101010",
  55572=>"111111111",
  55573=>"000000000",
  55574=>"000000000",
  55575=>"111011000",
  55576=>"011010110",
  55577=>"111001000",
  55578=>"010010010",
  55579=>"110111111",
  55580=>"100000000",
  55581=>"010110111",
  55582=>"011111111",
  55583=>"111101101",
  55584=>"101101000",
  55585=>"100000000",
  55586=>"111011001",
  55587=>"111111100",
  55588=>"010000000",
  55589=>"000100100",
  55590=>"100100000",
  55591=>"111000100",
  55592=>"111111000",
  55593=>"001101000",
  55594=>"101111111",
  55595=>"111111110",
  55596=>"111001000",
  55597=>"001011111",
  55598=>"000000101",
  55599=>"000000000",
  55600=>"000000000",
  55601=>"000000001",
  55602=>"111110000",
  55603=>"000000000",
  55604=>"111111000",
  55605=>"111101101",
  55606=>"100100000",
  55607=>"001000000",
  55608=>"000000100",
  55609=>"000000001",
  55610=>"000000001",
  55611=>"101111111",
  55612=>"100100000",
  55613=>"110000000",
  55614=>"000000000",
  55615=>"110110111",
  55616=>"111000000",
  55617=>"110111111",
  55618=>"100000000",
  55619=>"011111111",
  55620=>"010111111",
  55621=>"000000110",
  55622=>"000001001",
  55623=>"111111111",
  55624=>"000000000",
  55625=>"000100111",
  55626=>"111111111",
  55627=>"010010000",
  55628=>"110110000",
  55629=>"000001000",
  55630=>"000000110",
  55631=>"010000000",
  55632=>"000001000",
  55633=>"111111111",
  55634=>"000000010",
  55635=>"000000000",
  55636=>"011111100",
  55637=>"111111011",
  55638=>"111111111",
  55639=>"000100100",
  55640=>"111111111",
  55641=>"111111111",
  55642=>"110000111",
  55643=>"100111110",
  55644=>"111111111",
  55645=>"000001011",
  55646=>"111111111",
  55647=>"110000100",
  55648=>"100100101",
  55649=>"011001101",
  55650=>"001001001",
  55651=>"110111111",
  55652=>"111111111",
  55653=>"000011111",
  55654=>"000000000",
  55655=>"010110000",
  55656=>"100011011",
  55657=>"111111000",
  55658=>"111111110",
  55659=>"010111111",
  55660=>"111100100",
  55661=>"111111111",
  55662=>"011111111",
  55663=>"000000000",
  55664=>"000000000",
  55665=>"101001001",
  55666=>"111110000",
  55667=>"011011011",
  55668=>"111111111",
  55669=>"111001000",
  55670=>"000000000",
  55671=>"000000000",
  55672=>"111111111",
  55673=>"111111110",
  55674=>"111010010",
  55675=>"110111011",
  55676=>"111111011",
  55677=>"010010010",
  55678=>"110010111",
  55679=>"111111111",
  55680=>"100100110",
  55681=>"100110010",
  55682=>"000000111",
  55683=>"001000001",
  55684=>"111011000",
  55685=>"110111111",
  55686=>"100110110",
  55687=>"000001000",
  55688=>"000110110",
  55689=>"001000000",
  55690=>"111110111",
  55691=>"011111000",
  55692=>"111111111",
  55693=>"000000011",
  55694=>"111111111",
  55695=>"111111100",
  55696=>"001001100",
  55697=>"000111111",
  55698=>"111011010",
  55699=>"001001000",
  55700=>"000000000",
  55701=>"000110111",
  55702=>"100000000",
  55703=>"001001001",
  55704=>"111111101",
  55705=>"111110111",
  55706=>"000111000",
  55707=>"111111111",
  55708=>"010000000",
  55709=>"110111110",
  55710=>"111111111",
  55711=>"111111111",
  55712=>"100100000",
  55713=>"110110110",
  55714=>"000000000",
  55715=>"111011111",
  55716=>"000110110",
  55717=>"000000000",
  55718=>"101111111",
  55719=>"000011011",
  55720=>"111111000",
  55721=>"000110110",
  55722=>"001001111",
  55723=>"111111011",
  55724=>"001111111",
  55725=>"000000010",
  55726=>"000000000",
  55727=>"101101001",
  55728=>"000000000",
  55729=>"010000000",
  55730=>"000000000",
  55731=>"100110110",
  55732=>"000000111",
  55733=>"101001000",
  55734=>"111010111",
  55735=>"000010000",
  55736=>"111110010",
  55737=>"111101111",
  55738=>"111111111",
  55739=>"000000000",
  55740=>"110110111",
  55741=>"000000000",
  55742=>"001001111",
  55743=>"110110110",
  55744=>"100000000",
  55745=>"111111000",
  55746=>"111111111",
  55747=>"000000000",
  55748=>"101111100",
  55749=>"001111111",
  55750=>"100110100",
  55751=>"101111111",
  55752=>"100100000",
  55753=>"000000001",
  55754=>"101111111",
  55755=>"000000000",
  55756=>"111111111",
  55757=>"111110000",
  55758=>"110110110",
  55759=>"010000000",
  55760=>"000000000",
  55761=>"000000000",
  55762=>"010000111",
  55763=>"111001001",
  55764=>"000110111",
  55765=>"100111111",
  55766=>"111011011",
  55767=>"011011011",
  55768=>"111000000",
  55769=>"111000010",
  55770=>"111101111",
  55771=>"100100111",
  55772=>"000001001",
  55773=>"111111111",
  55774=>"111110111",
  55775=>"010000110",
  55776=>"000000110",
  55777=>"000010001",
  55778=>"100000000",
  55779=>"000000000",
  55780=>"111111111",
  55781=>"101011000",
  55782=>"111011000",
  55783=>"001001111",
  55784=>"000010011",
  55785=>"100010000",
  55786=>"111011111",
  55787=>"000000000",
  55788=>"111111000",
  55789=>"000000000",
  55790=>"111100100",
  55791=>"111111111",
  55792=>"000001001",
  55793=>"001001001",
  55794=>"111100000",
  55795=>"111111111",
  55796=>"111000000",
  55797=>"110010000",
  55798=>"000000111",
  55799=>"110010000",
  55800=>"111111111",
  55801=>"110110110",
  55802=>"001001001",
  55803=>"010000000",
  55804=>"100000000",
  55805=>"000000000",
  55806=>"111111100",
  55807=>"111111111",
  55808=>"000000000",
  55809=>"111100100",
  55810=>"111111111",
  55811=>"011010000",
  55812=>"100000000",
  55813=>"100110110",
  55814=>"010011111",
  55815=>"111111111",
  55816=>"000001001",
  55817=>"000000000",
  55818=>"110111111",
  55819=>"110110110",
  55820=>"100100000",
  55821=>"111111111",
  55822=>"000001011",
  55823=>"000000100",
  55824=>"000000000",
  55825=>"000000000",
  55826=>"110100111",
  55827=>"000010111",
  55828=>"000000000",
  55829=>"000000000",
  55830=>"111100111",
  55831=>"010110110",
  55832=>"110100100",
  55833=>"110100000",
  55834=>"100100100",
  55835=>"100100101",
  55836=>"000000000",
  55837=>"111110000",
  55838=>"000000000",
  55839=>"000000000",
  55840=>"000000000",
  55841=>"111111111",
  55842=>"000111111",
  55843=>"000000000",
  55844=>"101111111",
  55845=>"011000000",
  55846=>"111111110",
  55847=>"111111111",
  55848=>"101111111",
  55849=>"100100000",
  55850=>"111111111",
  55851=>"000100000",
  55852=>"110110000",
  55853=>"000000000",
  55854=>"000110100",
  55855=>"011010011",
  55856=>"000111111",
  55857=>"111000000",
  55858=>"000000000",
  55859=>"010011001",
  55860=>"010110100",
  55861=>"111001100",
  55862=>"110100111",
  55863=>"100110001",
  55864=>"000000000",
  55865=>"111111101",
  55866=>"000000000",
  55867=>"000000000",
  55868=>"101111111",
  55869=>"100100000",
  55870=>"111111111",
  55871=>"110000000",
  55872=>"000000000",
  55873=>"011001001",
  55874=>"111110111",
  55875=>"111011011",
  55876=>"100100110",
  55877=>"110100000",
  55878=>"001001001",
  55879=>"000000000",
  55880=>"000000000",
  55881=>"111111111",
  55882=>"000000000",
  55883=>"111011111",
  55884=>"111111111",
  55885=>"001111000",
  55886=>"111111110",
  55887=>"111111111",
  55888=>"000001111",
  55889=>"011111110",
  55890=>"000000000",
  55891=>"111111111",
  55892=>"000100111",
  55893=>"000000000",
  55894=>"110111011",
  55895=>"000010100",
  55896=>"000000100",
  55897=>"000001000",
  55898=>"011111111",
  55899=>"100111111",
  55900=>"000001001",
  55901=>"000000000",
  55902=>"000000000",
  55903=>"000000000",
  55904=>"111000100",
  55905=>"111111111",
  55906=>"100011111",
  55907=>"111111010",
  55908=>"111111100",
  55909=>"000000000",
  55910=>"111010000",
  55911=>"101100101",
  55912=>"011111111",
  55913=>"001011011",
  55914=>"110111111",
  55915=>"000000000",
  55916=>"111111111",
  55917=>"000000101",
  55918=>"110111111",
  55919=>"111111111",
  55920=>"000000000",
  55921=>"100111001",
  55922=>"111111101",
  55923=>"000000001",
  55924=>"000000100",
  55925=>"111011011",
  55926=>"000000000",
  55927=>"111111110",
  55928=>"111111111",
  55929=>"111101010",
  55930=>"101000000",
  55931=>"000000001",
  55932=>"100100110",
  55933=>"111011111",
  55934=>"000001111",
  55935=>"000010010",
  55936=>"000000000",
  55937=>"100100000",
  55938=>"000000000",
  55939=>"010000000",
  55940=>"111100000",
  55941=>"111111111",
  55942=>"000110100",
  55943=>"111111111",
  55944=>"111000000",
  55945=>"000000000",
  55946=>"011011011",
  55947=>"111111011",
  55948=>"111111111",
  55949=>"110111111",
  55950=>"101001111",
  55951=>"000000000",
  55952=>"111111111",
  55953=>"111111111",
  55954=>"111111111",
  55955=>"100000000",
  55956=>"000000000",
  55957=>"111011010",
  55958=>"111111111",
  55959=>"111111111",
  55960=>"010000111",
  55961=>"000001011",
  55962=>"000000000",
  55963=>"000000000",
  55964=>"000000111",
  55965=>"101101001",
  55966=>"111111111",
  55967=>"111111111",
  55968=>"100011000",
  55969=>"000011011",
  55970=>"000000000",
  55971=>"001001000",
  55972=>"101001000",
  55973=>"100111000",
  55974=>"000000011",
  55975=>"111111111",
  55976=>"111111110",
  55977=>"111100000",
  55978=>"001011001",
  55979=>"000000000",
  55980=>"100001000",
  55981=>"101100100",
  55982=>"111111111",
  55983=>"000000000",
  55984=>"111111100",
  55985=>"011011011",
  55986=>"110110110",
  55987=>"111000100",
  55988=>"011000000",
  55989=>"111111111",
  55990=>"111111110",
  55991=>"000000011",
  55992=>"000001011",
  55993=>"001110111",
  55994=>"111111000",
  55995=>"000000000",
  55996=>"111111111",
  55997=>"000001001",
  55998=>"111111111",
  55999=>"111000110",
  56000=>"100100100",
  56001=>"101000001",
  56002=>"000001001",
  56003=>"000000000",
  56004=>"111111111",
  56005=>"000000000",
  56006=>"000000101",
  56007=>"110011111",
  56008=>"111111111",
  56009=>"000000010",
  56010=>"101100000",
  56011=>"111101111",
  56012=>"110010110",
  56013=>"100100100",
  56014=>"011000000",
  56015=>"110110111",
  56016=>"010000000",
  56017=>"111100100",
  56018=>"111110100",
  56019=>"000000001",
  56020=>"000000111",
  56021=>"111111111",
  56022=>"001001111",
  56023=>"111111111",
  56024=>"000000000",
  56025=>"100100111",
  56026=>"111111101",
  56027=>"000011111",
  56028=>"110111111",
  56029=>"110000000",
  56030=>"110111111",
  56031=>"001111111",
  56032=>"001111111",
  56033=>"011011110",
  56034=>"001000000",
  56035=>"000000000",
  56036=>"001111111",
  56037=>"111111100",
  56038=>"010111111",
  56039=>"111111111",
  56040=>"011000001",
  56041=>"111111011",
  56042=>"000001111",
  56043=>"111111111",
  56044=>"010000000",
  56045=>"000000000",
  56046=>"111111111",
  56047=>"101101111",
  56048=>"111111111",
  56049=>"011000111",
  56050=>"011111000",
  56051=>"000000111",
  56052=>"011111111",
  56053=>"000000001",
  56054=>"111001011",
  56055=>"000000000",
  56056=>"110000000",
  56057=>"110110111",
  56058=>"110111110",
  56059=>"111111110",
  56060=>"111110110",
  56061=>"000000110",
  56062=>"111110000",
  56063=>"101101001",
  56064=>"111111011",
  56065=>"000001001",
  56066=>"000000000",
  56067=>"101000000",
  56068=>"000111111",
  56069=>"000001111",
  56070=>"000000110",
  56071=>"110111110",
  56072=>"000010010",
  56073=>"010000000",
  56074=>"100110110",
  56075=>"000000000",
  56076=>"110100100",
  56077=>"100110110",
  56078=>"000000001",
  56079=>"111111111",
  56080=>"111111111",
  56081=>"111011011",
  56082=>"000000000",
  56083=>"001011111",
  56084=>"101101000",
  56085=>"100000000",
  56086=>"100000000",
  56087=>"011111110",
  56088=>"111011010",
  56089=>"011000110",
  56090=>"000000100",
  56091=>"110110111",
  56092=>"110110111",
  56093=>"111111111",
  56094=>"111111111",
  56095=>"111111111",
  56096=>"111111001",
  56097=>"001111111",
  56098=>"000001111",
  56099=>"000111111",
  56100=>"000010001",
  56101=>"000000000",
  56102=>"000000000",
  56103=>"100111111",
  56104=>"110110000",
  56105=>"110111111",
  56106=>"110110110",
  56107=>"000000100",
  56108=>"000000000",
  56109=>"111111111",
  56110=>"110000000",
  56111=>"010110110",
  56112=>"101101000",
  56113=>"000110111",
  56114=>"110110010",
  56115=>"000100100",
  56116=>"000000000",
  56117=>"101001101",
  56118=>"000000001",
  56119=>"111111111",
  56120=>"000000000",
  56121=>"101101001",
  56122=>"111111100",
  56123=>"011010111",
  56124=>"011011000",
  56125=>"110110000",
  56126=>"110110100",
  56127=>"111011011",
  56128=>"111000000",
  56129=>"011110000",
  56130=>"001001000",
  56131=>"000000000",
  56132=>"100010110",
  56133=>"010011001",
  56134=>"111011000",
  56135=>"110111111",
  56136=>"110110111",
  56137=>"001111111",
  56138=>"101001000",
  56139=>"110110110",
  56140=>"100000000",
  56141=>"001011000",
  56142=>"000000000",
  56143=>"110100000",
  56144=>"100100100",
  56145=>"110001111",
  56146=>"111111110",
  56147=>"000000000",
  56148=>"000000000",
  56149=>"001001001",
  56150=>"000000111",
  56151=>"111000000",
  56152=>"111101111",
  56153=>"111010111",
  56154=>"000101111",
  56155=>"000000000",
  56156=>"000100000",
  56157=>"110000000",
  56158=>"000000111",
  56159=>"010000000",
  56160=>"001111111",
  56161=>"111100000",
  56162=>"000000001",
  56163=>"000000000",
  56164=>"111101011",
  56165=>"111111111",
  56166=>"111111111",
  56167=>"111111111",
  56168=>"111011011",
  56169=>"111111111",
  56170=>"100000000",
  56171=>"000000000",
  56172=>"100100110",
  56173=>"001111000",
  56174=>"111111001",
  56175=>"111111000",
  56176=>"010011111",
  56177=>"001000000",
  56178=>"111111111",
  56179=>"111110010",
  56180=>"000000010",
  56181=>"100000001",
  56182=>"111111111",
  56183=>"111010000",
  56184=>"000000101",
  56185=>"011000001",
  56186=>"111111111",
  56187=>"111000000",
  56188=>"000000000",
  56189=>"000110111",
  56190=>"111000000",
  56191=>"111111111",
  56192=>"101001101",
  56193=>"111111111",
  56194=>"000000000",
  56195=>"000000000",
  56196=>"111111111",
  56197=>"011111111",
  56198=>"000100000",
  56199=>"101111011",
  56200=>"111000000",
  56201=>"000000000",
  56202=>"000100100",
  56203=>"011111011",
  56204=>"000111000",
  56205=>"000000000",
  56206=>"111101111",
  56207=>"011110000",
  56208=>"001011111",
  56209=>"010001111",
  56210=>"110110111",
  56211=>"110111110",
  56212=>"000000000",
  56213=>"000000000",
  56214=>"100100111",
  56215=>"001001110",
  56216=>"000000000",
  56217=>"001100110",
  56218=>"000000111",
  56219=>"111011111",
  56220=>"110000000",
  56221=>"100000000",
  56222=>"111110111",
  56223=>"111111110",
  56224=>"111111111",
  56225=>"111111111",
  56226=>"100100001",
  56227=>"000011010",
  56228=>"111111001",
  56229=>"111111111",
  56230=>"111111111",
  56231=>"111111111",
  56232=>"000000000",
  56233=>"000000000",
  56234=>"000000000",
  56235=>"001001111",
  56236=>"000000000",
  56237=>"000001001",
  56238=>"010011001",
  56239=>"011011000",
  56240=>"011001000",
  56241=>"111111111",
  56242=>"011111111",
  56243=>"000000000",
  56244=>"000000000",
  56245=>"010011011",
  56246=>"111001001",
  56247=>"000001000",
  56248=>"000001000",
  56249=>"000001000",
  56250=>"011111111",
  56251=>"111111000",
  56252=>"000000000",
  56253=>"100100011",
  56254=>"100010110",
  56255=>"110010110",
  56256=>"000000000",
  56257=>"111111111",
  56258=>"000111110",
  56259=>"001000111",
  56260=>"000000000",
  56261=>"100110100",
  56262=>"000001000",
  56263=>"010000000",
  56264=>"000000010",
  56265=>"010111100",
  56266=>"110110010",
  56267=>"111100000",
  56268=>"111111110",
  56269=>"000000000",
  56270=>"111111111",
  56271=>"000000011",
  56272=>"101000000",
  56273=>"010010000",
  56274=>"010111111",
  56275=>"111111000",
  56276=>"111111111",
  56277=>"111111101",
  56278=>"000000000",
  56279=>"111100110",
  56280=>"110010000",
  56281=>"000000100",
  56282=>"111110000",
  56283=>"110010011",
  56284=>"111110110",
  56285=>"100000000",
  56286=>"111111111",
  56287=>"101000101",
  56288=>"110000000",
  56289=>"100111111",
  56290=>"000000000",
  56291=>"111111001",
  56292=>"000110111",
  56293=>"011001000",
  56294=>"100110111",
  56295=>"001000000",
  56296=>"110111111",
  56297=>"000000000",
  56298=>"001000111",
  56299=>"110010000",
  56300=>"000111111",
  56301=>"010010011",
  56302=>"011111111",
  56303=>"110110111",
  56304=>"111111000",
  56305=>"111111110",
  56306=>"000000000",
  56307=>"100000100",
  56308=>"111111111",
  56309=>"001001111",
  56310=>"000100110",
  56311=>"111111111",
  56312=>"010110000",
  56313=>"000000100",
  56314=>"100100000",
  56315=>"000000000",
  56316=>"110000000",
  56317=>"000000101",
  56318=>"001111111",
  56319=>"111111111",
  56320=>"111011001",
  56321=>"111000000",
  56322=>"111111111",
  56323=>"000001000",
  56324=>"000001111",
  56325=>"001111111",
  56326=>"000000000",
  56327=>"111111111",
  56328=>"110111111",
  56329=>"000000000",
  56330=>"111110000",
  56331=>"111111000",
  56332=>"000100110",
  56333=>"001000000",
  56334=>"000100111",
  56335=>"000000000",
  56336=>"000000000",
  56337=>"000010000",
  56338=>"110111111",
  56339=>"000000111",
  56340=>"000000000",
  56341=>"110111111",
  56342=>"100111101",
  56343=>"000001011",
  56344=>"000001111",
  56345=>"000001001",
  56346=>"000000000",
  56347=>"111010000",
  56348=>"111111111",
  56349=>"000000000",
  56350=>"011010010",
  56351=>"001000000",
  56352=>"000000000",
  56353=>"100000000",
  56354=>"000000000",
  56355=>"001111111",
  56356=>"000000000",
  56357=>"100000000",
  56358=>"000000000",
  56359=>"111111000",
  56360=>"000011111",
  56361=>"000110110",
  56362=>"110111010",
  56363=>"110111111",
  56364=>"000001000",
  56365=>"000000000",
  56366=>"001011000",
  56367=>"000000000",
  56368=>"011111111",
  56369=>"000001111",
  56370=>"000010010",
  56371=>"100000011",
  56372=>"000001010",
  56373=>"011111111",
  56374=>"011001111",
  56375=>"000000101",
  56376=>"111111011",
  56377=>"000000001",
  56378=>"100111111",
  56379=>"100100000",
  56380=>"111111000",
  56381=>"111111111",
  56382=>"000000111",
  56383=>"111111111",
  56384=>"111101111",
  56385=>"111111110",
  56386=>"000111111",
  56387=>"111111111",
  56388=>"110111000",
  56389=>"000111011",
  56390=>"011000000",
  56391=>"101000100",
  56392=>"111110100",
  56393=>"000000000",
  56394=>"000000000",
  56395=>"100000000",
  56396=>"001001001",
  56397=>"000000000",
  56398=>"110111111",
  56399=>"101101101",
  56400=>"000000000",
  56401=>"111111000",
  56402=>"010110100",
  56403=>"000011001",
  56404=>"111111111",
  56405=>"001001001",
  56406=>"111100100",
  56407=>"000100100",
  56408=>"001001111",
  56409=>"101000101",
  56410=>"000000000",
  56411=>"001001001",
  56412=>"000000000",
  56413=>"100100000",
  56414=>"101111101",
  56415=>"100110110",
  56416=>"111100000",
  56417=>"000000111",
  56418=>"111111100",
  56419=>"000000111",
  56420=>"111001111",
  56421=>"111111101",
  56422=>"110000000",
  56423=>"101111111",
  56424=>"111101111",
  56425=>"111110000",
  56426=>"111011111",
  56427=>"110110110",
  56428=>"100000111",
  56429=>"000111010",
  56430=>"000000000",
  56431=>"000111111",
  56432=>"111111000",
  56433=>"000000011",
  56434=>"000000101",
  56435=>"001000000",
  56436=>"011000000",
  56437=>"111111111",
  56438=>"110000000",
  56439=>"000000000",
  56440=>"000110111",
  56441=>"001111111",
  56442=>"000000000",
  56443=>"000000000",
  56444=>"110000001",
  56445=>"000000000",
  56446=>"100110100",
  56447=>"111111111",
  56448=>"011111111",
  56449=>"000000111",
  56450=>"000000100",
  56451=>"011001000",
  56452=>"100100111",
  56453=>"000000000",
  56454=>"111111111",
  56455=>"101001001",
  56456=>"111111111",
  56457=>"001001010",
  56458=>"000000001",
  56459=>"000011111",
  56460=>"110111111",
  56461=>"110110111",
  56462=>"100001001",
  56463=>"000000000",
  56464=>"111111011",
  56465=>"111111111",
  56466=>"000000000",
  56467=>"010110110",
  56468=>"001001111",
  56469=>"000000000",
  56470=>"000001111",
  56471=>"111111000",
  56472=>"000111000",
  56473=>"100111111",
  56474=>"000000000",
  56475=>"010111111",
  56476=>"011111111",
  56477=>"111111000",
  56478=>"111001111",
  56479=>"110111010",
  56480=>"011111111",
  56481=>"000000111",
  56482=>"111111100",
  56483=>"111111111",
  56484=>"100100110",
  56485=>"000001111",
  56486=>"111111010",
  56487=>"011111101",
  56488=>"111111111",
  56489=>"011111111",
  56490=>"000000111",
  56491=>"111111111",
  56492=>"111111110",
  56493=>"100110110",
  56494=>"111111111",
  56495=>"101111111",
  56496=>"001000111",
  56497=>"100100000",
  56498=>"011011111",
  56499=>"111111111",
  56500=>"110000000",
  56501=>"100111111",
  56502=>"100111111",
  56503=>"111111101",
  56504=>"000011111",
  56505=>"000001000",
  56506=>"000000000",
  56507=>"000001001",
  56508=>"000000000",
  56509=>"111111000",
  56510=>"000000000",
  56511=>"111110110",
  56512=>"010011011",
  56513=>"011010000",
  56514=>"110110110",
  56515=>"111111111",
  56516=>"000000000",
  56517=>"000101111",
  56518=>"111111111",
  56519=>"111111111",
  56520=>"111111111",
  56521=>"100100000",
  56522=>"001100101",
  56523=>"000000000",
  56524=>"111111000",
  56525=>"101011000",
  56526=>"000000000",
  56527=>"000000000",
  56528=>"111011000",
  56529=>"111111000",
  56530=>"000000101",
  56531=>"000001010",
  56532=>"001000000",
  56533=>"000001111",
  56534=>"111111000",
  56535=>"110110111",
  56536=>"000101111",
  56537=>"111011111",
  56538=>"001000100",
  56539=>"000000000",
  56540=>"111001000",
  56541=>"111111111",
  56542=>"001111000",
  56543=>"000000000",
  56544=>"000011111",
  56545=>"111110000",
  56546=>"111111111",
  56547=>"100110110",
  56548=>"111111111",
  56549=>"000000000",
  56550=>"000000001",
  56551=>"100000000",
  56552=>"111111111",
  56553=>"111111111",
  56554=>"110100111",
  56555=>"000000000",
  56556=>"000000000",
  56557=>"000111111",
  56558=>"100111010",
  56559=>"111111111",
  56560=>"000001001",
  56561=>"000111111",
  56562=>"000000000",
  56563=>"111011000",
  56564=>"000000000",
  56565=>"001000100",
  56566=>"000001001",
  56567=>"001111111",
  56568=>"101101001",
  56569=>"000001001",
  56570=>"111111111",
  56571=>"101111111",
  56572=>"100100000",
  56573=>"110111001",
  56574=>"000000000",
  56575=>"000000010",
  56576=>"000000000",
  56577=>"111111001",
  56578=>"000000111",
  56579=>"000000000",
  56580=>"000000111",
  56581=>"000000011",
  56582=>"111110000",
  56583=>"000000001",
  56584=>"110100100",
  56585=>"000010110",
  56586=>"000000000",
  56587=>"000100100",
  56588=>"001000111",
  56589=>"111111011",
  56590=>"111111111",
  56591=>"111100000",
  56592=>"000000101",
  56593=>"000001011",
  56594=>"111001001",
  56595=>"000000011",
  56596=>"110000000",
  56597=>"000000000",
  56598=>"100110000",
  56599=>"000000001",
  56600=>"000000001",
  56601=>"011111110",
  56602=>"111111111",
  56603=>"000100000",
  56604=>"001001000",
  56605=>"000000000",
  56606=>"010111111",
  56607=>"000000000",
  56608=>"111111111",
  56609=>"001000000",
  56610=>"000000000",
  56611=>"000111111",
  56612=>"000010111",
  56613=>"000000000",
  56614=>"011000000",
  56615=>"110110000",
  56616=>"000000000",
  56617=>"000000000",
  56618=>"011011000",
  56619=>"111111000",
  56620=>"000000000",
  56621=>"100111111",
  56622=>"000111100",
  56623=>"000000001",
  56624=>"011111111",
  56625=>"000000111",
  56626=>"001111111",
  56627=>"000001111",
  56628=>"100000111",
  56629=>"111111000",
  56630=>"000001111",
  56631=>"000011110",
  56632=>"111100100",
  56633=>"111111000",
  56634=>"010010000",
  56635=>"000000000",
  56636=>"001111111",
  56637=>"101001101",
  56638=>"000100100",
  56639=>"101111111",
  56640=>"000100111",
  56641=>"101000111",
  56642=>"100100001",
  56643=>"000000100",
  56644=>"000000000",
  56645=>"111011000",
  56646=>"111000000",
  56647=>"000000000",
  56648=>"111111111",
  56649=>"111001101",
  56650=>"011111111",
  56651=>"100101111",
  56652=>"111111111",
  56653=>"000000000",
  56654=>"000000000",
  56655=>"111111110",
  56656=>"000010111",
  56657=>"111111111",
  56658=>"101000111",
  56659=>"000000000",
  56660=>"111111100",
  56661=>"011011011",
  56662=>"111111111",
  56663=>"111111111",
  56664=>"011011001",
  56665=>"001010111",
  56666=>"111111111",
  56667=>"111110111",
  56668=>"111111111",
  56669=>"000000111",
  56670=>"111100100",
  56671=>"110111111",
  56672=>"000000111",
  56673=>"000000000",
  56674=>"000001111",
  56675=>"000000000",
  56676=>"000000111",
  56677=>"111001001",
  56678=>"010000000",
  56679=>"111111110",
  56680=>"011111101",
  56681=>"001000000",
  56682=>"110110111",
  56683=>"111101001",
  56684=>"011000000",
  56685=>"111001100",
  56686=>"000000000",
  56687=>"111111111",
  56688=>"000111100",
  56689=>"111111111",
  56690=>"110111111",
  56691=>"000000000",
  56692=>"000110010",
  56693=>"101101101",
  56694=>"000000000",
  56695=>"000000000",
  56696=>"111111110",
  56697=>"000000000",
  56698=>"000101111",
  56699=>"011111110",
  56700=>"111111111",
  56701=>"111110111",
  56702=>"000000000",
  56703=>"000000111",
  56704=>"000001000",
  56705=>"000000001",
  56706=>"000110110",
  56707=>"000000111",
  56708=>"110000111",
  56709=>"000111000",
  56710=>"000000000",
  56711=>"111010000",
  56712=>"111111111",
  56713=>"110100100",
  56714=>"110001000",
  56715=>"111111000",
  56716=>"111111111",
  56717=>"000000000",
  56718=>"000000001",
  56719=>"000111101",
  56720=>"111111111",
  56721=>"100000000",
  56722=>"100001001",
  56723=>"111111111",
  56724=>"111000100",
  56725=>"000011000",
  56726=>"111001000",
  56727=>"111100011",
  56728=>"000000101",
  56729=>"111001000",
  56730=>"100100101",
  56731=>"000000000",
  56732=>"100101111",
  56733=>"100100000",
  56734=>"000000000",
  56735=>"011110111",
  56736=>"000000000",
  56737=>"111111001",
  56738=>"000000001",
  56739=>"000000000",
  56740=>"101101100",
  56741=>"100101100",
  56742=>"111111111",
  56743=>"001000000",
  56744=>"011101000",
  56745=>"011011110",
  56746=>"000000000",
  56747=>"000111011",
  56748=>"011100000",
  56749=>"111111111",
  56750=>"111111111",
  56751=>"111111000",
  56752=>"111111111",
  56753=>"001000000",
  56754=>"000000000",
  56755=>"111111011",
  56756=>"000111101",
  56757=>"101001000",
  56758=>"000101111",
  56759=>"111011000",
  56760=>"100001111",
  56761=>"111000111",
  56762=>"110110000",
  56763=>"000000111",
  56764=>"111001111",
  56765=>"111100111",
  56766=>"011111000",
  56767=>"000001000",
  56768=>"001000000",
  56769=>"111111111",
  56770=>"111111111",
  56771=>"111111101",
  56772=>"000000111",
  56773=>"111111111",
  56774=>"000000000",
  56775=>"111111100",
  56776=>"111111111",
  56777=>"000111111",
  56778=>"000000001",
  56779=>"110111000",
  56780=>"000111111",
  56781=>"111001101",
  56782=>"111111001",
  56783=>"000000100",
  56784=>"000111111",
  56785=>"111111110",
  56786=>"000000000",
  56787=>"111111111",
  56788=>"011001000",
  56789=>"111110110",
  56790=>"111111111",
  56791=>"001011011",
  56792=>"111000000",
  56793=>"111110011",
  56794=>"111110000",
  56795=>"001100111",
  56796=>"010111111",
  56797=>"110000000",
  56798=>"100000000",
  56799=>"000001011",
  56800=>"111111111",
  56801=>"000000000",
  56802=>"000000000",
  56803=>"000000000",
  56804=>"011111111",
  56805=>"101101001",
  56806=>"001000000",
  56807=>"000000000",
  56808=>"110000000",
  56809=>"111111111",
  56810=>"111111111",
  56811=>"000001111",
  56812=>"010111101",
  56813=>"011001001",
  56814=>"111111111",
  56815=>"000001101",
  56816=>"000000001",
  56817=>"000001111",
  56818=>"111000000",
  56819=>"000111100",
  56820=>"110000100",
  56821=>"011111111",
  56822=>"111111101",
  56823=>"111011111",
  56824=>"001000000",
  56825=>"101111111",
  56826=>"000000000",
  56827=>"101111111",
  56828=>"100000000",
  56829=>"111111111",
  56830=>"001100111",
  56831=>"111111111",
  56832=>"000010000",
  56833=>"010110111",
  56834=>"000100111",
  56835=>"000000000",
  56836=>"000010111",
  56837=>"111011000",
  56838=>"000000111",
  56839=>"111000000",
  56840=>"111001001",
  56841=>"000000000",
  56842=>"001000011",
  56843=>"111110110",
  56844=>"110111011",
  56845=>"111011111",
  56846=>"110100000",
  56847=>"110110111",
  56848=>"000111111",
  56849=>"000011000",
  56850=>"000000100",
  56851=>"000001011",
  56852=>"001000000",
  56853=>"111111000",
  56854=>"000000000",
  56855=>"110011011",
  56856=>"000000000",
  56857=>"000000000",
  56858=>"111111000",
  56859=>"001000110",
  56860=>"000110111",
  56861=>"111111001",
  56862=>"011000111",
  56863=>"000000111",
  56864=>"111110000",
  56865=>"100111000",
  56866=>"111111111",
  56867=>"000010110",
  56868=>"001001111",
  56869=>"111001001",
  56870=>"010011111",
  56871=>"000000111",
  56872=>"110111010",
  56873=>"000001111",
  56874=>"111111111",
  56875=>"111001111",
  56876=>"111111001",
  56877=>"000001000",
  56878=>"111111111",
  56879=>"011000001",
  56880=>"000011000",
  56881=>"000111111",
  56882=>"000100000",
  56883=>"010000001",
  56884=>"000000000",
  56885=>"111111111",
  56886=>"000000000",
  56887=>"000101001",
  56888=>"000000000",
  56889=>"000100000",
  56890=>"000000000",
  56891=>"011111000",
  56892=>"000000111",
  56893=>"011000100",
  56894=>"001000000",
  56895=>"100000001",
  56896=>"100110111",
  56897=>"111111101",
  56898=>"100000000",
  56899=>"111011111",
  56900=>"011000001",
  56901=>"111111110",
  56902=>"111001111",
  56903=>"000011000",
  56904=>"011111111",
  56905=>"111111000",
  56906=>"111001000",
  56907=>"000000000",
  56908=>"111000000",
  56909=>"100111000",
  56910=>"111010111",
  56911=>"111111111",
  56912=>"100000000",
  56913=>"111111011",
  56914=>"000000000",
  56915=>"111101001",
  56916=>"000000111",
  56917=>"000000100",
  56918=>"001000101",
  56919=>"000000000",
  56920=>"111100000",
  56921=>"000000101",
  56922=>"101000000",
  56923=>"111000000",
  56924=>"000000101",
  56925=>"111100101",
  56926=>"011000000",
  56927=>"100110110",
  56928=>"110000000",
  56929=>"101000000",
  56930=>"000000000",
  56931=>"000000000",
  56932=>"000000111",
  56933=>"110000111",
  56934=>"111110000",
  56935=>"110111111",
  56936=>"111111001",
  56937=>"000000000",
  56938=>"111110000",
  56939=>"000000110",
  56940=>"000001111",
  56941=>"001111011",
  56942=>"111111110",
  56943=>"111111011",
  56944=>"001011001",
  56945=>"110000000",
  56946=>"011111110",
  56947=>"111000111",
  56948=>"011000000",
  56949=>"000001000",
  56950=>"000000001",
  56951=>"000000110",
  56952=>"010111111",
  56953=>"000000101",
  56954=>"011111111",
  56955=>"111011010",
  56956=>"001111001",
  56957=>"000110000",
  56958=>"011111111",
  56959=>"011001000",
  56960=>"110100110",
  56961=>"111111001",
  56962=>"000000001",
  56963=>"111000000",
  56964=>"110000110",
  56965=>"000111001",
  56966=>"110010110",
  56967=>"000000000",
  56968=>"011000000",
  56969=>"000000000",
  56970=>"111110110",
  56971=>"000000111",
  56972=>"111111101",
  56973=>"111000000",
  56974=>"000000000",
  56975=>"000000100",
  56976=>"000111111",
  56977=>"011111111",
  56978=>"111000100",
  56979=>"111001000",
  56980=>"000110110",
  56981=>"001111000",
  56982=>"111100111",
  56983=>"011111111",
  56984=>"111111000",
  56985=>"011010000",
  56986=>"001111111",
  56987=>"111000000",
  56988=>"001000000",
  56989=>"110000100",
  56990=>"111111000",
  56991=>"111000110",
  56992=>"111111111",
  56993=>"000000111",
  56994=>"111001111",
  56995=>"011000000",
  56996=>"010111110",
  56997=>"001000111",
  56998=>"001011110",
  56999=>"111111000",
  57000=>"111110111",
  57001=>"000000001",
  57002=>"000000000",
  57003=>"111111111",
  57004=>"110000000",
  57005=>"101000000",
  57006=>"000000100",
  57007=>"010010111",
  57008=>"111111000",
  57009=>"000100111",
  57010=>"111111010",
  57011=>"000100101",
  57012=>"111000000",
  57013=>"100000001",
  57014=>"000110110",
  57015=>"000000000",
  57016=>"100111111",
  57017=>"000000000",
  57018=>"000000000",
  57019=>"001111011",
  57020=>"111101111",
  57021=>"111000000",
  57022=>"111111000",
  57023=>"111100000",
  57024=>"000111111",
  57025=>"000010111",
  57026=>"000000000",
  57027=>"011000000",
  57028=>"000011000",
  57029=>"011111111",
  57030=>"110000000",
  57031=>"000000011",
  57032=>"111111111",
  57033=>"000000111",
  57034=>"000000010",
  57035=>"000111111",
  57036=>"011000110",
  57037=>"111011111",
  57038=>"111000000",
  57039=>"000000100",
  57040=>"000000111",
  57041=>"111011110",
  57042=>"001000000",
  57043=>"000001101",
  57044=>"000000000",
  57045=>"111100000",
  57046=>"111000001",
  57047=>"000000111",
  57048=>"000000111",
  57049=>"111000111",
  57050=>"001000000",
  57051=>"101000000",
  57052=>"111000000",
  57053=>"000000000",
  57054=>"000110001",
  57055=>"100000000",
  57056=>"000000000",
  57057=>"111111111",
  57058=>"111111111",
  57059=>"101000111",
  57060=>"000001111",
  57061=>"000000010",
  57062=>"000000100",
  57063=>"001000111",
  57064=>"100000000",
  57065=>"000000011",
  57066=>"111000000",
  57067=>"000001001",
  57068=>"000000000",
  57069=>"111000001",
  57070=>"101000111",
  57071=>"000000010",
  57072=>"000000000",
  57073=>"000000000",
  57074=>"111100000",
  57075=>"111110000",
  57076=>"001000010",
  57077=>"001001001",
  57078=>"110100101",
  57079=>"000000000",
  57080=>"111111111",
  57081=>"111111000",
  57082=>"111100111",
  57083=>"001001010",
  57084=>"111111000",
  57085=>"010000001",
  57086=>"101000000",
  57087=>"001000000",
  57088=>"111110100",
  57089=>"000000110",
  57090=>"001001000",
  57091=>"111110111",
  57092=>"000000000",
  57093=>"000110111",
  57094=>"100010110",
  57095=>"000000111",
  57096=>"111100111",
  57097=>"000000000",
  57098=>"001001000",
  57099=>"111111111",
  57100=>"000010010",
  57101=>"000001000",
  57102=>"011011111",
  57103=>"000000000",
  57104=>"111101000",
  57105=>"111000011",
  57106=>"011011000",
  57107=>"010010010",
  57108=>"000111111",
  57109=>"000000000",
  57110=>"000000001",
  57111=>"000111111",
  57112=>"100101001",
  57113=>"100111111",
  57114=>"000000001",
  57115=>"100000000",
  57116=>"000111111",
  57117=>"111000000",
  57118=>"010000000",
  57119=>"000000100",
  57120=>"001000011",
  57121=>"100000000",
  57122=>"111110000",
  57123=>"101111100",
  57124=>"000111111",
  57125=>"110110100",
  57126=>"111111111",
  57127=>"111111000",
  57128=>"100111000",
  57129=>"000000000",
  57130=>"010110111",
  57131=>"000111100",
  57132=>"000000110",
  57133=>"000001101",
  57134=>"001001110",
  57135=>"000000111",
  57136=>"100111111",
  57137=>"001001000",
  57138=>"111111111",
  57139=>"000000000",
  57140=>"111000000",
  57141=>"111011011",
  57142=>"111000000",
  57143=>"111110000",
  57144=>"000000000",
  57145=>"001000111",
  57146=>"101001111",
  57147=>"111000001",
  57148=>"111111000",
  57149=>"000000010",
  57150=>"110000100",
  57151=>"000000111",
  57152=>"000000011",
  57153=>"101001000",
  57154=>"111000001",
  57155=>"000000111",
  57156=>"111111111",
  57157=>"100000000",
  57158=>"010111110",
  57159=>"011011011",
  57160=>"111000111",
  57161=>"001000000",
  57162=>"111111111",
  57163=>"110100111",
  57164=>"111111000",
  57165=>"010010111",
  57166=>"101000011",
  57167=>"100100111",
  57168=>"001000001",
  57169=>"111011001",
  57170=>"100111101",
  57171=>"111111111",
  57172=>"000000001",
  57173=>"001111101",
  57174=>"000111111",
  57175=>"111110101",
  57176=>"111100111",
  57177=>"111000000",
  57178=>"111111011",
  57179=>"000000110",
  57180=>"100000111",
  57181=>"011110100",
  57182=>"011111111",
  57183=>"001000000",
  57184=>"000000111",
  57185=>"111111010",
  57186=>"000000000",
  57187=>"111000000",
  57188=>"111111111",
  57189=>"000000000",
  57190=>"111111010",
  57191=>"100111011",
  57192=>"001001101",
  57193=>"000011011",
  57194=>"000001001",
  57195=>"000111111",
  57196=>"111111111",
  57197=>"011111000",
  57198=>"111110100",
  57199=>"001000000",
  57200=>"111001010",
  57201=>"111001001",
  57202=>"011000000",
  57203=>"111011110",
  57204=>"111001000",
  57205=>"000110000",
  57206=>"111111111",
  57207=>"000111111",
  57208=>"000000100",
  57209=>"111000000",
  57210=>"001000000",
  57211=>"111001000",
  57212=>"000001111",
  57213=>"001001000",
  57214=>"111111000",
  57215=>"000000000",
  57216=>"110010000",
  57217=>"000010010",
  57218=>"111111001",
  57219=>"000000100",
  57220=>"111000001",
  57221=>"000110110",
  57222=>"111101000",
  57223=>"000010000",
  57224=>"000011100",
  57225=>"111111111",
  57226=>"000000000",
  57227=>"000000100",
  57228=>"000000001",
  57229=>"001000111",
  57230=>"000100100",
  57231=>"010010000",
  57232=>"000111101",
  57233=>"111111000",
  57234=>"111000111",
  57235=>"111110000",
  57236=>"111111000",
  57237=>"111011000",
  57238=>"000000000",
  57239=>"110000011",
  57240=>"000000111",
  57241=>"000001011",
  57242=>"001000010",
  57243=>"111010000",
  57244=>"111111011",
  57245=>"111110111",
  57246=>"000111111",
  57247=>"001000000",
  57248=>"111000000",
  57249=>"111110110",
  57250=>"000001001",
  57251=>"111000000",
  57252=>"000000000",
  57253=>"111111111",
  57254=>"000000111",
  57255=>"101111111",
  57256=>"111000000",
  57257=>"000111111",
  57258=>"111001111",
  57259=>"000111111",
  57260=>"111111111",
  57261=>"111000000",
  57262=>"111000111",
  57263=>"111010000",
  57264=>"100110100",
  57265=>"100111111",
  57266=>"000101111",
  57267=>"111000000",
  57268=>"000110111",
  57269=>"011011111",
  57270=>"110111111",
  57271=>"111111000",
  57272=>"000000011",
  57273=>"111000000",
  57274=>"000000000",
  57275=>"110000000",
  57276=>"111000111",
  57277=>"000000011",
  57278=>"001001000",
  57279=>"001011111",
  57280=>"111111111",
  57281=>"000000000",
  57282=>"111111110",
  57283=>"111000111",
  57284=>"000000101",
  57285=>"011111110",
  57286=>"000000001",
  57287=>"000001000",
  57288=>"111000100",
  57289=>"000111111",
  57290=>"111000000",
  57291=>"000110111",
  57292=>"000000100",
  57293=>"111111111",
  57294=>"000100111",
  57295=>"011000011",
  57296=>"000000111",
  57297=>"111011001",
  57298=>"000111111",
  57299=>"101000111",
  57300=>"110110110",
  57301=>"100111000",
  57302=>"111111000",
  57303=>"000100110",
  57304=>"111000111",
  57305=>"111111001",
  57306=>"000111001",
  57307=>"001000100",
  57308=>"110111111",
  57309=>"111111001",
  57310=>"000001010",
  57311=>"011000000",
  57312=>"000001111",
  57313=>"110000111",
  57314=>"111111100",
  57315=>"111111011",
  57316=>"111111111",
  57317=>"100001001",
  57318=>"000001111",
  57319=>"101100111",
  57320=>"000000000",
  57321=>"111011001",
  57322=>"100111000",
  57323=>"000000101",
  57324=>"111111111",
  57325=>"110111000",
  57326=>"000111111",
  57327=>"000000000",
  57328=>"000111111",
  57329=>"100111111",
  57330=>"111000000",
  57331=>"111000000",
  57332=>"111111111",
  57333=>"001001000",
  57334=>"000000000",
  57335=>"111001001",
  57336=>"000110000",
  57337=>"000110110",
  57338=>"110000000",
  57339=>"111000000",
  57340=>"000110011",
  57341=>"011001001",
  57342=>"000000111",
  57343=>"100111111",
  57344=>"011000000",
  57345=>"100111000",
  57346=>"101100100",
  57347=>"010110011",
  57348=>"000000101",
  57349=>"110111000",
  57350=>"000000000",
  57351=>"111111000",
  57352=>"111011111",
  57353=>"111110111",
  57354=>"000000000",
  57355=>"111010010",
  57356=>"100100110",
  57357=>"101000001",
  57358=>"000000000",
  57359=>"000000000",
  57360=>"111000100",
  57361=>"000010001",
  57362=>"001111111",
  57363=>"111101111",
  57364=>"100000000",
  57365=>"000000000",
  57366=>"111111111",
  57367=>"001000000",
  57368=>"001000111",
  57369=>"000100100",
  57370=>"000011000",
  57371=>"000111010",
  57372=>"111111111",
  57373=>"111001111",
  57374=>"100111010",
  57375=>"110111111",
  57376=>"011010000",
  57377=>"101111100",
  57378=>"010110001",
  57379=>"111111110",
  57380=>"111111011",
  57381=>"111111011",
  57382=>"000011000",
  57383=>"001101011",
  57384=>"000011000",
  57385=>"000101000",
  57386=>"111111111",
  57387=>"111110111",
  57388=>"000000100",
  57389=>"111110110",
  57390=>"101000000",
  57391=>"111111011",
  57392=>"111111100",
  57393=>"000000010",
  57394=>"001001001",
  57395=>"011000000",
  57396=>"000000111",
  57397=>"001001111",
  57398=>"000100000",
  57399=>"111111111",
  57400=>"000000101",
  57401=>"000000000",
  57402=>"000000000",
  57403=>"000000000",
  57404=>"111000111",
  57405=>"000000111",
  57406=>"111111111",
  57407=>"111000000",
  57408=>"111010100",
  57409=>"110000111",
  57410=>"111100111",
  57411=>"111111111",
  57412=>"000000000",
  57413=>"100111011",
  57414=>"111001000",
  57415=>"111000000",
  57416=>"100100100",
  57417=>"000000111",
  57418=>"111011011",
  57419=>"000110111",
  57420=>"000011100",
  57421=>"010000100",
  57422=>"101000000",
  57423=>"010000111",
  57424=>"000001101",
  57425=>"111111111",
  57426=>"001000000",
  57427=>"010011011",
  57428=>"111000010",
  57429=>"111110010",
  57430=>"001001001",
  57431=>"111111111",
  57432=>"000000000",
  57433=>"111101111",
  57434=>"111111111",
  57435=>"001110111",
  57436=>"000000000",
  57437=>"111111111",
  57438=>"000110000",
  57439=>"000101111",
  57440=>"000111111",
  57441=>"000000101",
  57442=>"111110000",
  57443=>"000110110",
  57444=>"001111000",
  57445=>"010110011",
  57446=>"000100111",
  57447=>"110100000",
  57448=>"111000000",
  57449=>"000000000",
  57450=>"111110000",
  57451=>"001001000",
  57452=>"111111000",
  57453=>"000000000",
  57454=>"011111111",
  57455=>"001000000",
  57456=>"000000001",
  57457=>"000000000",
  57458=>"111000111",
  57459=>"010111011",
  57460=>"011011111",
  57461=>"000111111",
  57462=>"010111000",
  57463=>"001000000",
  57464=>"110000001",
  57465=>"010000111",
  57466=>"000100111",
  57467=>"111000111",
  57468=>"001001100",
  57469=>"000111011",
  57470=>"100100110",
  57471=>"011101000",
  57472=>"000000000",
  57473=>"000000011",
  57474=>"000000000",
  57475=>"001000011",
  57476=>"011111111",
  57477=>"111000101",
  57478=>"001001111",
  57479=>"000111111",
  57480=>"001001111",
  57481=>"110000000",
  57482=>"000100100",
  57483=>"111111011",
  57484=>"000001111",
  57485=>"000000000",
  57486=>"100000100",
  57487=>"000000001",
  57488=>"111000111",
  57489=>"111110111",
  57490=>"000000001",
  57491=>"001000000",
  57492=>"010010000",
  57493=>"000111001",
  57494=>"111000000",
  57495=>"001000111",
  57496=>"011000011",
  57497=>"001000001",
  57498=>"111111111",
  57499=>"101011000",
  57500=>"101111111",
  57501=>"011011001",
  57502=>"111000110",
  57503=>"000000000",
  57504=>"010111111",
  57505=>"001000001",
  57506=>"111111001",
  57507=>"111001111",
  57508=>"000000000",
  57509=>"000111000",
  57510=>"111111110",
  57511=>"010010111",
  57512=>"111011011",
  57513=>"011110000",
  57514=>"111100000",
  57515=>"111000001",
  57516=>"000000111",
  57517=>"110110001",
  57518=>"001000100",
  57519=>"000100000",
  57520=>"000001111",
  57521=>"000111001",
  57522=>"010111000",
  57523=>"000001111",
  57524=>"011111010",
  57525=>"111000111",
  57526=>"011000000",
  57527=>"101100000",
  57528=>"000000000",
  57529=>"101000101",
  57530=>"000000111",
  57531=>"000000000",
  57532=>"011000000",
  57533=>"001001111",
  57534=>"111000111",
  57535=>"110000011",
  57536=>"011111111",
  57537=>"001011000",
  57538=>"001000000",
  57539=>"111111111",
  57540=>"111000001",
  57541=>"000111111",
  57542=>"011000000",
  57543=>"010111000",
  57544=>"001111000",
  57545=>"111001000",
  57546=>"000000011",
  57547=>"100111111",
  57548=>"000000101",
  57549=>"000100000",
  57550=>"000000000",
  57551=>"110000110",
  57552=>"010111011",
  57553=>"001110000",
  57554=>"000000000",
  57555=>"001000010",
  57556=>"000000101",
  57557=>"111111001",
  57558=>"100000100",
  57559=>"110010000",
  57560=>"110110000",
  57561=>"111010100",
  57562=>"111000111",
  57563=>"000111001",
  57564=>"000010010",
  57565=>"001001001",
  57566=>"111011000",
  57567=>"010000000",
  57568=>"001000010",
  57569=>"000111000",
  57570=>"110011000",
  57571=>"000111000",
  57572=>"111001111",
  57573=>"000110111",
  57574=>"000110000",
  57575=>"000000000",
  57576=>"111000001",
  57577=>"000000100",
  57578=>"111011111",
  57579=>"111110000",
  57580=>"111101000",
  57581=>"101101000",
  57582=>"111010111",
  57583=>"111001000",
  57584=>"111111111",
  57585=>"100000000",
  57586=>"000001111",
  57587=>"000101111",
  57588=>"000000000",
  57589=>"000110010",
  57590=>"011011000",
  57591=>"010110000",
  57592=>"000000001",
  57593=>"010010110",
  57594=>"111111011",
  57595=>"101111111",
  57596=>"011101111",
  57597=>"011011011",
  57598=>"001111111",
  57599=>"111010010",
  57600=>"010010011",
  57601=>"101000101",
  57602=>"100100100",
  57603=>"010000111",
  57604=>"111110010",
  57605=>"001001111",
  57606=>"111111111",
  57607=>"001011010",
  57608=>"000011001",
  57609=>"000000101",
  57610=>"111000000",
  57611=>"111111111",
  57612=>"101110000",
  57613=>"111000000",
  57614=>"001111000",
  57615=>"000000000",
  57616=>"011111111",
  57617=>"111111111",
  57618=>"111000001",
  57619=>"000111111",
  57620=>"100000001",
  57621=>"010000000",
  57622=>"001001001",
  57623=>"000000000",
  57624=>"011010111",
  57625=>"000000100",
  57626=>"000010011",
  57627=>"001001000",
  57628=>"000111110",
  57629=>"101111000",
  57630=>"111111111",
  57631=>"000100000",
  57632=>"100111011",
  57633=>"010010000",
  57634=>"011011111",
  57635=>"111111000",
  57636=>"111111000",
  57637=>"000000000",
  57638=>"111001000",
  57639=>"101001011",
  57640=>"000000111",
  57641=>"000000000",
  57642=>"000001000",
  57643=>"101111100",
  57644=>"001001001",
  57645=>"011001011",
  57646=>"001000000",
  57647=>"001111000",
  57648=>"111111011",
  57649=>"111011111",
  57650=>"111110000",
  57651=>"010011000",
  57652=>"000000000",
  57653=>"011000000",
  57654=>"010110101",
  57655=>"001000100",
  57656=>"000111000",
  57657=>"111111111",
  57658=>"000000001",
  57659=>"000010111",
  57660=>"111101100",
  57661=>"110110101",
  57662=>"111010000",
  57663=>"000000001",
  57664=>"111011001",
  57665=>"111100111",
  57666=>"000111000",
  57667=>"111000000",
  57668=>"111111100",
  57669=>"001011111",
  57670=>"111000000",
  57671=>"000110100",
  57672=>"000001000",
  57673=>"000111000",
  57674=>"000000101",
  57675=>"001101110",
  57676=>"110000000",
  57677=>"010010000",
  57678=>"000000100",
  57679=>"001001100",
  57680=>"101111100",
  57681=>"000000011",
  57682=>"000000000",
  57683=>"111011000",
  57684=>"011000000",
  57685=>"100110011",
  57686=>"001111111",
  57687=>"010111110",
  57688=>"100000101",
  57689=>"000111000",
  57690=>"000000111",
  57691=>"111000011",
  57692=>"011000011",
  57693=>"000000001",
  57694=>"001001001",
  57695=>"111111100",
  57696=>"010000000",
  57697=>"111110111",
  57698=>"001111000",
  57699=>"101000000",
  57700=>"000100111",
  57701=>"001001000",
  57702=>"010111110",
  57703=>"110110000",
  57704=>"011001001",
  57705=>"110100111",
  57706=>"000000000",
  57707=>"111111101",
  57708=>"001111000",
  57709=>"101110000",
  57710=>"000000000",
  57711=>"111001111",
  57712=>"001000000",
  57713=>"000110000",
  57714=>"000011010",
  57715=>"100000000",
  57716=>"010001000",
  57717=>"001000000",
  57718=>"000100111",
  57719=>"101000000",
  57720=>"100000000",
  57721=>"010110000",
  57722=>"000000000",
  57723=>"001001111",
  57724=>"111111010",
  57725=>"111111000",
  57726=>"000010111",
  57727=>"111000001",
  57728=>"000000111",
  57729=>"010010000",
  57730=>"011011011",
  57731=>"111001000",
  57732=>"000111111",
  57733=>"100100101",
  57734=>"000000111",
  57735=>"000001000",
  57736=>"111000000",
  57737=>"111101101",
  57738=>"011000001",
  57739=>"111111000",
  57740=>"111111111",
  57741=>"111011011",
  57742=>"000000000",
  57743=>"110010001",
  57744=>"111111010",
  57745=>"111100111",
  57746=>"000000000",
  57747=>"111111111",
  57748=>"101111111",
  57749=>"000000000",
  57750=>"111111111",
  57751=>"100100101",
  57752=>"110111101",
  57753=>"010010111",
  57754=>"000000000",
  57755=>"000100001",
  57756=>"111010111",
  57757=>"011111110",
  57758=>"111000111",
  57759=>"000000000",
  57760=>"011000110",
  57761=>"100110001",
  57762=>"000110010",
  57763=>"111101001",
  57764=>"100000000",
  57765=>"111000000",
  57766=>"001001000",
  57767=>"000110000",
  57768=>"001110110",
  57769=>"110111000",
  57770=>"011111111",
  57771=>"001101111",
  57772=>"000001000",
  57773=>"100111001",
  57774=>"000000000",
  57775=>"001111111",
  57776=>"000001101",
  57777=>"000000000",
  57778=>"001010000",
  57779=>"000111010",
  57780=>"111111110",
  57781=>"000111111",
  57782=>"110000000",
  57783=>"001000000",
  57784=>"111011000",
  57785=>"000000100",
  57786=>"111101000",
  57787=>"111000111",
  57788=>"101101001",
  57789=>"111000000",
  57790=>"110111111",
  57791=>"100100100",
  57792=>"101101011",
  57793=>"001001000",
  57794=>"111100000",
  57795=>"111000000",
  57796=>"111111111",
  57797=>"101111100",
  57798=>"010110010",
  57799=>"000110110",
  57800=>"100000010",
  57801=>"111000100",
  57802=>"011111000",
  57803=>"111000000",
  57804=>"110000000",
  57805=>"111110000",
  57806=>"110110110",
  57807=>"001000000",
  57808=>"101001001",
  57809=>"000101001",
  57810=>"000101100",
  57811=>"010000001",
  57812=>"111111000",
  57813=>"100100000",
  57814=>"010100111",
  57815=>"000000001",
  57816=>"000000111",
  57817=>"111110111",
  57818=>"101111000",
  57819=>"000000111",
  57820=>"101101111",
  57821=>"000110000",
  57822=>"000100000",
  57823=>"001011111",
  57824=>"111111000",
  57825=>"000111111",
  57826=>"100000111",
  57827=>"000000010",
  57828=>"111011000",
  57829=>"011011011",
  57830=>"101101000",
  57831=>"111000000",
  57832=>"110100100",
  57833=>"111010010",
  57834=>"000011001",
  57835=>"000110000",
  57836=>"101111111",
  57837=>"011011111",
  57838=>"111110111",
  57839=>"111111111",
  57840=>"000000101",
  57841=>"000000111",
  57842=>"111100001",
  57843=>"000011011",
  57844=>"000110111",
  57845=>"111000000",
  57846=>"110101111",
  57847=>"011001001",
  57848=>"100000000",
  57849=>"011000100",
  57850=>"000000011",
  57851=>"000001000",
  57852=>"110111111",
  57853=>"111111000",
  57854=>"100111110",
  57855=>"101000101",
  57856=>"000000000",
  57857=>"000000000",
  57858=>"101111111",
  57859=>"111011001",
  57860=>"000110101",
  57861=>"001001001",
  57862=>"000000111",
  57863=>"111111111",
  57864=>"111111111",
  57865=>"000000001",
  57866=>"111111111",
  57867=>"000000111",
  57868=>"110010010",
  57869=>"011111110",
  57870=>"000000110",
  57871=>"111111111",
  57872=>"001111111",
  57873=>"000000000",
  57874=>"001111101",
  57875=>"111111111",
  57876=>"100100000",
  57877=>"000000111",
  57878=>"111011001",
  57879=>"001011011",
  57880=>"110110010",
  57881=>"000000000",
  57882=>"001001111",
  57883=>"001000000",
  57884=>"000111111",
  57885=>"110111111",
  57886=>"001011011",
  57887=>"011000100",
  57888=>"111111111",
  57889=>"100000000",
  57890=>"000000000",
  57891=>"111100000",
  57892=>"000110110",
  57893=>"111111111",
  57894=>"111001001",
  57895=>"000000000",
  57896=>"111111111",
  57897=>"111011010",
  57898=>"000111111",
  57899=>"111111111",
  57900=>"100101101",
  57901=>"111111010",
  57902=>"111111111",
  57903=>"111101000",
  57904=>"000000000",
  57905=>"000000000",
  57906=>"000000000",
  57907=>"100000000",
  57908=>"111111111",
  57909=>"100000110",
  57910=>"011111111",
  57911=>"000000000",
  57912=>"010000111",
  57913=>"000000000",
  57914=>"000000111",
  57915=>"111111111",
  57916=>"101000000",
  57917=>"111111111",
  57918=>"001011000",
  57919=>"111000111",
  57920=>"111111110",
  57921=>"000000000",
  57922=>"000000111",
  57923=>"000011000",
  57924=>"111011000",
  57925=>"000001011",
  57926=>"000000111",
  57927=>"111000000",
  57928=>"111111110",
  57929=>"000000101",
  57930=>"111111111",
  57931=>"000000000",
  57932=>"111111101",
  57933=>"011000000",
  57934=>"000000000",
  57935=>"111111111",
  57936=>"111111000",
  57937=>"101100101",
  57938=>"000010011",
  57939=>"110111111",
  57940=>"000000000",
  57941=>"000111111",
  57942=>"000000000",
  57943=>"000001000",
  57944=>"011010011",
  57945=>"000000111",
  57946=>"101101011",
  57947=>"000000010",
  57948=>"010000000",
  57949=>"000000111",
  57950=>"000000100",
  57951=>"110100000",
  57952=>"100000000",
  57953=>"111100100",
  57954=>"000100000",
  57955=>"000000000",
  57956=>"111111111",
  57957=>"000110110",
  57958=>"111111110",
  57959=>"000000000",
  57960=>"000000111",
  57961=>"111000000",
  57962=>"000100111",
  57963=>"000000000",
  57964=>"100000000",
  57965=>"000010010",
  57966=>"000000000",
  57967=>"000000111",
  57968=>"111111111",
  57969=>"000000000",
  57970=>"100100100",
  57971=>"000000000",
  57972=>"000000000",
  57973=>"111111011",
  57974=>"011111111",
  57975=>"000000000",
  57976=>"111110000",
  57977=>"111111111",
  57978=>"001011000",
  57979=>"000111111",
  57980=>"000110110",
  57981=>"000000000",
  57982=>"000111111",
  57983=>"001011001",
  57984=>"000000000",
  57985=>"100000000",
  57986=>"100000000",
  57987=>"100110111",
  57988=>"111111100",
  57989=>"111101101",
  57990=>"100100000",
  57991=>"111110111",
  57992=>"000000000",
  57993=>"000000111",
  57994=>"110000000",
  57995=>"111111111",
  57996=>"000000100",
  57997=>"001011011",
  57998=>"000000000",
  57999=>"000000000",
  58000=>"000000000",
  58001=>"010010000",
  58002=>"000001000",
  58003=>"100110110",
  58004=>"100100000",
  58005=>"000000110",
  58006=>"001111111",
  58007=>"111111111",
  58008=>"111000000",
  58009=>"111111111",
  58010=>"011001000",
  58011=>"100000000",
  58012=>"000000010",
  58013=>"000000100",
  58014=>"000000111",
  58015=>"111111111",
  58016=>"111111111",
  58017=>"111011000",
  58018=>"000000001",
  58019=>"000000000",
  58020=>"011011000",
  58021=>"000000001",
  58022=>"111100000",
  58023=>"001001011",
  58024=>"000100111",
  58025=>"001001000",
  58026=>"000000000",
  58027=>"001001001",
  58028=>"000000000",
  58029=>"110110110",
  58030=>"111111111",
  58031=>"010000000",
  58032=>"000000000",
  58033=>"000110110",
  58034=>"111111111",
  58035=>"000000000",
  58036=>"001001000",
  58037=>"000000100",
  58038=>"000000011",
  58039=>"000000000",
  58040=>"111111111",
  58041=>"000000000",
  58042=>"110010011",
  58043=>"111011111",
  58044=>"100000000",
  58045=>"000011111",
  58046=>"101111111",
  58047=>"111101111",
  58048=>"000011111",
  58049=>"111011100",
  58050=>"001111111",
  58051=>"000000111",
  58052=>"100000000",
  58053=>"111111111",
  58054=>"111111111",
  58055=>"011011111",
  58056=>"001000000",
  58057=>"000000000",
  58058=>"000000011",
  58059=>"111111011",
  58060=>"000000111",
  58061=>"000000000",
  58062=>"111111111",
  58063=>"000000000",
  58064=>"101000000",
  58065=>"001111111",
  58066=>"000000000",
  58067=>"011000000",
  58068=>"110011011",
  58069=>"110111110",
  58070=>"000000000",
  58071=>"000000000",
  58072=>"111001001",
  58073=>"011111111",
  58074=>"000010111",
  58075=>"000011011",
  58076=>"001001001",
  58077=>"010010000",
  58078=>"100000111",
  58079=>"111111111",
  58080=>"000000000",
  58081=>"000000111",
  58082=>"000000110",
  58083=>"000000000",
  58084=>"011111111",
  58085=>"000000001",
  58086=>"000000111",
  58087=>"111101000",
  58088=>"111111000",
  58089=>"110000010",
  58090=>"000000000",
  58091=>"110000110",
  58092=>"011111010",
  58093=>"000000000",
  58094=>"100110111",
  58095=>"111111111",
  58096=>"111110100",
  58097=>"000001111",
  58098=>"111111111",
  58099=>"110000000",
  58100=>"000100100",
  58101=>"011001000",
  58102=>"000000001",
  58103=>"100000000",
  58104=>"110101111",
  58105=>"111111111",
  58106=>"000000000",
  58107=>"101101101",
  58108=>"011000000",
  58109=>"000000111",
  58110=>"010000000",
  58111=>"000001000",
  58112=>"111000000",
  58113=>"100000000",
  58114=>"110110110",
  58115=>"111111000",
  58116=>"110111111",
  58117=>"000000000",
  58118=>"111001000",
  58119=>"011110000",
  58120=>"000000100",
  58121=>"000000000",
  58122=>"100001111",
  58123=>"111111111",
  58124=>"101001101",
  58125=>"010110110",
  58126=>"111111111",
  58127=>"111111001",
  58128=>"000001011",
  58129=>"000000011",
  58130=>"000000000",
  58131=>"000000000",
  58132=>"000110111",
  58133=>"000000000",
  58134=>"110110110",
  58135=>"010011110",
  58136=>"110111111",
  58137=>"000111111",
  58138=>"000100000",
  58139=>"000111111",
  58140=>"000110100",
  58141=>"011001000",
  58142=>"111111111",
  58143=>"111111100",
  58144=>"000000000",
  58145=>"111011111",
  58146=>"001111100",
  58147=>"000000100",
  58148=>"100111111",
  58149=>"000000000",
  58150=>"111111111",
  58151=>"111110000",
  58152=>"000000000",
  58153=>"111011011",
  58154=>"111000000",
  58155=>"110100000",
  58156=>"110110111",
  58157=>"111111000",
  58158=>"000000000",
  58159=>"000000000",
  58160=>"110100110",
  58161=>"000000010",
  58162=>"111000000",
  58163=>"111111111",
  58164=>"111101101",
  58165=>"000110000",
  58166=>"111001000",
  58167=>"110110111",
  58168=>"110010000",
  58169=>"101110111",
  58170=>"010000000",
  58171=>"100000000",
  58172=>"000011011",
  58173=>"000000011",
  58174=>"111100101",
  58175=>"011011011",
  58176=>"000010000",
  58177=>"111111000",
  58178=>"000000111",
  58179=>"000000000",
  58180=>"000000000",
  58181=>"000000111",
  58182=>"000000000",
  58183=>"000001001",
  58184=>"000000011",
  58185=>"111111111",
  58186=>"111111100",
  58187=>"111111111",
  58188=>"000000000",
  58189=>"000000100",
  58190=>"000000111",
  58191=>"111111111",
  58192=>"011001111",
  58193=>"111111111",
  58194=>"101111111",
  58195=>"111111111",
  58196=>"110110000",
  58197=>"011011011",
  58198=>"111111111",
  58199=>"011111111",
  58200=>"000101111",
  58201=>"000000000",
  58202=>"000000000",
  58203=>"110000000",
  58204=>"001011011",
  58205=>"000010011",
  58206=>"000100100",
  58207=>"010011010",
  58208=>"010000000",
  58209=>"111111111",
  58210=>"010010000",
  58211=>"100000100",
  58212=>"011111111",
  58213=>"000000000",
  58214=>"101101111",
  58215=>"011111111",
  58216=>"001001001",
  58217=>"100111110",
  58218=>"000000000",
  58219=>"000000000",
  58220=>"000010011",
  58221=>"111111111",
  58222=>"010110010",
  58223=>"000000000",
  58224=>"000000010",
  58225=>"111111011",
  58226=>"110110111",
  58227=>"011001011",
  58228=>"011000000",
  58229=>"111111111",
  58230=>"100010010",
  58231=>"000000100",
  58232=>"000000000",
  58233=>"000000000",
  58234=>"000000100",
  58235=>"111110111",
  58236=>"000000010",
  58237=>"111111111",
  58238=>"000000001",
  58239=>"000000000",
  58240=>"000000000",
  58241=>"010000100",
  58242=>"010010010",
  58243=>"100100100",
  58244=>"000000110",
  58245=>"111111111",
  58246=>"000100110",
  58247=>"001011000",
  58248=>"000010110",
  58249=>"100100000",
  58250=>"011111111",
  58251=>"111111111",
  58252=>"100100100",
  58253=>"111111111",
  58254=>"111111111",
  58255=>"000110000",
  58256=>"111000000",
  58257=>"111111111",
  58258=>"001000000",
  58259=>"010000000",
  58260=>"011001001",
  58261=>"010000000",
  58262=>"000000000",
  58263=>"110010110",
  58264=>"111001000",
  58265=>"000110111",
  58266=>"111111111",
  58267=>"111111110",
  58268=>"110111000",
  58269=>"000001000",
  58270=>"000000001",
  58271=>"001000000",
  58272=>"011111111",
  58273=>"100110111",
  58274=>"000000001",
  58275=>"111101101",
  58276=>"111100000",
  58277=>"111111111",
  58278=>"001000000",
  58279=>"000111111",
  58280=>"000000000",
  58281=>"001001001",
  58282=>"000000000",
  58283=>"111111011",
  58284=>"000000110",
  58285=>"001001100",
  58286=>"000110111",
  58287=>"000011111",
  58288=>"000000011",
  58289=>"111000000",
  58290=>"111111111",
  58291=>"111111000",
  58292=>"100100111",
  58293=>"111111101",
  58294=>"000000000",
  58295=>"111111111",
  58296=>"111000000",
  58297=>"111111110",
  58298=>"111110110",
  58299=>"000000000",
  58300=>"001001111",
  58301=>"000000000",
  58302=>"000000000",
  58303=>"111110110",
  58304=>"011011000",
  58305=>"111111111",
  58306=>"111111111",
  58307=>"001000001",
  58308=>"111111111",
  58309=>"000000101",
  58310=>"000000001",
  58311=>"111001000",
  58312=>"111000001",
  58313=>"100100100",
  58314=>"000000001",
  58315=>"111111011",
  58316=>"000000010",
  58317=>"111111111",
  58318=>"111001001",
  58319=>"110111111",
  58320=>"000000000",
  58321=>"011111111",
  58322=>"111001010",
  58323=>"111111111",
  58324=>"100100110",
  58325=>"000000111",
  58326=>"011011000",
  58327=>"111111111",
  58328=>"000000000",
  58329=>"011000111",
  58330=>"000000000",
  58331=>"000000000",
  58332=>"000000000",
  58333=>"111110000",
  58334=>"110000000",
  58335=>"000111111",
  58336=>"000100111",
  58337=>"111111111",
  58338=>"111111001",
  58339=>"000000001",
  58340=>"000110100",
  58341=>"000000000",
  58342=>"100000010",
  58343=>"111000000",
  58344=>"000000000",
  58345=>"000001001",
  58346=>"110000000",
  58347=>"000000111",
  58348=>"111111111",
  58349=>"111111111",
  58350=>"111111111",
  58351=>"111111111",
  58352=>"000000000",
  58353=>"011010000",
  58354=>"010110010",
  58355=>"001000001",
  58356=>"011000000",
  58357=>"000000000",
  58358=>"100000000",
  58359=>"111111111",
  58360=>"001000100",
  58361=>"101101111",
  58362=>"111110000",
  58363=>"101111011",
  58364=>"000000111",
  58365=>"111001100",
  58366=>"000000011",
  58367=>"000000000",
  58368=>"111011011",
  58369=>"111111111",
  58370=>"101000000",
  58371=>"000011001",
  58372=>"011011011",
  58373=>"000001101",
  58374=>"110110110",
  58375=>"000000001",
  58376=>"001111001",
  58377=>"110110001",
  58378=>"000000000",
  58379=>"011011011",
  58380=>"100110110",
  58381=>"111010010",
  58382=>"101101000",
  58383=>"000000001",
  58384=>"000000000",
  58385=>"000011111",
  58386=>"010110110",
  58387=>"111111110",
  58388=>"111001001",
  58389=>"010111110",
  58390=>"111101000",
  58391=>"110011011",
  58392=>"100100000",
  58393=>"001011100",
  58394=>"000000000",
  58395=>"110111111",
  58396=>"000100011",
  58397=>"000000110",
  58398=>"001001001",
  58399=>"000000001",
  58400=>"000110111",
  58401=>"001100000",
  58402=>"110110000",
  58403=>"000000000",
  58404=>"011111111",
  58405=>"000000000",
  58406=>"000000001",
  58407=>"000001000",
  58408=>"000001001",
  58409=>"110111111",
  58410=>"100100111",
  58411=>"000000000",
  58412=>"000000111",
  58413=>"011111111",
  58414=>"001000111",
  58415=>"111001000",
  58416=>"001001001",
  58417=>"000000100",
  58418=>"011111001",
  58419=>"110111100",
  58420=>"000000000",
  58421=>"000000000",
  58422=>"000000000",
  58423=>"001001001",
  58424=>"111111011",
  58425=>"000000110",
  58426=>"010110111",
  58427=>"101101111",
  58428=>"111111011",
  58429=>"000000101",
  58430=>"000111000",
  58431=>"101000101",
  58432=>"110111100",
  58433=>"100110110",
  58434=>"111000001",
  58435=>"111111111",
  58436=>"110110011",
  58437=>"001001111",
  58438=>"111010000",
  58439=>"111101101",
  58440=>"111111111",
  58441=>"010110010",
  58442=>"111110000",
  58443=>"001000001",
  58444=>"100000101",
  58445=>"111111101",
  58446=>"101000000",
  58447=>"000100111",
  58448=>"110111110",
  58449=>"011111111",
  58450=>"111011000",
  58451=>"010010000",
  58452=>"001101101",
  58453=>"000010000",
  58454=>"111001010",
  58455=>"011111000",
  58456=>"111111001",
  58457=>"101101101",
  58458=>"111111111",
  58459=>"001001000",
  58460=>"101001001",
  58461=>"101000000",
  58462=>"110110111",
  58463=>"100100000",
  58464=>"000000000",
  58465=>"111000000",
  58466=>"000000111",
  58467=>"100110111",
  58468=>"111110000",
  58469=>"000000000",
  58470=>"111010000",
  58471=>"110110010",
  58472=>"100111111",
  58473=>"001000000",
  58474=>"110110110",
  58475=>"000011111",
  58476=>"001001001",
  58477=>"000000101",
  58478=>"111111111",
  58479=>"000110000",
  58480=>"111000000",
  58481=>"000011011",
  58482=>"000110000",
  58483=>"001001111",
  58484=>"000010010",
  58485=>"001001001",
  58486=>"100000000",
  58487=>"000100101",
  58488=>"000000111",
  58489=>"111101111",
  58490=>"001000000",
  58491=>"000000001",
  58492=>"001001001",
  58493=>"001001000",
  58494=>"010001000",
  58495=>"000101111",
  58496=>"011111111",
  58497=>"001111110",
  58498=>"111101101",
  58499=>"111010000",
  58500=>"000000000",
  58501=>"000000111",
  58502=>"110011001",
  58503=>"111110010",
  58504=>"010000000",
  58505=>"111111111",
  58506=>"111000000",
  58507=>"111111000",
  58508=>"010000000",
  58509=>"111111110",
  58510=>"110110010",
  58511=>"010110010",
  58512=>"101101101",
  58513=>"111111110",
  58514=>"111101001",
  58515=>"111111111",
  58516=>"100000000",
  58517=>"100100111",
  58518=>"110110110",
  58519=>"000000000",
  58520=>"000000101",
  58521=>"111111011",
  58522=>"010110111",
  58523=>"000000000",
  58524=>"110110110",
  58525=>"000001001",
  58526=>"101101111",
  58527=>"000000000",
  58528=>"000111111",
  58529=>"001110110",
  58530=>"111111111",
  58531=>"100000000",
  58532=>"001001001",
  58533=>"111000100",
  58534=>"000000000",
  58535=>"000000000",
  58536=>"100000000",
  58537=>"000000000",
  58538=>"000000000",
  58539=>"001101100",
  58540=>"011010010",
  58541=>"001000000",
  58542=>"111111111",
  58543=>"001001001",
  58544=>"010111111",
  58545=>"100100000",
  58546=>"111111110",
  58547=>"000000000",
  58548=>"111111111",
  58549=>"001000001",
  58550=>"001011000",
  58551=>"000000000",
  58552=>"010011111",
  58553=>"111111110",
  58554=>"000000001",
  58555=>"001000000",
  58556=>"000000100",
  58557=>"001101111",
  58558=>"000100101",
  58559=>"000000000",
  58560=>"000010000",
  58561=>"111111011",
  58562=>"000000100",
  58563=>"110010000",
  58564=>"111111111",
  58565=>"111001000",
  58566=>"000000000",
  58567=>"000011010",
  58568=>"101111000",
  58569=>"111110001",
  58570=>"001000001",
  58571=>"111111101",
  58572=>"010010000",
  58573=>"101100000",
  58574=>"111100111",
  58575=>"111111111",
  58576=>"000000100",
  58577=>"000000001",
  58578=>"101000110",
  58579=>"110111111",
  58580=>"111111000",
  58581=>"111101101",
  58582=>"101100000",
  58583=>"110000001",
  58584=>"000000000",
  58585=>"111111111",
  58586=>"111111111",
  58587=>"000011111",
  58588=>"111001001",
  58589=>"010000000",
  58590=>"001001001",
  58591=>"011000000",
  58592=>"000000001",
  58593=>"000010000",
  58594=>"000100100",
  58595=>"101001111",
  58596=>"111111101",
  58597=>"000000000",
  58598=>"110111010",
  58599=>"111111111",
  58600=>"001001001",
  58601=>"011011111",
  58602=>"011111111",
  58603=>"000000011",
  58604=>"111111111",
  58605=>"000000000",
  58606=>"111000000",
  58607=>"001000000",
  58608=>"011000000",
  58609=>"111111111",
  58610=>"010111110",
  58611=>"001001001",
  58612=>"000000010",
  58613=>"000000000",
  58614=>"100101111",
  58615=>"000010000",
  58616=>"110110010",
  58617=>"010010010",
  58618=>"001001001",
  58619=>"111111111",
  58620=>"110110110",
  58621=>"010000000",
  58622=>"000000000",
  58623=>"100110111",
  58624=>"000001101",
  58625=>"010000000",
  58626=>"111111110",
  58627=>"111100000",
  58628=>"101101111",
  58629=>"000110110",
  58630=>"101000000",
  58631=>"100000101",
  58632=>"000000001",
  58633=>"111101001",
  58634=>"101001111",
  58635=>"111111111",
  58636=>"000010010",
  58637=>"100111111",
  58638=>"111111111",
  58639=>"100110110",
  58640=>"111111111",
  58641=>"001000000",
  58642=>"000001111",
  58643=>"001101111",
  58644=>"010111110",
  58645=>"011011111",
  58646=>"110110110",
  58647=>"111001011",
  58648=>"001001001",
  58649=>"111111001",
  58650=>"000000000",
  58651=>"101001000",
  58652=>"111111111",
  58653=>"010100100",
  58654=>"010010000",
  58655=>"111101100",
  58656=>"100000100",
  58657=>"111110010",
  58658=>"110111111",
  58659=>"000000001",
  58660=>"000000001",
  58661=>"000000101",
  58662=>"111111011",
  58663=>"111111011",
  58664=>"111011001",
  58665=>"111111111",
  58666=>"000001110",
  58667=>"100100111",
  58668=>"100100111",
  58669=>"001001001",
  58670=>"100100000",
  58671=>"100100000",
  58672=>"000000010",
  58673=>"100111000",
  58674=>"001101111",
  58675=>"111111010",
  58676=>"000000101",
  58677=>"000111011",
  58678=>"000010010",
  58679=>"010011011",
  58680=>"110000000",
  58681=>"110110111",
  58682=>"101100100",
  58683=>"000010011",
  58684=>"100100111",
  58685=>"000000001",
  58686=>"111000000",
  58687=>"000000000",
  58688=>"111110010",
  58689=>"111110101",
  58690=>"001001000",
  58691=>"000000000",
  58692=>"000011011",
  58693=>"111111111",
  58694=>"000010111",
  58695=>"110110110",
  58696=>"101111111",
  58697=>"000000000",
  58698=>"000111111",
  58699=>"100110110",
  58700=>"000000000",
  58701=>"011011111",
  58702=>"100111111",
  58703=>"000010000",
  58704=>"000000001",
  58705=>"111000001",
  58706=>"111111111",
  58707=>"000111111",
  58708=>"010011111",
  58709=>"011011011",
  58710=>"001011110",
  58711=>"110000010",
  58712=>"000000000",
  58713=>"000000000",
  58714=>"111111101",
  58715=>"000000000",
  58716=>"110011001",
  58717=>"000000001",
  58718=>"000000000",
  58719=>"111111111",
  58720=>"111101111",
  58721=>"111101101",
  58722=>"100100110",
  58723=>"111110000",
  58724=>"000000000",
  58725=>"001000001",
  58726=>"000111111",
  58727=>"111111111",
  58728=>"001111110",
  58729=>"111110000",
  58730=>"000010000",
  58731=>"110010000",
  58732=>"000011011",
  58733=>"000111001",
  58734=>"000000000",
  58735=>"111100000",
  58736=>"110110010",
  58737=>"101101111",
  58738=>"110110110",
  58739=>"101000000",
  58740=>"000000001",
  58741=>"101001001",
  58742=>"111000001",
  58743=>"111111000",
  58744=>"000010011",
  58745=>"000001111",
  58746=>"001000111",
  58747=>"100000000",
  58748=>"001000011",
  58749=>"001001101",
  58750=>"000001011",
  58751=>"101001101",
  58752=>"000000000",
  58753=>"111111111",
  58754=>"111101110",
  58755=>"000000000",
  58756=>"011011111",
  58757=>"101001000",
  58758=>"000000110",
  58759=>"010011000",
  58760=>"011011000",
  58761=>"011011011",
  58762=>"000010010",
  58763=>"010110110",
  58764=>"111111111",
  58765=>"000100100",
  58766=>"111101111",
  58767=>"000000001",
  58768=>"111111111",
  58769=>"110111111",
  58770=>"100101111",
  58771=>"011011111",
  58772=>"010110110",
  58773=>"110000000",
  58774=>"000000000",
  58775=>"001001101",
  58776=>"000110111",
  58777=>"111110000",
  58778=>"111111000",
  58779=>"110110010",
  58780=>"000000000",
  58781=>"000000001",
  58782=>"111000000",
  58783=>"000001000",
  58784=>"101000100",
  58785=>"100100000",
  58786=>"111011001",
  58787=>"111111111",
  58788=>"001001111",
  58789=>"110000000",
  58790=>"000000000",
  58791=>"001000100",
  58792=>"111111011",
  58793=>"111111101",
  58794=>"110111010",
  58795=>"001000000",
  58796=>"001011111",
  58797=>"000000101",
  58798=>"000000111",
  58799=>"000000000",
  58800=>"000000111",
  58801=>"101111111",
  58802=>"110111110",
  58803=>"010111111",
  58804=>"000000000",
  58805=>"111111111",
  58806=>"100111100",
  58807=>"111110000",
  58808=>"000000000",
  58809=>"111111111",
  58810=>"000000111",
  58811=>"000000000",
  58812=>"000000001",
  58813=>"001000001",
  58814=>"111111100",
  58815=>"100100001",
  58816=>"111111011",
  58817=>"000000000",
  58818=>"000111111",
  58819=>"010010000",
  58820=>"111111110",
  58821=>"001011001",
  58822=>"111110110",
  58823=>"000000001",
  58824=>"110111111",
  58825=>"000000110",
  58826=>"111000000",
  58827=>"001101111",
  58828=>"011001000",
  58829=>"000010111",
  58830=>"100000000",
  58831=>"000000000",
  58832=>"100000101",
  58833=>"001000001",
  58834=>"000110110",
  58835=>"111111111",
  58836=>"000100111",
  58837=>"111111111",
  58838=>"001000000",
  58839=>"011111011",
  58840=>"000000000",
  58841=>"100111111",
  58842=>"111011011",
  58843=>"111111010",
  58844=>"000000000",
  58845=>"110000000",
  58846=>"001000000",
  58847=>"000110000",
  58848=>"001001000",
  58849=>"111010000",
  58850=>"000000011",
  58851=>"000000000",
  58852=>"111111111",
  58853=>"000000000",
  58854=>"000100000",
  58855=>"000000000",
  58856=>"100011011",
  58857=>"111111011",
  58858=>"000000000",
  58859=>"011101001",
  58860=>"010010010",
  58861=>"000100100",
  58862=>"101101101",
  58863=>"001000110",
  58864=>"111001001",
  58865=>"000011111",
  58866=>"011111111",
  58867=>"000100000",
  58868=>"000000000",
  58869=>"000000000",
  58870=>"000000000",
  58871=>"111111111",
  58872=>"000000000",
  58873=>"011011011",
  58874=>"110110110",
  58875=>"100100100",
  58876=>"110111111",
  58877=>"000110111",
  58878=>"000000001",
  58879=>"001000011",
  58880=>"100100100",
  58881=>"000000000",
  58882=>"111111000",
  58883=>"000111111",
  58884=>"111111111",
  58885=>"000000000",
  58886=>"110111110",
  58887=>"111111001",
  58888=>"011000000",
  58889=>"111111100",
  58890=>"011011011",
  58891=>"000100111",
  58892=>"000000000",
  58893=>"000111111",
  58894=>"100000101",
  58895=>"101111111",
  58896=>"111100010",
  58897=>"111111000",
  58898=>"111100000",
  58899=>"111101000",
  58900=>"000000000",
  58901=>"011011001",
  58902=>"000111111",
  58903=>"001111111",
  58904=>"000111111",
  58905=>"111111111",
  58906=>"111111110",
  58907=>"000100000",
  58908=>"111110000",
  58909=>"111011000",
  58910=>"000000111",
  58911=>"000111111",
  58912=>"000111110",
  58913=>"000111111",
  58914=>"111000110",
  58915=>"111111111",
  58916=>"000010110",
  58917=>"100111111",
  58918=>"000000000",
  58919=>"000000111",
  58920=>"100100000",
  58921=>"011000000",
  58922=>"011000000",
  58923=>"011000011",
  58924=>"111111111",
  58925=>"100000000",
  58926=>"011000110",
  58927=>"000000111",
  58928=>"100000000",
  58929=>"000000000",
  58930=>"001111111",
  58931=>"100111001",
  58932=>"000000111",
  58933=>"000110110",
  58934=>"000101111",
  58935=>"000001111",
  58936=>"000000000",
  58937=>"111011111",
  58938=>"111000000",
  58939=>"011000000",
  58940=>"111111111",
  58941=>"111111011",
  58942=>"011001000",
  58943=>"111111111",
  58944=>"001101111",
  58945=>"000000010",
  58946=>"000111111",
  58947=>"111000111",
  58948=>"000000101",
  58949=>"000001111",
  58950=>"000110101",
  58951=>"110111000",
  58952=>"001001011",
  58953=>"000000000",
  58954=>"111000011",
  58955=>"100000000",
  58956=>"000011011",
  58957=>"000000000",
  58958=>"000100110",
  58959=>"100100000",
  58960=>"110110010",
  58961=>"111111000",
  58962=>"111101111",
  58963=>"000100101",
  58964=>"111111110",
  58965=>"111001000",
  58966=>"101000111",
  58967=>"001111011",
  58968=>"000000010",
  58969=>"111110100",
  58970=>"111111000",
  58971=>"000100110",
  58972=>"000000111",
  58973=>"000000101",
  58974=>"000000000",
  58975=>"000000111",
  58976=>"111110110",
  58977=>"000000000",
  58978=>"111000100",
  58979=>"001011111",
  58980=>"000000000",
  58981=>"000111111",
  58982=>"111000110",
  58983=>"000000000",
  58984=>"000000111",
  58985=>"000010111",
  58986=>"111111101",
  58987=>"111111001",
  58988=>"101000001",
  58989=>"000000000",
  58990=>"000111111",
  58991=>"001111101",
  58992=>"000000111",
  58993=>"100111111",
  58994=>"000000000",
  58995=>"011011000",
  58996=>"111001000",
  58997=>"111111000",
  58998=>"111000000",
  58999=>"000011001",
  59000=>"111101000",
  59001=>"001000000",
  59002=>"000000000",
  59003=>"111011000",
  59004=>"000110111",
  59005=>"000100100",
  59006=>"000010000",
  59007=>"000000111",
  59008=>"000101111",
  59009=>"110110110",
  59010=>"110111000",
  59011=>"110110001",
  59012=>"111001000",
  59013=>"011011011",
  59014=>"000001000",
  59015=>"000000000",
  59016=>"111111000",
  59017=>"101101111",
  59018=>"000000010",
  59019=>"111001000",
  59020=>"111111000",
  59021=>"100110000",
  59022=>"111111001",
  59023=>"000000000",
  59024=>"111111001",
  59025=>"111011000",
  59026=>"010111111",
  59027=>"010111111",
  59028=>"000000110",
  59029=>"000000011",
  59030=>"000111001",
  59031=>"001101000",
  59032=>"000000001",
  59033=>"111111111",
  59034=>"000000000",
  59035=>"000111111",
  59036=>"100101000",
  59037=>"111000000",
  59038=>"000111111",
  59039=>"000010000",
  59040=>"111111000",
  59041=>"000000001",
  59042=>"111000000",
  59043=>"000000000",
  59044=>"000000000",
  59045=>"110000001",
  59046=>"000011011",
  59047=>"011111111",
  59048=>"000000000",
  59049=>"110111100",
  59050=>"000111111",
  59051=>"111111111",
  59052=>"001001111",
  59053=>"000110111",
  59054=>"111111001",
  59055=>"000111111",
  59056=>"000000111",
  59057=>"111000100",
  59058=>"111011010",
  59059=>"011000001",
  59060=>"000000000",
  59061=>"000011011",
  59062=>"000000101",
  59063=>"101111000",
  59064=>"110111111",
  59065=>"111010000",
  59066=>"000000111",
  59067=>"100000000",
  59068=>"110000000",
  59069=>"111111001",
  59070=>"111000111",
  59071=>"111111111",
  59072=>"001001011",
  59073=>"000001011",
  59074=>"000000000",
  59075=>"000000010",
  59076=>"111000111",
  59077=>"000000000",
  59078=>"110011111",
  59079=>"100000000",
  59080=>"111111100",
  59081=>"000000000",
  59082=>"000011011",
  59083=>"100000000",
  59084=>"111001000",
  59085=>"011111111",
  59086=>"000000000",
  59087=>"100000000",
  59088=>"011111000",
  59089=>"000001111",
  59090=>"111000000",
  59091=>"000000000",
  59092=>"111100111",
  59093=>"000010010",
  59094=>"111111000",
  59095=>"000000001",
  59096=>"000000000",
  59097=>"101000000",
  59098=>"111001000",
  59099=>"000000111",
  59100=>"001111111",
  59101=>"111111101",
  59102=>"111111011",
  59103=>"000000000",
  59104=>"111111111",
  59105=>"000111011",
  59106=>"000000000",
  59107=>"111000000",
  59108=>"111111000",
  59109=>"000110111",
  59110=>"000110111",
  59111=>"001000110",
  59112=>"000000111",
  59113=>"011011101",
  59114=>"000000000",
  59115=>"000101111",
  59116=>"000100111",
  59117=>"011001111",
  59118=>"010110111",
  59119=>"111100111",
  59120=>"100001000",
  59121=>"000000000",
  59122=>"111000000",
  59123=>"000100011",
  59124=>"000000000",
  59125=>"000100111",
  59126=>"111000000",
  59127=>"111000000",
  59128=>"000111111",
  59129=>"111111000",
  59130=>"000000011",
  59131=>"111110010",
  59132=>"000111111",
  59133=>"111111111",
  59134=>"000000000",
  59135=>"001011001",
  59136=>"111111011",
  59137=>"111111111",
  59138=>"111000000",
  59139=>"111111111",
  59140=>"000000000",
  59141=>"000000111",
  59142=>"000000000",
  59143=>"001010000",
  59144=>"111000000",
  59145=>"000000100",
  59146=>"000100111",
  59147=>"000000000",
  59148=>"111110001",
  59149=>"111000000",
  59150=>"000110111",
  59151=>"111100111",
  59152=>"000000000",
  59153=>"000101111",
  59154=>"111001000",
  59155=>"000000000",
  59156=>"111111011",
  59157=>"111110111",
  59158=>"011011110",
  59159=>"000000000",
  59160=>"111111000",
  59161=>"000111111",
  59162=>"000111010",
  59163=>"000010010",
  59164=>"000000111",
  59165=>"110001000",
  59166=>"000000111",
  59167=>"000001101",
  59168=>"111011111",
  59169=>"000011000",
  59170=>"111111000",
  59171=>"110000001",
  59172=>"000000111",
  59173=>"000110000",
  59174=>"110111111",
  59175=>"111111011",
  59176=>"000111111",
  59177=>"101000000",
  59178=>"111111000",
  59179=>"111000000",
  59180=>"110111111",
  59181=>"111111000",
  59182=>"000000000",
  59183=>"000000110",
  59184=>"111001011",
  59185=>"111111010",
  59186=>"111111000",
  59187=>"011001001",
  59188=>"111001000",
  59189=>"000000100",
  59190=>"110000000",
  59191=>"010100111",
  59192=>"000111010",
  59193=>"111001000",
  59194=>"000111111",
  59195=>"000000010",
  59196=>"111000000",
  59197=>"111000101",
  59198=>"000110111",
  59199=>"111110000",
  59200=>"111111000",
  59201=>"111111000",
  59202=>"000000000",
  59203=>"000100101",
  59204=>"111111110",
  59205=>"100101111",
  59206=>"110110110",
  59207=>"000000011",
  59208=>"000000000",
  59209=>"000000000",
  59210=>"101100111",
  59211=>"100000100",
  59212=>"000111011",
  59213=>"000011001",
  59214=>"000000001",
  59215=>"110000000",
  59216=>"000000111",
  59217=>"100000011",
  59218=>"000101101",
  59219=>"001001000",
  59220=>"111001111",
  59221=>"111001001",
  59222=>"000000000",
  59223=>"001001011",
  59224=>"111000000",
  59225=>"111111111",
  59226=>"100000100",
  59227=>"100111010",
  59228=>"011001000",
  59229=>"000000000",
  59230=>"111111000",
  59231=>"001001001",
  59232=>"110000000",
  59233=>"111111111",
  59234=>"000111110",
  59235=>"000111111",
  59236=>"111011011",
  59237=>"111111110",
  59238=>"000111111",
  59239=>"011000001",
  59240=>"000000101",
  59241=>"110111111",
  59242=>"000011111",
  59243=>"111111001",
  59244=>"001000000",
  59245=>"000010000",
  59246=>"111111110",
  59247=>"000011111",
  59248=>"000000000",
  59249=>"100011111",
  59250=>"110110100",
  59251=>"000000001",
  59252=>"111111000",
  59253=>"011111100",
  59254=>"111000000",
  59255=>"000111001",
  59256=>"000111111",
  59257=>"001111111",
  59258=>"000100000",
  59259=>"000111000",
  59260=>"110000000",
  59261=>"000000100",
  59262=>"000011111",
  59263=>"000000000",
  59264=>"101100000",
  59265=>"000000111",
  59266=>"100111000",
  59267=>"100110000",
  59268=>"111111111",
  59269=>"000000111",
  59270=>"110110000",
  59271=>"011111111",
  59272=>"000000100",
  59273=>"111111111",
  59274=>"111100110",
  59275=>"111111000",
  59276=>"101100100",
  59277=>"011011111",
  59278=>"110110000",
  59279=>"010001111",
  59280=>"000000000",
  59281=>"111000000",
  59282=>"111000000",
  59283=>"111011001",
  59284=>"101000011",
  59285=>"000000010",
  59286=>"111111000",
  59287=>"111000000",
  59288=>"000000000",
  59289=>"000110111",
  59290=>"110111111",
  59291=>"011000000",
  59292=>"111111111",
  59293=>"000011000",
  59294=>"111111111",
  59295=>"000000011",
  59296=>"111111011",
  59297=>"001111000",
  59298=>"001011011",
  59299=>"000111111",
  59300=>"101111101",
  59301=>"110111000",
  59302=>"111111010",
  59303=>"000000011",
  59304=>"000000001",
  59305=>"000000000",
  59306=>"111000000",
  59307=>"000000111",
  59308=>"100000000",
  59309=>"111100111",
  59310=>"000000000",
  59311=>"111011000",
  59312=>"000000100",
  59313=>"000110111",
  59314=>"000100000",
  59315=>"000000111",
  59316=>"100111010",
  59317=>"000001111",
  59318=>"111011011",
  59319=>"111111111",
  59320=>"111000000",
  59321=>"111001000",
  59322=>"000000100",
  59323=>"000111100",
  59324=>"001000111",
  59325=>"111000000",
  59326=>"000000000",
  59327=>"000101111",
  59328=>"000000111",
  59329=>"000000000",
  59330=>"111111000",
  59331=>"111111101",
  59332=>"111111100",
  59333=>"111001101",
  59334=>"000000011",
  59335=>"011011111",
  59336=>"000000000",
  59337=>"011011000",
  59338=>"000111111",
  59339=>"111111000",
  59340=>"111111010",
  59341=>"000111000",
  59342=>"000000111",
  59343=>"000000010",
  59344=>"001001111",
  59345=>"000111111",
  59346=>"111110111",
  59347=>"111111000",
  59348=>"111111011",
  59349=>"111110000",
  59350=>"011001111",
  59351=>"000011111",
  59352=>"000100110",
  59353=>"111111011",
  59354=>"000000011",
  59355=>"101111111",
  59356=>"000001011",
  59357=>"000100011",
  59358=>"100100111",
  59359=>"000000001",
  59360=>"000100100",
  59361=>"100110110",
  59362=>"001000111",
  59363=>"111111111",
  59364=>"000000011",
  59365=>"111001000",
  59366=>"000000110",
  59367=>"000111111",
  59368=>"101111100",
  59369=>"000000110",
  59370=>"000000000",
  59371=>"000100111",
  59372=>"100000001",
  59373=>"110011011",
  59374=>"111111101",
  59375=>"000000001",
  59376=>"000000000",
  59377=>"111111011",
  59378=>"000000111",
  59379=>"000111111",
  59380=>"111000000",
  59381=>"100001001",
  59382=>"000000000",
  59383=>"010011001",
  59384=>"000001111",
  59385=>"000000111",
  59386=>"000000000",
  59387=>"111111111",
  59388=>"000000111",
  59389=>"000000001",
  59390=>"000000000",
  59391=>"000111111",
  59392=>"110111111",
  59393=>"000111111",
  59394=>"000000001",
  59395=>"000000000",
  59396=>"000000001",
  59397=>"001011010",
  59398=>"111111111",
  59399=>"111101111",
  59400=>"111111000",
  59401=>"000000000",
  59402=>"000000000",
  59403=>"111111111",
  59404=>"000110001",
  59405=>"000000000",
  59406=>"000000000",
  59407=>"000000000",
  59408=>"000000000",
  59409=>"011111011",
  59410=>"000000101",
  59411=>"000000100",
  59412=>"111000100",
  59413=>"111111111",
  59414=>"000010010",
  59415=>"110111011",
  59416=>"000000000",
  59417=>"000100000",
  59418=>"101011111",
  59419=>"100100100",
  59420=>"111001001",
  59421=>"010111100",
  59422=>"001001101",
  59423=>"000100110",
  59424=>"000000000",
  59425=>"110110000",
  59426=>"111100110",
  59427=>"100100001",
  59428=>"111111001",
  59429=>"111111011",
  59430=>"110110110",
  59431=>"111111111",
  59432=>"000100111",
  59433=>"101101111",
  59434=>"111111011",
  59435=>"111111111",
  59436=>"111101000",
  59437=>"000000000",
  59438=>"001011000",
  59439=>"000000111",
  59440=>"101001001",
  59441=>"000000000",
  59442=>"000001001",
  59443=>"000000000",
  59444=>"000000000",
  59445=>"000001001",
  59446=>"101111111",
  59447=>"111111000",
  59448=>"001000000",
  59449=>"111001111",
  59450=>"000000001",
  59451=>"000000000",
  59452=>"111100111",
  59453=>"110000110",
  59454=>"111111110",
  59455=>"111111111",
  59456=>"000110111",
  59457=>"000000001",
  59458=>"010111010",
  59459=>"000001010",
  59460=>"000010011",
  59461=>"111111111",
  59462=>"111111111",
  59463=>"111111111",
  59464=>"000101111",
  59465=>"000000000",
  59466=>"000001011",
  59467=>"010000000",
  59468=>"000000000",
  59469=>"011111100",
  59470=>"111011011",
  59471=>"111111100",
  59472=>"111111110",
  59473=>"111111111",
  59474=>"111111110",
  59475=>"000001001",
  59476=>"000000000",
  59477=>"111010000",
  59478=>"000000000",
  59479=>"000000100",
  59480=>"000000011",
  59481=>"000000111",
  59482=>"000000100",
  59483=>"110110110",
  59484=>"000100111",
  59485=>"000101101",
  59486=>"000000000",
  59487=>"100000011",
  59488=>"000000000",
  59489=>"001000000",
  59490=>"110111111",
  59491=>"111000000",
  59492=>"000111110",
  59493=>"011011111",
  59494=>"111111000",
  59495=>"000011011",
  59496=>"000001111",
  59497=>"011000000",
  59498=>"111111111",
  59499=>"000000001",
  59500=>"111111111",
  59501=>"100100111",
  59502=>"110110000",
  59503=>"111000000",
  59504=>"000000000",
  59505=>"000000000",
  59506=>"011011000",
  59507=>"111000011",
  59508=>"000000000",
  59509=>"100000111",
  59510=>"011111000",
  59511=>"000000000",
  59512=>"111000000",
  59513=>"011111111",
  59514=>"000000000",
  59515=>"000000011",
  59516=>"100110110",
  59517=>"111111111",
  59518=>"111110001",
  59519=>"000010000",
  59520=>"111100000",
  59521=>"111111101",
  59522=>"110000000",
  59523=>"100110111",
  59524=>"110100100",
  59525=>"000000000",
  59526=>"111111011",
  59527=>"010111000",
  59528=>"000000111",
  59529=>"000001100",
  59530=>"000000111",
  59531=>"001000000",
  59532=>"000000110",
  59533=>"000000000",
  59534=>"100000000",
  59535=>"000000000",
  59536=>"111111111",
  59537=>"111111111",
  59538=>"000000000",
  59539=>"111111110",
  59540=>"100100110",
  59541=>"000000000",
  59542=>"111000000",
  59543=>"000011111",
  59544=>"000000000",
  59545=>"111111110",
  59546=>"000000100",
  59547=>"000000010",
  59548=>"111111111",
  59549=>"000011000",
  59550=>"111111111",
  59551=>"000000000",
  59552=>"111101101",
  59553=>"100100100",
  59554=>"100000000",
  59555=>"101000001",
  59556=>"000000000",
  59557=>"000000100",
  59558=>"101101111",
  59559=>"111001001",
  59560=>"111111111",
  59561=>"000000000",
  59562=>"111110000",
  59563=>"000000000",
  59564=>"111011111",
  59565=>"101101111",
  59566=>"111111111",
  59567=>"011100100",
  59568=>"001111111",
  59569=>"100000000",
  59570=>"011011010",
  59571=>"000000111",
  59572=>"111001111",
  59573=>"111111011",
  59574=>"101111100",
  59575=>"000000000",
  59576=>"100100000",
  59577=>"110000000",
  59578=>"000000000",
  59579=>"001001001",
  59580=>"011001011",
  59581=>"111010000",
  59582=>"100000000",
  59583=>"011111111",
  59584=>"000000100",
  59585=>"000000000",
  59586=>"001111111",
  59587=>"000000000",
  59588=>"000000000",
  59589=>"011000000",
  59590=>"000000010",
  59591=>"000001000",
  59592=>"111111111",
  59593=>"111111101",
  59594=>"000000001",
  59595=>"000111110",
  59596=>"001100000",
  59597=>"111111110",
  59598=>"000000001",
  59599=>"000000000",
  59600=>"001000000",
  59601=>"011111110",
  59602=>"000011011",
  59603=>"000000000",
  59604=>"110110000",
  59605=>"111111111",
  59606=>"000100000",
  59607=>"001111111",
  59608=>"001001111",
  59609=>"001111111",
  59610=>"000000000",
  59611=>"111111111",
  59612=>"110110111",
  59613=>"111111001",
  59614=>"001111101",
  59615=>"111111110",
  59616=>"111111011",
  59617=>"000010000",
  59618=>"000000011",
  59619=>"101100100",
  59620=>"000000000",
  59621=>"111111011",
  59622=>"000000111",
  59623=>"000000000",
  59624=>"111111111",
  59625=>"000001111",
  59626=>"111000000",
  59627=>"000100111",
  59628=>"010000111",
  59629=>"000010011",
  59630=>"111000110",
  59631=>"000011111",
  59632=>"110000000",
  59633=>"000000000",
  59634=>"111101100",
  59635=>"011011111",
  59636=>"000000000",
  59637=>"100000110",
  59638=>"111100000",
  59639=>"000000000",
  59640=>"000000000",
  59641=>"111000001",
  59642=>"100111111",
  59643=>"000001011",
  59644=>"110110110",
  59645=>"000001011",
  59646=>"111110100",
  59647=>"100000000",
  59648=>"111111111",
  59649=>"000000100",
  59650=>"000000000",
  59651=>"000001000",
  59652=>"100100100",
  59653=>"111111000",
  59654=>"000100101",
  59655=>"100110011",
  59656=>"101001001",
  59657=>"110011000",
  59658=>"000001011",
  59659=>"111111001",
  59660=>"000000000",
  59661=>"000110110",
  59662=>"000000000",
  59663=>"110010011",
  59664=>"001000100",
  59665=>"111111011",
  59666=>"111111111",
  59667=>"011111000",
  59668=>"000001011",
  59669=>"000000111",
  59670=>"001001001",
  59671=>"000000000",
  59672=>"000111111",
  59673=>"111111111",
  59674=>"111111111",
  59675=>"110111111",
  59676=>"111111100",
  59677=>"111111111",
  59678=>"111111111",
  59679=>"000000000",
  59680=>"010010000",
  59681=>"000111001",
  59682=>"011011111",
  59683=>"000100101",
  59684=>"001011011",
  59685=>"100100000",
  59686=>"001011100",
  59687=>"000000100",
  59688=>"000010000",
  59689=>"111111111",
  59690=>"000111011",
  59691=>"000011111",
  59692=>"001011000",
  59693=>"101111111",
  59694=>"001111111",
  59695=>"000000100",
  59696=>"011011000",
  59697=>"111111111",
  59698=>"000000100",
  59699=>"111111011",
  59700=>"000000000",
  59701=>"000110111",
  59702=>"111111101",
  59703=>"000000001",
  59704=>"000000000",
  59705=>"000000000",
  59706=>"000000000",
  59707=>"000100100",
  59708=>"001100110",
  59709=>"111111111",
  59710=>"011010000",
  59711=>"000111111",
  59712=>"000000000",
  59713=>"100000000",
  59714=>"111111111",
  59715=>"000111111",
  59716=>"111111100",
  59717=>"100111111",
  59718=>"111111111",
  59719=>"000000011",
  59720=>"100000010",
  59721=>"111111111",
  59722=>"111111111",
  59723=>"110110111",
  59724=>"000001001",
  59725=>"011001001",
  59726=>"100110110",
  59727=>"001001111",
  59728=>"001001100",
  59729=>"011000000",
  59730=>"000000000",
  59731=>"111111111",
  59732=>"000000011",
  59733=>"011000000",
  59734=>"111111111",
  59735=>"000001000",
  59736=>"110111011",
  59737=>"111111111",
  59738=>"001101011",
  59739=>"000100111",
  59740=>"111000110",
  59741=>"000011010",
  59742=>"000001111",
  59743=>"111011001",
  59744=>"101111000",
  59745=>"111111001",
  59746=>"000000100",
  59747=>"000000111",
  59748=>"100000000",
  59749=>"000000000",
  59750=>"000001001",
  59751=>"000001001",
  59752=>"111111111",
  59753=>"011011111",
  59754=>"111111010",
  59755=>"011000000",
  59756=>"000001011",
  59757=>"000010111",
  59758=>"000000000",
  59759=>"000110000",
  59760=>"001001111",
  59761=>"111001001",
  59762=>"000100111",
  59763=>"100110111",
  59764=>"111111111",
  59765=>"100100110",
  59766=>"000000000",
  59767=>"000000000",
  59768=>"000000000",
  59769=>"001000000",
  59770=>"000000000",
  59771=>"111111111",
  59772=>"100000000",
  59773=>"000000100",
  59774=>"111111001",
  59775=>"000000000",
  59776=>"110110110",
  59777=>"110100100",
  59778=>"111111011",
  59779=>"011001000",
  59780=>"001000000",
  59781=>"000110111",
  59782=>"111111111",
  59783=>"001011111",
  59784=>"000000000",
  59785=>"001001011",
  59786=>"010011111",
  59787=>"000110111",
  59788=>"000000101",
  59789=>"000000000",
  59790=>"000000000",
  59791=>"000000000",
  59792=>"100100000",
  59793=>"111100000",
  59794=>"111011010",
  59795=>"011011011",
  59796=>"111011011",
  59797=>"000000000",
  59798=>"100100000",
  59799=>"010010111",
  59800=>"111101101",
  59801=>"100111010",
  59802=>"000000000",
  59803=>"101101111",
  59804=>"111111111",
  59805=>"110000000",
  59806=>"000000100",
  59807=>"111111101",
  59808=>"011001000",
  59809=>"100100111",
  59810=>"000000110",
  59811=>"000000000",
  59812=>"110110111",
  59813=>"000000000",
  59814=>"000000000",
  59815=>"111011000",
  59816=>"000000000",
  59817=>"010111001",
  59818=>"111111111",
  59819=>"000000000",
  59820=>"100100100",
  59821=>"100000100",
  59822=>"000000001",
  59823=>"111111111",
  59824=>"000111111",
  59825=>"000000010",
  59826=>"011000000",
  59827=>"000011111",
  59828=>"111111111",
  59829=>"111111111",
  59830=>"111100010",
  59831=>"111111000",
  59832=>"000001011",
  59833=>"001011000",
  59834=>"111100111",
  59835=>"000000001",
  59836=>"011000000",
  59837=>"000000000",
  59838=>"100100100",
  59839=>"100101101",
  59840=>"110110001",
  59841=>"111111111",
  59842=>"010010111",
  59843=>"111111111",
  59844=>"000000000",
  59845=>"001001011",
  59846=>"000111111",
  59847=>"000100101",
  59848=>"001001001",
  59849=>"000100111",
  59850=>"000000000",
  59851=>"000000000",
  59852=>"000000000",
  59853=>"100100110",
  59854=>"000001000",
  59855=>"111011011",
  59856=>"000111111",
  59857=>"000000000",
  59858=>"011111111",
  59859=>"111000111",
  59860=>"000111101",
  59861=>"010110000",
  59862=>"000001001",
  59863=>"000111111",
  59864=>"110111111",
  59865=>"000000100",
  59866=>"000000001",
  59867=>"001000000",
  59868=>"000111111",
  59869=>"110001011",
  59870=>"111111111",
  59871=>"111111111",
  59872=>"000000000",
  59873=>"000000110",
  59874=>"000011101",
  59875=>"000000011",
  59876=>"000000000",
  59877=>"111100000",
  59878=>"100000000",
  59879=>"011010011",
  59880=>"011011001",
  59881=>"000000000",
  59882=>"111011110",
  59883=>"010111110",
  59884=>"011111010",
  59885=>"000100100",
  59886=>"000000000",
  59887=>"000000100",
  59888=>"001001000",
  59889=>"000000000",
  59890=>"111111111",
  59891=>"000000000",
  59892=>"000001111",
  59893=>"000001001",
  59894=>"111111111",
  59895=>"001001011",
  59896=>"000111111",
  59897=>"000000100",
  59898=>"000000001",
  59899=>"111111110",
  59900=>"111111000",
  59901=>"111111111",
  59902=>"100111111",
  59903=>"000100110",
  59904=>"000000000",
  59905=>"111111111",
  59906=>"101000000",
  59907=>"111111111",
  59908=>"111111111",
  59909=>"111111110",
  59910=>"000000000",
  59911=>"000000000",
  59912=>"111111011",
  59913=>"111000000",
  59914=>"111111111",
  59915=>"000000001",
  59916=>"000001001",
  59917=>"110110110",
  59918=>"000000100",
  59919=>"000000000",
  59920=>"110001000",
  59921=>"000010000",
  59922=>"000000000",
  59923=>"000000000",
  59924=>"111111111",
  59925=>"000000011",
  59926=>"000000000",
  59927=>"101100110",
  59928=>"111110111",
  59929=>"100000001",
  59930=>"111001000",
  59931=>"111100101",
  59932=>"111000111",
  59933=>"111111111",
  59934=>"111111010",
  59935=>"000011111",
  59936=>"000000000",
  59937=>"111111111",
  59938=>"000001000",
  59939=>"111111111",
  59940=>"011111011",
  59941=>"110000000",
  59942=>"111001001",
  59943=>"100111111",
  59944=>"001000000",
  59945=>"111111111",
  59946=>"110100111",
  59947=>"100000000",
  59948=>"111111111",
  59949=>"000000110",
  59950=>"100110111",
  59951=>"111111111",
  59952=>"000000000",
  59953=>"000001000",
  59954=>"000000100",
  59955=>"000000111",
  59956=>"111111100",
  59957=>"000000000",
  59958=>"000001001",
  59959=>"101101011",
  59960=>"000111111",
  59961=>"000111111",
  59962=>"111111111",
  59963=>"000000010",
  59964=>"101000101",
  59965=>"111111111",
  59966=>"011011110",
  59967=>"110000111",
  59968=>"100100100",
  59969=>"000100010",
  59970=>"111111100",
  59971=>"111111111",
  59972=>"111001001",
  59973=>"001001011",
  59974=>"000000000",
  59975=>"001000000",
  59976=>"111111111",
  59977=>"000000000",
  59978=>"000000000",
  59979=>"000001111",
  59980=>"111011010",
  59981=>"001001100",
  59982=>"111111111",
  59983=>"000000000",
  59984=>"101011111",
  59985=>"111111111",
  59986=>"000000000",
  59987=>"101101100",
  59988=>"000000000",
  59989=>"111111001",
  59990=>"111111111",
  59991=>"111101101",
  59992=>"000000000",
  59993=>"000000111",
  59994=>"001001111",
  59995=>"001011011",
  59996=>"000000000",
  59997=>"111111111",
  59998=>"111111110",
  59999=>"111111011",
  60000=>"000000000",
  60001=>"111110111",
  60002=>"000001011",
  60003=>"001100000",
  60004=>"111111110",
  60005=>"011000100",
  60006=>"000000000",
  60007=>"000011111",
  60008=>"111111110",
  60009=>"110111111",
  60010=>"100001000",
  60011=>"000111011",
  60012=>"101101100",
  60013=>"000000100",
  60014=>"111111111",
  60015=>"111011000",
  60016=>"111111100",
  60017=>"000110000",
  60018=>"001011000",
  60019=>"111000000",
  60020=>"000000000",
  60021=>"101011111",
  60022=>"000000000",
  60023=>"111111111",
  60024=>"000111111",
  60025=>"100100000",
  60026=>"000000000",
  60027=>"000000000",
  60028=>"110110110",
  60029=>"100101111",
  60030=>"010010000",
  60031=>"001001000",
  60032=>"100100000",
  60033=>"111001101",
  60034=>"111111111",
  60035=>"111111111",
  60036=>"000001111",
  60037=>"111111101",
  60038=>"111111000",
  60039=>"000000000",
  60040=>"111110000",
  60041=>"111111111",
  60042=>"111000000",
  60043=>"100100000",
  60044=>"111111111",
  60045=>"111111111",
  60046=>"011000000",
  60047=>"000000010",
  60048=>"111111111",
  60049=>"111111011",
  60050=>"111111110",
  60051=>"111111110",
  60052=>"000000000",
  60053=>"111111111",
  60054=>"000011011",
  60055=>"000000000",
  60056=>"100000100",
  60057=>"000000000",
  60058=>"111101000",
  60059=>"011011000",
  60060=>"100010000",
  60061=>"010111111",
  60062=>"000000111",
  60063=>"000000000",
  60064=>"000111000",
  60065=>"000000111",
  60066=>"000000000",
  60067=>"110111111",
  60068=>"000000000",
  60069=>"110100100",
  60070=>"000000000",
  60071=>"011011111",
  60072=>"000110111",
  60073=>"000000000",
  60074=>"111000000",
  60075=>"000000100",
  60076=>"110111101",
  60077=>"010001011",
  60078=>"100000011",
  60079=>"111110100",
  60080=>"111110110",
  60081=>"001011110",
  60082=>"000101000",
  60083=>"111111111",
  60084=>"000001101",
  60085=>"111111100",
  60086=>"001000000",
  60087=>"111111111",
  60088=>"101001011",
  60089=>"001001011",
  60090=>"000000000",
  60091=>"111011000",
  60092=>"111111111",
  60093=>"111111111",
  60094=>"000000000",
  60095=>"001000000",
  60096=>"000000000",
  60097=>"000000000",
  60098=>"111011011",
  60099=>"000010010",
  60100=>"111111111",
  60101=>"000000000",
  60102=>"000110111",
  60103=>"001001011",
  60104=>"110000111",
  60105=>"000111111",
  60106=>"110000001",
  60107=>"111111111",
  60108=>"000000000",
  60109=>"001111000",
  60110=>"111111111",
  60111=>"000111111",
  60112=>"111111101",
  60113=>"110100000",
  60114=>"000000100",
  60115=>"111111111",
  60116=>"000000000",
  60117=>"000010000",
  60118=>"000000000",
  60119=>"111111111",
  60120=>"000000000",
  60121=>"111111111",
  60122=>"001000000",
  60123=>"011000000",
  60124=>"000000111",
  60125=>"000000000",
  60126=>"000001011",
  60127=>"111111111",
  60128=>"000000000",
  60129=>"000010111",
  60130=>"000111110",
  60131=>"000000111",
  60132=>"000000000",
  60133=>"110100110",
  60134=>"111111111",
  60135=>"111111111",
  60136=>"111111110",
  60137=>"100110110",
  60138=>"111111010",
  60139=>"000000000",
  60140=>"000111111",
  60141=>"000000000",
  60142=>"000111111",
  60143=>"111110000",
  60144=>"111111111",
  60145=>"101001001",
  60146=>"000111000",
  60147=>"000000000",
  60148=>"000000000",
  60149=>"111111000",
  60150=>"000000000",
  60151=>"111111110",
  60152=>"001001001",
  60153=>"000000000",
  60154=>"100100000",
  60155=>"011000100",
  60156=>"000000001",
  60157=>"111001011",
  60158=>"000001111",
  60159=>"111111011",
  60160=>"000000000",
  60161=>"001011011",
  60162=>"111111111",
  60163=>"000011111",
  60164=>"000011001",
  60165=>"000000000",
  60166=>"000000000",
  60167=>"111111111",
  60168=>"000000000",
  60169=>"100000000",
  60170=>"111100111",
  60171=>"110000000",
  60172=>"100100000",
  60173=>"110100111",
  60174=>"000000000",
  60175=>"001001000",
  60176=>"000000011",
  60177=>"000000110",
  60178=>"000000000",
  60179=>"000001101",
  60180=>"000111111",
  60181=>"111111000",
  60182=>"100111111",
  60183=>"100100000",
  60184=>"000000001",
  60185=>"001001001",
  60186=>"000000000",
  60187=>"111111111",
  60188=>"111111111",
  60189=>"000010111",
  60190=>"000000100",
  60191=>"100110111",
  60192=>"111111111",
  60193=>"011001001",
  60194=>"100000000",
  60195=>"110111101",
  60196=>"110000000",
  60197=>"000000000",
  60198=>"000000000",
  60199=>"111111111",
  60200=>"000000111",
  60201=>"000000100",
  60202=>"100100101",
  60203=>"000001000",
  60204=>"111011111",
  60205=>"011001001",
  60206=>"111111010",
  60207=>"000000000",
  60208=>"000000000",
  60209=>"111011111",
  60210=>"111111111",
  60211=>"000000000",
  60212=>"000100110",
  60213=>"000000100",
  60214=>"111001000",
  60215=>"000000000",
  60216=>"000000000",
  60217=>"101000000",
  60218=>"010000000",
  60219=>"101111111",
  60220=>"000000000",
  60221=>"100100000",
  60222=>"011111111",
  60223=>"000000000",
  60224=>"000011000",
  60225=>"000000000",
  60226=>"100001111",
  60227=>"000000101",
  60228=>"000111111",
  60229=>"111111111",
  60230=>"000000000",
  60231=>"100000000",
  60232=>"000000000",
  60233=>"000110111",
  60234=>"111111011",
  60235=>"111101001",
  60236=>"111001111",
  60237=>"111001000",
  60238=>"000000000",
  60239=>"111111100",
  60240=>"000100111",
  60241=>"111111000",
  60242=>"111111111",
  60243=>"000000000",
  60244=>"000000000",
  60245=>"001001011",
  60246=>"000111111",
  60247=>"111111111",
  60248=>"111111111",
  60249=>"111111001",
  60250=>"111111110",
  60251=>"000000000",
  60252=>"000000000",
  60253=>"000000000",
  60254=>"000000000",
  60255=>"111111111",
  60256=>"000111000",
  60257=>"111111111",
  60258=>"001000000",
  60259=>"100100111",
  60260=>"111111000",
  60261=>"000000000",
  60262=>"000000000",
  60263=>"111111111",
  60264=>"001001001",
  60265=>"010010000",
  60266=>"011111000",
  60267=>"111111111",
  60268=>"000000000",
  60269=>"000111111",
  60270=>"110111111",
  60271=>"111100110",
  60272=>"110111000",
  60273=>"000000000",
  60274=>"000000000",
  60275=>"111001001",
  60276=>"000010010",
  60277=>"100000001",
  60278=>"111111011",
  60279=>"111111111",
  60280=>"000000000",
  60281=>"111011010",
  60282=>"001000001",
  60283=>"111111111",
  60284=>"000000000",
  60285=>"111111111",
  60286=>"111000011",
  60287=>"111111111",
  60288=>"100100000",
  60289=>"110110110",
  60290=>"000000000",
  60291=>"000000111",
  60292=>"000101111",
  60293=>"100100100",
  60294=>"111111001",
  60295=>"000000000",
  60296=>"111111000",
  60297=>"111111110",
  60298=>"100110110",
  60299=>"000000110",
  60300=>"111111111",
  60301=>"100110010",
  60302=>"101101111",
  60303=>"111111111",
  60304=>"000000000",
  60305=>"111111111",
  60306=>"000000000",
  60307=>"000000000",
  60308=>"110110010",
  60309=>"000000000",
  60310=>"000000000",
  60311=>"000001110",
  60312=>"001101000",
  60313=>"110110110",
  60314=>"000000000",
  60315=>"000000000",
  60316=>"000100111",
  60317=>"001111111",
  60318=>"111000000",
  60319=>"000000000",
  60320=>"100000000",
  60321=>"011011011",
  60322=>"100000100",
  60323=>"001011111",
  60324=>"101101101",
  60325=>"000010110",
  60326=>"111111110",
  60327=>"001111111",
  60328=>"111111100",
  60329=>"100111111",
  60330=>"000000000",
  60331=>"000000110",
  60332=>"000000000",
  60333=>"011111111",
  60334=>"011010000",
  60335=>"000000000",
  60336=>"011111001",
  60337=>"000000001",
  60338=>"110111111",
  60339=>"001000000",
  60340=>"111111111",
  60341=>"000000000",
  60342=>"000110110",
  60343=>"111011011",
  60344=>"001001111",
  60345=>"011001000",
  60346=>"111111011",
  60347=>"100101001",
  60348=>"111111111",
  60349=>"000000000",
  60350=>"111111110",
  60351=>"000000000",
  60352=>"000100110",
  60353=>"000000000",
  60354=>"000000000",
  60355=>"111111110",
  60356=>"111111000",
  60357=>"010010000",
  60358=>"011011000",
  60359=>"100111111",
  60360=>"010000000",
  60361=>"000000000",
  60362=>"000000000",
  60363=>"000000000",
  60364=>"000111000",
  60365=>"010000100",
  60366=>"111100100",
  60367=>"000000000",
  60368=>"000010000",
  60369=>"000000111",
  60370=>"011000000",
  60371=>"111010011",
  60372=>"000000000",
  60373=>"111110010",
  60374=>"000000000",
  60375=>"101110111",
  60376=>"111011000",
  60377=>"111111111",
  60378=>"111111011",
  60379=>"111111111",
  60380=>"110100000",
  60381=>"000000000",
  60382=>"011001000",
  60383=>"000011111",
  60384=>"110110000",
  60385=>"111011001",
  60386=>"011011111",
  60387=>"001101001",
  60388=>"100111111",
  60389=>"000110100",
  60390=>"011000000",
  60391=>"111111111",
  60392=>"111001001",
  60393=>"001000000",
  60394=>"000011011",
  60395=>"111100000",
  60396=>"100100101",
  60397=>"000000000",
  60398=>"000000000",
  60399=>"000000000",
  60400=>"000000000",
  60401=>"000000000",
  60402=>"111111111",
  60403=>"000000000",
  60404=>"000000000",
  60405=>"111011011",
  60406=>"000000000",
  60407=>"110100100",
  60408=>"110111111",
  60409=>"000111110",
  60410=>"111111000",
  60411=>"111000000",
  60412=>"000000111",
  60413=>"000000000",
  60414=>"110100101",
  60415=>"111111111",
  60416=>"000000000",
  60417=>"101011111",
  60418=>"101101111",
  60419=>"111100000",
  60420=>"011011011",
  60421=>"111111111",
  60422=>"000001111",
  60423=>"111100000",
  60424=>"111111111",
  60425=>"111111000",
  60426=>"110000000",
  60427=>"000000111",
  60428=>"000000101",
  60429=>"111111100",
  60430=>"111001100",
  60431=>"001111011",
  60432=>"000000000",
  60433=>"000000000",
  60434=>"010111111",
  60435=>"110010000",
  60436=>"000000000",
  60437=>"111000000",
  60438=>"000000100",
  60439=>"011011110",
  60440=>"000100111",
  60441=>"111111101",
  60442=>"111001000",
  60443=>"111110000",
  60444=>"111110000",
  60445=>"000000000",
  60446=>"111111100",
  60447=>"111111100",
  60448=>"000101000",
  60449=>"001111001",
  60450=>"001001001",
  60451=>"000000000",
  60452=>"000000000",
  60453=>"110111111",
  60454=>"100000101",
  60455=>"000101000",
  60456=>"111100000",
  60457=>"000000000",
  60458=>"111000001",
  60459=>"100000000",
  60460=>"111110111",
  60461=>"000000111",
  60462=>"000001111",
  60463=>"101111000",
  60464=>"111110000",
  60465=>"000001000",
  60466=>"100001001",
  60467=>"000111000",
  60468=>"000000101",
  60469=>"000111011",
  60470=>"000000000",
  60471=>"111111100",
  60472=>"000000111",
  60473=>"111101011",
  60474=>"000001001",
  60475=>"000000000",
  60476=>"000000000",
  60477=>"011000000",
  60478=>"000000000",
  60479=>"101000001",
  60480=>"100110011",
  60481=>"000000111",
  60482=>"000000000",
  60483=>"111011000",
  60484=>"111111111",
  60485=>"000000011",
  60486=>"000000100",
  60487=>"111111111",
  60488=>"110110001",
  60489=>"000000111",
  60490=>"111111111",
  60491=>"011000111",
  60492=>"111111001",
  60493=>"000000100",
  60494=>"000000000",
  60495=>"000110000",
  60496=>"110111000",
  60497=>"110111111",
  60498=>"111011111",
  60499=>"110111000",
  60500=>"000001111",
  60501=>"111101100",
  60502=>"111101101",
  60503=>"000000000",
  60504=>"001000001",
  60505=>"111100000",
  60506=>"000000000",
  60507=>"000000110",
  60508=>"111111010",
  60509=>"111100000",
  60510=>"000000101",
  60511=>"110111000",
  60512=>"111000000",
  60513=>"000011001",
  60514=>"000000110",
  60515=>"111111101",
  60516=>"101001001",
  60517=>"011111111",
  60518=>"111001000",
  60519=>"000111111",
  60520=>"111111000",
  60521=>"111000000",
  60522=>"111111000",
  60523=>"000000111",
  60524=>"000001011",
  60525=>"111111111",
  60526=>"101000111",
  60527=>"000000000",
  60528=>"000000000",
  60529=>"000000111",
  60530=>"111111111",
  60531=>"101001111",
  60532=>"000000111",
  60533=>"010111111",
  60534=>"000000000",
  60535=>"000000000",
  60536=>"001001001",
  60537=>"001000011",
  60538=>"000110000",
  60539=>"100000000",
  60540=>"111111000",
  60541=>"110100000",
  60542=>"000000111",
  60543=>"000011000",
  60544=>"111010111",
  60545=>"000000000",
  60546=>"010110111",
  60547=>"111111111",
  60548=>"011011111",
  60549=>"100100111",
  60550=>"100000000",
  60551=>"111111111",
  60552=>"110000110",
  60553=>"101000100",
  60554=>"111111000",
  60555=>"000000111",
  60556=>"111100111",
  60557=>"000101111",
  60558=>"111111000",
  60559=>"000000000",
  60560=>"000000011",
  60561=>"000011000",
  60562=>"000000111",
  60563=>"000111010",
  60564=>"000000000",
  60565=>"010110111",
  60566=>"111111111",
  60567=>"110000000",
  60568=>"000000000",
  60569=>"111110110",
  60570=>"001001101",
  60571=>"000000000",
  60572=>"000000000",
  60573=>"000000111",
  60574=>"111111101",
  60575=>"011011111",
  60576=>"000000110",
  60577=>"000111111",
  60578=>"001111011",
  60579=>"111111111",
  60580=>"000111001",
  60581=>"000011111",
  60582=>"110111111",
  60583=>"000111100",
  60584=>"000000000",
  60585=>"000000000",
  60586=>"011111001",
  60587=>"000011011",
  60588=>"001001011",
  60589=>"100110110",
  60590=>"111111001",
  60591=>"000000101",
  60592=>"000000101",
  60593=>"000111111",
  60594=>"000111111",
  60595=>"000000000",
  60596=>"011111111",
  60597=>"111000111",
  60598=>"000111110",
  60599=>"110111111",
  60600=>"111111101",
  60601=>"111111111",
  60602=>"000111100",
  60603=>"100100111",
  60604=>"000000000",
  60605=>"100000000",
  60606=>"111111111",
  60607=>"000000001",
  60608=>"101111111",
  60609=>"001111101",
  60610=>"001011011",
  60611=>"010111011",
  60612=>"000111000",
  60613=>"000000100",
  60614=>"111111000",
  60615=>"111111000",
  60616=>"000000000",
  60617=>"111111111",
  60618=>"000000000",
  60619=>"000000110",
  60620=>"111111000",
  60621=>"010111000",
  60622=>"111111000",
  60623=>"000001000",
  60624=>"100110111",
  60625=>"000000000",
  60626=>"100000111",
  60627=>"000111111",
  60628=>"111111111",
  60629=>"101001001",
  60630=>"110110001",
  60631=>"111111111",
  60632=>"111111001",
  60633=>"000001001",
  60634=>"000000000",
  60635=>"001001001",
  60636=>"111010110",
  60637=>"100001111",
  60638=>"110111111",
  60639=>"000000001",
  60640=>"100000000",
  60641=>"000000000",
  60642=>"111111111",
  60643=>"111111101",
  60644=>"000000001",
  60645=>"110111110",
  60646=>"000000111",
  60647=>"111111000",
  60648=>"111111111",
  60649=>"001000000",
  60650=>"000000111",
  60651=>"000000000",
  60652=>"111111111",
  60653=>"000000001",
  60654=>"111101111",
  60655=>"000000000",
  60656=>"111111010",
  60657=>"000000111",
  60658=>"011111000",
  60659=>"010111000",
  60660=>"000000000",
  60661=>"111111000",
  60662=>"000000111",
  60663=>"111000111",
  60664=>"000111111",
  60665=>"000001100",
  60666=>"111111000",
  60667=>"111111110",
  60668=>"110110101",
  60669=>"000000000",
  60670=>"111011111",
  60671=>"000000000",
  60672=>"000000000",
  60673=>"111000000",
  60674=>"111111111",
  60675=>"100110000",
  60676=>"000000000",
  60677=>"101111111",
  60678=>"111110100",
  60679=>"101000000",
  60680=>"111111000",
  60681=>"111111111",
  60682=>"000000001",
  60683=>"000000000",
  60684=>"101000101",
  60685=>"011000001",
  60686=>"111111000",
  60687=>"000000111",
  60688=>"111010000",
  60689=>"000000000",
  60690=>"011000011",
  60691=>"001011111",
  60692=>"000000101",
  60693=>"000100100",
  60694=>"111111000",
  60695=>"000000111",
  60696=>"111111011",
  60697=>"111111110",
  60698=>"000000000",
  60699=>"000000010",
  60700=>"100110000",
  60701=>"111111010",
  60702=>"111111000",
  60703=>"000011111",
  60704=>"100111111",
  60705=>"111111111",
  60706=>"000000000",
  60707=>"110110000",
  60708=>"111000111",
  60709=>"001000000",
  60710=>"000110000",
  60711=>"111111110",
  60712=>"111111111",
  60713=>"000000000",
  60714=>"111111000",
  60715=>"100000000",
  60716=>"000001001",
  60717=>"110111000",
  60718=>"000111111",
  60719=>"000000000",
  60720=>"000000001",
  60721=>"000000100",
  60722=>"111111000",
  60723=>"111111111",
  60724=>"000000000",
  60725=>"000001011",
  60726=>"000110000",
  60727=>"111111111",
  60728=>"110111100",
  60729=>"111000000",
  60730=>"000000111",
  60731=>"111000000",
  60732=>"000000111",
  60733=>"111111100",
  60734=>"000011011",
  60735=>"000000000",
  60736=>"111011000",
  60737=>"100000000",
  60738=>"111101011",
  60739=>"000000000",
  60740=>"111111001",
  60741=>"100000011",
  60742=>"000011111",
  60743=>"100100111",
  60744=>"111101000",
  60745=>"000000000",
  60746=>"110110000",
  60747=>"000000011",
  60748=>"000010011",
  60749=>"111111111",
  60750=>"000000000",
  60751=>"000000111",
  60752=>"000100111",
  60753=>"001000011",
  60754=>"111001001",
  60755=>"000000001",
  60756=>"000111001",
  60757=>"011011111",
  60758=>"111111001",
  60759=>"111111000",
  60760=>"001011111",
  60761=>"111111111",
  60762=>"000000111",
  60763=>"011111000",
  60764=>"111000000",
  60765=>"001000001",
  60766=>"000000110",
  60767=>"001001000",
  60768=>"100110000",
  60769=>"000000000",
  60770=>"111011001",
  60771=>"111000000",
  60772=>"010011011",
  60773=>"000000011",
  60774=>"000001111",
  60775=>"111111000",
  60776=>"000000110",
  60777=>"110111001",
  60778=>"111111000",
  60779=>"110111111",
  60780=>"000110111",
  60781=>"000011010",
  60782=>"110111110",
  60783=>"111000000",
  60784=>"111000000",
  60785=>"100111011",
  60786=>"001011011",
  60787=>"111110100",
  60788=>"001001001",
  60789=>"011011001",
  60790=>"111100110",
  60791=>"111011111",
  60792=>"111000001",
  60793=>"111111000",
  60794=>"111000001",
  60795=>"000000000",
  60796=>"001111111",
  60797=>"001000000",
  60798=>"000000011",
  60799=>"011111111",
  60800=>"110110110",
  60801=>"001001111",
  60802=>"000000010",
  60803=>"111001001",
  60804=>"000000000",
  60805=>"110100110",
  60806=>"111001000",
  60807=>"110111110",
  60808=>"001011111",
  60809=>"000110100",
  60810=>"001000000",
  60811=>"000000000",
  60812=>"001001001",
  60813=>"100111100",
  60814=>"110000000",
  60815=>"011011101",
  60816=>"000000000",
  60817=>"111101001",
  60818=>"000000000",
  60819=>"000000001",
  60820=>"000001111",
  60821=>"000010111",
  60822=>"000111111",
  60823=>"110111111",
  60824=>"000000110",
  60825=>"000000001",
  60826=>"000000011",
  60827=>"111011111",
  60828=>"111111111",
  60829=>"000000000",
  60830=>"000000111",
  60831=>"000000000",
  60832=>"000111000",
  60833=>"111011011",
  60834=>"001111001",
  60835=>"100101101",
  60836=>"101111000",
  60837=>"000111110",
  60838=>"000000000",
  60839=>"000000000",
  60840=>"001111111",
  60841=>"111111111",
  60842=>"111111000",
  60843=>"000000001",
  60844=>"000000110",
  60845=>"000111111",
  60846=>"111101000",
  60847=>"111000000",
  60848=>"000100111",
  60849=>"111011001",
  60850=>"000000000",
  60851=>"111111001",
  60852=>"000000000",
  60853=>"110111110",
  60854=>"111111111",
  60855=>"100110111",
  60856=>"111000000",
  60857=>"111111111",
  60858=>"011100101",
  60859=>"000000000",
  60860=>"000000100",
  60861=>"101111111",
  60862=>"000000000",
  60863=>"100100000",
  60864=>"111111111",
  60865=>"000000000",
  60866=>"000000000",
  60867=>"000000000",
  60868=>"001001111",
  60869=>"101001011",
  60870=>"010111001",
  60871=>"000111111",
  60872=>"000000111",
  60873=>"011000111",
  60874=>"000000000",
  60875=>"000000000",
  60876=>"110000111",
  60877=>"111111000",
  60878=>"100110000",
  60879=>"011111011",
  60880=>"100000000",
  60881=>"111011000",
  60882=>"000000110",
  60883=>"001011001",
  60884=>"111000000",
  60885=>"101111111",
  60886=>"000000111",
  60887=>"001001001",
  60888=>"100100000",
  60889=>"010000000",
  60890=>"111111000",
  60891=>"111111111",
  60892=>"010111011",
  60893=>"111111110",
  60894=>"111111101",
  60895=>"010000000",
  60896=>"000000100",
  60897=>"111111111",
  60898=>"000000100",
  60899=>"111111111",
  60900=>"001001111",
  60901=>"000111000",
  60902=>"100100111",
  60903=>"001000001",
  60904=>"000000000",
  60905=>"111111000",
  60906=>"010110000",
  60907=>"000001111",
  60908=>"111111111",
  60909=>"000001111",
  60910=>"000101111",
  60911=>"111000000",
  60912=>"000001011",
  60913=>"001011011",
  60914=>"100111111",
  60915=>"000000101",
  60916=>"110111011",
  60917=>"000000001",
  60918=>"000011111",
  60919=>"001000110",
  60920=>"111100111",
  60921=>"100010000",
  60922=>"100111101",
  60923=>"000000001",
  60924=>"111010111",
  60925=>"000001001",
  60926=>"000000001",
  60927=>"100000111",
  60928=>"101111111",
  60929=>"011000001",
  60930=>"000000111",
  60931=>"000000000",
  60932=>"111001101",
  60933=>"000000000",
  60934=>"010000000",
  60935=>"111111111",
  60936=>"111111000",
  60937=>"000011111",
  60938=>"111111110",
  60939=>"000110111",
  60940=>"000000000",
  60941=>"111100000",
  60942=>"000001001",
  60943=>"111111000",
  60944=>"011111111",
  60945=>"000010110",
  60946=>"111111111",
  60947=>"111111000",
  60948=>"111111111",
  60949=>"000000100",
  60950=>"111111111",
  60951=>"011011011",
  60952=>"000000111",
  60953=>"000000000",
  60954=>"111110111",
  60955=>"000000111",
  60956=>"110110110",
  60957=>"010110100",
  60958=>"111000000",
  60959=>"000000111",
  60960=>"111111011",
  60961=>"111110110",
  60962=>"111111100",
  60963=>"000000000",
  60964=>"111110000",
  60965=>"000000000",
  60966=>"111100000",
  60967=>"111111111",
  60968=>"000000111",
  60969=>"000000000",
  60970=>"110110000",
  60971=>"100000100",
  60972=>"111111100",
  60973=>"111111000",
  60974=>"100110111",
  60975=>"111111111",
  60976=>"100000000",
  60977=>"000000000",
  60978=>"000000000",
  60979=>"111010000",
  60980=>"011011111",
  60981=>"010011000",
  60982=>"111110111",
  60983=>"010010011",
  60984=>"000000011",
  60985=>"111101111",
  60986=>"000000000",
  60987=>"011111111",
  60988=>"000001000",
  60989=>"111111111",
  60990=>"000000110",
  60991=>"111111011",
  60992=>"000000101",
  60993=>"111111111",
  60994=>"000000011",
  60995=>"111111000",
  60996=>"010000000",
  60997=>"000000011",
  60998=>"000000100",
  60999=>"111111111",
  61000=>"100000000",
  61001=>"000000111",
  61002=>"111111110",
  61003=>"000000000",
  61004=>"011011111",
  61005=>"110100100",
  61006=>"000000000",
  61007=>"111111100",
  61008=>"000111111",
  61009=>"011011101",
  61010=>"110100000",
  61011=>"000000000",
  61012=>"111111111",
  61013=>"111111111",
  61014=>"111000111",
  61015=>"110110110",
  61016=>"111101101",
  61017=>"101000000",
  61018=>"111111111",
  61019=>"111111001",
  61020=>"000001111",
  61021=>"111110000",
  61022=>"011001001",
  61023=>"111000000",
  61024=>"111111110",
  61025=>"011000100",
  61026=>"000000000",
  61027=>"111101000",
  61028=>"001001100",
  61029=>"000000000",
  61030=>"100000000",
  61031=>"111111000",
  61032=>"111111000",
  61033=>"111100000",
  61034=>"111111111",
  61035=>"000000010",
  61036=>"001011111",
  61037=>"111111111",
  61038=>"010111111",
  61039=>"010011011",
  61040=>"111111001",
  61041=>"000000100",
  61042=>"101111111",
  61043=>"000001111",
  61044=>"110110111",
  61045=>"111111111",
  61046=>"101111110",
  61047=>"011100111",
  61048=>"000000100",
  61049=>"000000000",
  61050=>"101101000",
  61051=>"000000100",
  61052=>"010000000",
  61053=>"000110011",
  61054=>"001001001",
  61055=>"010100111",
  61056=>"000011000",
  61057=>"111111111",
  61058=>"011001000",
  61059=>"000000000",
  61060=>"111011110",
  61061=>"001000000",
  61062=>"000000000",
  61063=>"110100100",
  61064=>"111111111",
  61065=>"000010111",
  61066=>"000000000",
  61067=>"100110111",
  61068=>"000000000",
  61069=>"011000000",
  61070=>"111111111",
  61071=>"000000000",
  61072=>"000000000",
  61073=>"100111111",
  61074=>"000100111",
  61075=>"010010111",
  61076=>"110000111",
  61077=>"000010000",
  61078=>"000000000",
  61079=>"111111111",
  61080=>"111000000",
  61081=>"111101100",
  61082=>"111111111",
  61083=>"000000000",
  61084=>"111110000",
  61085=>"111111111",
  61086=>"010000000",
  61087=>"000000000",
  61088=>"000000000",
  61089=>"011000000",
  61090=>"100110111",
  61091=>"111111111",
  61092=>"000000001",
  61093=>"010000001",
  61094=>"000000100",
  61095=>"101111111",
  61096=>"100000111",
  61097=>"000000111",
  61098=>"100000000",
  61099=>"111110100",
  61100=>"011111111",
  61101=>"000000000",
  61102=>"000000000",
  61103=>"000000001",
  61104=>"000011111",
  61105=>"000000000",
  61106=>"110110111",
  61107=>"000000000",
  61108=>"111101100",
  61109=>"111111111",
  61110=>"110000000",
  61111=>"000010000",
  61112=>"111101111",
  61113=>"000000110",
  61114=>"000000000",
  61115=>"111111000",
  61116=>"001001111",
  61117=>"111111111",
  61118=>"110000101",
  61119=>"100000000",
  61120=>"000110000",
  61121=>"010000000",
  61122=>"011001111",
  61123=>"000000000",
  61124=>"111101100",
  61125=>"111000000",
  61126=>"000000000",
  61127=>"100100100",
  61128=>"111111000",
  61129=>"000000011",
  61130=>"100111111",
  61131=>"000000000",
  61132=>"001000111",
  61133=>"011000100",
  61134=>"010000000",
  61135=>"000000111",
  61136=>"101100100",
  61137=>"000010001",
  61138=>"000000000",
  61139=>"000000000",
  61140=>"000000000",
  61141=>"111001000",
  61142=>"000000000",
  61143=>"000000110",
  61144=>"111101100",
  61145=>"000100100",
  61146=>"000000110",
  61147=>"111111111",
  61148=>"111111000",
  61149=>"000000000",
  61150=>"011001000",
  61151=>"011000111",
  61152=>"001000100",
  61153=>"111111000",
  61154=>"110111111",
  61155=>"111000100",
  61156=>"101001000",
  61157=>"111111010",
  61158=>"110111011",
  61159=>"111111101",
  61160=>"000110111",
  61161=>"111111111",
  61162=>"000001111",
  61163=>"111111111",
  61164=>"000001001",
  61165=>"010110111",
  61166=>"111111001",
  61167=>"000000000",
  61168=>"010000111",
  61169=>"110010010",
  61170=>"011001001",
  61171=>"000000000",
  61172=>"111111111",
  61173=>"111111000",
  61174=>"011010011",
  61175=>"011000000",
  61176=>"000010010",
  61177=>"110000110",
  61178=>"011001000",
  61179=>"111111111",
  61180=>"000000000",
  61181=>"111111111",
  61182=>"111011010",
  61183=>"000000000",
  61184=>"000000000",
  61185=>"111111100",
  61186=>"111111111",
  61187=>"000011011",
  61188=>"111111111",
  61189=>"001000000",
  61190=>"000100000",
  61191=>"000011111",
  61192=>"111011011",
  61193=>"111000000",
  61194=>"000000000",
  61195=>"000000111",
  61196=>"111111111",
  61197=>"000000110",
  61198=>"000000000",
  61199=>"100111000",
  61200=>"111110100",
  61201=>"111100000",
  61202=>"000000110",
  61203=>"001001000",
  61204=>"000000111",
  61205=>"111111111",
  61206=>"001000001",
  61207=>"010000110",
  61208=>"000011111",
  61209=>"000000000",
  61210=>"000000111",
  61211=>"110011011",
  61212=>"000000000",
  61213=>"000000000",
  61214=>"011111111",
  61215=>"111000001",
  61216=>"110111111",
  61217=>"001000000",
  61218=>"001000000",
  61219=>"110000000",
  61220=>"000000110",
  61221=>"111111001",
  61222=>"001000000",
  61223=>"001000111",
  61224=>"100110100",
  61225=>"000000000",
  61226=>"000111000",
  61227=>"100110000",
  61228=>"000000111",
  61229=>"000000111",
  61230=>"100110111",
  61231=>"000010000",
  61232=>"111110111",
  61233=>"110000100",
  61234=>"000000000",
  61235=>"111111111",
  61236=>"001000000",
  61237=>"111111111",
  61238=>"111001000",
  61239=>"000000000",
  61240=>"110100110",
  61241=>"111101000",
  61242=>"100100100",
  61243=>"000000111",
  61244=>"000000001",
  61245=>"110111000",
  61246=>"110101101",
  61247=>"111111111",
  61248=>"000000001",
  61249=>"011011000",
  61250=>"111001001",
  61251=>"000110111",
  61252=>"000000010",
  61253=>"000000000",
  61254=>"000000100",
  61255=>"111111110",
  61256=>"011010000",
  61257=>"000110111",
  61258=>"111111001",
  61259=>"000011001",
  61260=>"011000001",
  61261=>"000001001",
  61262=>"111111111",
  61263=>"111111111",
  61264=>"010000111",
  61265=>"000000101",
  61266=>"111111011",
  61267=>"000100100",
  61268=>"011000000",
  61269=>"000010000",
  61270=>"110111111",
  61271=>"111110000",
  61272=>"111011011",
  61273=>"000000000",
  61274=>"111111111",
  61275=>"000000101",
  61276=>"000000000",
  61277=>"000000111",
  61278=>"111010111",
  61279=>"001111111",
  61280=>"000000001",
  61281=>"000000100",
  61282=>"010001000",
  61283=>"111111111",
  61284=>"000000000",
  61285=>"110000000",
  61286=>"111111111",
  61287=>"000000000",
  61288=>"001110111",
  61289=>"000100000",
  61290=>"100111111",
  61291=>"000110111",
  61292=>"000000000",
  61293=>"000000111",
  61294=>"000000000",
  61295=>"111101111",
  61296=>"111111001",
  61297=>"000111110",
  61298=>"000000000",
  61299=>"111111111",
  61300=>"110111111",
  61301=>"000000100",
  61302=>"111111111",
  61303=>"001101101",
  61304=>"110110110",
  61305=>"000000000",
  61306=>"111101011",
  61307=>"111100100",
  61308=>"000000000",
  61309=>"000000100",
  61310=>"000000000",
  61311=>"011000000",
  61312=>"000000000",
  61313=>"010000111",
  61314=>"000111110",
  61315=>"000000000",
  61316=>"000000111",
  61317=>"000000100",
  61318=>"111111111",
  61319=>"111110111",
  61320=>"000000111",
  61321=>"111111011",
  61322=>"011000000",
  61323=>"111111111",
  61324=>"000001001",
  61325=>"000000000",
  61326=>"000000111",
  61327=>"011000011",
  61328=>"111111000",
  61329=>"001001101",
  61330=>"001011111",
  61331=>"000000000",
  61332=>"000000110",
  61333=>"110111000",
  61334=>"001000000",
  61335=>"011000000",
  61336=>"111101000",
  61337=>"000000000",
  61338=>"111111111",
  61339=>"000111111",
  61340=>"000000000",
  61341=>"000000000",
  61342=>"000000000",
  61343=>"000000000",
  61344=>"000000000",
  61345=>"000000101",
  61346=>"000011000",
  61347=>"111111111",
  61348=>"000011001",
  61349=>"111111111",
  61350=>"000101111",
  61351=>"000000011",
  61352=>"111111111",
  61353=>"111111111",
  61354=>"111010101",
  61355=>"010010000",
  61356=>"010000111",
  61357=>"111011111",
  61358=>"000000001",
  61359=>"111111111",
  61360=>"000000000",
  61361=>"000000000",
  61362=>"011001000",
  61363=>"000000000",
  61364=>"111111111",
  61365=>"000000000",
  61366=>"111111111",
  61367=>"100000000",
  61368=>"111100000",
  61369=>"111111111",
  61370=>"000000000",
  61371=>"110111100",
  61372=>"111111110",
  61373=>"110111111",
  61374=>"000000000",
  61375=>"000000000",
  61376=>"111111000",
  61377=>"110000000",
  61378=>"000000000",
  61379=>"010000001",
  61380=>"010111111",
  61381=>"111010010",
  61382=>"111111000",
  61383=>"111100100",
  61384=>"111011111",
  61385=>"111111111",
  61386=>"111000000",
  61387=>"111111111",
  61388=>"100001111",
  61389=>"001011011",
  61390=>"000001111",
  61391=>"111111111",
  61392=>"000000000",
  61393=>"111111011",
  61394=>"011111111",
  61395=>"000101000",
  61396=>"100000000",
  61397=>"111111000",
  61398=>"111111111",
  61399=>"000000000",
  61400=>"000000000",
  61401=>"011010011",
  61402=>"100000000",
  61403=>"010010111",
  61404=>"110111111",
  61405=>"111111111",
  61406=>"011000111",
  61407=>"000000100",
  61408=>"111000000",
  61409=>"100100000",
  61410=>"111111000",
  61411=>"111111111",
  61412=>"111111111",
  61413=>"001011000",
  61414=>"111111111",
  61415=>"010000000",
  61416=>"000000111",
  61417=>"000000000",
  61418=>"100000000",
  61419=>"000101111",
  61420=>"000000000",
  61421=>"000000000",
  61422=>"111011111",
  61423=>"011011001",
  61424=>"000000000",
  61425=>"111111111",
  61426=>"000001001",
  61427=>"110110111",
  61428=>"000000000",
  61429=>"111111111",
  61430=>"111010000",
  61431=>"000000000",
  61432=>"011011000",
  61433=>"010000010",
  61434=>"111111111",
  61435=>"110110100",
  61436=>"110111111",
  61437=>"111111111",
  61438=>"111001011",
  61439=>"111111111",
  61440=>"001001011",
  61441=>"111111100",
  61442=>"111111111",
  61443=>"111111111",
  61444=>"111111111",
  61445=>"010010111",
  61446=>"000000000",
  61447=>"111111111",
  61448=>"000110110",
  61449=>"100100101",
  61450=>"000100111",
  61451=>"110111000",
  61452=>"001000011",
  61453=>"000000101",
  61454=>"111000000",
  61455=>"000000000",
  61456=>"111110000",
  61457=>"000000011",
  61458=>"000010010",
  61459=>"000000101",
  61460=>"000000000",
  61461=>"000000000",
  61462=>"000000000",
  61463=>"000000000",
  61464=>"111111110",
  61465=>"111111000",
  61466=>"111111111",
  61467=>"011000000",
  61468=>"111100100",
  61469=>"000000000",
  61470=>"001001001",
  61471=>"000001000",
  61472=>"000010000",
  61473=>"111111111",
  61474=>"001011010",
  61475=>"111111111",
  61476=>"111111111",
  61477=>"000000001",
  61478=>"000000000",
  61479=>"000000000",
  61480=>"100101100",
  61481=>"000000000",
  61482=>"000000000",
  61483=>"111111100",
  61484=>"111111111",
  61485=>"110111111",
  61486=>"000010000",
  61487=>"110110011",
  61488=>"000000000",
  61489=>"000000000",
  61490=>"110110010",
  61491=>"000000101",
  61492=>"000000000",
  61493=>"110001000",
  61494=>"000000000",
  61495=>"000000000",
  61496=>"100000110",
  61497=>"111111111",
  61498=>"111001000",
  61499=>"000000011",
  61500=>"000000000",
  61501=>"000000000",
  61502=>"011010110",
  61503=>"100000000",
  61504=>"111111111",
  61505=>"000111100",
  61506=>"111111111",
  61507=>"110000111",
  61508=>"100111111",
  61509=>"000000001",
  61510=>"111111111",
  61511=>"111111111",
  61512=>"110111111",
  61513=>"111111111",
  61514=>"000110000",
  61515=>"110110000",
  61516=>"000000000",
  61517=>"100100111",
  61518=>"000000000",
  61519=>"111111111",
  61520=>"111111111",
  61521=>"111110000",
  61522=>"001001000",
  61523=>"111111111",
  61524=>"111111000",
  61525=>"000000100",
  61526=>"111000001",
  61527=>"111111111",
  61528=>"100000000",
  61529=>"001000101",
  61530=>"111111000",
  61531=>"001000000",
  61532=>"111111111",
  61533=>"000111111",
  61534=>"001001000",
  61535=>"000000000",
  61536=>"000000010",
  61537=>"010111010",
  61538=>"000111111",
  61539=>"000011111",
  61540=>"000000000",
  61541=>"000000010",
  61542=>"111100111",
  61543=>"000000000",
  61544=>"111111110",
  61545=>"111111010",
  61546=>"000111111",
  61547=>"000000000",
  61548=>"000001001",
  61549=>"100111000",
  61550=>"000000000",
  61551=>"000000101",
  61552=>"000010000",
  61553=>"111010101",
  61554=>"000111000",
  61555=>"000000000",
  61556=>"111111111",
  61557=>"000000001",
  61558=>"111111000",
  61559=>"000000000",
  61560=>"000000010",
  61561=>"111111111",
  61562=>"000000000",
  61563=>"000000000",
  61564=>"100000100",
  61565=>"000000000",
  61566=>"000000000",
  61567=>"111111000",
  61568=>"000000111",
  61569=>"000000100",
  61570=>"000000000",
  61571=>"001001111",
  61572=>"000000000",
  61573=>"011101111",
  61574=>"011111001",
  61575=>"000100000",
  61576=>"000000000",
  61577=>"000000000",
  61578=>"000111111",
  61579=>"110000000",
  61580=>"000010000",
  61581=>"111111111",
  61582=>"100000000",
  61583=>"000000000",
  61584=>"000101000",
  61585=>"111111110",
  61586=>"000000000",
  61587=>"110110100",
  61588=>"000110110",
  61589=>"000111111",
  61590=>"111111111",
  61591=>"111111111",
  61592=>"000000000",
  61593=>"111111110",
  61594=>"000000000",
  61595=>"100101000",
  61596=>"100000000",
  61597=>"100100100",
  61598=>"100000000",
  61599=>"000000000",
  61600=>"111101001",
  61601=>"111111110",
  61602=>"111111111",
  61603=>"000000001",
  61604=>"111001011",
  61605=>"111111111",
  61606=>"000111111",
  61607=>"001001000",
  61608=>"110110000",
  61609=>"000000111",
  61610=>"000000000",
  61611=>"111111100",
  61612=>"000000000",
  61613=>"001001110",
  61614=>"100000000",
  61615=>"110111011",
  61616=>"000000000",
  61617=>"110111111",
  61618=>"111111100",
  61619=>"111111111",
  61620=>"000000000",
  61621=>"111111001",
  61622=>"110111111",
  61623=>"000000000",
  61624=>"100000001",
  61625=>"000000111",
  61626=>"111000000",
  61627=>"100101111",
  61628=>"011000000",
  61629=>"111111111",
  61630=>"000000000",
  61631=>"000001001",
  61632=>"111111111",
  61633=>"110110111",
  61634=>"111111111",
  61635=>"011000000",
  61636=>"111111111",
  61637=>"011011011",
  61638=>"000000000",
  61639=>"111111111",
  61640=>"100110111",
  61641=>"100101011",
  61642=>"000000000",
  61643=>"011111111",
  61644=>"110111111",
  61645=>"111111110",
  61646=>"000000110",
  61647=>"100000000",
  61648=>"010000011",
  61649=>"000000101",
  61650=>"001000100",
  61651=>"111111111",
  61652=>"100000000",
  61653=>"110111111",
  61654=>"000000000",
  61655=>"000011000",
  61656=>"000000000",
  61657=>"111111111",
  61658=>"001000000",
  61659=>"000100010",
  61660=>"111110101",
  61661=>"011010000",
  61662=>"011111111",
  61663=>"111000111",
  61664=>"111111111",
  61665=>"011001111",
  61666=>"110000000",
  61667=>"000000000",
  61668=>"111110111",
  61669=>"100100000",
  61670=>"111111111",
  61671=>"101000000",
  61672=>"111111111",
  61673=>"111010100",
  61674=>"110010000",
  61675=>"110010010",
  61676=>"111111111",
  61677=>"111111111",
  61678=>"111111111",
  61679=>"010110111",
  61680=>"101100100",
  61681=>"111101100",
  61682=>"000000000",
  61683=>"111001000",
  61684=>"000100001",
  61685=>"111001000",
  61686=>"001011100",
  61687=>"110000000",
  61688=>"000001000",
  61689=>"111110000",
  61690=>"111000000",
  61691=>"011111111",
  61692=>"100110110",
  61693=>"111111001",
  61694=>"000000000",
  61695=>"000000100",
  61696=>"101111000",
  61697=>"001000000",
  61698=>"001111111",
  61699=>"100111111",
  61700=>"000000111",
  61701=>"100100101",
  61702=>"000000000",
  61703=>"111000100",
  61704=>"000000101",
  61705=>"000000000",
  61706=>"000110111",
  61707=>"011000111",
  61708=>"111111000",
  61709=>"000000000",
  61710=>"000000011",
  61711=>"000111000",
  61712=>"000000011",
  61713=>"111111111",
  61714=>"111100100",
  61715=>"100100110",
  61716=>"111111111",
  61717=>"111111111",
  61718=>"001001001",
  61719=>"110110000",
  61720=>"111111111",
  61721=>"111111111",
  61722=>"000000000",
  61723=>"111111111",
  61724=>"110111101",
  61725=>"111111111",
  61726=>"000000000",
  61727=>"111111111",
  61728=>"111011011",
  61729=>"000001001",
  61730=>"111000000",
  61731=>"110110111",
  61732=>"000000100",
  61733=>"000000000",
  61734=>"110111111",
  61735=>"000000000",
  61736=>"000000000",
  61737=>"100101111",
  61738=>"110110111",
  61739=>"000000001",
  61740=>"111111000",
  61741=>"100000000",
  61742=>"000000110",
  61743=>"000000000",
  61744=>"110111110",
  61745=>"110111001",
  61746=>"000000000",
  61747=>"000010011",
  61748=>"010010000",
  61749=>"010010000",
  61750=>"000000000",
  61751=>"111001111",
  61752=>"000000000",
  61753=>"111111101",
  61754=>"010010000",
  61755=>"001000111",
  61756=>"001001000",
  61757=>"000000010",
  61758=>"100110111",
  61759=>"000111111",
  61760=>"101101000",
  61761=>"111111101",
  61762=>"000000000",
  61763=>"000000000",
  61764=>"011111000",
  61765=>"000110110",
  61766=>"111111111",
  61767=>"000000000",
  61768=>"000000000",
  61769=>"000000000",
  61770=>"111111111",
  61771=>"100000100",
  61772=>"111111111",
  61773=>"111111110",
  61774=>"110101111",
  61775=>"110100110",
  61776=>"000110110",
  61777=>"110000011",
  61778=>"111111101",
  61779=>"000000111",
  61780=>"000000000",
  61781=>"001011001",
  61782=>"111100111",
  61783=>"110100111",
  61784=>"000001111",
  61785=>"000000000",
  61786=>"100111111",
  61787=>"110011000",
  61788=>"000000111",
  61789=>"100101101",
  61790=>"000010111",
  61791=>"100000000",
  61792=>"100000101",
  61793=>"011111111",
  61794=>"101000000",
  61795=>"000111111",
  61796=>"100000000",
  61797=>"111000000",
  61798=>"111111111",
  61799=>"000000100",
  61800=>"001001001",
  61801=>"111010000",
  61802=>"000000000",
  61803=>"100001001",
  61804=>"000100111",
  61805=>"111111111",
  61806=>"000000111",
  61807=>"101100100",
  61808=>"011110111",
  61809=>"111110111",
  61810=>"111110111",
  61811=>"111110110",
  61812=>"111111111",
  61813=>"001000100",
  61814=>"000000000",
  61815=>"000000000",
  61816=>"011111111",
  61817=>"001000000",
  61818=>"000000000",
  61819=>"110100000",
  61820=>"111101111",
  61821=>"110111111",
  61822=>"000000000",
  61823=>"100111111",
  61824=>"111111000",
  61825=>"111010010",
  61826=>"000111110",
  61827=>"000111111",
  61828=>"111111111",
  61829=>"000000000",
  61830=>"000000000",
  61831=>"110000000",
  61832=>"000000000",
  61833=>"100110111",
  61834=>"110000111",
  61835=>"111111111",
  61836=>"111111111",
  61837=>"111111111",
  61838=>"111111110",
  61839=>"000000000",
  61840=>"111000000",
  61841=>"100001001",
  61842=>"110110100",
  61843=>"110110111",
  61844=>"011000000",
  61845=>"011111000",
  61846=>"000000001",
  61847=>"111111000",
  61848=>"000111100",
  61849=>"000000000",
  61850=>"000000000",
  61851=>"110001000",
  61852=>"100111011",
  61853=>"000000000",
  61854=>"111101100",
  61855=>"111110100",
  61856=>"101000110",
  61857=>"011011011",
  61858=>"110000000",
  61859=>"000000000",
  61860=>"110110100",
  61861=>"111111100",
  61862=>"000000000",
  61863=>"011011011",
  61864=>"011001000",
  61865=>"000000111",
  61866=>"000000111",
  61867=>"111011011",
  61868=>"000000000",
  61869=>"000000000",
  61870=>"111111111",
  61871=>"111111000",
  61872=>"110100111",
  61873=>"000000001",
  61874=>"100100100",
  61875=>"000000000",
  61876=>"111111111",
  61877=>"000111111",
  61878=>"000001111",
  61879=>"110100000",
  61880=>"100111100",
  61881=>"000000000",
  61882=>"000011111",
  61883=>"110100100",
  61884=>"111111111",
  61885=>"101111100",
  61886=>"100111000",
  61887=>"111000000",
  61888=>"011011111",
  61889=>"000000000",
  61890=>"111111011",
  61891=>"111101000",
  61892=>"111111111",
  61893=>"100000101",
  61894=>"000011011",
  61895=>"000000111",
  61896=>"000000000",
  61897=>"111111111",
  61898=>"110000000",
  61899=>"111111111",
  61900=>"000110000",
  61901=>"111111111",
  61902=>"000000000",
  61903=>"111010110",
  61904=>"000000010",
  61905=>"000000000",
  61906=>"111111011",
  61907=>"011111011",
  61908=>"001101001",
  61909=>"111111111",
  61910=>"110000000",
  61911=>"000000011",
  61912=>"100001001",
  61913=>"110110011",
  61914=>"111111111",
  61915=>"001001000",
  61916=>"001000000",
  61917=>"000000000",
  61918=>"111111011",
  61919=>"001001001",
  61920=>"111110111",
  61921=>"011011000",
  61922=>"111111111",
  61923=>"101000000",
  61924=>"100101001",
  61925=>"010110100",
  61926=>"000111100",
  61927=>"111111111",
  61928=>"111111111",
  61929=>"000000000",
  61930=>"111111011",
  61931=>"111111100",
  61932=>"111011111",
  61933=>"111011000",
  61934=>"000000000",
  61935=>"100011111",
  61936=>"100100000",
  61937=>"100100101",
  61938=>"000000000",
  61939=>"000000000",
  61940=>"111111011",
  61941=>"000000000",
  61942=>"000000010",
  61943=>"000101111",
  61944=>"011011010",
  61945=>"100100000",
  61946=>"111111100",
  61947=>"000001000",
  61948=>"111000000",
  61949=>"111000000",
  61950=>"111011000",
  61951=>"000000110",
  61952=>"001100110",
  61953=>"000000000",
  61954=>"110000000",
  61955=>"111001000",
  61956=>"000101100",
  61957=>"000000100",
  61958=>"011001111",
  61959=>"111111110",
  61960=>"111111001",
  61961=>"000001000",
  61962=>"111111111",
  61963=>"101000000",
  61964=>"111011111",
  61965=>"110111111",
  61966=>"000000000",
  61967=>"000000110",
  61968=>"111011001",
  61969=>"000000000",
  61970=>"001010110",
  61971=>"001111111",
  61972=>"000000000",
  61973=>"111111000",
  61974=>"000000000",
  61975=>"111111111",
  61976=>"101111010",
  61977=>"101000100",
  61978=>"000000000",
  61979=>"000000000",
  61980=>"000000000",
  61981=>"111111111",
  61982=>"100000100",
  61983=>"001000000",
  61984=>"000000000",
  61985=>"111111111",
  61986=>"000001001",
  61987=>"111111111",
  61988=>"000111111",
  61989=>"110110101",
  61990=>"011011010",
  61991=>"000001000",
  61992=>"000000110",
  61993=>"000000000",
  61994=>"111111111",
  61995=>"111111010",
  61996=>"010011111",
  61997=>"111000000",
  61998=>"000000111",
  61999=>"111111010",
  62000=>"000000000",
  62001=>"000000100",
  62002=>"001000100",
  62003=>"110010000",
  62004=>"001001111",
  62005=>"011010000",
  62006=>"001000000",
  62007=>"110011111",
  62008=>"111111111",
  62009=>"110011011",
  62010=>"111000000",
  62011=>"000001101",
  62012=>"000111111",
  62013=>"111111111",
  62014=>"001001001",
  62015=>"000000100",
  62016=>"010010111",
  62017=>"110111011",
  62018=>"111100101",
  62019=>"111111111",
  62020=>"100000000",
  62021=>"001000000",
  62022=>"000001001",
  62023=>"000000111",
  62024=>"000100101",
  62025=>"111111101",
  62026=>"111011001",
  62027=>"000000000",
  62028=>"100000000",
  62029=>"111111000",
  62030=>"000000011",
  62031=>"011000000",
  62032=>"100100111",
  62033=>"000000011",
  62034=>"000000000",
  62035=>"011011001",
  62036=>"111111111",
  62037=>"000000111",
  62038=>"100001000",
  62039=>"000000000",
  62040=>"111111111",
  62041=>"000001111",
  62042=>"000000000",
  62043=>"110101101",
  62044=>"000000010",
  62045=>"110101001",
  62046=>"000000000",
  62047=>"111111111",
  62048=>"111111111",
  62049=>"011111111",
  62050=>"111111011",
  62051=>"010000010",
  62052=>"100111011",
  62053=>"110111000",
  62054=>"000001000",
  62055=>"000000000",
  62056=>"111110000",
  62057=>"110111110",
  62058=>"110111110",
  62059=>"000000000",
  62060=>"000000100",
  62061=>"000001011",
  62062=>"100100111",
  62063=>"111111111",
  62064=>"000010000",
  62065=>"000000100",
  62066=>"100111111",
  62067=>"000000000",
  62068=>"011001000",
  62069=>"010100100",
  62070=>"000000000",
  62071=>"111111110",
  62072=>"111111111",
  62073=>"111111111",
  62074=>"000000000",
  62075=>"000000000",
  62076=>"111111111",
  62077=>"100101111",
  62078=>"000110111",
  62079=>"011001000",
  62080=>"111111111",
  62081=>"000111111",
  62082=>"000000000",
  62083=>"000110000",
  62084=>"101110110",
  62085=>"100100111",
  62086=>"111111110",
  62087=>"000000000",
  62088=>"111111111",
  62089=>"000000100",
  62090=>"011001000",
  62091=>"010000000",
  62092=>"111111000",
  62093=>"001000000",
  62094=>"000010000",
  62095=>"000000000",
  62096=>"000000000",
  62097=>"011000000",
  62098=>"000000000",
  62099=>"110000000",
  62100=>"111111111",
  62101=>"101000000",
  62102=>"111111111",
  62103=>"111111111",
  62104=>"111000111",
  62105=>"111111110",
  62106=>"000000000",
  62107=>"000000010",
  62108=>"111111111",
  62109=>"000000000",
  62110=>"000000011",
  62111=>"110000000",
  62112=>"011010010",
  62113=>"111110110",
  62114=>"111111111",
  62115=>"100000000",
  62116=>"011010000",
  62117=>"001111101",
  62118=>"011111111",
  62119=>"111001111",
  62120=>"110111111",
  62121=>"000001111",
  62122=>"111111000",
  62123=>"001000000",
  62124=>"110010011",
  62125=>"100011110",
  62126=>"111011110",
  62127=>"000100111",
  62128=>"000000111",
  62129=>"111110100",
  62130=>"000000100",
  62131=>"111111111",
  62132=>"000001111",
  62133=>"111111111",
  62134=>"111111111",
  62135=>"111111011",
  62136=>"100100000",
  62137=>"110110110",
  62138=>"100000011",
  62139=>"111001011",
  62140=>"111111111",
  62141=>"110001000",
  62142=>"011000000",
  62143=>"100000111",
  62144=>"000000011",
  62145=>"011000000",
  62146=>"010010111",
  62147=>"111101000",
  62148=>"100111111",
  62149=>"111011000",
  62150=>"000000000",
  62151=>"000000000",
  62152=>"000000000",
  62153=>"111111011",
  62154=>"000000011",
  62155=>"110000000",
  62156=>"000000000",
  62157=>"111011111",
  62158=>"011000011",
  62159=>"000000000",
  62160=>"111111011",
  62161=>"000000010",
  62162=>"000000111",
  62163=>"000000100",
  62164=>"000000000",
  62165=>"000000000",
  62166=>"000110110",
  62167=>"000001111",
  62168=>"101111111",
  62169=>"110111001",
  62170=>"111111111",
  62171=>"001001111",
  62172=>"111111111",
  62173=>"111111111",
  62174=>"000000111",
  62175=>"000000000",
  62176=>"110110111",
  62177=>"000000111",
  62178=>"111111100",
  62179=>"000000000",
  62180=>"001111111",
  62181=>"000000000",
  62182=>"111011110",
  62183=>"100100111",
  62184=>"101011000",
  62185=>"001000000",
  62186=>"111011001",
  62187=>"000011111",
  62188=>"000000000",
  62189=>"110010110",
  62190=>"000000100",
  62191=>"100000000",
  62192=>"000000111",
  62193=>"111111111",
  62194=>"000000000",
  62195=>"001001000",
  62196=>"100000000",
  62197=>"111111111",
  62198=>"000000010",
  62199=>"001000000",
  62200=>"111111111",
  62201=>"111000000",
  62202=>"000000000",
  62203=>"111011000",
  62204=>"011000100",
  62205=>"000000010",
  62206=>"011011011",
  62207=>"111001100",
  62208=>"111011011",
  62209=>"111101001",
  62210=>"000000000",
  62211=>"100100101",
  62212=>"000001011",
  62213=>"100010011",
  62214=>"111111111",
  62215=>"000100100",
  62216=>"011100011",
  62217=>"000000000",
  62218=>"011001001",
  62219=>"000100000",
  62220=>"000000000",
  62221=>"011011111",
  62222=>"111100000",
  62223=>"000000101",
  62224=>"000000111",
  62225=>"111111111",
  62226=>"111011001",
  62227=>"111111001",
  62228=>"000010111",
  62229=>"011011000",
  62230=>"100100110",
  62231=>"111111111",
  62232=>"000110100",
  62233=>"111111000",
  62234=>"100111110",
  62235=>"100000001",
  62236=>"100001011",
  62237=>"011000000",
  62238=>"111111000",
  62239=>"110000000",
  62240=>"011010110",
  62241=>"000000000",
  62242=>"111000000",
  62243=>"000100101",
  62244=>"100011010",
  62245=>"000111111",
  62246=>"000100000",
  62247=>"000000111",
  62248=>"000000011",
  62249=>"111111111",
  62250=>"010100101",
  62251=>"111000000",
  62252=>"100000000",
  62253=>"110110010",
  62254=>"000011111",
  62255=>"100111111",
  62256=>"000000000",
  62257=>"000000111",
  62258=>"000001111",
  62259=>"111111000",
  62260=>"000000000",
  62261=>"111110000",
  62262=>"111111111",
  62263=>"011000000",
  62264=>"000000100",
  62265=>"110100000",
  62266=>"000000000",
  62267=>"000000100",
  62268=>"111111111",
  62269=>"111111110",
  62270=>"111101111",
  62271=>"001000000",
  62272=>"000000000",
  62273=>"111111110",
  62274=>"001001000",
  62275=>"111111110",
  62276=>"000000000",
  62277=>"111111111",
  62278=>"111100111",
  62279=>"000000000",
  62280=>"000000010",
  62281=>"010000000",
  62282=>"101000110",
  62283=>"111111111",
  62284=>"100111111",
  62285=>"111111110",
  62286=>"000000011",
  62287=>"110000110",
  62288=>"111111100",
  62289=>"011011000",
  62290=>"111111110",
  62291=>"111111111",
  62292=>"000000111",
  62293=>"011011111",
  62294=>"111000000",
  62295=>"111000000",
  62296=>"000000000",
  62297=>"001011111",
  62298=>"000000000",
  62299=>"000001011",
  62300=>"000000000",
  62301=>"111111011",
  62302=>"100000110",
  62303=>"000100101",
  62304=>"111111100",
  62305=>"111001111",
  62306=>"000000001",
  62307=>"000100110",
  62308=>"001000000",
  62309=>"111111111",
  62310=>"110110100",
  62311=>"111111111",
  62312=>"111111111",
  62313=>"000000000",
  62314=>"000000000",
  62315=>"010011111",
  62316=>"111110100",
  62317=>"001111011",
  62318=>"001001111",
  62319=>"111111011",
  62320=>"110010010",
  62321=>"001001011",
  62322=>"000010010",
  62323=>"000100110",
  62324=>"111000000",
  62325=>"000000000",
  62326=>"110111111",
  62327=>"111111000",
  62328=>"111111111",
  62329=>"000100100",
  62330=>"111011111",
  62331=>"101101000",
  62332=>"110000000",
  62333=>"000000000",
  62334=>"111111111",
  62335=>"111111111",
  62336=>"001000000",
  62337=>"000000110",
  62338=>"111010000",
  62339=>"111111111",
  62340=>"111111011",
  62341=>"111001001",
  62342=>"000000111",
  62343=>"001110100",
  62344=>"111111111",
  62345=>"000000111",
  62346=>"000010110",
  62347=>"100000000",
  62348=>"000000000",
  62349=>"100001001",
  62350=>"111100000",
  62351=>"111111111",
  62352=>"000000001",
  62353=>"110111010",
  62354=>"100100100",
  62355=>"111111111",
  62356=>"111101001",
  62357=>"000110111",
  62358=>"111110000",
  62359=>"010011010",
  62360=>"100100000",
  62361=>"000000010",
  62362=>"100100110",
  62363=>"111110110",
  62364=>"111111111",
  62365=>"011011111",
  62366=>"110110111",
  62367=>"111111111",
  62368=>"000010100",
  62369=>"001011011",
  62370=>"000100111",
  62371=>"000111000",
  62372=>"101111111",
  62373=>"000010111",
  62374=>"111111111",
  62375=>"111111110",
  62376=>"011011111",
  62377=>"111111111",
  62378=>"000000001",
  62379=>"000000000",
  62380=>"000000000",
  62381=>"001000110",
  62382=>"000000011",
  62383=>"000110000",
  62384=>"000000000",
  62385=>"000111111",
  62386=>"111111111",
  62387=>"010011111",
  62388=>"000010000",
  62389=>"001100000",
  62390=>"111111111",
  62391=>"111110000",
  62392=>"000110110",
  62393=>"000111011",
  62394=>"111011000",
  62395=>"011001001",
  62396=>"000001001",
  62397=>"110100100",
  62398=>"111111111",
  62399=>"100101111",
  62400=>"000001100",
  62401=>"000000111",
  62402=>"001111111",
  62403=>"111011011",
  62404=>"110110000",
  62405=>"001000100",
  62406=>"000000111",
  62407=>"001101100",
  62408=>"111100011",
  62409=>"000000000",
  62410=>"000001000",
  62411=>"000000101",
  62412=>"000101000",
  62413=>"000000000",
  62414=>"111100110",
  62415=>"111111010",
  62416=>"110111111",
  62417=>"100000100",
  62418=>"100110111",
  62419=>"111111110",
  62420=>"000000001",
  62421=>"111111000",
  62422=>"000000000",
  62423=>"111111110",
  62424=>"000011110",
  62425=>"000001100",
  62426=>"100000010",
  62427=>"111111010",
  62428=>"011111011",
  62429=>"000000110",
  62430=>"000000000",
  62431=>"100101111",
  62432=>"111111000",
  62433=>"000000000",
  62434=>"000000000",
  62435=>"010010110",
  62436=>"110111111",
  62437=>"111111000",
  62438=>"111111101",
  62439=>"110110111",
  62440=>"111101100",
  62441=>"011011000",
  62442=>"100100110",
  62443=>"000110111",
  62444=>"001000000",
  62445=>"000000100",
  62446=>"111001000",
  62447=>"111111111",
  62448=>"100000001",
  62449=>"000001111",
  62450=>"000000000",
  62451=>"110111111",
  62452=>"111111100",
  62453=>"011001001",
  62454=>"001000000",
  62455=>"111111111",
  62456=>"111111100",
  62457=>"000110110",
  62458=>"111111000",
  62459=>"000000000",
  62460=>"011011011",
  62461=>"111111111",
  62462=>"000000011",
  62463=>"000111111",
  62464=>"000000000",
  62465=>"000111111",
  62466=>"111100100",
  62467=>"110111111",
  62468=>"111101000",
  62469=>"111011001",
  62470=>"000000000",
  62471=>"111111111",
  62472=>"111111111",
  62473=>"010010000",
  62474=>"110111111",
  62475=>"110111111",
  62476=>"000000000",
  62477=>"111001000",
  62478=>"000110001",
  62479=>"001000000",
  62480=>"111111111",
  62481=>"111111001",
  62482=>"000000000",
  62483=>"111001000",
  62484=>"000100111",
  62485=>"000000000",
  62486=>"000000000",
  62487=>"001001100",
  62488=>"001001011",
  62489=>"101111111",
  62490=>"000010000",
  62491=>"111011000",
  62492=>"000111011",
  62493=>"000000000",
  62494=>"111110000",
  62495=>"111111111",
  62496=>"000010010",
  62497=>"000001111",
  62498=>"111000000",
  62499=>"000100000",
  62500=>"110100111",
  62501=>"011111011",
  62502=>"010010000",
  62503=>"001111110",
  62504=>"000000000",
  62505=>"000000000",
  62506=>"111111111",
  62507=>"001111110",
  62508=>"101000011",
  62509=>"111110110",
  62510=>"000000100",
  62511=>"010110111",
  62512=>"111111111",
  62513=>"000000000",
  62514=>"001001011",
  62515=>"110110000",
  62516=>"111111110",
  62517=>"001000000",
  62518=>"100111000",
  62519=>"001100100",
  62520=>"000000111",
  62521=>"000000000",
  62522=>"000000000",
  62523=>"111111000",
  62524=>"111111111",
  62525=>"111000000",
  62526=>"100100100",
  62527=>"000000000",
  62528=>"000000000",
  62529=>"001000000",
  62530=>"111111111",
  62531=>"010110111",
  62532=>"011000000",
  62533=>"001011011",
  62534=>"000000000",
  62535=>"000000100",
  62536=>"101110100",
  62537=>"000000101",
  62538=>"110100110",
  62539=>"111100000",
  62540=>"000111111",
  62541=>"111111111",
  62542=>"000000000",
  62543=>"001000000",
  62544=>"111111000",
  62545=>"100110110",
  62546=>"111111000",
  62547=>"001100000",
  62548=>"111000000",
  62549=>"111000000",
  62550=>"000111000",
  62551=>"111111111",
  62552=>"111110110",
  62553=>"000000000",
  62554=>"000000000",
  62555=>"111111000",
  62556=>"000110111",
  62557=>"111101111",
  62558=>"000000111",
  62559=>"100100100",
  62560=>"000000001",
  62561=>"000011111",
  62562=>"111111111",
  62563=>"000000000",
  62564=>"110111110",
  62565=>"011001000",
  62566=>"001000111",
  62567=>"101000000",
  62568=>"111000101",
  62569=>"000111111",
  62570=>"001111111",
  62571=>"001001000",
  62572=>"001011110",
  62573=>"110000000",
  62574=>"000110011",
  62575=>"111111111",
  62576=>"001011111",
  62577=>"111111110",
  62578=>"001000001",
  62579=>"001001111",
  62580=>"111000000",
  62581=>"000000011",
  62582=>"010010010",
  62583=>"000000000",
  62584=>"000111111",
  62585=>"000110000",
  62586=>"000000000",
  62587=>"100000000",
  62588=>"011111110",
  62589=>"000000000",
  62590=>"000000000",
  62591=>"000100000",
  62592=>"000000000",
  62593=>"000111110",
  62594=>"110110111",
  62595=>"111100100",
  62596=>"111111111",
  62597=>"000100101",
  62598=>"110110110",
  62599=>"000000011",
  62600=>"000001000",
  62601=>"001000100",
  62602=>"111010000",
  62603=>"000001001",
  62604=>"111100001",
  62605=>"001000000",
  62606=>"110000000",
  62607=>"111111111",
  62608=>"000000000",
  62609=>"111101100",
  62610=>"111000000",
  62611=>"010111001",
  62612=>"000000001",
  62613=>"111111111",
  62614=>"001001011",
  62615=>"110100110",
  62616=>"000001111",
  62617=>"100111111",
  62618=>"110000000",
  62619=>"001000000",
  62620=>"111110100",
  62621=>"000000001",
  62622=>"111111111",
  62623=>"000000000",
  62624=>"000111111",
  62625=>"000000000",
  62626=>"110111111",
  62627=>"101101101",
  62628=>"000000001",
  62629=>"111111111",
  62630=>"001111111",
  62631=>"111011111",
  62632=>"000000011",
  62633=>"000000001",
  62634=>"111000000",
  62635=>"111011100",
  62636=>"000000011",
  62637=>"100110010",
  62638=>"011111111",
  62639=>"110100110",
  62640=>"000000100",
  62641=>"111111111",
  62642=>"111111111",
  62643=>"000000111",
  62644=>"111111111",
  62645=>"111111111",
  62646=>"111101011",
  62647=>"000111101",
  62648=>"000010010",
  62649=>"111111111",
  62650=>"000000111",
  62651=>"011111110",
  62652=>"000000000",
  62653=>"000000000",
  62654=>"111111111",
  62655=>"111111111",
  62656=>"000010011",
  62657=>"111110000",
  62658=>"000000000",
  62659=>"111111111",
  62660=>"111111110",
  62661=>"000111111",
  62662=>"011111011",
  62663=>"001000001",
  62664=>"111111111",
  62665=>"001111111",
  62666=>"111100011",
  62667=>"110100001",
  62668=>"100100001",
  62669=>"100000000",
  62670=>"110111110",
  62671=>"000011000",
  62672=>"000111111",
  62673=>"000111010",
  62674=>"000111011",
  62675=>"000000000",
  62676=>"000000000",
  62677=>"000100001",
  62678=>"000000000",
  62679=>"100110010",
  62680=>"111111011",
  62681=>"100001000",
  62682=>"011111111",
  62683=>"111111111",
  62684=>"001000001",
  62685=>"100111111",
  62686=>"111000010",
  62687=>"010110111",
  62688=>"010000000",
  62689=>"000000000",
  62690=>"111111111",
  62691=>"001000000",
  62692=>"000000100",
  62693=>"111111010",
  62694=>"000111111",
  62695=>"110110101",
  62696=>"100000110",
  62697=>"000001111",
  62698=>"111111111",
  62699=>"000000000",
  62700=>"001011001",
  62701=>"001000110",
  62702=>"111100000",
  62703=>"000000000",
  62704=>"011001001",
  62705=>"000000000",
  62706=>"000000111",
  62707=>"000100111",
  62708=>"111111000",
  62709=>"000001011",
  62710=>"011111000",
  62711=>"100100000",
  62712=>"110111111",
  62713=>"011111111",
  62714=>"111111000",
  62715=>"101110111",
  62716=>"100100110",
  62717=>"000000001",
  62718=>"111001001",
  62719=>"110000000",
  62720=>"000000001",
  62721=>"011000000",
  62722=>"000000100",
  62723=>"111111001",
  62724=>"111010000",
  62725=>"000000000",
  62726=>"111111111",
  62727=>"000111100",
  62728=>"101111011",
  62729=>"111111111",
  62730=>"000000000",
  62731=>"100000111",
  62732=>"101101001",
  62733=>"111100100",
  62734=>"100111110",
  62735=>"110110000",
  62736=>"011011001",
  62737=>"010111011",
  62738=>"100000101",
  62739=>"111101000",
  62740=>"100000000",
  62741=>"111111000",
  62742=>"111111011",
  62743=>"001001000",
  62744=>"111111110",
  62745=>"101110000",
  62746=>"100001001",
  62747=>"100000001",
  62748=>"000111111",
  62749=>"000000000",
  62750=>"000000000",
  62751=>"011011011",
  62752=>"000000000",
  62753=>"111111000",
  62754=>"000000110",
  62755=>"111111111",
  62756=>"011111011",
  62757=>"001011000",
  62758=>"111111111",
  62759=>"100110111",
  62760=>"001001001",
  62761=>"011111111",
  62762=>"100100111",
  62763=>"111110110",
  62764=>"001000111",
  62765=>"000000000",
  62766=>"000000000",
  62767=>"000000000",
  62768=>"111111111",
  62769=>"111111110",
  62770=>"111111111",
  62771=>"111111110",
  62772=>"111111111",
  62773=>"001001001",
  62774=>"111111000",
  62775=>"001000100",
  62776=>"000010100",
  62777=>"111010111",
  62778=>"000000000",
  62779=>"000000000",
  62780=>"000000000",
  62781=>"100110111",
  62782=>"111011011",
  62783=>"110111111",
  62784=>"000000010",
  62785=>"111111111",
  62786=>"111111111",
  62787=>"000000000",
  62788=>"001000000",
  62789=>"111001000",
  62790=>"000000000",
  62791=>"000000001",
  62792=>"101000000",
  62793=>"111011000",
  62794=>"000011111",
  62795=>"001111111",
  62796=>"010000000",
  62797=>"000000000",
  62798=>"000000100",
  62799=>"000000110",
  62800=>"111110110",
  62801=>"000111111",
  62802=>"001001011",
  62803=>"101001001",
  62804=>"111000000",
  62805=>"000110110",
  62806=>"000001111",
  62807=>"000111111",
  62808=>"111010000",
  62809=>"111000000",
  62810=>"110010111",
  62811=>"001101001",
  62812=>"000000000",
  62813=>"000000001",
  62814=>"000000000",
  62815=>"011111111",
  62816=>"000000000",
  62817=>"111000110",
  62818=>"111111101",
  62819=>"000000100",
  62820=>"111111110",
  62821=>"000000000",
  62822=>"000000111",
  62823=>"101111001",
  62824=>"100111111",
  62825=>"111110000",
  62826=>"001000001",
  62827=>"010110100",
  62828=>"001011001",
  62829=>"000011111",
  62830=>"000110111",
  62831=>"000000011",
  62832=>"001001101",
  62833=>"001000000",
  62834=>"111101111",
  62835=>"111011011",
  62836=>"111110011",
  62837=>"000000000",
  62838=>"000010111",
  62839=>"111111111",
  62840=>"000000000",
  62841=>"111111010",
  62842=>"000100100",
  62843=>"000000001",
  62844=>"010110000",
  62845=>"111111001",
  62846=>"111111001",
  62847=>"000000000",
  62848=>"110110110",
  62849=>"111001011",
  62850=>"000000000",
  62851=>"000000010",
  62852=>"100111001",
  62853=>"000000000",
  62854=>"011111111",
  62855=>"111001110",
  62856=>"000000000",
  62857=>"111011000",
  62858=>"000000001",
  62859=>"111111000",
  62860=>"111101000",
  62861=>"111111111",
  62862=>"110100111",
  62863=>"000000111",
  62864=>"111100000",
  62865=>"111000000",
  62866=>"101111111",
  62867=>"000000000",
  62868=>"000000110",
  62869=>"000011110",
  62870=>"100000000",
  62871=>"011110010",
  62872=>"000000010",
  62873=>"001011011",
  62874=>"110110000",
  62875=>"000000011",
  62876=>"011000001",
  62877=>"110110111",
  62878=>"101000000",
  62879=>"000111111",
  62880=>"111111111",
  62881=>"001011011",
  62882=>"110111111",
  62883=>"111000000",
  62884=>"110000001",
  62885=>"111111000",
  62886=>"101000110",
  62887=>"111000000",
  62888=>"010000000",
  62889=>"110000000",
  62890=>"011010011",
  62891=>"000000100",
  62892=>"001001000",
  62893=>"000000111",
  62894=>"000000000",
  62895=>"001101001",
  62896=>"000000111",
  62897=>"000100110",
  62898=>"001000000",
  62899=>"110010000",
  62900=>"000000000",
  62901=>"110110000",
  62902=>"111111000",
  62903=>"111000000",
  62904=>"000000000",
  62905=>"111111111",
  62906=>"111111000",
  62907=>"111100111",
  62908=>"111101110",
  62909=>"110111111",
  62910=>"000000000",
  62911=>"011001000",
  62912=>"000000111",
  62913=>"110110000",
  62914=>"111111111",
  62915=>"000000000",
  62916=>"000000110",
  62917=>"000100000",
  62918=>"011111000",
  62919=>"101000000",
  62920=>"000000101",
  62921=>"101111111",
  62922=>"100001001",
  62923=>"000000000",
  62924=>"010110110",
  62925=>"111111000",
  62926=>"000000010",
  62927=>"001111111",
  62928=>"111111111",
  62929=>"001000100",
  62930=>"111111000",
  62931=>"000111110",
  62932=>"111111011",
  62933=>"111111111",
  62934=>"000000111",
  62935=>"000000000",
  62936=>"000000111",
  62937=>"111000100",
  62938=>"101111110",
  62939=>"000000000",
  62940=>"111111111",
  62941=>"111111000",
  62942=>"111111110",
  62943=>"001001111",
  62944=>"000000100",
  62945=>"101111111",
  62946=>"111111111",
  62947=>"111110111",
  62948=>"101111110",
  62949=>"000000000",
  62950=>"000111000",
  62951=>"000000000",
  62952=>"110110010",
  62953=>"111111000",
  62954=>"000000111",
  62955=>"111111100",
  62956=>"000111111",
  62957=>"011111101",
  62958=>"001001011",
  62959=>"111001001",
  62960=>"000000001",
  62961=>"011011111",
  62962=>"000000001",
  62963=>"000000111",
  62964=>"111110000",
  62965=>"111101000",
  62966=>"111111011",
  62967=>"010110111",
  62968=>"100100110",
  62969=>"000011101",
  62970=>"111111111",
  62971=>"000000000",
  62972=>"000000000",
  62973=>"111101111",
  62974=>"000000000",
  62975=>"000000000",
  62976=>"111111111",
  62977=>"011000000",
  62978=>"000001000",
  62979=>"000000000",
  62980=>"001000000",
  62981=>"110111111",
  62982=>"101001001",
  62983=>"000000000",
  62984=>"111110100",
  62985=>"000000000",
  62986=>"111111111",
  62987=>"101100111",
  62988=>"111011011",
  62989=>"110110100",
  62990=>"111110111",
  62991=>"111100101",
  62992=>"000000011",
  62993=>"111000000",
  62994=>"101000000",
  62995=>"000001000",
  62996=>"111000000",
  62997=>"000000111",
  62998=>"111100000",
  62999=>"110110111",
  63000=>"001000000",
  63001=>"111111111",
  63002=>"000000111",
  63003=>"001000100",
  63004=>"000000000",
  63005=>"000000000",
  63006=>"111111111",
  63007=>"000110000",
  63008=>"011010000",
  63009=>"111111111",
  63010=>"011011011",
  63011=>"000000000",
  63012=>"111111111",
  63013=>"111111111",
  63014=>"000111110",
  63015=>"000001101",
  63016=>"111111111",
  63017=>"010111110",
  63018=>"011101111",
  63019=>"111111111",
  63020=>"111000111",
  63021=>"000000000",
  63022=>"001101111",
  63023=>"111111111",
  63024=>"001000000",
  63025=>"001000000",
  63026=>"100111111",
  63027=>"000000000",
  63028=>"111111000",
  63029=>"000000001",
  63030=>"111111111",
  63031=>"111111111",
  63032=>"111111111",
  63033=>"100000000",
  63034=>"111001111",
  63035=>"000110111",
  63036=>"000000000",
  63037=>"000000000",
  63038=>"101111000",
  63039=>"000000111",
  63040=>"111110100",
  63041=>"110110110",
  63042=>"111111111",
  63043=>"100010011",
  63044=>"010000101",
  63045=>"000000000",
  63046=>"110111111",
  63047=>"000000000",
  63048=>"000100000",
  63049=>"111111011",
  63050=>"000001011",
  63051=>"000000000",
  63052=>"111111000",
  63053=>"111011001",
  63054=>"111111010",
  63055=>"000000100",
  63056=>"000000000",
  63057=>"000110011",
  63058=>"011010000",
  63059=>"011110111",
  63060=>"111001001",
  63061=>"111111111",
  63062=>"000000000",
  63063=>"000000000",
  63064=>"111101111",
  63065=>"111111111",
  63066=>"011111111",
  63067=>"111110110",
  63068=>"111111101",
  63069=>"111111111",
  63070=>"010001000",
  63071=>"000111111",
  63072=>"001111111",
  63073=>"100000000",
  63074=>"111011000",
  63075=>"100000100",
  63076=>"111111111",
  63077=>"001111011",
  63078=>"000011000",
  63079=>"000110111",
  63080=>"111111111",
  63081=>"000111111",
  63082=>"111111111",
  63083=>"001001001",
  63084=>"110110110",
  63085=>"000000000",
  63086=>"000011000",
  63087=>"111111100",
  63088=>"111111110",
  63089=>"000000111",
  63090=>"000000000",
  63091=>"001001011",
  63092=>"001000000",
  63093=>"111000000",
  63094=>"000000000",
  63095=>"111111011",
  63096=>"000111011",
  63097=>"111111111",
  63098=>"111111001",
  63099=>"111111111",
  63100=>"111111111",
  63101=>"111001111",
  63102=>"111111010",
  63103=>"000000000",
  63104=>"111011011",
  63105=>"100111001",
  63106=>"111111110",
  63107=>"011001001",
  63108=>"000000000",
  63109=>"111111001",
  63110=>"001001001",
  63111=>"111111111",
  63112=>"001001000",
  63113=>"000000000",
  63114=>"010111111",
  63115=>"000000100",
  63116=>"111100111",
  63117=>"010000000",
  63118=>"000000000",
  63119=>"011000000",
  63120=>"000000000",
  63121=>"000000010",
  63122=>"000010110",
  63123=>"000000000",
  63124=>"001000000",
  63125=>"000000000",
  63126=>"111111011",
  63127=>"000000001",
  63128=>"110110110",
  63129=>"000000000",
  63130=>"111111111",
  63131=>"000000000",
  63132=>"111110000",
  63133=>"001111111",
  63134=>"111111111",
  63135=>"000000000",
  63136=>"111111110",
  63137=>"111111111",
  63138=>"111111111",
  63139=>"000110111",
  63140=>"011111111",
  63141=>"011111111",
  63142=>"111100100",
  63143=>"011001011",
  63144=>"111111111",
  63145=>"000000000",
  63146=>"111110110",
  63147=>"111111111",
  63148=>"000000000",
  63149=>"000000100",
  63150=>"000000111",
  63151=>"000000000",
  63152=>"111111111",
  63153=>"011011011",
  63154=>"100000000",
  63155=>"111100000",
  63156=>"001000011",
  63157=>"111111111",
  63158=>"101000101",
  63159=>"111001000",
  63160=>"000110110",
  63161=>"000000110",
  63162=>"000001111",
  63163=>"100100000",
  63164=>"000110111",
  63165=>"000000000",
  63166=>"111111110",
  63167=>"000000100",
  63168=>"000000000",
  63169=>"001111011",
  63170=>"000001001",
  63171=>"111000000",
  63172=>"111111111",
  63173=>"000000000",
  63174=>"000000000",
  63175=>"110000000",
  63176=>"000000110",
  63177=>"111111111",
  63178=>"010111000",
  63179=>"111000000",
  63180=>"110011111",
  63181=>"111110111",
  63182=>"111111111",
  63183=>"111101101",
  63184=>"000000100",
  63185=>"111111111",
  63186=>"111100111",
  63187=>"111111111",
  63188=>"000000000",
  63189=>"000000000",
  63190=>"000011111",
  63191=>"000110110",
  63192=>"111111111",
  63193=>"111111111",
  63194=>"000000000",
  63195=>"101000001",
  63196=>"001001001",
  63197=>"111111111",
  63198=>"111111111",
  63199=>"001000000",
  63200=>"111100100",
  63201=>"000000000",
  63202=>"000000000",
  63203=>"111111011",
  63204=>"101100001",
  63205=>"100110110",
  63206=>"111110111",
  63207=>"111111111",
  63208=>"000010000",
  63209=>"001001000",
  63210=>"011000000",
  63211=>"111111101",
  63212=>"000000001",
  63213=>"111111111",
  63214=>"000000000",
  63215=>"000000000",
  63216=>"000000000",
  63217=>"000000000",
  63218=>"111111111",
  63219=>"000000000",
  63220=>"000000000",
  63221=>"000000010",
  63222=>"000000001",
  63223=>"001000111",
  63224=>"000110000",
  63225=>"111111111",
  63226=>"000100111",
  63227=>"111111110",
  63228=>"101100100",
  63229=>"011111111",
  63230=>"111111011",
  63231=>"001011001",
  63232=>"111111111",
  63233=>"011011001",
  63234=>"000100000",
  63235=>"111111000",
  63236=>"000000000",
  63237=>"010011001",
  63238=>"000000000",
  63239=>"001001001",
  63240=>"000000000",
  63241=>"000000000",
  63242=>"000000100",
  63243=>"111111111",
  63244=>"000000110",
  63245=>"000101111",
  63246=>"111001100",
  63247=>"000011100",
  63248=>"100111111",
  63249=>"000000000",
  63250=>"000000000",
  63251=>"001011100",
  63252=>"011000000",
  63253=>"111110111",
  63254=>"111000000",
  63255=>"111111100",
  63256=>"110011111",
  63257=>"000001111",
  63258=>"111100000",
  63259=>"111100000",
  63260=>"011001001",
  63261=>"011100001",
  63262=>"111111111",
  63263=>"000011111",
  63264=>"001111111",
  63265=>"101111111",
  63266=>"000000011",
  63267=>"000000000",
  63268=>"001011111",
  63269=>"000000000",
  63270=>"111110000",
  63271=>"111111011",
  63272=>"001000000",
  63273=>"000000000",
  63274=>"111000000",
  63275=>"111101100",
  63276=>"000000000",
  63277=>"000101110",
  63278=>"000000111",
  63279=>"100100000",
  63280=>"000000110",
  63281=>"000000000",
  63282=>"001001001",
  63283=>"111111111",
  63284=>"100000100",
  63285=>"001111111",
  63286=>"000010010",
  63287=>"111111111",
  63288=>"000000000",
  63289=>"000110111",
  63290=>"111000000",
  63291=>"000000000",
  63292=>"000111001",
  63293=>"100000111",
  63294=>"011011000",
  63295=>"111110101",
  63296=>"000000000",
  63297=>"000000000",
  63298=>"011000110",
  63299=>"010000000",
  63300=>"000000000",
  63301=>"110111010",
  63302=>"101111111",
  63303=>"000000000",
  63304=>"000000010",
  63305=>"111000100",
  63306=>"111111000",
  63307=>"011011111",
  63308=>"111101111",
  63309=>"000111111",
  63310=>"000000001",
  63311=>"110110100",
  63312=>"100101111",
  63313=>"111111111",
  63314=>"111111111",
  63315=>"111111111",
  63316=>"111100110",
  63317=>"001011011",
  63318=>"111111111",
  63319=>"111111111",
  63320=>"000000000",
  63321=>"000000000",
  63322=>"000000001",
  63323=>"100000011",
  63324=>"111101100",
  63325=>"100000000",
  63326=>"001001000",
  63327=>"011011111",
  63328=>"100100000",
  63329=>"000000000",
  63330=>"111110010",
  63331=>"111000000",
  63332=>"001001001",
  63333=>"000010010",
  63334=>"000000000",
  63335=>"001000000",
  63336=>"110110110",
  63337=>"000000000",
  63338=>"111111100",
  63339=>"111111111",
  63340=>"000000000",
  63341=>"000000000",
  63342=>"000000000",
  63343=>"011111011",
  63344=>"000000000",
  63345=>"011000010",
  63346=>"000111011",
  63347=>"111100110",
  63348=>"111111111",
  63349=>"111111101",
  63350=>"000000110",
  63351=>"010000000",
  63352=>"000000000",
  63353=>"000000000",
  63354=>"010111111",
  63355=>"111100100",
  63356=>"000111111",
  63357=>"111000000",
  63358=>"110110110",
  63359=>"111111111",
  63360=>"111111111",
  63361=>"110000000",
  63362=>"111000000",
  63363=>"010010000",
  63364=>"100100000",
  63365=>"111111000",
  63366=>"111111111",
  63367=>"111011111",
  63368=>"000010000",
  63369=>"001000000",
  63370=>"000100100",
  63371=>"111111111",
  63372=>"001111111",
  63373=>"000000010",
  63374=>"010111100",
  63375=>"000000000",
  63376=>"111111000",
  63377=>"001001001",
  63378=>"000100000",
  63379=>"001011000",
  63380=>"111101000",
  63381=>"011000000",
  63382=>"111101111",
  63383=>"000001000",
  63384=>"000000110",
  63385=>"111001111",
  63386=>"000000100",
  63387=>"000000010",
  63388=>"100111100",
  63389=>"000100111",
  63390=>"000011001",
  63391=>"111111000",
  63392=>"111111111",
  63393=>"000000000",
  63394=>"111011111",
  63395=>"110111011",
  63396=>"010111111",
  63397=>"111111100",
  63398=>"000000000",
  63399=>"000100111",
  63400=>"111010000",
  63401=>"110111111",
  63402=>"011111111",
  63403=>"010010000",
  63404=>"000000000",
  63405=>"100110110",
  63406=>"110010000",
  63407=>"000110010",
  63408=>"110111111",
  63409=>"111111111",
  63410=>"111111111",
  63411=>"100000000",
  63412=>"100001111",
  63413=>"000000000",
  63414=>"110110110",
  63415=>"111111111",
  63416=>"111111111",
  63417=>"111011111",
  63418=>"111011000",
  63419=>"111111111",
  63420=>"000111111",
  63421=>"111111011",
  63422=>"000000010",
  63423=>"010000000",
  63424=>"000110111",
  63425=>"000100100",
  63426=>"111111000",
  63427=>"111011000",
  63428=>"010000000",
  63429=>"000010010",
  63430=>"000000010",
  63431=>"100101000",
  63432=>"000000000",
  63433=>"110110111",
  63434=>"111111111",
  63435=>"000000000",
  63436=>"000010011",
  63437=>"000000000",
  63438=>"100000000",
  63439=>"000100110",
  63440=>"000000000",
  63441=>"110111111",
  63442=>"111111111",
  63443=>"011001111",
  63444=>"111111111",
  63445=>"110000000",
  63446=>"010110111",
  63447=>"100001000",
  63448=>"000001001",
  63449=>"101110000",
  63450=>"000000000",
  63451=>"100000100",
  63452=>"110100111",
  63453=>"001000001",
  63454=>"000000000",
  63455=>"001000000",
  63456=>"100000000",
  63457=>"110111111",
  63458=>"000001000",
  63459=>"111111111",
  63460=>"110111010",
  63461=>"111111111",
  63462=>"001011011",
  63463=>"101111101",
  63464=>"111111111",
  63465=>"001011011",
  63466=>"110000000",
  63467=>"111111111",
  63468=>"010000111",
  63469=>"000000000",
  63470=>"000000000",
  63471=>"000000000",
  63472=>"000001001",
  63473=>"111111000",
  63474=>"111111110",
  63475=>"000000000",
  63476=>"011111111",
  63477=>"111111011",
  63478=>"111111111",
  63479=>"100000000",
  63480=>"111110110",
  63481=>"100110000",
  63482=>"011000000",
  63483=>"000110111",
  63484=>"111111111",
  63485=>"011110100",
  63486=>"111000000",
  63487=>"111111111",
  63488=>"100000000",
  63489=>"000000000",
  63490=>"000000000",
  63491=>"111111100",
  63492=>"000001000",
  63493=>"110100100",
  63494=>"001001001",
  63495=>"111111111",
  63496=>"011000000",
  63497=>"000000111",
  63498=>"110010011",
  63499=>"001100101",
  63500=>"100110110",
  63501=>"111111100",
  63502=>"100000100",
  63503=>"000000000",
  63504=>"001000000",
  63505=>"111100100",
  63506=>"111000000",
  63507=>"110110100",
  63508=>"000000111",
  63509=>"101010110",
  63510=>"000000011",
  63511=>"000100101",
  63512=>"100101001",
  63513=>"010011011",
  63514=>"111111000",
  63515=>"110100100",
  63516=>"011000000",
  63517=>"111111111",
  63518=>"111110110",
  63519=>"000000000",
  63520=>"000000000",
  63521=>"010000000",
  63522=>"111111111",
  63523=>"110100111",
  63524=>"100000000",
  63525=>"101000111",
  63526=>"101000000",
  63527=>"011000000",
  63528=>"111111011",
  63529=>"110111000",
  63530=>"000000000",
  63531=>"111111111",
  63532=>"000111111",
  63533=>"111100100",
  63534=>"011011001",
  63535=>"000100111",
  63536=>"000000000",
  63537=>"001001001",
  63538=>"110110110",
  63539=>"000110001",
  63540=>"011111111",
  63541=>"000000100",
  63542=>"100001001",
  63543=>"110110000",
  63544=>"001011111",
  63545=>"111111111",
  63546=>"101111101",
  63547=>"111111000",
  63548=>"111110111",
  63549=>"000000101",
  63550=>"010110100",
  63551=>"100000011",
  63552=>"001000000",
  63553=>"111011011",
  63554=>"111111100",
  63555=>"100110110",
  63556=>"000100000",
  63557=>"100000000",
  63558=>"011111111",
  63559=>"000000000",
  63560=>"011011010",
  63561=>"000000111",
  63562=>"000111110",
  63563=>"111011011",
  63564=>"110111111",
  63565=>"001001101",
  63566=>"000000000",
  63567=>"000000000",
  63568=>"000110101",
  63569=>"011111111",
  63570=>"111111111",
  63571=>"110110100",
  63572=>"111010110",
  63573=>"010000000",
  63574=>"000100110",
  63575=>"111100111",
  63576=>"000000000",
  63577=>"111101111",
  63578=>"011001110",
  63579=>"000000000",
  63580=>"110110111",
  63581=>"111111111",
  63582=>"000110111",
  63583=>"000000000",
  63584=>"111111001",
  63585=>"000000000",
  63586=>"000000000",
  63587=>"000111111",
  63588=>"111000110",
  63589=>"000000111",
  63590=>"100111111",
  63591=>"101000000",
  63592=>"000000111",
  63593=>"111100000",
  63594=>"000111001",
  63595=>"111111111",
  63596=>"000110010",
  63597=>"000000000",
  63598=>"111111111",
  63599=>"011001111",
  63600=>"001011111",
  63601=>"001110111",
  63602=>"001100111",
  63603=>"011011000",
  63604=>"111111111",
  63605=>"111111000",
  63606=>"110111000",
  63607=>"000000000",
  63608=>"000000001",
  63609=>"101001001",
  63610=>"110110110",
  63611=>"000000001",
  63612=>"100000000",
  63613=>"110110111",
  63614=>"111100000",
  63615=>"111111000",
  63616=>"111111010",
  63617=>"000000000",
  63618=>"110111111",
  63619=>"111011011",
  63620=>"111111111",
  63621=>"111000000",
  63622=>"100100110",
  63623=>"111000000",
  63624=>"011000000",
  63625=>"000000000",
  63626=>"101000111",
  63627=>"111111111",
  63628=>"111111111",
  63629=>"000000000",
  63630=>"100000111",
  63631=>"000000001",
  63632=>"111111111",
  63633=>"000000000",
  63634=>"000000000",
  63635=>"000000001",
  63636=>"111111110",
  63637=>"111111111",
  63638=>"111000000",
  63639=>"000001001",
  63640=>"111111111",
  63641=>"111111111",
  63642=>"110011111",
  63643=>"000000000",
  63644=>"000011011",
  63645=>"001001000",
  63646=>"000100100",
  63647=>"000101111",
  63648=>"100000101",
  63649=>"111000000",
  63650=>"010000000",
  63651=>"000000111",
  63652=>"111000000",
  63653=>"010001000",
  63654=>"111111000",
  63655=>"000111111",
  63656=>"111111111",
  63657=>"000000000",
  63658=>"100000111",
  63659=>"000000000",
  63660=>"111100110",
  63661=>"000000011",
  63662=>"111111111",
  63663=>"000011111",
  63664=>"111111010",
  63665=>"000000000",
  63666=>"010011000",
  63667=>"111111010",
  63668=>"000000000",
  63669=>"001111011",
  63670=>"000000000",
  63671=>"111001000",
  63672=>"001011111",
  63673=>"000000111",
  63674=>"111001000",
  63675=>"001000001",
  63676=>"110111011",
  63677=>"011000000",
  63678=>"111111111",
  63679=>"111111111",
  63680=>"111111001",
  63681=>"001000000",
  63682=>"001000111",
  63683=>"111111111",
  63684=>"111111111",
  63685=>"000001000",
  63686=>"111001000",
  63687=>"000000000",
  63688=>"001001000",
  63689=>"011111111",
  63690=>"110000000",
  63691=>"000000001",
  63692=>"011000011",
  63693=>"000111111",
  63694=>"111011000",
  63695=>"000100000",
  63696=>"000000000",
  63697=>"111111110",
  63698=>"111111111",
  63699=>"111110000",
  63700=>"000000000",
  63701=>"100110111",
  63702=>"111010111",
  63703=>"000100110",
  63704=>"111111000",
  63705=>"111011011",
  63706=>"000000000",
  63707=>"000010111",
  63708=>"110111111",
  63709=>"111110010",
  63710=>"111111100",
  63711=>"111111110",
  63712=>"001000001",
  63713=>"111000000",
  63714=>"111001010",
  63715=>"100000000",
  63716=>"100000001",
  63717=>"001001000",
  63718=>"111111111",
  63719=>"000000000",
  63720=>"000000111",
  63721=>"111111010",
  63722=>"111001000",
  63723=>"011001111",
  63724=>"011011000",
  63725=>"001111111",
  63726=>"110111101",
  63727=>"111111100",
  63728=>"100111111",
  63729=>"000000000",
  63730=>"111111111",
  63731=>"110110000",
  63732=>"101000000",
  63733=>"000000000",
  63734=>"000001000",
  63735=>"111111111",
  63736=>"000000000",
  63737=>"110111111",
  63738=>"111111110",
  63739=>"000000000",
  63740=>"011001001",
  63741=>"010011001",
  63742=>"111111111",
  63743=>"000000000",
  63744=>"000100111",
  63745=>"110110110",
  63746=>"111111111",
  63747=>"111111111",
  63748=>"000000000",
  63749=>"100000100",
  63750=>"011000000",
  63751=>"000000010",
  63752=>"000101111",
  63753=>"001000000",
  63754=>"111111111",
  63755=>"111111111",
  63756=>"111001111",
  63757=>"000000000",
  63758=>"111001000",
  63759=>"000000000",
  63760=>"100111111",
  63761=>"001111111",
  63762=>"000000000",
  63763=>"000011011",
  63764=>"100000000",
  63765=>"111110110",
  63766=>"011111010",
  63767=>"000000111",
  63768=>"100110110",
  63769=>"000000000",
  63770=>"011111111",
  63771=>"111000000",
  63772=>"110110111",
  63773=>"111111110",
  63774=>"111101111",
  63775=>"111011000",
  63776=>"101111101",
  63777=>"000001000",
  63778=>"000000101",
  63779=>"111000011",
  63780=>"111111111",
  63781=>"000000000",
  63782=>"111111000",
  63783=>"000000000",
  63784=>"110000000",
  63785=>"000000000",
  63786=>"111111111",
  63787=>"100111111",
  63788=>"000000000",
  63789=>"011010000",
  63790=>"000000010",
  63791=>"000001000",
  63792=>"100101111",
  63793=>"000000000",
  63794=>"000000111",
  63795=>"000100111",
  63796=>"000010010",
  63797=>"111110100",
  63798=>"111111111",
  63799=>"111111101",
  63800=>"000000000",
  63801=>"000000001",
  63802=>"101101111",
  63803=>"011111111",
  63804=>"111111111",
  63805=>"100110000",
  63806=>"000000000",
  63807=>"000100100",
  63808=>"100000000",
  63809=>"111111111",
  63810=>"000000000",
  63811=>"000000000",
  63812=>"000001000",
  63813=>"110111111",
  63814=>"000000000",
  63815=>"001101100",
  63816=>"000110011",
  63817=>"110110000",
  63818=>"000100111",
  63819=>"000100000",
  63820=>"000000000",
  63821=>"111111000",
  63822=>"000001011",
  63823=>"000100000",
  63824=>"111111001",
  63825=>"111111000",
  63826=>"100100000",
  63827=>"111011001",
  63828=>"000000000",
  63829=>"011001011",
  63830=>"111111000",
  63831=>"101001101",
  63832=>"110000111",
  63833=>"010110010",
  63834=>"111111001",
  63835=>"000000000",
  63836=>"111111110",
  63837=>"111111111",
  63838=>"000000000",
  63839=>"001011111",
  63840=>"000000001",
  63841=>"111001000",
  63842=>"011111111",
  63843=>"011011111",
  63844=>"111111111",
  63845=>"000000000",
  63846=>"111111111",
  63847=>"110111001",
  63848=>"001001001",
  63849=>"111111111",
  63850=>"111111111",
  63851=>"000111000",
  63852=>"000100110",
  63853=>"111111111",
  63854=>"000000001",
  63855=>"000000001",
  63856=>"111111111",
  63857=>"111111011",
  63858=>"111111111",
  63859=>"111111011",
  63860=>"000001111",
  63861=>"010000000",
  63862=>"111111111",
  63863=>"000000000",
  63864=>"000111111",
  63865=>"111111111",
  63866=>"000000000",
  63867=>"000000000",
  63868=>"000111111",
  63869=>"111111111",
  63870=>"110111111",
  63871=>"101101111",
  63872=>"100000000",
  63873=>"111101111",
  63874=>"000000000",
  63875=>"111010000",
  63876=>"001111111",
  63877=>"000000000",
  63878=>"000000000",
  63879=>"000110110",
  63880=>"000000000",
  63881=>"011111101",
  63882=>"000000000",
  63883=>"000001000",
  63884=>"101111111",
  63885=>"000000010",
  63886=>"111111111",
  63887=>"011111111",
  63888=>"010111111",
  63889=>"010111111",
  63890=>"111111111",
  63891=>"010111111",
  63892=>"000000000",
  63893=>"011011000",
  63894=>"100100111",
  63895=>"011011000",
  63896=>"000000110",
  63897=>"000000000",
  63898=>"000000000",
  63899=>"011010011",
  63900=>"000100001",
  63901=>"000000000",
  63902=>"101101101",
  63903=>"101111111",
  63904=>"111001001",
  63905=>"000100000",
  63906=>"000110111",
  63907=>"111111000",
  63908=>"110110110",
  63909=>"010000000",
  63910=>"000011111",
  63911=>"000000000",
  63912=>"000000010",
  63913=>"000001011",
  63914=>"000110111",
  63915=>"011001000",
  63916=>"000000000",
  63917=>"111110000",
  63918=>"000001111",
  63919=>"001001011",
  63920=>"111100011",
  63921=>"000000000",
  63922=>"101100111",
  63923=>"000000011",
  63924=>"000000000",
  63925=>"010000001",
  63926=>"110111111",
  63927=>"000011111",
  63928=>"000000100",
  63929=>"110011001",
  63930=>"010010110",
  63931=>"100000000",
  63932=>"000000000",
  63933=>"111111111",
  63934=>"101100100",
  63935=>"100101101",
  63936=>"111111011",
  63937=>"000000000",
  63938=>"000000000",
  63939=>"000001001",
  63940=>"111010011",
  63941=>"110110100",
  63942=>"111111111",
  63943=>"000000000",
  63944=>"100100110",
  63945=>"000011011",
  63946=>"000111011",
  63947=>"000000000",
  63948=>"000000000",
  63949=>"011111011",
  63950=>"010110111",
  63951=>"110000111",
  63952=>"101101110",
  63953=>"111111000",
  63954=>"111111000",
  63955=>"000111111",
  63956=>"100010011",
  63957=>"100100101",
  63958=>"000000000",
  63959=>"011011011",
  63960=>"001101001",
  63961=>"110111111",
  63962=>"111111111",
  63963=>"000000010",
  63964=>"111011011",
  63965=>"101111000",
  63966=>"111111110",
  63967=>"111111111",
  63968=>"111111000",
  63969=>"001011011",
  63970=>"000000000",
  63971=>"001001000",
  63972=>"000000000",
  63973=>"000000011",
  63974=>"111001000",
  63975=>"110111101",
  63976=>"001000000",
  63977=>"000000000",
  63978=>"000111111",
  63979=>"111111000",
  63980=>"100000011",
  63981=>"100100110",
  63982=>"111111111",
  63983=>"111011011",
  63984=>"000100111",
  63985=>"000100100",
  63986=>"000000110",
  63987=>"000000000",
  63988=>"000000000",
  63989=>"000000000",
  63990=>"111011000",
  63991=>"000000000",
  63992=>"000010011",
  63993=>"001111111",
  63994=>"100111111",
  63995=>"000001111",
  63996=>"100000000",
  63997=>"110100000",
  63998=>"000000111",
  63999=>"000111111",
  64000=>"111100100",
  64001=>"011000111",
  64002=>"111111111",
  64003=>"000111111",
  64004=>"011000001",
  64005=>"111111110",
  64006=>"111111000",
  64007=>"100100101",
  64008=>"000000000",
  64009=>"100000100",
  64010=>"011000000",
  64011=>"000101111",
  64012=>"000111111",
  64013=>"000111111",
  64014=>"000000011",
  64015=>"111000000",
  64016=>"001000101",
  64017=>"111110111",
  64018=>"111111000",
  64019=>"111100111",
  64020=>"000001001",
  64021=>"111111111",
  64022=>"000001000",
  64023=>"110110111",
  64024=>"111111010",
  64025=>"000110111",
  64026=>"010111111",
  64027=>"000000000",
  64028=>"111011001",
  64029=>"101000000",
  64030=>"010110100",
  64031=>"000000101",
  64032=>"001111111",
  64033=>"111111111",
  64034=>"111000000",
  64035=>"111111111",
  64036=>"000000000",
  64037=>"010100000",
  64038=>"011000000",
  64039=>"111111000",
  64040=>"001011011",
  64041=>"101000000",
  64042=>"011000101",
  64043=>"100000000",
  64044=>"111000000",
  64045=>"000010111",
  64046=>"000000000",
  64047=>"111111001",
  64048=>"011101001",
  64049=>"111111000",
  64050=>"000000000",
  64051=>"000111111",
  64052=>"000000000",
  64053=>"111111000",
  64054=>"111111111",
  64055=>"000100111",
  64056=>"000111000",
  64057=>"001000000",
  64058=>"000000000",
  64059=>"001101111",
  64060=>"011011000",
  64061=>"111100000",
  64062=>"110110110",
  64063=>"111110000",
  64064=>"000000111",
  64065=>"000100001",
  64066=>"000000000",
  64067=>"000000001",
  64068=>"111111001",
  64069=>"111111000",
  64070=>"111111111",
  64071=>"000000000",
  64072=>"001111011",
  64073=>"110111101",
  64074=>"011001000",
  64075=>"000000001",
  64076=>"000110111",
  64077=>"000000000",
  64078=>"111000000",
  64079=>"000000000",
  64080=>"000000000",
  64081=>"111111000",
  64082=>"001001111",
  64083=>"000111111",
  64084=>"111000000",
  64085=>"100000000",
  64086=>"000000000",
  64087=>"101100000",
  64088=>"000111011",
  64089=>"111111101",
  64090=>"000000000",
  64091=>"111001011",
  64092=>"111111111",
  64093=>"001001001",
  64094=>"000000100",
  64095=>"111111110",
  64096=>"110111000",
  64097=>"000000000",
  64098=>"001011111",
  64099=>"111000000",
  64100=>"001001000",
  64101=>"000000111",
  64102=>"000100111",
  64103=>"100000111",
  64104=>"011000000",
  64105=>"000111111",
  64106=>"000000011",
  64107=>"001111111",
  64108=>"111111111",
  64109=>"111000010",
  64110=>"111111101",
  64111=>"111111001",
  64112=>"000000000",
  64113=>"000100100",
  64114=>"010001000",
  64115=>"010111111",
  64116=>"111000000",
  64117=>"011011111",
  64118=>"111111000",
  64119=>"110100000",
  64120=>"000000000",
  64121=>"111111101",
  64122=>"000000000",
  64123=>"101000000",
  64124=>"000000110",
  64125=>"000111111",
  64126=>"110111111",
  64127=>"000000111",
  64128=>"111111111",
  64129=>"000010101",
  64130=>"000000000",
  64131=>"000100111",
  64132=>"000000000",
  64133=>"101101111",
  64134=>"001111000",
  64135=>"111011011",
  64136=>"000000011",
  64137=>"111000100",
  64138=>"010101000",
  64139=>"000000001",
  64140=>"000001111",
  64141=>"000000000",
  64142=>"111111111",
  64143=>"000000000",
  64144=>"000000011",
  64145=>"000110111",
  64146=>"000000000",
  64147=>"000000011",
  64148=>"010110111",
  64149=>"000001111",
  64150=>"011111100",
  64151=>"001000011",
  64152=>"101000000",
  64153=>"000000000",
  64154=>"111000000",
  64155=>"000000011",
  64156=>"001001000",
  64157=>"000111111",
  64158=>"000000111",
  64159=>"111110000",
  64160=>"001111101",
  64161=>"000000111",
  64162=>"110110010",
  64163=>"111111111",
  64164=>"111111000",
  64165=>"110110001",
  64166=>"000000000",
  64167=>"000000000",
  64168=>"100110011",
  64169=>"111111011",
  64170=>"000111111",
  64171=>"000110110",
  64172=>"011111101",
  64173=>"101111111",
  64174=>"111000000",
  64175=>"101111110",
  64176=>"000000111",
  64177=>"111111101",
  64178=>"010111111",
  64179=>"111111000",
  64180=>"110000100",
  64181=>"000000000",
  64182=>"011011000",
  64183=>"100110000",
  64184=>"001111111",
  64185=>"000111000",
  64186=>"111011100",
  64187=>"000000001",
  64188=>"011000000",
  64189=>"111000000",
  64190=>"111111101",
  64191=>"111111111",
  64192=>"000000000",
  64193=>"111000000",
  64194=>"000000111",
  64195=>"111111000",
  64196=>"100000110",
  64197=>"000111111",
  64198=>"000000000",
  64199=>"000000111",
  64200=>"000000001",
  64201=>"111111000",
  64202=>"000000111",
  64203=>"111111010",
  64204=>"000000111",
  64205=>"110000000",
  64206=>"111111111",
  64207=>"111110000",
  64208=>"110111111",
  64209=>"000000110",
  64210=>"001000111",
  64211=>"100110111",
  64212=>"000000000",
  64213=>"111110110",
  64214=>"111000000",
  64215=>"000000111",
  64216=>"111110110",
  64217=>"111011111",
  64218=>"000110111",
  64219=>"111101001",
  64220=>"000000000",
  64221=>"000110111",
  64222=>"110111111",
  64223=>"000000101",
  64224=>"110000010",
  64225=>"111111111",
  64226=>"011101001",
  64227=>"111111001",
  64228=>"010000000",
  64229=>"111101111",
  64230=>"100000000",
  64231=>"000011111",
  64232=>"000111111",
  64233=>"111111111",
  64234=>"000000000",
  64235=>"000100100",
  64236=>"011000000",
  64237=>"111000000",
  64238=>"111000000",
  64239=>"010000000",
  64240=>"011001111",
  64241=>"000111110",
  64242=>"000000111",
  64243=>"100101000",
  64244=>"001111111",
  64245=>"011111111",
  64246=>"111011000",
  64247=>"000000111",
  64248=>"000001100",
  64249=>"111001001",
  64250=>"000000000",
  64251=>"110111111",
  64252=>"000000001",
  64253=>"111100000",
  64254=>"000000001",
  64255=>"111111111",
  64256=>"111111100",
  64257=>"011001001",
  64258=>"110000111",
  64259=>"111111111",
  64260=>"111000000",
  64261=>"000100110",
  64262=>"111101101",
  64263=>"000000000",
  64264=>"000100011",
  64265=>"000000000",
  64266=>"001000011",
  64267=>"000000111",
  64268=>"100100000",
  64269=>"000111000",
  64270=>"111111111",
  64271=>"010000111",
  64272=>"000000000",
  64273=>"001101111",
  64274=>"000000110",
  64275=>"100000010",
  64276=>"111000001",
  64277=>"001001111",
  64278=>"000011111",
  64279=>"111111000",
  64280=>"000000110",
  64281=>"000000000",
  64282=>"010111000",
  64283=>"110000111",
  64284=>"000000110",
  64285=>"000000000",
  64286=>"111111100",
  64287=>"111111111",
  64288=>"100111111",
  64289=>"000110110",
  64290=>"000111111",
  64291=>"000000011",
  64292=>"110111111",
  64293=>"000111111",
  64294=>"001111111",
  64295=>"000000000",
  64296=>"111111000",
  64297=>"111001000",
  64298=>"000011111",
  64299=>"000000000",
  64300=>"000000000",
  64301=>"000001111",
  64302=>"000000000",
  64303=>"000000111",
  64304=>"000101111",
  64305=>"000000000",
  64306=>"111111110",
  64307=>"111111111",
  64308=>"111111000",
  64309=>"000110111",
  64310=>"000000000",
  64311=>"000000111",
  64312=>"111111010",
  64313=>"111001000",
  64314=>"111000000",
  64315=>"111111111",
  64316=>"110110100",
  64317=>"100010000",
  64318=>"011111110",
  64319=>"000000000",
  64320=>"000111011",
  64321=>"111111111",
  64322=>"000000111",
  64323=>"000000000",
  64324=>"000100000",
  64325=>"000000000",
  64326=>"111000000",
  64327=>"111100000",
  64328=>"011111111",
  64329=>"111111101",
  64330=>"111111111",
  64331=>"011011111",
  64332=>"000000111",
  64333=>"000000000",
  64334=>"000000111",
  64335=>"111101000",
  64336=>"011111111",
  64337=>"100000100",
  64338=>"111111111",
  64339=>"001000000",
  64340=>"110111111",
  64341=>"000000001",
  64342=>"000111111",
  64343=>"000000000",
  64344=>"111111000",
  64345=>"000000001",
  64346=>"111001000",
  64347=>"111000000",
  64348=>"111100111",
  64349=>"100100100",
  64350=>"000000001",
  64351=>"010000000",
  64352=>"100111111",
  64353=>"000000111",
  64354=>"100001011",
  64355=>"000100011",
  64356=>"111111110",
  64357=>"000000111",
  64358=>"000000111",
  64359=>"011011000",
  64360=>"100000000",
  64361=>"101001111",
  64362=>"000000111",
  64363=>"000000111",
  64364=>"011001111",
  64365=>"111000100",
  64366=>"000000000",
  64367=>"011000000",
  64368=>"000000100",
  64369=>"000011000",
  64370=>"101111111",
  64371=>"100001000",
  64372=>"111111111",
  64373=>"111011000",
  64374=>"000000000",
  64375=>"000001111",
  64376=>"111100000",
  64377=>"011010111",
  64378=>"111111111",
  64379=>"011111111",
  64380=>"011111111",
  64381=>"111001001",
  64382=>"000000101",
  64383=>"111000000",
  64384=>"011101001",
  64385=>"100111111",
  64386=>"100100000",
  64387=>"111111111",
  64388=>"000000000",
  64389=>"111100100",
  64390=>"010000110",
  64391=>"110111011",
  64392=>"111110000",
  64393=>"111000000",
  64394=>"011000000",
  64395=>"100110111",
  64396=>"110111111",
  64397=>"000000000",
  64398=>"111111000",
  64399=>"100100000",
  64400=>"111111111",
  64401=>"111011000",
  64402=>"000110111",
  64403=>"111111000",
  64404=>"111111111",
  64405=>"110010000",
  64406=>"010111111",
  64407=>"011000000",
  64408=>"110111111",
  64409=>"000011011",
  64410=>"100011000",
  64411=>"000001111",
  64412=>"000001111",
  64413=>"000000000",
  64414=>"111000000",
  64415=>"100111110",
  64416=>"000000000",
  64417=>"000000110",
  64418=>"000101111",
  64419=>"100100000",
  64420=>"111101000",
  64421=>"000111011",
  64422=>"000000001",
  64423=>"000111110",
  64424=>"110000000",
  64425=>"000111111",
  64426=>"111111011",
  64427=>"011010000",
  64428=>"000000111",
  64429=>"000000000",
  64430=>"000001000",
  64431=>"000010000",
  64432=>"000000000",
  64433=>"111111001",
  64434=>"000110111",
  64435=>"111001011",
  64436=>"000000111",
  64437=>"110000000",
  64438=>"111111000",
  64439=>"111111111",
  64440=>"000111011",
  64441=>"011111111",
  64442=>"011000111",
  64443=>"000001001",
  64444=>"111111011",
  64445=>"111111000",
  64446=>"000010011",
  64447=>"111100010",
  64448=>"000111111",
  64449=>"111100111",
  64450=>"110111000",
  64451=>"111111111",
  64452=>"111111111",
  64453=>"000000001",
  64454=>"000000111",
  64455=>"000000000",
  64456=>"100100000",
  64457=>"111000000",
  64458=>"000011111",
  64459=>"010111000",
  64460=>"110111010",
  64461=>"001111111",
  64462=>"101110111",
  64463=>"000000100",
  64464=>"111101000",
  64465=>"001100100",
  64466=>"111111111",
  64467=>"000011111",
  64468=>"111111011",
  64469=>"111110000",
  64470=>"000100111",
  64471=>"110111111",
  64472=>"000000000",
  64473=>"000000000",
  64474=>"111111111",
  64475=>"000000110",
  64476=>"000000111",
  64477=>"000000011",
  64478=>"100111111",
  64479=>"011011000",
  64480=>"100000111",
  64481=>"000001100",
  64482=>"111111010",
  64483=>"011000000",
  64484=>"000000101",
  64485=>"111111001",
  64486=>"111111111",
  64487=>"110000000",
  64488=>"000110111",
  64489=>"111111101",
  64490=>"000001001",
  64491=>"100110110",
  64492=>"011000101",
  64493=>"111111111",
  64494=>"111111111",
  64495=>"111001000",
  64496=>"111000000",
  64497=>"111111101",
  64498=>"001011110",
  64499=>"000000111",
  64500=>"111111011",
  64501=>"110000000",
  64502=>"001000111",
  64503=>"001001000",
  64504=>"000000011",
  64505=>"001001110",
  64506=>"111111101",
  64507=>"110110111",
  64508=>"001000011",
  64509=>"000001101",
  64510=>"000000111",
  64511=>"100000100",
  64512=>"000000000",
  64513=>"000110111",
  64514=>"000000111",
  64515=>"111000000",
  64516=>"000000000",
  64517=>"110100000",
  64518=>"000000111",
  64519=>"111111111",
  64520=>"111100110",
  64521=>"000110000",
  64522=>"011100111",
  64523=>"111110010",
  64524=>"000000100",
  64525=>"111001000",
  64526=>"100000000",
  64527=>"000111110",
  64528=>"010001000",
  64529=>"111111110",
  64530=>"000000111",
  64531=>"000000000",
  64532=>"000000000",
  64533=>"111000000",
  64534=>"101111100",
  64535=>"100001001",
  64536=>"111111011",
  64537=>"000111000",
  64538=>"000000000",
  64539=>"111100101",
  64540=>"000000001",
  64541=>"111111111",
  64542=>"000110111",
  64543=>"000000111",
  64544=>"000000000",
  64545=>"111111100",
  64546=>"000000000",
  64547=>"111111111",
  64548=>"111111111",
  64549=>"111111111",
  64550=>"101100000",
  64551=>"000101111",
  64552=>"001011000",
  64553=>"000000001",
  64554=>"111111000",
  64555=>"111111110",
  64556=>"111000000",
  64557=>"111000000",
  64558=>"000000011",
  64559=>"011010010",
  64560=>"111111111",
  64561=>"000010000",
  64562=>"000000000",
  64563=>"111111000",
  64564=>"000000110",
  64565=>"000110111",
  64566=>"000111111",
  64567=>"000000000",
  64568=>"111000000",
  64569=>"000000000",
  64570=>"000000000",
  64571=>"111111111",
  64572=>"000100111",
  64573=>"000111111",
  64574=>"100110111",
  64575=>"111101000",
  64576=>"110000000",
  64577=>"111011000",
  64578=>"111111111",
  64579=>"110111111",
  64580=>"000000010",
  64581=>"111110110",
  64582=>"000110110",
  64583=>"000000000",
  64584=>"111111011",
  64585=>"000000101",
  64586=>"100111000",
  64587=>"111011011",
  64588=>"111111111",
  64589=>"001101110",
  64590=>"000000000",
  64591=>"111111111",
  64592=>"111111000",
  64593=>"001110000",
  64594=>"000110111",
  64595=>"000000010",
  64596=>"000000000",
  64597=>"100000100",
  64598=>"111100000",
  64599=>"111001101",
  64600=>"111000000",
  64601=>"100110000",
  64602=>"000000111",
  64603=>"011001000",
  64604=>"000000000",
  64605=>"111100000",
  64606=>"000111111",
  64607=>"100100101",
  64608=>"000110000",
  64609=>"001000000",
  64610=>"111111111",
  64611=>"000110110",
  64612=>"000000000",
  64613=>"000011111",
  64614=>"000000000",
  64615=>"101111111",
  64616=>"111111000",
  64617=>"000000000",
  64618=>"111111000",
  64619=>"000001011",
  64620=>"111111111",
  64621=>"000000000",
  64622=>"111111001",
  64623=>"111111111",
  64624=>"111110000",
  64625=>"110111111",
  64626=>"001001000",
  64627=>"000001000",
  64628=>"111111100",
  64629=>"000000000",
  64630=>"110010000",
  64631=>"000000001",
  64632=>"000000000",
  64633=>"111101000",
  64634=>"010011000",
  64635=>"000000000",
  64636=>"111111111",
  64637=>"110110000",
  64638=>"001000000",
  64639=>"000000100",
  64640=>"111111100",
  64641=>"000100111",
  64642=>"000000111",
  64643=>"000000000",
  64644=>"111111111",
  64645=>"000101111",
  64646=>"110111100",
  64647=>"000000111",
  64648=>"000001111",
  64649=>"110000000",
  64650=>"000001111",
  64651=>"000000000",
  64652=>"100100111",
  64653=>"111111010",
  64654=>"000000000",
  64655=>"000000000",
  64656=>"111111111",
  64657=>"111110000",
  64658=>"111110110",
  64659=>"110000001",
  64660=>"111000000",
  64661=>"111111000",
  64662=>"111111001",
  64663=>"111111110",
  64664=>"000100000",
  64665=>"001111111",
  64666=>"111001000",
  64667=>"000011000",
  64668=>"100111111",
  64669=>"110110010",
  64670=>"111001111",
  64671=>"001000111",
  64672=>"110000000",
  64673=>"000000100",
  64674=>"110100110",
  64675=>"101111100",
  64676=>"000011000",
  64677=>"110111111",
  64678=>"111111111",
  64679=>"111111110",
  64680=>"001001001",
  64681=>"111010110",
  64682=>"111111100",
  64683=>"111110000",
  64684=>"001000000",
  64685=>"110111111",
  64686=>"111111000",
  64687=>"100000000",
  64688=>"000000100",
  64689=>"101111111",
  64690=>"111111111",
  64691=>"000000000",
  64692=>"000000000",
  64693=>"110010000",
  64694=>"111101111",
  64695=>"000100100",
  64696=>"111111011",
  64697=>"000000001",
  64698=>"000001111",
  64699=>"000000000",
  64700=>"100100000",
  64701=>"111000000",
  64702=>"000000000",
  64703=>"111001001",
  64704=>"111000000",
  64705=>"000111111",
  64706=>"000000001",
  64707=>"111111111",
  64708=>"101101111",
  64709=>"111000111",
  64710=>"000010000",
  64711=>"011111111",
  64712=>"000000000",
  64713=>"011001100",
  64714=>"111111111",
  64715=>"000000100",
  64716=>"111011001",
  64717=>"111111000",
  64718=>"000111111",
  64719=>"010100000",
  64720=>"011011111",
  64721=>"110000000",
  64722=>"111010000",
  64723=>"001001111",
  64724=>"000010000",
  64725=>"110000000",
  64726=>"111000000",
  64727=>"110110000",
  64728=>"000000100",
  64729=>"111110011",
  64730=>"000011111",
  64731=>"110000000",
  64732=>"001001000",
  64733=>"111001000",
  64734=>"000000000",
  64735=>"111111111",
  64736=>"111000000",
  64737=>"101000000",
  64738=>"100100111",
  64739=>"000000000",
  64740=>"011011110",
  64741=>"000110110",
  64742=>"000000000",
  64743=>"111111111",
  64744=>"111111011",
  64745=>"111111111",
  64746=>"101001111",
  64747=>"111000000",
  64748=>"000011011",
  64749=>"111111000",
  64750=>"000000000",
  64751=>"001000000",
  64752=>"001000000",
  64753=>"000111010",
  64754=>"100001111",
  64755=>"101000111",
  64756=>"100000000",
  64757=>"001001011",
  64758=>"000111111",
  64759=>"111111111",
  64760=>"000000000",
  64761=>"111111011",
  64762=>"010000100",
  64763=>"000000111",
  64764=>"011000001",
  64765=>"011111111",
  64766=>"000000000",
  64767=>"001111111",
  64768=>"000111111",
  64769=>"011000000",
  64770=>"111000000",
  64771=>"111111000",
  64772=>"000000000",
  64773=>"111001001",
  64774=>"111111111",
  64775=>"000001111",
  64776=>"111111111",
  64777=>"111000000",
  64778=>"000000001",
  64779=>"000000000",
  64780=>"000011111",
  64781=>"001000000",
  64782=>"000000111",
  64783=>"110100000",
  64784=>"100000000",
  64785=>"000000000",
  64786=>"000000000",
  64787=>"011111111",
  64788=>"000111111",
  64789=>"000000111",
  64790=>"001011011",
  64791=>"001100100",
  64792=>"110110110",
  64793=>"111111000",
  64794=>"100110111",
  64795=>"000000000",
  64796=>"111111111",
  64797=>"001000111",
  64798=>"111111111",
  64799=>"101000000",
  64800=>"111100011",
  64801=>"000011011",
  64802=>"111111110",
  64803=>"111111000",
  64804=>"001111101",
  64805=>"111111111",
  64806=>"100101000",
  64807=>"010000000",
  64808=>"000001011",
  64809=>"000000111",
  64810=>"100100101",
  64811=>"100111111",
  64812=>"111111111",
  64813=>"000111000",
  64814=>"000111000",
  64815=>"000101111",
  64816=>"111111111",
  64817=>"000111111",
  64818=>"111111111",
  64819=>"000000011",
  64820=>"011111111",
  64821=>"000000001",
  64822=>"111100000",
  64823=>"100100111",
  64824=>"000110100",
  64825=>"111111001",
  64826=>"000000000",
  64827=>"110000000",
  64828=>"111111100",
  64829=>"111111000",
  64830=>"111000000",
  64831=>"001111111",
  64832=>"010000000",
  64833=>"000100000",
  64834=>"100111111",
  64835=>"000001001",
  64836=>"111111010",
  64837=>"111000000",
  64838=>"000000000",
  64839=>"000000000",
  64840=>"111000100",
  64841=>"111000100",
  64842=>"000100000",
  64843=>"110111111",
  64844=>"010000000",
  64845=>"100000000",
  64846=>"110110101",
  64847=>"100001001",
  64848=>"101100111",
  64849=>"000000000",
  64850=>"011111000",
  64851=>"111110111",
  64852=>"111000000",
  64853=>"001111111",
  64854=>"111111000",
  64855=>"111100110",
  64856=>"001001111",
  64857=>"000110111",
  64858=>"000000000",
  64859=>"011111111",
  64860=>"000000000",
  64861=>"000000100",
  64862=>"000000000",
  64863=>"111111111",
  64864=>"000000000",
  64865=>"001000000",
  64866=>"000010111",
  64867=>"111000000",
  64868=>"111111111",
  64869=>"000000000",
  64870=>"110000000",
  64871=>"000111111",
  64872=>"010111111",
  64873=>"110111111",
  64874=>"000111111",
  64875=>"001001001",
  64876=>"000111011",
  64877=>"000111111",
  64878=>"000000000",
  64879=>"000000000",
  64880=>"111111111",
  64881=>"000101010",
  64882=>"111011000",
  64883=>"111001000",
  64884=>"111111111",
  64885=>"111111100",
  64886=>"000000011",
  64887=>"110101111",
  64888=>"000000011",
  64889=>"111000000",
  64890=>"000000000",
  64891=>"110000011",
  64892=>"110111111",
  64893=>"000000000",
  64894=>"111000010",
  64895=>"111000011",
  64896=>"111100110",
  64897=>"111000111",
  64898=>"111111111",
  64899=>"000000000",
  64900=>"000100111",
  64901=>"110000111",
  64902=>"000000000",
  64903=>"001000000",
  64904=>"000000000",
  64905=>"001111111",
  64906=>"000000000",
  64907=>"001011111",
  64908=>"100110111",
  64909=>"000111111",
  64910=>"001001001",
  64911=>"000000000",
  64912=>"000000100",
  64913=>"111101111",
  64914=>"110110000",
  64915=>"111011011",
  64916=>"000011000",
  64917=>"000000000",
  64918=>"100000000",
  64919=>"100111011",
  64920=>"111111111",
  64921=>"000000000",
  64922=>"011000000",
  64923=>"100111111",
  64924=>"110010010",
  64925=>"111111111",
  64926=>"000000000",
  64927=>"111011111",
  64928=>"111101111",
  64929=>"000000000",
  64930=>"000001000",
  64931=>"111100000",
  64932=>"111111001",
  64933=>"110111000",
  64934=>"000000000",
  64935=>"000111111",
  64936=>"000000110",
  64937=>"110111111",
  64938=>"111001011",
  64939=>"000000000",
  64940=>"010100111",
  64941=>"111000000",
  64942=>"111111100",
  64943=>"100000000",
  64944=>"000111111",
  64945=>"111111111",
  64946=>"000000000",
  64947=>"111111110",
  64948=>"010111111",
  64949=>"111111011",
  64950=>"111111000",
  64951=>"111000000",
  64952=>"111000000",
  64953=>"111001000",
  64954=>"000000110",
  64955=>"111111001",
  64956=>"011111111",
  64957=>"001000000",
  64958=>"000000000",
  64959=>"111111001",
  64960=>"000101000",
  64961=>"011001000",
  64962=>"111110110",
  64963=>"111111100",
  64964=>"111111111",
  64965=>"000000000",
  64966=>"010000000",
  64967=>"001011011",
  64968=>"000011111",
  64969=>"000000111",
  64970=>"111100000",
  64971=>"111111000",
  64972=>"000000110",
  64973=>"111111111",
  64974=>"000110111",
  64975=>"000000000",
  64976=>"000010111",
  64977=>"111000000",
  64978=>"000000000",
  64979=>"110111111",
  64980=>"000110111",
  64981=>"111111000",
  64982=>"000101111",
  64983=>"001011001",
  64984=>"000000000",
  64985=>"000000110",
  64986=>"000000000",
  64987=>"000000000",
  64988=>"111011011",
  64989=>"111111000",
  64990=>"111111000",
  64991=>"000001011",
  64992=>"000000000",
  64993=>"000111111",
  64994=>"111110111",
  64995=>"111011000",
  64996=>"111111111",
  64997=>"010000000",
  64998=>"111111000",
  64999=>"111111111",
  65000=>"100000000",
  65001=>"111000000",
  65002=>"000000000",
  65003=>"000000000",
  65004=>"000000111",
  65005=>"011111100",
  65006=>"000000000",
  65007=>"000010111",
  65008=>"000000000",
  65009=>"111111111",
  65010=>"100000001",
  65011=>"010111111",
  65012=>"111100000",
  65013=>"100010010",
  65014=>"110110111",
  65015=>"000000000",
  65016=>"000111111",
  65017=>"010111110",
  65018=>"100000000",
  65019=>"111111110",
  65020=>"000000000",
  65021=>"111011001",
  65022=>"101111111",
  65023=>"110000000",
  65024=>"111111111",
  65025=>"000000101",
  65026=>"111111111",
  65027=>"110000000",
  65028=>"011001001",
  65029=>"000000111",
  65030=>"100000000",
  65031=>"111111111",
  65032=>"000111111",
  65033=>"111111001",
  65034=>"111111110",
  65035=>"111111111",
  65036=>"000000110",
  65037=>"110110111",
  65038=>"100100100",
  65039=>"000111111",
  65040=>"110110111",
  65041=>"111111000",
  65042=>"111111111",
  65043=>"110000000",
  65044=>"110111111",
  65045=>"000100110",
  65046=>"000000111",
  65047=>"011010111",
  65048=>"111001001",
  65049=>"011011000",
  65050=>"000000000",
  65051=>"010000100",
  65052=>"000001011",
  65053=>"110000111",
  65054=>"110100110",
  65055=>"111111111",
  65056=>"111111111",
  65057=>"111110110",
  65058=>"111111111",
  65059=>"111111000",
  65060=>"000000000",
  65061=>"111111110",
  65062=>"011010010",
  65063=>"000110111",
  65064=>"111111111",
  65065=>"000000000",
  65066=>"000110100",
  65067=>"001111111",
  65068=>"110110010",
  65069=>"111111000",
  65070=>"111111011",
  65071=>"000001000",
  65072=>"000111111",
  65073=>"111111110",
  65074=>"111001001",
  65075=>"000000111",
  65076=>"111000111",
  65077=>"111101000",
  65078=>"100001101",
  65079=>"000000000",
  65080=>"001000000",
  65081=>"000000000",
  65082=>"000100100",
  65083=>"111101111",
  65084=>"111111001",
  65085=>"111001000",
  65086=>"111111011",
  65087=>"001000000",
  65088=>"111111111",
  65089=>"000000000",
  65090=>"001000110",
  65091=>"000110111",
  65092=>"000100100",
  65093=>"111011000",
  65094=>"000000000",
  65095=>"000010011",
  65096=>"000000000",
  65097=>"000000000",
  65098=>"111111111",
  65099=>"001001000",
  65100=>"000000000",
  65101=>"110000000",
  65102=>"101100011",
  65103=>"000111011",
  65104=>"110111111",
  65105=>"111101001",
  65106=>"111111000",
  65107=>"111101110",
  65108=>"111111000",
  65109=>"000000111",
  65110=>"000011000",
  65111=>"111111101",
  65112=>"000100111",
  65113=>"001111111",
  65114=>"000001001",
  65115=>"100100110",
  65116=>"000001111",
  65117=>"000111111",
  65118=>"001111101",
  65119=>"001000011",
  65120=>"000000001",
  65121=>"000110000",
  65122=>"111000111",
  65123=>"111001001",
  65124=>"111111111",
  65125=>"111111100",
  65126=>"111111000",
  65127=>"111000000",
  65128=>"111111111",
  65129=>"000000111",
  65130=>"000010000",
  65131=>"010010011",
  65132=>"011011111",
  65133=>"000000001",
  65134=>"111111001",
  65135=>"000010110",
  65136=>"000000111",
  65137=>"000000000",
  65138=>"100111001",
  65139=>"101111111",
  65140=>"001011001",
  65141=>"100000110",
  65142=>"001001001",
  65143=>"101111111",
  65144=>"100101100",
  65145=>"110111111",
  65146=>"111000000",
  65147=>"111111111",
  65148=>"101111111",
  65149=>"000111000",
  65150=>"111111111",
  65151=>"000001001",
  65152=>"111111000",
  65153=>"000100000",
  65154=>"000000000",
  65155=>"100111111",
  65156=>"000111111",
  65157=>"111100110",
  65158=>"111111111",
  65159=>"000010111",
  65160=>"111111111",
  65161=>"111000111",
  65162=>"111111111",
  65163=>"111111111",
  65164=>"001001011",
  65165=>"111111111",
  65166=>"001000000",
  65167=>"110000000",
  65168=>"000001111",
  65169=>"001111111",
  65170=>"000000000",
  65171=>"111111111",
  65172=>"111111111",
  65173=>"000000100",
  65174=>"111111111",
  65175=>"000000000",
  65176=>"000000000",
  65177=>"111101000",
  65178=>"000000000",
  65179=>"111111111",
  65180=>"000000111",
  65181=>"111111111",
  65182=>"000000101",
  65183=>"010011000",
  65184=>"000000011",
  65185=>"000101111",
  65186=>"000000000",
  65187=>"000000000",
  65188=>"111000000",
  65189=>"000000101",
  65190=>"111001000",
  65191=>"111111000",
  65192=>"000000000",
  65193=>"001011111",
  65194=>"100111100",
  65195=>"000000000",
  65196=>"000101000",
  65197=>"100111111",
  65198=>"000000011",
  65199=>"100111111",
  65200=>"000000110",
  65201=>"000000000",
  65202=>"100100111",
  65203=>"111111111",
  65204=>"000010111",
  65205=>"000111010",
  65206=>"000000111",
  65207=>"111100000",
  65208=>"100000011",
  65209=>"110110100",
  65210=>"111000000",
  65211=>"000010111",
  65212=>"111111111",
  65213=>"001111111",
  65214=>"010011111",
  65215=>"000000000",
  65216=>"111101111",
  65217=>"100000111",
  65218=>"000000111",
  65219=>"011111111",
  65220=>"000000100",
  65221=>"000000001",
  65222=>"110100000",
  65223=>"111001100",
  65224=>"000000010",
  65225=>"001000000",
  65226=>"001000111",
  65227=>"111100000",
  65228=>"000111111",
  65229=>"000010000",
  65230=>"000000111",
  65231=>"000100100",
  65232=>"000111111",
  65233=>"000000000",
  65234=>"111111111",
  65235=>"010000000",
  65236=>"111111000",
  65237=>"111110110",
  65238=>"111000000",
  65239=>"000111111",
  65240=>"110000000",
  65241=>"001010000",
  65242=>"000000000",
  65243=>"000000001",
  65244=>"000000000",
  65245=>"000111111",
  65246=>"001000111",
  65247=>"000000000",
  65248=>"000000111",
  65249=>"010010010",
  65250=>"000011111",
  65251=>"111111111",
  65252=>"000000000",
  65253=>"000000011",
  65254=>"000000000",
  65255=>"111111000",
  65256=>"101000000",
  65257=>"111001001",
  65258=>"111000111",
  65259=>"111111111",
  65260=>"111111010",
  65261=>"111000111",
  65262=>"000000001",
  65263=>"100110111",
  65264=>"100110100",
  65265=>"011010000",
  65266=>"000010000",
  65267=>"000000000",
  65268=>"110100110",
  65269=>"101101100",
  65270=>"000000001",
  65271=>"101100111",
  65272=>"110000111",
  65273=>"000111111",
  65274=>"000000000",
  65275=>"000110110",
  65276=>"111111111",
  65277=>"000000000",
  65278=>"100000000",
  65279=>"111111000",
  65280=>"011111111",
  65281=>"111110100",
  65282=>"111000100",
  65283=>"000000000",
  65284=>"000000000",
  65285=>"110111111",
  65286=>"111101000",
  65287=>"000000111",
  65288=>"001001000",
  65289=>"111111111",
  65290=>"111111111",
  65291=>"000000000",
  65292=>"111110111",
  65293=>"011001001",
  65294=>"111011011",
  65295=>"000000000",
  65296=>"110100111",
  65297=>"000000001",
  65298=>"100111111",
  65299=>"100000000",
  65300=>"110000111",
  65301=>"000001111",
  65302=>"111000100",
  65303=>"100100111",
  65304=>"111111111",
  65305=>"000000000",
  65306=>"111111000",
  65307=>"000000111",
  65308=>"000000000",
  65309=>"000000000",
  65310=>"000100100",
  65311=>"000000111",
  65312=>"100111011",
  65313=>"000000000",
  65314=>"000001011",
  65315=>"101111111",
  65316=>"100000000",
  65317=>"100000111",
  65318=>"111000100",
  65319=>"000000111",
  65320=>"111111111",
  65321=>"000000000",
  65322=>"001000010",
  65323=>"000000000",
  65324=>"000111011",
  65325=>"001100101",
  65326=>"001001111",
  65327=>"111111111",
  65328=>"100000110",
  65329=>"010000000",
  65330=>"000000110",
  65331=>"111111111",
  65332=>"011111111",
  65333=>"011111111",
  65334=>"000000000",
  65335=>"000000111",
  65336=>"111101100",
  65337=>"000000000",
  65338=>"000000000",
  65339=>"100100111",
  65340=>"000000010",
  65341=>"000000100",
  65342=>"000100110",
  65343=>"111001111",
  65344=>"001000100",
  65345=>"110000111",
  65346=>"000000000",
  65347=>"111111111",
  65348=>"111001000",
  65349=>"111001110",
  65350=>"100100000",
  65351=>"111001001",
  65352=>"111100000",
  65353=>"111000111",
  65354=>"111111111",
  65355=>"000000010",
  65356=>"000110110",
  65357=>"000100100",
  65358=>"000000000",
  65359=>"111111000",
  65360=>"111111111",
  65361=>"100110110",
  65362=>"111111111",
  65363=>"111100100",
  65364=>"111111110",
  65365=>"001001011",
  65366=>"111111111",
  65367=>"001001000",
  65368=>"000000111",
  65369=>"000000111",
  65370=>"111111111",
  65371=>"111001001",
  65372=>"000100000",
  65373=>"111111100",
  65374=>"111111111",
  65375=>"000000000",
  65376=>"111111111",
  65377=>"111001000",
  65378=>"001011011",
  65379=>"110001001",
  65380=>"001101011",
  65381=>"110000000",
  65382=>"010000111",
  65383=>"111000000",
  65384=>"001000100",
  65385=>"001000001",
  65386=>"111111111",
  65387=>"111001001",
  65388=>"011011111",
  65389=>"000111000",
  65390=>"000000000",
  65391=>"000000001",
  65392=>"001111111",
  65393=>"110110000",
  65394=>"111000000",
  65395=>"000000000",
  65396=>"000010010",
  65397=>"011111111",
  65398=>"000110110",
  65399=>"111000000",
  65400=>"111001000",
  65401=>"000000000",
  65402=>"111111111",
  65403=>"111000000",
  65404=>"110111001",
  65405=>"111111101",
  65406=>"100111111",
  65407=>"000000000",
  65408=>"101111111",
  65409=>"100000000",
  65410=>"111101000",
  65411=>"010000000",
  65412=>"110111111",
  65413=>"000000000",
  65414=>"000000010",
  65415=>"000000110",
  65416=>"111111000",
  65417=>"001111001",
  65418=>"000000111",
  65419=>"000000000",
  65420=>"111111111",
  65421=>"000000000",
  65422=>"101000000",
  65423=>"011010010",
  65424=>"000000000",
  65425=>"111111111",
  65426=>"100100100",
  65427=>"001011001",
  65428=>"001001111",
  65429=>"000000000",
  65430=>"111110110",
  65431=>"001000000",
  65432=>"000000000",
  65433=>"100000000",
  65434=>"100111000",
  65435=>"111101001",
  65436=>"111111101",
  65437=>"001010110",
  65438=>"111111000",
  65439=>"000000000",
  65440=>"010111111",
  65441=>"001011001",
  65442=>"000000000",
  65443=>"000000000",
  65444=>"001111111",
  65445=>"000001111",
  65446=>"111000001",
  65447=>"000000111",
  65448=>"100101111",
  65449=>"000000000",
  65450=>"111111100",
  65451=>"011000000",
  65452=>"011000000",
  65453=>"000000111",
  65454=>"001111101",
  65455=>"000000000",
  65456=>"000111111",
  65457=>"111000000",
  65458=>"110110000",
  65459=>"000010000",
  65460=>"011000010",
  65461=>"111111111",
  65462=>"001000000",
  65463=>"011111111",
  65464=>"000000000",
  65465=>"100100110",
  65466=>"000000001",
  65467=>"111110110",
  65468=>"000000000",
  65469=>"111111111",
  65470=>"111000000",
  65471=>"110110000",
  65472=>"001000000",
  65473=>"011000000",
  65474=>"000000111",
  65475=>"000011011",
  65476=>"000000000",
  65477=>"001011010",
  65478=>"000000000",
  65479=>"111101000",
  65480=>"000000000",
  65481=>"111111111",
  65482=>"000001011",
  65483=>"111110111",
  65484=>"000000111",
  65485=>"000111111",
  65486=>"101001000",
  65487=>"000010110",
  65488=>"011000000",
  65489=>"000000100",
  65490=>"110100110",
  65491=>"111111111",
  65492=>"101101011",
  65493=>"000000111",
  65494=>"000000100",
  65495=>"000001111",
  65496=>"000111111",
  65497=>"110100111",
  65498=>"001000110",
  65499=>"001000000",
  65500=>"111111111",
  65501=>"000000111",
  65502=>"111001111",
  65503=>"000111111",
  65504=>"000000000",
  65505=>"111001000",
  65506=>"000000111",
  65507=>"101111001",
  65508=>"111111111",
  65509=>"000111000",
  65510=>"001000110",
  65511=>"111000000",
  65512=>"111111111",
  65513=>"111111111",
  65514=>"000000000",
  65515=>"111000111",
  65516=>"000000110",
  65517=>"001000000",
  65518=>"111111111",
  65519=>"111000010",
  65520=>"111111110",
  65521=>"000001111",
  65522=>"111101111",
  65523=>"000001101",
  65524=>"000100100",
  65525=>"000000000",
  65526=>"111111111",
  65527=>"000101111",
  65528=>"000111111",
  65529=>"111100100",
  65530=>"001111111",
  65531=>"000000000",
  65532=>"010000100",
  65533=>"001111111",
  65534=>"110111111",
  65535=>"000000000");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;